module rompcm352(
	input clk,//45m
	input reset_n,
	output signed [31:0]addrout
);

wire signed [31:0]addr[0:65535];
reg [6:0]k;
wire lrck;
always @(posedge clk or negedge reset_n)begin
	if(reset_n ==0) 
	k = 0;
	
	else
	k <= k+1;

end
assign lrck = k[6];
reg [15:0]i;
always @(posedge lrck or negedge reset_n)begin
	if(reset_n ==0)begin
		i <= 0;
	//	addrout <= 32'd0;
		end
	
	else begin
		i <= i+1;
	//	addrout <= addr[i];
		end
end

assign addrout = addr[i];
assign addr[0]= 0;
assign addr[1]= 38243550;
assign addr[2]= 76474970;
assign addr[3]= 114682135;
assign addr[4]= 152852926;
assign addr[5]= 190975237;
assign addr[6]= 229036977;
assign addr[7]= 267026072;
assign addr[8]= 304930476;
assign addr[9]= 342738165;
assign addr[10]= 380437148;
assign addr[11]= 418015468;
assign addr[12]= 455461206;
assign addr[13]= 492762486;
assign addr[14]= 529907477;
assign addr[15]= 566884397;
assign addr[16]= 603681519;
assign addr[17]= 640287172;
assign addr[18]= 676689746;
assign addr[19]= 712877694;
assign addr[20]= 748839539;
assign addr[21]= 784563876;
assign addr[22]= 820039373;
assign addr[23]= 855254778;
assign addr[24]= 890198924;
assign addr[25]= 924860725;
assign addr[26]= 959229189;
assign addr[27]= 993293415;
assign addr[28]= 1027042599;
assign addr[29]= 1060466036;
assign addr[30]= 1093553126;
assign addr[31]= 1126293375;
assign addr[32]= 1158676398;
assign addr[33]= 1190691925;
assign addr[34]= 1222329801;
assign addr[35]= 1253579991;
assign addr[36]= 1284432584;
assign addr[37]= 1314877795;
assign addr[38]= 1344905966;
assign addr[39]= 1374507575;
assign addr[40]= 1403673233;
assign addr[41]= 1432393688;
assign addr[42]= 1460659832;
assign addr[43]= 1488462700;
assign addr[44]= 1515793473;
assign addr[45]= 1542643483;
assign addr[46]= 1569004214;
assign addr[47]= 1594867305;
assign addr[48]= 1620224553;
assign addr[49]= 1645067915;
assign addr[50]= 1669389513;
assign addr[51]= 1693181631;
assign addr[52]= 1716436725;
assign addr[53]= 1739147417;
assign addr[54]= 1761306505;
assign addr[55]= 1782906961;
assign addr[56]= 1803941934;
assign addr[57]= 1824404752;
assign addr[58]= 1844288924;
assign addr[59]= 1863588145;
assign addr[60]= 1882296293;
assign addr[61]= 1900407434;
assign addr[62]= 1917915825;
assign addr[63]= 1934815911;
assign addr[64]= 1951102334;
assign addr[65]= 1966769926;
assign addr[66]= 1981813720;
assign addr[67]= 1996228943;
assign addr[68]= 2010011024;
assign addr[69]= 2023155591;
assign addr[70]= 2035658475;
assign addr[71]= 2047515711;
assign addr[72]= 2058723538;
assign addr[73]= 2069278401;
assign addr[74]= 2079176953;
assign addr[75]= 2088416053;
assign addr[76]= 2096992772;
assign addr[77]= 2104904390;
assign addr[78]= 2112148396;
assign addr[79]= 2118722494;
assign addr[80]= 2124624598;
assign addr[81]= 2129852837;
assign addr[82]= 2134405552;
assign addr[83]= 2138281298;
assign addr[84]= 2141478848;
assign addr[85]= 2143997187;
assign addr[86]= 2145835515;
assign addr[87]= 2146993250;
assign addr[88]= 2147470025;
assign addr[89]= 2147265689;
assign addr[90]= 2146380306;
assign addr[91]= 2144814157;
assign addr[92]= 2142567738;
assign addr[93]= 2139641764;
assign addr[94]= 2136037160;
assign addr[95]= 2131755071;
assign addr[96]= 2126796855;
assign addr[97]= 2121164085;
assign addr[98]= 2114858546;
assign addr[99]= 2107882239;
assign addr[100]= 2100237377;
assign addr[101]= 2091926384;
assign addr[102]= 2082951896;
assign addr[103]= 2073316760;
assign addr[104]= 2063024031;
assign addr[105]= 2052076975;
assign addr[106]= 2040479063;
assign addr[107]= 2028233973;
assign addr[108]= 2015345591;
assign addr[109]= 2001818002;
assign addr[110]= 1987655498;
assign addr[111]= 1972862571;
assign addr[112]= 1957443913;
assign addr[113]= 1941404413;
assign addr[114]= 1924749160;
assign addr[115]= 1907483436;
assign addr[116]= 1889612716;
assign addr[117]= 1871142669;
assign addr[118]= 1852079154;
assign addr[119]= 1832428215;
assign addr[120]= 1812196087;
assign addr[121]= 1791389186;
assign addr[122]= 1770014111;
assign addr[123]= 1748077642;
assign addr[124]= 1725586737;
assign addr[125]= 1702548529;
assign addr[126]= 1678970324;
assign addr[127]= 1654859602;
assign addr[128]= 1630224009;
assign addr[129]= 1605071359;
assign addr[130]= 1579409630;
assign addr[131]= 1553246960;
assign addr[132]= 1526591649;
assign addr[133]= 1499452149;
assign addr[134]= 1471837070;
assign addr[135]= 1443755168;
assign addr[136]= 1415215352;
assign addr[137]= 1386226674;
assign addr[138]= 1356798326;
assign addr[139]= 1326939644;
assign addr[140]= 1296660098;
assign addr[141]= 1265969291;
assign addr[142]= 1234876957;
assign addr[143]= 1203392958;
assign addr[144]= 1171527280;
assign addr[145]= 1139290029;
assign addr[146]= 1106691431;
assign addr[147]= 1073741824;
assign addr[148]= 1040451659;
assign addr[149]= 1006831495;
assign addr[150]= 972891995;
assign addr[151]= 938643924;
assign addr[152]= 904098143;
assign addr[153]= 869265610;
assign addr[154]= 834157373;
assign addr[155]= 798784567;
assign addr[156]= 763158411;
assign addr[157]= 727290205;
assign addr[158]= 691191324;
assign addr[159]= 654873219;
assign addr[160]= 618347408;
assign addr[161]= 581625477;
assign addr[162]= 544719071;
assign addr[163]= 507639898;
assign addr[164]= 470399716;
assign addr[165]= 433010339;
assign addr[166]= 395483624;
assign addr[167]= 357831473;
assign addr[168]= 320065829;
assign addr[169]= 282198671;
assign addr[170]= 244242007;
assign addr[171]= 206207878;
assign addr[172]= 168108346;
assign addr[173]= 129955495;
assign addr[174]= 91761426;
assign addr[175]= 53538253;
assign addr[176]= 15298099;
assign addr[177]= -22946906;
assign addr[178]= -61184634;
assign addr[179]= -99402956;
assign addr[180]= -137589750;
assign addr[181]= -175732905;
assign addr[182]= -213820322;
assign addr[183]= -251839923;
assign addr[184]= -289779648;
assign addr[185]= -327627463;
assign addr[186]= -365371365;
assign addr[187]= -402999383;
assign addr[188]= -440499581;
assign addr[189]= -477860067;
assign addr[190]= -515068990;
assign addr[191]= -552114549;
assign addr[192]= -588984994;
assign addr[193]= -625668632;
assign addr[194]= -662153826;
assign addr[195]= -698429006;
assign addr[196]= -734482665;
assign addr[197]= -770303369;
assign addr[198]= -805879757;
assign addr[199]= -841200544;
assign addr[200]= -876254528;
assign addr[201]= -911030591;
assign addr[202]= -945517704;
assign addr[203]= -979704927;
assign addr[204]= -1013581418;
assign addr[205]= -1047136432;
assign addr[206]= -1080359326;
assign addr[207]= -1113239564;
assign addr[208]= -1145766716;
assign addr[209]= -1177930466;
assign addr[210]= -1209720613;
assign addr[211]= -1241127074;
assign addr[212]= -1272139887;
assign addr[213]= -1302749217;
assign addr[214]= -1332945355;
assign addr[215]= -1362718723;
assign addr[216]= -1392059879;
assign addr[217]= -1420959516;
assign addr[218]= -1449408469;
assign addr[219]= -1477397714;
assign addr[220]= -1504918373;
assign addr[221]= -1531961719;
assign addr[222]= -1558519173;
assign addr[223]= -1584582314;
assign addr[224]= -1610142873;
assign addr[225]= -1635192744;
assign addr[226]= -1659723983;
assign addr[227]= -1683728808;
assign addr[228]= -1707199606;
assign addr[229]= -1730128933;
assign addr[230]= -1752509516;
assign addr[231]= -1774334257;
assign addr[232]= -1795596234;
assign addr[233]= -1816288703;
assign addr[234]= -1836405100;
assign addr[235]= -1855939047;
assign addr[236]= -1874884346;
assign addr[237]= -1893234990;
assign addr[238]= -1910985158;
assign addr[239]= -1928129220;
assign addr[240]= -1944661739;
assign addr[241]= -1960577471;
assign addr[242]= -1975871368;
assign addr[243]= -1990538579;
assign addr[244]= -2004574453;
assign addr[245]= -2017974537;
assign addr[246]= -2030734582;
assign addr[247]= -2042850540;
assign addr[248]= -2054318569;
assign addr[249]= -2065135031;
assign addr[250]= -2075296495;
assign addr[251]= -2084799740;
assign addr[252]= -2093641749;
assign addr[253]= -2101819720;
assign addr[254]= -2109331059;
assign addr[255]= -2116173382;
assign addr[256]= -2122344521;
assign addr[257]= -2127842516;
assign addr[258]= -2132665626;
assign addr[259]= -2136812319;
assign addr[260]= -2140281282;
assign addr[261]= -2143071413;
assign addr[262]= -2145181827;
assign addr[263]= -2146611856;
assign addr[264]= -2147361045;
assign addr[265]= -2147429158;
assign addr[266]= -2146816171;
assign addr[267]= -2145522281;
assign addr[268]= -2143547897;
assign addr[269]= -2140893646;
assign addr[270]= -2137560369;
assign addr[271]= -2133549123;
assign addr[272]= -2128861181;
assign addr[273]= -2123498030;
assign addr[274]= -2117461370;
assign addr[275]= -2110753117;
assign addr[276]= -2103375398;
assign addr[277]= -2095330553;
assign addr[278]= -2086621133;
assign addr[279]= -2077249901;
assign addr[280]= -2067219829;
assign addr[281]= -2056534099;
assign addr[282]= -2045196100;
assign addr[283]= -2033209426;
assign addr[284]= -2020577882;
assign addr[285]= -2007305472;
assign addr[286]= -1993396407;
assign addr[287]= -1978855097;
assign addr[288]= -1963686155;
assign addr[289]= -1947894393;
assign addr[290]= -1931484818;
assign addr[291]= -1914462636;
assign addr[292]= -1896833245;
assign addr[293]= -1878602237;
assign addr[294]= -1859775393;
assign addr[295]= -1840358687;
assign addr[296]= -1820358275;
assign addr[297]= -1799780501;
assign addr[298]= -1778631892;
assign addr[299]= -1756919156;
assign addr[300]= -1734649179;
assign addr[301]= -1711829025;
assign addr[302]= -1688465931;
assign addr[303]= -1664567307;
assign addr[304]= -1640140734;
assign addr[305]= -1615193959;
assign addr[306]= -1589734894;
assign addr[307]= -1563771613;
assign addr[308]= -1537312353;
assign addr[309]= -1510365504;
assign addr[310]= -1482939614;
assign addr[311]= -1455043381;
assign addr[312]= -1426685652;
assign addr[313]= -1397875423;
assign addr[314]= -1368621831;
assign addr[315]= -1338934154;
assign addr[316]= -1308821808;
assign addr[317]= -1278294345;
assign addr[318]= -1247361445;
assign addr[319]= -1216032921;
assign addr[320]= -1184318708;
assign addr[321]= -1152228866;
assign addr[322]= -1119773573;
assign addr[323]= -1086963121;
assign addr[324]= -1053807919;
assign addr[325]= -1020318481;
assign addr[326]= -986505429;
assign addr[327]= -952379488;
assign addr[328]= -917951481;
assign addr[329]= -883232329;
assign addr[330]= -848233042;
assign addr[331]= -812964722;
assign addr[332]= -777438554;
assign addr[333]= -741665807;
assign addr[334]= -705657826;
assign addr[335]= -669426032;
assign addr[336]= -632981917;
assign addr[337]= -596337040;
assign addr[338]= -559503022;
assign addr[339]= -522491548;
assign addr[340]= -485314355;
assign addr[341]= -447983235;
assign addr[342]= -410510029;
assign addr[343]= -372906622;
assign addr[344]= -335184940;
assign addr[345]= -297356948;
assign addr[346]= -259434643;
assign addr[347]= -221430054;
assign addr[348]= -183355234;
assign addr[349]= -145222259;
assign addr[350]= -107043224;
assign addr[351]= -68830239;
assign addr[352]= -30595422;
assign addr[353]= 7649098;
assign addr[354]= 45891193;
assign addr[355]= 84118732;
assign addr[356]= 122319591;
assign addr[357]= 160481654;
assign addr[358]= 198592817;
assign addr[359]= 236640993;
assign addr[360]= 274614114;
assign addr[361]= 312500135;
assign addr[362]= 350287041;
assign addr[363]= 387962847;
assign addr[364]= 425515602;
assign addr[365]= 462933398;
assign addr[366]= 500204365;
assign addr[367]= 537316682;
assign addr[368]= 574258580;
assign addr[369]= 611018340;
assign addr[370]= 647584304;
assign addr[371]= 683944874;
assign addr[372]= 720088517;
assign addr[373]= 756003771;
assign addr[374]= 791679244;
assign addr[375]= 827103620;
assign addr[376]= 862265664;
assign addr[377]= 897154224;
assign addr[378]= 931758235;
assign addr[379]= 966066720;
assign addr[380]= 1000068799;
assign addr[381]= 1033753687;
assign addr[382]= 1067110699;
assign addr[383]= 1100129257;
assign addr[384]= 1132798888;
assign addr[385]= 1165109230;
assign addr[386]= 1197050035;
assign addr[387]= 1228611172;
assign addr[388]= 1259782632;
assign addr[389]= 1290554528;
assign addr[390]= 1320917099;
assign addr[391]= 1350860716;
assign addr[392]= 1380375881;
assign addr[393]= 1409453233;
assign addr[394]= 1438083551;
assign addr[395]= 1466257752;
assign addr[396]= 1493966902;
assign addr[397]= 1521202211;
assign addr[398]= 1547955041;
assign addr[399]= 1574216908;
assign addr[400]= 1599979481;
assign addr[401]= 1625234591;
assign addr[402]= 1649974225;
assign addr[403]= 1674190539;
assign addr[404]= 1697875851;
assign addr[405]= 1721022648;
assign addr[406]= 1743623590;
assign addr[407]= 1765671509;
assign addr[408]= 1787159411;
assign addr[409]= 1808080480;
assign addr[410]= 1828428082;
assign addr[411]= 1848195763;
assign addr[412]= 1867377253;
assign addr[413]= 1885966468;
assign addr[414]= 1903957513;
assign addr[415]= 1921344681;
assign addr[416]= 1938122457;
assign addr[417]= 1954285520;
assign addr[418]= 1969828744;
assign addr[419]= 1984747199;
assign addr[420]= 1999036154;
assign addr[421]= 2012691075;
assign addr[422]= 2025707632;
assign addr[423]= 2038081698;
assign addr[424]= 2049809346;
assign addr[425]= 2060886858;
assign addr[426]= 2071310720;
assign addr[427]= 2081077626;
assign addr[428]= 2090184478;
assign addr[429]= 2098628387;
assign addr[430]= 2106406677;
assign addr[431]= 2113516878;
assign addr[432]= 2119956737;
assign addr[433]= 2125724211;
assign addr[434]= 2130817471;
assign addr[435]= 2135234901;
assign addr[436]= 2138975100;
assign addr[437]= 2142036881;
assign addr[438]= 2144419275;
assign addr[439]= 2146121524;
assign addr[440]= 2147143090;
assign addr[441]= 2147483648;
assign addr[442]= 2147143090;
assign addr[443]= 2146121524;
assign addr[444]= 2144419275;
assign addr[445]= 2142036881;
assign addr[446]= 2138975100;
assign addr[447]= 2135234901;
assign addr[448]= 2130817471;
assign addr[449]= 2125724211;
assign addr[450]= 2119956737;
assign addr[451]= 2113516878;
assign addr[452]= 2106406677;
assign addr[453]= 2098628387;
assign addr[454]= 2090184478;
assign addr[455]= 2081077626;
assign addr[456]= 2071310720;
assign addr[457]= 2060886858;
assign addr[458]= 2049809346;
assign addr[459]= 2038081698;
assign addr[460]= 2025707632;
assign addr[461]= 2012691075;
assign addr[462]= 1999036154;
assign addr[463]= 1984747199;
assign addr[464]= 1969828744;
assign addr[465]= 1954285520;
assign addr[466]= 1938122457;
assign addr[467]= 1921344681;
assign addr[468]= 1903957513;
assign addr[469]= 1885966468;
assign addr[470]= 1867377253;
assign addr[471]= 1848195763;
assign addr[472]= 1828428082;
assign addr[473]= 1808080480;
assign addr[474]= 1787159411;
assign addr[475]= 1765671509;
assign addr[476]= 1743623590;
assign addr[477]= 1721022648;
assign addr[478]= 1697875851;
assign addr[479]= 1674190539;
assign addr[480]= 1649974225;
assign addr[481]= 1625234591;
assign addr[482]= 1599979481;
assign addr[483]= 1574216908;
assign addr[484]= 1547955041;
assign addr[485]= 1521202211;
assign addr[486]= 1493966902;
assign addr[487]= 1466257752;
assign addr[488]= 1438083551;
assign addr[489]= 1409453233;
assign addr[490]= 1380375881;
assign addr[491]= 1350860716;
assign addr[492]= 1320917099;
assign addr[493]= 1290554528;
assign addr[494]= 1259782632;
assign addr[495]= 1228611172;
assign addr[496]= 1197050035;
assign addr[497]= 1165109230;
assign addr[498]= 1132798888;
assign addr[499]= 1100129257;
assign addr[500]= 1067110699;
assign addr[501]= 1033753687;
assign addr[502]= 1000068799;
assign addr[503]= 966066720;
assign addr[504]= 931758235;
assign addr[505]= 897154224;
assign addr[506]= 862265664;
assign addr[507]= 827103620;
assign addr[508]= 791679244;
assign addr[509]= 756003771;
assign addr[510]= 720088517;
assign addr[511]= 683944874;
assign addr[512]= 647584304;
assign addr[513]= 611018340;
assign addr[514]= 574258580;
assign addr[515]= 537316682;
assign addr[516]= 500204365;
assign addr[517]= 462933398;
assign addr[518]= 425515602;
assign addr[519]= 387962847;
assign addr[520]= 350287041;
assign addr[521]= 312500135;
assign addr[522]= 274614114;
assign addr[523]= 236640993;
assign addr[524]= 198592817;
assign addr[525]= 160481654;
assign addr[526]= 122319591;
assign addr[527]= 84118732;
assign addr[528]= 45891193;
assign addr[529]= 7649098;
assign addr[530]= -30595422;
assign addr[531]= -68830239;
assign addr[532]= -107043224;
assign addr[533]= -145222259;
assign addr[534]= -183355234;
assign addr[535]= -221430054;
assign addr[536]= -259434643;
assign addr[537]= -297356948;
assign addr[538]= -335184940;
assign addr[539]= -372906622;
assign addr[540]= -410510029;
assign addr[541]= -447983235;
assign addr[542]= -485314355;
assign addr[543]= -522491548;
assign addr[544]= -559503022;
assign addr[545]= -596337040;
assign addr[546]= -632981917;
assign addr[547]= -669426032;
assign addr[548]= -705657826;
assign addr[549]= -741665807;
assign addr[550]= -777438554;
assign addr[551]= -812964722;
assign addr[552]= -848233042;
assign addr[553]= -883232329;
assign addr[554]= -917951481;
assign addr[555]= -952379488;
assign addr[556]= -986505429;
assign addr[557]= -1020318481;
assign addr[558]= -1053807919;
assign addr[559]= -1086963121;
assign addr[560]= -1119773573;
assign addr[561]= -1152228866;
assign addr[562]= -1184318708;
assign addr[563]= -1216032921;
assign addr[564]= -1247361445;
assign addr[565]= -1278294345;
assign addr[566]= -1308821808;
assign addr[567]= -1338934154;
assign addr[568]= -1368621831;
assign addr[569]= -1397875423;
assign addr[570]= -1426685652;
assign addr[571]= -1455043381;
assign addr[572]= -1482939614;
assign addr[573]= -1510365504;
assign addr[574]= -1537312353;
assign addr[575]= -1563771613;
assign addr[576]= -1589734894;
assign addr[577]= -1615193959;
assign addr[578]= -1640140734;
assign addr[579]= -1664567307;
assign addr[580]= -1688465931;
assign addr[581]= -1711829025;
assign addr[582]= -1734649179;
assign addr[583]= -1756919156;
assign addr[584]= -1778631892;
assign addr[585]= -1799780501;
assign addr[586]= -1820358275;
assign addr[587]= -1840358687;
assign addr[588]= -1859775393;
assign addr[589]= -1878602237;
assign addr[590]= -1896833245;
assign addr[591]= -1914462636;
assign addr[592]= -1931484818;
assign addr[593]= -1947894393;
assign addr[594]= -1963686155;
assign addr[595]= -1978855097;
assign addr[596]= -1993396407;
assign addr[597]= -2007305472;
assign addr[598]= -2020577882;
assign addr[599]= -2033209426;
assign addr[600]= -2045196100;
assign addr[601]= -2056534099;
assign addr[602]= -2067219829;
assign addr[603]= -2077249901;
assign addr[604]= -2086621133;
assign addr[605]= -2095330553;
assign addr[606]= -2103375398;
assign addr[607]= -2110753117;
assign addr[608]= -2117461370;
assign addr[609]= -2123498030;
assign addr[610]= -2128861181;
assign addr[611]= -2133549123;
assign addr[612]= -2137560369;
assign addr[613]= -2140893646;
assign addr[614]= -2143547897;
assign addr[615]= -2145522281;
assign addr[616]= -2146816171;
assign addr[617]= -2147429158;
assign addr[618]= -2147361045;
assign addr[619]= -2146611856;
assign addr[620]= -2145181827;
assign addr[621]= -2143071413;
assign addr[622]= -2140281282;
assign addr[623]= -2136812319;
assign addr[624]= -2132665626;
assign addr[625]= -2127842516;
assign addr[626]= -2122344521;
assign addr[627]= -2116173382;
assign addr[628]= -2109331059;
assign addr[629]= -2101819720;
assign addr[630]= -2093641749;
assign addr[631]= -2084799740;
assign addr[632]= -2075296495;
assign addr[633]= -2065135031;
assign addr[634]= -2054318569;
assign addr[635]= -2042850540;
assign addr[636]= -2030734582;
assign addr[637]= -2017974537;
assign addr[638]= -2004574453;
assign addr[639]= -1990538579;
assign addr[640]= -1975871368;
assign addr[641]= -1960577471;
assign addr[642]= -1944661739;
assign addr[643]= -1928129220;
assign addr[644]= -1910985158;
assign addr[645]= -1893234990;
assign addr[646]= -1874884346;
assign addr[647]= -1855939047;
assign addr[648]= -1836405100;
assign addr[649]= -1816288703;
assign addr[650]= -1795596234;
assign addr[651]= -1774334257;
assign addr[652]= -1752509516;
assign addr[653]= -1730128933;
assign addr[654]= -1707199606;
assign addr[655]= -1683728808;
assign addr[656]= -1659723983;
assign addr[657]= -1635192744;
assign addr[658]= -1610142873;
assign addr[659]= -1584582314;
assign addr[660]= -1558519173;
assign addr[661]= -1531961719;
assign addr[662]= -1504918373;
assign addr[663]= -1477397714;
assign addr[664]= -1449408469;
assign addr[665]= -1420959516;
assign addr[666]= -1392059879;
assign addr[667]= -1362718723;
assign addr[668]= -1332945355;
assign addr[669]= -1302749217;
assign addr[670]= -1272139887;
assign addr[671]= -1241127074;
assign addr[672]= -1209720613;
assign addr[673]= -1177930466;
assign addr[674]= -1145766716;
assign addr[675]= -1113239564;
assign addr[676]= -1080359326;
assign addr[677]= -1047136432;
assign addr[678]= -1013581418;
assign addr[679]= -979704927;
assign addr[680]= -945517704;
assign addr[681]= -911030591;
assign addr[682]= -876254528;
assign addr[683]= -841200544;
assign addr[684]= -805879757;
assign addr[685]= -770303369;
assign addr[686]= -734482665;
assign addr[687]= -698429006;
assign addr[688]= -662153826;
assign addr[689]= -625668632;
assign addr[690]= -588984994;
assign addr[691]= -552114549;
assign addr[692]= -515068990;
assign addr[693]= -477860067;
assign addr[694]= -440499581;
assign addr[695]= -402999383;
assign addr[696]= -365371365;
assign addr[697]= -327627463;
assign addr[698]= -289779648;
assign addr[699]= -251839923;
assign addr[700]= -213820322;
assign addr[701]= -175732905;
assign addr[702]= -137589750;
assign addr[703]= -99402956;
assign addr[704]= -61184634;
assign addr[705]= -22946906;
assign addr[706]= 15298099;
assign addr[707]= 53538253;
assign addr[708]= 91761426;
assign addr[709]= 129955495;
assign addr[710]= 168108346;
assign addr[711]= 206207878;
assign addr[712]= 244242007;
assign addr[713]= 282198671;
assign addr[714]= 320065829;
assign addr[715]= 357831473;
assign addr[716]= 395483624;
assign addr[717]= 433010339;
assign addr[718]= 470399716;
assign addr[719]= 507639898;
assign addr[720]= 544719071;
assign addr[721]= 581625477;
assign addr[722]= 618347408;
assign addr[723]= 654873219;
assign addr[724]= 691191324;
assign addr[725]= 727290205;
assign addr[726]= 763158411;
assign addr[727]= 798784567;
assign addr[728]= 834157373;
assign addr[729]= 869265610;
assign addr[730]= 904098143;
assign addr[731]= 938643924;
assign addr[732]= 972891995;
assign addr[733]= 1006831495;
assign addr[734]= 1040451659;
assign addr[735]= 1073741824;
assign addr[736]= 1106691431;
assign addr[737]= 1139290029;
assign addr[738]= 1171527280;
assign addr[739]= 1203392958;
assign addr[740]= 1234876957;
assign addr[741]= 1265969291;
assign addr[742]= 1296660098;
assign addr[743]= 1326939644;
assign addr[744]= 1356798326;
assign addr[745]= 1386226674;
assign addr[746]= 1415215352;
assign addr[747]= 1443755168;
assign addr[748]= 1471837070;
assign addr[749]= 1499452149;
assign addr[750]= 1526591649;
assign addr[751]= 1553246960;
assign addr[752]= 1579409630;
assign addr[753]= 1605071359;
assign addr[754]= 1630224009;
assign addr[755]= 1654859602;
assign addr[756]= 1678970324;
assign addr[757]= 1702548529;
assign addr[758]= 1725586737;
assign addr[759]= 1748077642;
assign addr[760]= 1770014111;
assign addr[761]= 1791389186;
assign addr[762]= 1812196087;
assign addr[763]= 1832428215;
assign addr[764]= 1852079154;
assign addr[765]= 1871142669;
assign addr[766]= 1889612716;
assign addr[767]= 1907483436;
assign addr[768]= 1924749160;
assign addr[769]= 1941404413;
assign addr[770]= 1957443913;
assign addr[771]= 1972862571;
assign addr[772]= 1987655498;
assign addr[773]= 2001818002;
assign addr[774]= 2015345591;
assign addr[775]= 2028233973;
assign addr[776]= 2040479063;
assign addr[777]= 2052076975;
assign addr[778]= 2063024031;
assign addr[779]= 2073316760;
assign addr[780]= 2082951896;
assign addr[781]= 2091926384;
assign addr[782]= 2100237377;
assign addr[783]= 2107882239;
assign addr[784]= 2114858546;
assign addr[785]= 2121164085;
assign addr[786]= 2126796855;
assign addr[787]= 2131755071;
assign addr[788]= 2136037160;
assign addr[789]= 2139641764;
assign addr[790]= 2142567738;
assign addr[791]= 2144814157;
assign addr[792]= 2146380306;
assign addr[793]= 2147265689;
assign addr[794]= 2147470025;
assign addr[795]= 2146993250;
assign addr[796]= 2145835515;
assign addr[797]= 2143997187;
assign addr[798]= 2141478848;
assign addr[799]= 2138281298;
assign addr[800]= 2134405552;
assign addr[801]= 2129852837;
assign addr[802]= 2124624598;
assign addr[803]= 2118722494;
assign addr[804]= 2112148396;
assign addr[805]= 2104904390;
assign addr[806]= 2096992772;
assign addr[807]= 2088416053;
assign addr[808]= 2079176953;
assign addr[809]= 2069278401;
assign addr[810]= 2058723538;
assign addr[811]= 2047515711;
assign addr[812]= 2035658475;
assign addr[813]= 2023155591;
assign addr[814]= 2010011024;
assign addr[815]= 1996228943;
assign addr[816]= 1981813720;
assign addr[817]= 1966769926;
assign addr[818]= 1951102334;
assign addr[819]= 1934815911;
assign addr[820]= 1917915825;
assign addr[821]= 1900407434;
assign addr[822]= 1882296293;
assign addr[823]= 1863588145;
assign addr[824]= 1844288924;
assign addr[825]= 1824404752;
assign addr[826]= 1803941934;
assign addr[827]= 1782906961;
assign addr[828]= 1761306505;
assign addr[829]= 1739147417;
assign addr[830]= 1716436725;
assign addr[831]= 1693181631;
assign addr[832]= 1669389513;
assign addr[833]= 1645067915;
assign addr[834]= 1620224553;
assign addr[835]= 1594867305;
assign addr[836]= 1569004214;
assign addr[837]= 1542643483;
assign addr[838]= 1515793473;
assign addr[839]= 1488462700;
assign addr[840]= 1460659832;
assign addr[841]= 1432393688;
assign addr[842]= 1403673233;
assign addr[843]= 1374507575;
assign addr[844]= 1344905966;
assign addr[845]= 1314877795;
assign addr[846]= 1284432584;
assign addr[847]= 1253579991;
assign addr[848]= 1222329801;
assign addr[849]= 1190691925;
assign addr[850]= 1158676398;
assign addr[851]= 1126293375;
assign addr[852]= 1093553126;
assign addr[853]= 1060466036;
assign addr[854]= 1027042599;
assign addr[855]= 993293415;
assign addr[856]= 959229189;
assign addr[857]= 924860725;
assign addr[858]= 890198924;
assign addr[859]= 855254778;
assign addr[860]= 820039373;
assign addr[861]= 784563876;
assign addr[862]= 748839539;
assign addr[863]= 712877694;
assign addr[864]= 676689746;
assign addr[865]= 640287172;
assign addr[866]= 603681519;
assign addr[867]= 566884397;
assign addr[868]= 529907477;
assign addr[869]= 492762486;
assign addr[870]= 455461206;
assign addr[871]= 418015468;
assign addr[872]= 380437148;
assign addr[873]= 342738165;
assign addr[874]= 304930476;
assign addr[875]= 267026072;
assign addr[876]= 229036977;
assign addr[877]= 190975237;
assign addr[878]= 152852926;
assign addr[879]= 114682135;
assign addr[880]= 76474970;
assign addr[881]= 38243550;
assign addr[882]= 0;
assign addr[883]= -38243550;
assign addr[884]= -76474970;
assign addr[885]= -114682135;
assign addr[886]= -152852926;
assign addr[887]= -190975237;
assign addr[888]= -229036977;
assign addr[889]= -267026072;
assign addr[890]= -304930476;
assign addr[891]= -342738165;
assign addr[892]= -380437148;
assign addr[893]= -418015468;
assign addr[894]= -455461206;
assign addr[895]= -492762486;
assign addr[896]= -529907477;
assign addr[897]= -566884397;
assign addr[898]= -603681519;
assign addr[899]= -640287172;
assign addr[900]= -676689746;
assign addr[901]= -712877694;
assign addr[902]= -748839539;
assign addr[903]= -784563876;
assign addr[904]= -820039373;
assign addr[905]= -855254778;
assign addr[906]= -890198924;
assign addr[907]= -924860725;
assign addr[908]= -959229189;
assign addr[909]= -993293415;
assign addr[910]= -1027042599;
assign addr[911]= -1060466036;
assign addr[912]= -1093553126;
assign addr[913]= -1126293375;
assign addr[914]= -1158676398;
assign addr[915]= -1190691925;
assign addr[916]= -1222329801;
assign addr[917]= -1253579991;
assign addr[918]= -1284432584;
assign addr[919]= -1314877795;
assign addr[920]= -1344905966;
assign addr[921]= -1374507575;
assign addr[922]= -1403673233;
assign addr[923]= -1432393688;
assign addr[924]= -1460659832;
assign addr[925]= -1488462700;
assign addr[926]= -1515793473;
assign addr[927]= -1542643483;
assign addr[928]= -1569004214;
assign addr[929]= -1594867305;
assign addr[930]= -1620224553;
assign addr[931]= -1645067915;
assign addr[932]= -1669389513;
assign addr[933]= -1693181631;
assign addr[934]= -1716436725;
assign addr[935]= -1739147417;
assign addr[936]= -1761306505;
assign addr[937]= -1782906961;
assign addr[938]= -1803941934;
assign addr[939]= -1824404752;
assign addr[940]= -1844288924;
assign addr[941]= -1863588145;
assign addr[942]= -1882296293;
assign addr[943]= -1900407434;
assign addr[944]= -1917915825;
assign addr[945]= -1934815911;
assign addr[946]= -1951102334;
assign addr[947]= -1966769926;
assign addr[948]= -1981813720;
assign addr[949]= -1996228943;
assign addr[950]= -2010011024;
assign addr[951]= -2023155591;
assign addr[952]= -2035658475;
assign addr[953]= -2047515711;
assign addr[954]= -2058723538;
assign addr[955]= -2069278401;
assign addr[956]= -2079176953;
assign addr[957]= -2088416053;
assign addr[958]= -2096992772;
assign addr[959]= -2104904390;
assign addr[960]= -2112148396;
assign addr[961]= -2118722494;
assign addr[962]= -2124624598;
assign addr[963]= -2129852837;
assign addr[964]= -2134405552;
assign addr[965]= -2138281298;
assign addr[966]= -2141478848;
assign addr[967]= -2143997187;
assign addr[968]= -2145835515;
assign addr[969]= -2146993250;
assign addr[970]= -2147470025;
assign addr[971]= -2147265689;
assign addr[972]= -2146380306;
assign addr[973]= -2144814157;
assign addr[974]= -2142567738;
assign addr[975]= -2139641764;
assign addr[976]= -2136037160;
assign addr[977]= -2131755071;
assign addr[978]= -2126796855;
assign addr[979]= -2121164085;
assign addr[980]= -2114858546;
assign addr[981]= -2107882239;
assign addr[982]= -2100237377;
assign addr[983]= -2091926384;
assign addr[984]= -2082951896;
assign addr[985]= -2073316760;
assign addr[986]= -2063024031;
assign addr[987]= -2052076975;
assign addr[988]= -2040479063;
assign addr[989]= -2028233973;
assign addr[990]= -2015345591;
assign addr[991]= -2001818002;
assign addr[992]= -1987655498;
assign addr[993]= -1972862571;
assign addr[994]= -1957443913;
assign addr[995]= -1941404413;
assign addr[996]= -1924749160;
assign addr[997]= -1907483436;
assign addr[998]= -1889612716;
assign addr[999]= -1871142669;
assign addr[1000]= -1852079154;
assign addr[1001]= -1832428215;
assign addr[1002]= -1812196087;
assign addr[1003]= -1791389186;
assign addr[1004]= -1770014111;
assign addr[1005]= -1748077642;
assign addr[1006]= -1725586737;
assign addr[1007]= -1702548529;
assign addr[1008]= -1678970324;
assign addr[1009]= -1654859602;
assign addr[1010]= -1630224009;
assign addr[1011]= -1605071359;
assign addr[1012]= -1579409630;
assign addr[1013]= -1553246960;
assign addr[1014]= -1526591649;
assign addr[1015]= -1499452149;
assign addr[1016]= -1471837070;
assign addr[1017]= -1443755168;
assign addr[1018]= -1415215352;
assign addr[1019]= -1386226674;
assign addr[1020]= -1356798326;
assign addr[1021]= -1326939644;
assign addr[1022]= -1296660098;
assign addr[1023]= -1265969291;
assign addr[1024]= -1234876957;
assign addr[1025]= -1203392958;
assign addr[1026]= -1171527280;
assign addr[1027]= -1139290029;
assign addr[1028]= -1106691431;
assign addr[1029]= -1073741824;
assign addr[1030]= -1040451659;
assign addr[1031]= -1006831495;
assign addr[1032]= -972891995;
assign addr[1033]= -938643924;
assign addr[1034]= -904098143;
assign addr[1035]= -869265610;
assign addr[1036]= -834157373;
assign addr[1037]= -798784567;
assign addr[1038]= -763158411;
assign addr[1039]= -727290205;
assign addr[1040]= -691191324;
assign addr[1041]= -654873219;
assign addr[1042]= -618347408;
assign addr[1043]= -581625477;
assign addr[1044]= -544719071;
assign addr[1045]= -507639898;
assign addr[1046]= -470399716;
assign addr[1047]= -433010339;
assign addr[1048]= -395483624;
assign addr[1049]= -357831473;
assign addr[1050]= -320065829;
assign addr[1051]= -282198671;
assign addr[1052]= -244242007;
assign addr[1053]= -206207878;
assign addr[1054]= -168108346;
assign addr[1055]= -129955495;
assign addr[1056]= -91761426;
assign addr[1057]= -53538253;
assign addr[1058]= -15298099;
assign addr[1059]= 22946906;
assign addr[1060]= 61184634;
assign addr[1061]= 99402956;
assign addr[1062]= 137589750;
assign addr[1063]= 175732905;
assign addr[1064]= 213820322;
assign addr[1065]= 251839923;
assign addr[1066]= 289779648;
assign addr[1067]= 327627463;
assign addr[1068]= 365371365;
assign addr[1069]= 402999383;
assign addr[1070]= 440499581;
assign addr[1071]= 477860067;
assign addr[1072]= 515068990;
assign addr[1073]= 552114549;
assign addr[1074]= 588984994;
assign addr[1075]= 625668632;
assign addr[1076]= 662153826;
assign addr[1077]= 698429006;
assign addr[1078]= 734482665;
assign addr[1079]= 770303369;
assign addr[1080]= 805879757;
assign addr[1081]= 841200544;
assign addr[1082]= 876254528;
assign addr[1083]= 911030591;
assign addr[1084]= 945517704;
assign addr[1085]= 979704927;
assign addr[1086]= 1013581418;
assign addr[1087]= 1047136432;
assign addr[1088]= 1080359326;
assign addr[1089]= 1113239564;
assign addr[1090]= 1145766716;
assign addr[1091]= 1177930466;
assign addr[1092]= 1209720613;
assign addr[1093]= 1241127074;
assign addr[1094]= 1272139887;
assign addr[1095]= 1302749217;
assign addr[1096]= 1332945355;
assign addr[1097]= 1362718723;
assign addr[1098]= 1392059879;
assign addr[1099]= 1420959516;
assign addr[1100]= 1449408469;
assign addr[1101]= 1477397714;
assign addr[1102]= 1504918373;
assign addr[1103]= 1531961719;
assign addr[1104]= 1558519173;
assign addr[1105]= 1584582314;
assign addr[1106]= 1610142873;
assign addr[1107]= 1635192744;
assign addr[1108]= 1659723983;
assign addr[1109]= 1683728808;
assign addr[1110]= 1707199606;
assign addr[1111]= 1730128933;
assign addr[1112]= 1752509516;
assign addr[1113]= 1774334257;
assign addr[1114]= 1795596234;
assign addr[1115]= 1816288703;
assign addr[1116]= 1836405100;
assign addr[1117]= 1855939047;
assign addr[1118]= 1874884346;
assign addr[1119]= 1893234990;
assign addr[1120]= 1910985158;
assign addr[1121]= 1928129220;
assign addr[1122]= 1944661739;
assign addr[1123]= 1960577471;
assign addr[1124]= 1975871368;
assign addr[1125]= 1990538579;
assign addr[1126]= 2004574453;
assign addr[1127]= 2017974537;
assign addr[1128]= 2030734582;
assign addr[1129]= 2042850540;
assign addr[1130]= 2054318569;
assign addr[1131]= 2065135031;
assign addr[1132]= 2075296495;
assign addr[1133]= 2084799740;
assign addr[1134]= 2093641749;
assign addr[1135]= 2101819720;
assign addr[1136]= 2109331059;
assign addr[1137]= 2116173382;
assign addr[1138]= 2122344521;
assign addr[1139]= 2127842516;
assign addr[1140]= 2132665626;
assign addr[1141]= 2136812319;
assign addr[1142]= 2140281282;
assign addr[1143]= 2143071413;
assign addr[1144]= 2145181827;
assign addr[1145]= 2146611856;
assign addr[1146]= 2147361045;
assign addr[1147]= 2147429158;
assign addr[1148]= 2146816171;
assign addr[1149]= 2145522281;
assign addr[1150]= 2143547897;
assign addr[1151]= 2140893646;
assign addr[1152]= 2137560369;
assign addr[1153]= 2133549123;
assign addr[1154]= 2128861181;
assign addr[1155]= 2123498030;
assign addr[1156]= 2117461370;
assign addr[1157]= 2110753117;
assign addr[1158]= 2103375398;
assign addr[1159]= 2095330553;
assign addr[1160]= 2086621133;
assign addr[1161]= 2077249901;
assign addr[1162]= 2067219829;
assign addr[1163]= 2056534099;
assign addr[1164]= 2045196100;
assign addr[1165]= 2033209426;
assign addr[1166]= 2020577882;
assign addr[1167]= 2007305472;
assign addr[1168]= 1993396407;
assign addr[1169]= 1978855097;
assign addr[1170]= 1963686155;
assign addr[1171]= 1947894393;
assign addr[1172]= 1931484818;
assign addr[1173]= 1914462636;
assign addr[1174]= 1896833245;
assign addr[1175]= 1878602237;
assign addr[1176]= 1859775393;
assign addr[1177]= 1840358687;
assign addr[1178]= 1820358275;
assign addr[1179]= 1799780501;
assign addr[1180]= 1778631892;
assign addr[1181]= 1756919156;
assign addr[1182]= 1734649179;
assign addr[1183]= 1711829025;
assign addr[1184]= 1688465931;
assign addr[1185]= 1664567307;
assign addr[1186]= 1640140734;
assign addr[1187]= 1615193959;
assign addr[1188]= 1589734894;
assign addr[1189]= 1563771613;
assign addr[1190]= 1537312353;
assign addr[1191]= 1510365504;
assign addr[1192]= 1482939614;
assign addr[1193]= 1455043381;
assign addr[1194]= 1426685652;
assign addr[1195]= 1397875423;
assign addr[1196]= 1368621831;
assign addr[1197]= 1338934154;
assign addr[1198]= 1308821808;
assign addr[1199]= 1278294345;
assign addr[1200]= 1247361445;
assign addr[1201]= 1216032921;
assign addr[1202]= 1184318708;
assign addr[1203]= 1152228866;
assign addr[1204]= 1119773573;
assign addr[1205]= 1086963121;
assign addr[1206]= 1053807919;
assign addr[1207]= 1020318481;
assign addr[1208]= 986505429;
assign addr[1209]= 952379488;
assign addr[1210]= 917951481;
assign addr[1211]= 883232329;
assign addr[1212]= 848233042;
assign addr[1213]= 812964722;
assign addr[1214]= 777438554;
assign addr[1215]= 741665807;
assign addr[1216]= 705657826;
assign addr[1217]= 669426032;
assign addr[1218]= 632981917;
assign addr[1219]= 596337040;
assign addr[1220]= 559503022;
assign addr[1221]= 522491548;
assign addr[1222]= 485314355;
assign addr[1223]= 447983235;
assign addr[1224]= 410510029;
assign addr[1225]= 372906622;
assign addr[1226]= 335184940;
assign addr[1227]= 297356948;
assign addr[1228]= 259434643;
assign addr[1229]= 221430054;
assign addr[1230]= 183355234;
assign addr[1231]= 145222259;
assign addr[1232]= 107043224;
assign addr[1233]= 68830239;
assign addr[1234]= 30595422;
assign addr[1235]= -7649098;
assign addr[1236]= -45891193;
assign addr[1237]= -84118732;
assign addr[1238]= -122319591;
assign addr[1239]= -160481654;
assign addr[1240]= -198592817;
assign addr[1241]= -236640993;
assign addr[1242]= -274614114;
assign addr[1243]= -312500135;
assign addr[1244]= -350287041;
assign addr[1245]= -387962847;
assign addr[1246]= -425515602;
assign addr[1247]= -462933398;
assign addr[1248]= -500204365;
assign addr[1249]= -537316682;
assign addr[1250]= -574258580;
assign addr[1251]= -611018340;
assign addr[1252]= -647584304;
assign addr[1253]= -683944874;
assign addr[1254]= -720088517;
assign addr[1255]= -756003771;
assign addr[1256]= -791679244;
assign addr[1257]= -827103620;
assign addr[1258]= -862265664;
assign addr[1259]= -897154224;
assign addr[1260]= -931758235;
assign addr[1261]= -966066720;
assign addr[1262]= -1000068799;
assign addr[1263]= -1033753687;
assign addr[1264]= -1067110699;
assign addr[1265]= -1100129257;
assign addr[1266]= -1132798888;
assign addr[1267]= -1165109230;
assign addr[1268]= -1197050035;
assign addr[1269]= -1228611172;
assign addr[1270]= -1259782632;
assign addr[1271]= -1290554528;
assign addr[1272]= -1320917099;
assign addr[1273]= -1350860716;
assign addr[1274]= -1380375881;
assign addr[1275]= -1409453233;
assign addr[1276]= -1438083551;
assign addr[1277]= -1466257752;
assign addr[1278]= -1493966902;
assign addr[1279]= -1521202211;
assign addr[1280]= -1547955041;
assign addr[1281]= -1574216908;
assign addr[1282]= -1599979481;
assign addr[1283]= -1625234591;
assign addr[1284]= -1649974225;
assign addr[1285]= -1674190539;
assign addr[1286]= -1697875851;
assign addr[1287]= -1721022648;
assign addr[1288]= -1743623590;
assign addr[1289]= -1765671509;
assign addr[1290]= -1787159411;
assign addr[1291]= -1808080480;
assign addr[1292]= -1828428082;
assign addr[1293]= -1848195763;
assign addr[1294]= -1867377253;
assign addr[1295]= -1885966468;
assign addr[1296]= -1903957513;
assign addr[1297]= -1921344681;
assign addr[1298]= -1938122457;
assign addr[1299]= -1954285520;
assign addr[1300]= -1969828744;
assign addr[1301]= -1984747199;
assign addr[1302]= -1999036154;
assign addr[1303]= -2012691075;
assign addr[1304]= -2025707632;
assign addr[1305]= -2038081698;
assign addr[1306]= -2049809346;
assign addr[1307]= -2060886858;
assign addr[1308]= -2071310720;
assign addr[1309]= -2081077626;
assign addr[1310]= -2090184478;
assign addr[1311]= -2098628387;
assign addr[1312]= -2106406677;
assign addr[1313]= -2113516878;
assign addr[1314]= -2119956737;
assign addr[1315]= -2125724211;
assign addr[1316]= -2130817471;
assign addr[1317]= -2135234901;
assign addr[1318]= -2138975100;
assign addr[1319]= -2142036881;
assign addr[1320]= -2144419275;
assign addr[1321]= -2146121524;
assign addr[1322]= -2147143090;
assign addr[1323]= -2147483648;
assign addr[1324]= -2147143090;
assign addr[1325]= -2146121524;
assign addr[1326]= -2144419275;
assign addr[1327]= -2142036881;
assign addr[1328]= -2138975100;
assign addr[1329]= -2135234901;
assign addr[1330]= -2130817471;
assign addr[1331]= -2125724211;
assign addr[1332]= -2119956737;
assign addr[1333]= -2113516878;
assign addr[1334]= -2106406677;
assign addr[1335]= -2098628387;
assign addr[1336]= -2090184478;
assign addr[1337]= -2081077626;
assign addr[1338]= -2071310720;
assign addr[1339]= -2060886858;
assign addr[1340]= -2049809346;
assign addr[1341]= -2038081698;
assign addr[1342]= -2025707632;
assign addr[1343]= -2012691075;
assign addr[1344]= -1999036154;
assign addr[1345]= -1984747199;
assign addr[1346]= -1969828744;
assign addr[1347]= -1954285520;
assign addr[1348]= -1938122457;
assign addr[1349]= -1921344681;
assign addr[1350]= -1903957513;
assign addr[1351]= -1885966468;
assign addr[1352]= -1867377253;
assign addr[1353]= -1848195763;
assign addr[1354]= -1828428082;
assign addr[1355]= -1808080480;
assign addr[1356]= -1787159411;
assign addr[1357]= -1765671509;
assign addr[1358]= -1743623590;
assign addr[1359]= -1721022648;
assign addr[1360]= -1697875851;
assign addr[1361]= -1674190539;
assign addr[1362]= -1649974225;
assign addr[1363]= -1625234591;
assign addr[1364]= -1599979481;
assign addr[1365]= -1574216908;
assign addr[1366]= -1547955041;
assign addr[1367]= -1521202211;
assign addr[1368]= -1493966902;
assign addr[1369]= -1466257752;
assign addr[1370]= -1438083551;
assign addr[1371]= -1409453233;
assign addr[1372]= -1380375881;
assign addr[1373]= -1350860716;
assign addr[1374]= -1320917099;
assign addr[1375]= -1290554528;
assign addr[1376]= -1259782632;
assign addr[1377]= -1228611172;
assign addr[1378]= -1197050035;
assign addr[1379]= -1165109230;
assign addr[1380]= -1132798888;
assign addr[1381]= -1100129257;
assign addr[1382]= -1067110699;
assign addr[1383]= -1033753687;
assign addr[1384]= -1000068799;
assign addr[1385]= -966066720;
assign addr[1386]= -931758235;
assign addr[1387]= -897154224;
assign addr[1388]= -862265664;
assign addr[1389]= -827103620;
assign addr[1390]= -791679244;
assign addr[1391]= -756003771;
assign addr[1392]= -720088517;
assign addr[1393]= -683944874;
assign addr[1394]= -647584304;
assign addr[1395]= -611018340;
assign addr[1396]= -574258580;
assign addr[1397]= -537316682;
assign addr[1398]= -500204365;
assign addr[1399]= -462933398;
assign addr[1400]= -425515602;
assign addr[1401]= -387962847;
assign addr[1402]= -350287041;
assign addr[1403]= -312500135;
assign addr[1404]= -274614114;
assign addr[1405]= -236640993;
assign addr[1406]= -198592817;
assign addr[1407]= -160481654;
assign addr[1408]= -122319591;
assign addr[1409]= -84118732;
assign addr[1410]= -45891193;
assign addr[1411]= -7649098;
assign addr[1412]= 30595422;
assign addr[1413]= 68830239;
assign addr[1414]= 107043224;
assign addr[1415]= 145222259;
assign addr[1416]= 183355234;
assign addr[1417]= 221430054;
assign addr[1418]= 259434643;
assign addr[1419]= 297356948;
assign addr[1420]= 335184940;
assign addr[1421]= 372906622;
assign addr[1422]= 410510029;
assign addr[1423]= 447983235;
assign addr[1424]= 485314355;
assign addr[1425]= 522491548;
assign addr[1426]= 559503022;
assign addr[1427]= 596337040;
assign addr[1428]= 632981917;
assign addr[1429]= 669426032;
assign addr[1430]= 705657826;
assign addr[1431]= 741665807;
assign addr[1432]= 777438554;
assign addr[1433]= 812964722;
assign addr[1434]= 848233042;
assign addr[1435]= 883232329;
assign addr[1436]= 917951481;
assign addr[1437]= 952379488;
assign addr[1438]= 986505429;
assign addr[1439]= 1020318481;
assign addr[1440]= 1053807919;
assign addr[1441]= 1086963121;
assign addr[1442]= 1119773573;
assign addr[1443]= 1152228866;
assign addr[1444]= 1184318708;
assign addr[1445]= 1216032921;
assign addr[1446]= 1247361445;
assign addr[1447]= 1278294345;
assign addr[1448]= 1308821808;
assign addr[1449]= 1338934154;
assign addr[1450]= 1368621831;
assign addr[1451]= 1397875423;
assign addr[1452]= 1426685652;
assign addr[1453]= 1455043381;
assign addr[1454]= 1482939614;
assign addr[1455]= 1510365504;
assign addr[1456]= 1537312353;
assign addr[1457]= 1563771613;
assign addr[1458]= 1589734894;
assign addr[1459]= 1615193959;
assign addr[1460]= 1640140734;
assign addr[1461]= 1664567307;
assign addr[1462]= 1688465931;
assign addr[1463]= 1711829025;
assign addr[1464]= 1734649179;
assign addr[1465]= 1756919156;
assign addr[1466]= 1778631892;
assign addr[1467]= 1799780501;
assign addr[1468]= 1820358275;
assign addr[1469]= 1840358687;
assign addr[1470]= 1859775393;
assign addr[1471]= 1878602237;
assign addr[1472]= 1896833245;
assign addr[1473]= 1914462636;
assign addr[1474]= 1931484818;
assign addr[1475]= 1947894393;
assign addr[1476]= 1963686155;
assign addr[1477]= 1978855097;
assign addr[1478]= 1993396407;
assign addr[1479]= 2007305472;
assign addr[1480]= 2020577882;
assign addr[1481]= 2033209426;
assign addr[1482]= 2045196100;
assign addr[1483]= 2056534099;
assign addr[1484]= 2067219829;
assign addr[1485]= 2077249901;
assign addr[1486]= 2086621133;
assign addr[1487]= 2095330553;
assign addr[1488]= 2103375398;
assign addr[1489]= 2110753117;
assign addr[1490]= 2117461370;
assign addr[1491]= 2123498030;
assign addr[1492]= 2128861181;
assign addr[1493]= 2133549123;
assign addr[1494]= 2137560369;
assign addr[1495]= 2140893646;
assign addr[1496]= 2143547897;
assign addr[1497]= 2145522281;
assign addr[1498]= 2146816171;
assign addr[1499]= 2147429158;
assign addr[1500]= 2147361045;
assign addr[1501]= 2146611856;
assign addr[1502]= 2145181827;
assign addr[1503]= 2143071413;
assign addr[1504]= 2140281282;
assign addr[1505]= 2136812319;
assign addr[1506]= 2132665626;
assign addr[1507]= 2127842516;
assign addr[1508]= 2122344521;
assign addr[1509]= 2116173382;
assign addr[1510]= 2109331059;
assign addr[1511]= 2101819720;
assign addr[1512]= 2093641749;
assign addr[1513]= 2084799740;
assign addr[1514]= 2075296495;
assign addr[1515]= 2065135031;
assign addr[1516]= 2054318569;
assign addr[1517]= 2042850540;
assign addr[1518]= 2030734582;
assign addr[1519]= 2017974537;
assign addr[1520]= 2004574453;
assign addr[1521]= 1990538579;
assign addr[1522]= 1975871368;
assign addr[1523]= 1960577471;
assign addr[1524]= 1944661739;
assign addr[1525]= 1928129220;
assign addr[1526]= 1910985158;
assign addr[1527]= 1893234990;
assign addr[1528]= 1874884346;
assign addr[1529]= 1855939047;
assign addr[1530]= 1836405100;
assign addr[1531]= 1816288703;
assign addr[1532]= 1795596234;
assign addr[1533]= 1774334257;
assign addr[1534]= 1752509516;
assign addr[1535]= 1730128933;
assign addr[1536]= 1707199606;
assign addr[1537]= 1683728808;
assign addr[1538]= 1659723983;
assign addr[1539]= 1635192744;
assign addr[1540]= 1610142873;
assign addr[1541]= 1584582314;
assign addr[1542]= 1558519173;
assign addr[1543]= 1531961719;
assign addr[1544]= 1504918373;
assign addr[1545]= 1477397714;
assign addr[1546]= 1449408469;
assign addr[1547]= 1420959516;
assign addr[1548]= 1392059879;
assign addr[1549]= 1362718723;
assign addr[1550]= 1332945355;
assign addr[1551]= 1302749217;
assign addr[1552]= 1272139887;
assign addr[1553]= 1241127074;
assign addr[1554]= 1209720613;
assign addr[1555]= 1177930466;
assign addr[1556]= 1145766716;
assign addr[1557]= 1113239564;
assign addr[1558]= 1080359326;
assign addr[1559]= 1047136432;
assign addr[1560]= 1013581418;
assign addr[1561]= 979704927;
assign addr[1562]= 945517704;
assign addr[1563]= 911030591;
assign addr[1564]= 876254528;
assign addr[1565]= 841200544;
assign addr[1566]= 805879757;
assign addr[1567]= 770303369;
assign addr[1568]= 734482665;
assign addr[1569]= 698429006;
assign addr[1570]= 662153826;
assign addr[1571]= 625668632;
assign addr[1572]= 588984994;
assign addr[1573]= 552114549;
assign addr[1574]= 515068990;
assign addr[1575]= 477860067;
assign addr[1576]= 440499581;
assign addr[1577]= 402999383;
assign addr[1578]= 365371365;
assign addr[1579]= 327627463;
assign addr[1580]= 289779648;
assign addr[1581]= 251839923;
assign addr[1582]= 213820322;
assign addr[1583]= 175732905;
assign addr[1584]= 137589750;
assign addr[1585]= 99402956;
assign addr[1586]= 61184634;
assign addr[1587]= 22946906;
assign addr[1588]= -15298099;
assign addr[1589]= -53538253;
assign addr[1590]= -91761426;
assign addr[1591]= -129955495;
assign addr[1592]= -168108346;
assign addr[1593]= -206207878;
assign addr[1594]= -244242007;
assign addr[1595]= -282198671;
assign addr[1596]= -320065829;
assign addr[1597]= -357831473;
assign addr[1598]= -395483624;
assign addr[1599]= -433010339;
assign addr[1600]= -470399716;
assign addr[1601]= -507639898;
assign addr[1602]= -544719071;
assign addr[1603]= -581625477;
assign addr[1604]= -618347408;
assign addr[1605]= -654873219;
assign addr[1606]= -691191324;
assign addr[1607]= -727290205;
assign addr[1608]= -763158411;
assign addr[1609]= -798784567;
assign addr[1610]= -834157373;
assign addr[1611]= -869265610;
assign addr[1612]= -904098143;
assign addr[1613]= -938643924;
assign addr[1614]= -972891995;
assign addr[1615]= -1006831495;
assign addr[1616]= -1040451659;
assign addr[1617]= -1073741824;
assign addr[1618]= -1106691431;
assign addr[1619]= -1139290029;
assign addr[1620]= -1171527280;
assign addr[1621]= -1203392958;
assign addr[1622]= -1234876957;
assign addr[1623]= -1265969291;
assign addr[1624]= -1296660098;
assign addr[1625]= -1326939644;
assign addr[1626]= -1356798326;
assign addr[1627]= -1386226674;
assign addr[1628]= -1415215352;
assign addr[1629]= -1443755168;
assign addr[1630]= -1471837070;
assign addr[1631]= -1499452149;
assign addr[1632]= -1526591649;
assign addr[1633]= -1553246960;
assign addr[1634]= -1579409630;
assign addr[1635]= -1605071359;
assign addr[1636]= -1630224009;
assign addr[1637]= -1654859602;
assign addr[1638]= -1678970324;
assign addr[1639]= -1702548529;
assign addr[1640]= -1725586737;
assign addr[1641]= -1748077642;
assign addr[1642]= -1770014111;
assign addr[1643]= -1791389186;
assign addr[1644]= -1812196087;
assign addr[1645]= -1832428215;
assign addr[1646]= -1852079154;
assign addr[1647]= -1871142669;
assign addr[1648]= -1889612716;
assign addr[1649]= -1907483436;
assign addr[1650]= -1924749160;
assign addr[1651]= -1941404413;
assign addr[1652]= -1957443913;
assign addr[1653]= -1972862571;
assign addr[1654]= -1987655498;
assign addr[1655]= -2001818002;
assign addr[1656]= -2015345591;
assign addr[1657]= -2028233973;
assign addr[1658]= -2040479063;
assign addr[1659]= -2052076975;
assign addr[1660]= -2063024031;
assign addr[1661]= -2073316760;
assign addr[1662]= -2082951896;
assign addr[1663]= -2091926384;
assign addr[1664]= -2100237377;
assign addr[1665]= -2107882239;
assign addr[1666]= -2114858546;
assign addr[1667]= -2121164085;
assign addr[1668]= -2126796855;
assign addr[1669]= -2131755071;
assign addr[1670]= -2136037160;
assign addr[1671]= -2139641764;
assign addr[1672]= -2142567738;
assign addr[1673]= -2144814157;
assign addr[1674]= -2146380306;
assign addr[1675]= -2147265689;
assign addr[1676]= -2147470025;
assign addr[1677]= -2146993250;
assign addr[1678]= -2145835515;
assign addr[1679]= -2143997187;
assign addr[1680]= -2141478848;
assign addr[1681]= -2138281298;
assign addr[1682]= -2134405552;
assign addr[1683]= -2129852837;
assign addr[1684]= -2124624598;
assign addr[1685]= -2118722494;
assign addr[1686]= -2112148396;
assign addr[1687]= -2104904390;
assign addr[1688]= -2096992772;
assign addr[1689]= -2088416053;
assign addr[1690]= -2079176953;
assign addr[1691]= -2069278401;
assign addr[1692]= -2058723538;
assign addr[1693]= -2047515711;
assign addr[1694]= -2035658475;
assign addr[1695]= -2023155591;
assign addr[1696]= -2010011024;
assign addr[1697]= -1996228943;
assign addr[1698]= -1981813720;
assign addr[1699]= -1966769926;
assign addr[1700]= -1951102334;
assign addr[1701]= -1934815911;
assign addr[1702]= -1917915825;
assign addr[1703]= -1900407434;
assign addr[1704]= -1882296293;
assign addr[1705]= -1863588145;
assign addr[1706]= -1844288924;
assign addr[1707]= -1824404752;
assign addr[1708]= -1803941934;
assign addr[1709]= -1782906961;
assign addr[1710]= -1761306505;
assign addr[1711]= -1739147417;
assign addr[1712]= -1716436725;
assign addr[1713]= -1693181631;
assign addr[1714]= -1669389513;
assign addr[1715]= -1645067915;
assign addr[1716]= -1620224553;
assign addr[1717]= -1594867305;
assign addr[1718]= -1569004214;
assign addr[1719]= -1542643483;
assign addr[1720]= -1515793473;
assign addr[1721]= -1488462700;
assign addr[1722]= -1460659832;
assign addr[1723]= -1432393688;
assign addr[1724]= -1403673233;
assign addr[1725]= -1374507575;
assign addr[1726]= -1344905966;
assign addr[1727]= -1314877795;
assign addr[1728]= -1284432584;
assign addr[1729]= -1253579991;
assign addr[1730]= -1222329801;
assign addr[1731]= -1190691925;
assign addr[1732]= -1158676398;
assign addr[1733]= -1126293375;
assign addr[1734]= -1093553126;
assign addr[1735]= -1060466036;
assign addr[1736]= -1027042599;
assign addr[1737]= -993293415;
assign addr[1738]= -959229189;
assign addr[1739]= -924860725;
assign addr[1740]= -890198924;
assign addr[1741]= -855254778;
assign addr[1742]= -820039373;
assign addr[1743]= -784563876;
assign addr[1744]= -748839539;
assign addr[1745]= -712877694;
assign addr[1746]= -676689746;
assign addr[1747]= -640287172;
assign addr[1748]= -603681519;
assign addr[1749]= -566884397;
assign addr[1750]= -529907477;
assign addr[1751]= -492762486;
assign addr[1752]= -455461206;
assign addr[1753]= -418015468;
assign addr[1754]= -380437148;
assign addr[1755]= -342738165;
assign addr[1756]= -304930476;
assign addr[1757]= -267026072;
assign addr[1758]= -229036977;
assign addr[1759]= -190975237;
assign addr[1760]= -152852926;
assign addr[1761]= -114682135;
assign addr[1762]= -76474970;
assign addr[1763]= -38243550;
assign addr[1764]= 0;
assign addr[1765]= 38243550;
assign addr[1766]= 76474970;
assign addr[1767]= 114682135;
assign addr[1768]= 152852926;
assign addr[1769]= 190975237;
assign addr[1770]= 229036977;
assign addr[1771]= 267026072;
assign addr[1772]= 304930476;
assign addr[1773]= 342738165;
assign addr[1774]= 380437148;
assign addr[1775]= 418015468;
assign addr[1776]= 455461206;
assign addr[1777]= 492762486;
assign addr[1778]= 529907477;
assign addr[1779]= 566884397;
assign addr[1780]= 603681519;
assign addr[1781]= 640287172;
assign addr[1782]= 676689746;
assign addr[1783]= 712877694;
assign addr[1784]= 748839539;
assign addr[1785]= 784563876;
assign addr[1786]= 820039373;
assign addr[1787]= 855254778;
assign addr[1788]= 890198924;
assign addr[1789]= 924860725;
assign addr[1790]= 959229189;
assign addr[1791]= 993293415;
assign addr[1792]= 1027042599;
assign addr[1793]= 1060466036;
assign addr[1794]= 1093553126;
assign addr[1795]= 1126293375;
assign addr[1796]= 1158676398;
assign addr[1797]= 1190691925;
assign addr[1798]= 1222329801;
assign addr[1799]= 1253579991;
assign addr[1800]= 1284432584;
assign addr[1801]= 1314877795;
assign addr[1802]= 1344905966;
assign addr[1803]= 1374507575;
assign addr[1804]= 1403673233;
assign addr[1805]= 1432393688;
assign addr[1806]= 1460659832;
assign addr[1807]= 1488462700;
assign addr[1808]= 1515793473;
assign addr[1809]= 1542643483;
assign addr[1810]= 1569004214;
assign addr[1811]= 1594867305;
assign addr[1812]= 1620224553;
assign addr[1813]= 1645067915;
assign addr[1814]= 1669389513;
assign addr[1815]= 1693181631;
assign addr[1816]= 1716436725;
assign addr[1817]= 1739147417;
assign addr[1818]= 1761306505;
assign addr[1819]= 1782906961;
assign addr[1820]= 1803941934;
assign addr[1821]= 1824404752;
assign addr[1822]= 1844288924;
assign addr[1823]= 1863588145;
assign addr[1824]= 1882296293;
assign addr[1825]= 1900407434;
assign addr[1826]= 1917915825;
assign addr[1827]= 1934815911;
assign addr[1828]= 1951102334;
assign addr[1829]= 1966769926;
assign addr[1830]= 1981813720;
assign addr[1831]= 1996228943;
assign addr[1832]= 2010011024;
assign addr[1833]= 2023155591;
assign addr[1834]= 2035658475;
assign addr[1835]= 2047515711;
assign addr[1836]= 2058723538;
assign addr[1837]= 2069278401;
assign addr[1838]= 2079176953;
assign addr[1839]= 2088416053;
assign addr[1840]= 2096992772;
assign addr[1841]= 2104904390;
assign addr[1842]= 2112148396;
assign addr[1843]= 2118722494;
assign addr[1844]= 2124624598;
assign addr[1845]= 2129852837;
assign addr[1846]= 2134405552;
assign addr[1847]= 2138281298;
assign addr[1848]= 2141478848;
assign addr[1849]= 2143997187;
assign addr[1850]= 2145835515;
assign addr[1851]= 2146993250;
assign addr[1852]= 2147470025;
assign addr[1853]= 2147265689;
assign addr[1854]= 2146380306;
assign addr[1855]= 2144814157;
assign addr[1856]= 2142567738;
assign addr[1857]= 2139641764;
assign addr[1858]= 2136037160;
assign addr[1859]= 2131755071;
assign addr[1860]= 2126796855;
assign addr[1861]= 2121164085;
assign addr[1862]= 2114858546;
assign addr[1863]= 2107882239;
assign addr[1864]= 2100237377;
assign addr[1865]= 2091926384;
assign addr[1866]= 2082951896;
assign addr[1867]= 2073316760;
assign addr[1868]= 2063024031;
assign addr[1869]= 2052076975;
assign addr[1870]= 2040479063;
assign addr[1871]= 2028233973;
assign addr[1872]= 2015345591;
assign addr[1873]= 2001818002;
assign addr[1874]= 1987655498;
assign addr[1875]= 1972862571;
assign addr[1876]= 1957443913;
assign addr[1877]= 1941404413;
assign addr[1878]= 1924749160;
assign addr[1879]= 1907483436;
assign addr[1880]= 1889612716;
assign addr[1881]= 1871142669;
assign addr[1882]= 1852079154;
assign addr[1883]= 1832428215;
assign addr[1884]= 1812196087;
assign addr[1885]= 1791389186;
assign addr[1886]= 1770014111;
assign addr[1887]= 1748077642;
assign addr[1888]= 1725586737;
assign addr[1889]= 1702548529;
assign addr[1890]= 1678970324;
assign addr[1891]= 1654859602;
assign addr[1892]= 1630224009;
assign addr[1893]= 1605071359;
assign addr[1894]= 1579409630;
assign addr[1895]= 1553246960;
assign addr[1896]= 1526591649;
assign addr[1897]= 1499452149;
assign addr[1898]= 1471837070;
assign addr[1899]= 1443755168;
assign addr[1900]= 1415215352;
assign addr[1901]= 1386226674;
assign addr[1902]= 1356798326;
assign addr[1903]= 1326939644;
assign addr[1904]= 1296660098;
assign addr[1905]= 1265969291;
assign addr[1906]= 1234876957;
assign addr[1907]= 1203392958;
assign addr[1908]= 1171527280;
assign addr[1909]= 1139290029;
assign addr[1910]= 1106691431;
assign addr[1911]= 1073741824;
assign addr[1912]= 1040451659;
assign addr[1913]= 1006831495;
assign addr[1914]= 972891995;
assign addr[1915]= 938643924;
assign addr[1916]= 904098143;
assign addr[1917]= 869265610;
assign addr[1918]= 834157373;
assign addr[1919]= 798784567;
assign addr[1920]= 763158411;
assign addr[1921]= 727290205;
assign addr[1922]= 691191324;
assign addr[1923]= 654873219;
assign addr[1924]= 618347408;
assign addr[1925]= 581625477;
assign addr[1926]= 544719071;
assign addr[1927]= 507639898;
assign addr[1928]= 470399716;
assign addr[1929]= 433010339;
assign addr[1930]= 395483624;
assign addr[1931]= 357831473;
assign addr[1932]= 320065829;
assign addr[1933]= 282198671;
assign addr[1934]= 244242007;
assign addr[1935]= 206207878;
assign addr[1936]= 168108346;
assign addr[1937]= 129955495;
assign addr[1938]= 91761426;
assign addr[1939]= 53538253;
assign addr[1940]= 15298099;
assign addr[1941]= -22946906;
assign addr[1942]= -61184634;
assign addr[1943]= -99402956;
assign addr[1944]= -137589750;
assign addr[1945]= -175732905;
assign addr[1946]= -213820322;
assign addr[1947]= -251839923;
assign addr[1948]= -289779648;
assign addr[1949]= -327627463;
assign addr[1950]= -365371365;
assign addr[1951]= -402999383;
assign addr[1952]= -440499581;
assign addr[1953]= -477860067;
assign addr[1954]= -515068990;
assign addr[1955]= -552114549;
assign addr[1956]= -588984994;
assign addr[1957]= -625668632;
assign addr[1958]= -662153826;
assign addr[1959]= -698429006;
assign addr[1960]= -734482665;
assign addr[1961]= -770303369;
assign addr[1962]= -805879757;
assign addr[1963]= -841200544;
assign addr[1964]= -876254528;
assign addr[1965]= -911030591;
assign addr[1966]= -945517704;
assign addr[1967]= -979704927;
assign addr[1968]= -1013581418;
assign addr[1969]= -1047136432;
assign addr[1970]= -1080359326;
assign addr[1971]= -1113239564;
assign addr[1972]= -1145766716;
assign addr[1973]= -1177930466;
assign addr[1974]= -1209720613;
assign addr[1975]= -1241127074;
assign addr[1976]= -1272139887;
assign addr[1977]= -1302749217;
assign addr[1978]= -1332945355;
assign addr[1979]= -1362718723;
assign addr[1980]= -1392059879;
assign addr[1981]= -1420959516;
assign addr[1982]= -1449408469;
assign addr[1983]= -1477397714;
assign addr[1984]= -1504918373;
assign addr[1985]= -1531961719;
assign addr[1986]= -1558519173;
assign addr[1987]= -1584582314;
assign addr[1988]= -1610142873;
assign addr[1989]= -1635192744;
assign addr[1990]= -1659723983;
assign addr[1991]= -1683728808;
assign addr[1992]= -1707199606;
assign addr[1993]= -1730128933;
assign addr[1994]= -1752509516;
assign addr[1995]= -1774334257;
assign addr[1996]= -1795596234;
assign addr[1997]= -1816288703;
assign addr[1998]= -1836405100;
assign addr[1999]= -1855939047;
assign addr[2000]= -1874884346;
assign addr[2001]= -1893234990;
assign addr[2002]= -1910985158;
assign addr[2003]= -1928129220;
assign addr[2004]= -1944661739;
assign addr[2005]= -1960577471;
assign addr[2006]= -1975871368;
assign addr[2007]= -1990538579;
assign addr[2008]= -2004574453;
assign addr[2009]= -2017974537;
assign addr[2010]= -2030734582;
assign addr[2011]= -2042850540;
assign addr[2012]= -2054318569;
assign addr[2013]= -2065135031;
assign addr[2014]= -2075296495;
assign addr[2015]= -2084799740;
assign addr[2016]= -2093641749;
assign addr[2017]= -2101819720;
assign addr[2018]= -2109331059;
assign addr[2019]= -2116173382;
assign addr[2020]= -2122344521;
assign addr[2021]= -2127842516;
assign addr[2022]= -2132665626;
assign addr[2023]= -2136812319;
assign addr[2024]= -2140281282;
assign addr[2025]= -2143071413;
assign addr[2026]= -2145181827;
assign addr[2027]= -2146611856;
assign addr[2028]= -2147361045;
assign addr[2029]= -2147429158;
assign addr[2030]= -2146816171;
assign addr[2031]= -2145522281;
assign addr[2032]= -2143547897;
assign addr[2033]= -2140893646;
assign addr[2034]= -2137560369;
assign addr[2035]= -2133549123;
assign addr[2036]= -2128861181;
assign addr[2037]= -2123498030;
assign addr[2038]= -2117461370;
assign addr[2039]= -2110753117;
assign addr[2040]= -2103375398;
assign addr[2041]= -2095330553;
assign addr[2042]= -2086621133;
assign addr[2043]= -2077249901;
assign addr[2044]= -2067219829;
assign addr[2045]= -2056534099;
assign addr[2046]= -2045196100;
assign addr[2047]= -2033209426;
assign addr[2048]= -2020577882;
assign addr[2049]= -2007305472;
assign addr[2050]= -1993396407;
assign addr[2051]= -1978855097;
assign addr[2052]= -1963686155;
assign addr[2053]= -1947894393;
assign addr[2054]= -1931484818;
assign addr[2055]= -1914462636;
assign addr[2056]= -1896833245;
assign addr[2057]= -1878602237;
assign addr[2058]= -1859775393;
assign addr[2059]= -1840358687;
assign addr[2060]= -1820358275;
assign addr[2061]= -1799780501;
assign addr[2062]= -1778631892;
assign addr[2063]= -1756919156;
assign addr[2064]= -1734649179;
assign addr[2065]= -1711829025;
assign addr[2066]= -1688465931;
assign addr[2067]= -1664567307;
assign addr[2068]= -1640140734;
assign addr[2069]= -1615193959;
assign addr[2070]= -1589734894;
assign addr[2071]= -1563771613;
assign addr[2072]= -1537312353;
assign addr[2073]= -1510365504;
assign addr[2074]= -1482939614;
assign addr[2075]= -1455043381;
assign addr[2076]= -1426685652;
assign addr[2077]= -1397875423;
assign addr[2078]= -1368621831;
assign addr[2079]= -1338934154;
assign addr[2080]= -1308821808;
assign addr[2081]= -1278294345;
assign addr[2082]= -1247361445;
assign addr[2083]= -1216032921;
assign addr[2084]= -1184318708;
assign addr[2085]= -1152228866;
assign addr[2086]= -1119773573;
assign addr[2087]= -1086963121;
assign addr[2088]= -1053807919;
assign addr[2089]= -1020318481;
assign addr[2090]= -986505429;
assign addr[2091]= -952379488;
assign addr[2092]= -917951481;
assign addr[2093]= -883232329;
assign addr[2094]= -848233042;
assign addr[2095]= -812964722;
assign addr[2096]= -777438554;
assign addr[2097]= -741665807;
assign addr[2098]= -705657826;
assign addr[2099]= -669426032;
assign addr[2100]= -632981917;
assign addr[2101]= -596337040;
assign addr[2102]= -559503022;
assign addr[2103]= -522491548;
assign addr[2104]= -485314355;
assign addr[2105]= -447983235;
assign addr[2106]= -410510029;
assign addr[2107]= -372906622;
assign addr[2108]= -335184940;
assign addr[2109]= -297356948;
assign addr[2110]= -259434643;
assign addr[2111]= -221430054;
assign addr[2112]= -183355234;
assign addr[2113]= -145222259;
assign addr[2114]= -107043224;
assign addr[2115]= -68830239;
assign addr[2116]= -30595422;
assign addr[2117]= 7649098;
assign addr[2118]= 45891193;
assign addr[2119]= 84118732;
assign addr[2120]= 122319591;
assign addr[2121]= 160481654;
assign addr[2122]= 198592817;
assign addr[2123]= 236640993;
assign addr[2124]= 274614114;
assign addr[2125]= 312500135;
assign addr[2126]= 350287041;
assign addr[2127]= 387962847;
assign addr[2128]= 425515602;
assign addr[2129]= 462933398;
assign addr[2130]= 500204365;
assign addr[2131]= 537316682;
assign addr[2132]= 574258580;
assign addr[2133]= 611018340;
assign addr[2134]= 647584304;
assign addr[2135]= 683944874;
assign addr[2136]= 720088517;
assign addr[2137]= 756003771;
assign addr[2138]= 791679244;
assign addr[2139]= 827103620;
assign addr[2140]= 862265664;
assign addr[2141]= 897154224;
assign addr[2142]= 931758235;
assign addr[2143]= 966066720;
assign addr[2144]= 1000068799;
assign addr[2145]= 1033753687;
assign addr[2146]= 1067110699;
assign addr[2147]= 1100129257;
assign addr[2148]= 1132798888;
assign addr[2149]= 1165109230;
assign addr[2150]= 1197050035;
assign addr[2151]= 1228611172;
assign addr[2152]= 1259782632;
assign addr[2153]= 1290554528;
assign addr[2154]= 1320917099;
assign addr[2155]= 1350860716;
assign addr[2156]= 1380375881;
assign addr[2157]= 1409453233;
assign addr[2158]= 1438083551;
assign addr[2159]= 1466257752;
assign addr[2160]= 1493966902;
assign addr[2161]= 1521202211;
assign addr[2162]= 1547955041;
assign addr[2163]= 1574216908;
assign addr[2164]= 1599979481;
assign addr[2165]= 1625234591;
assign addr[2166]= 1649974225;
assign addr[2167]= 1674190539;
assign addr[2168]= 1697875851;
assign addr[2169]= 1721022648;
assign addr[2170]= 1743623590;
assign addr[2171]= 1765671509;
assign addr[2172]= 1787159411;
assign addr[2173]= 1808080480;
assign addr[2174]= 1828428082;
assign addr[2175]= 1848195763;
assign addr[2176]= 1867377253;
assign addr[2177]= 1885966468;
assign addr[2178]= 1903957513;
assign addr[2179]= 1921344681;
assign addr[2180]= 1938122457;
assign addr[2181]= 1954285520;
assign addr[2182]= 1969828744;
assign addr[2183]= 1984747199;
assign addr[2184]= 1999036154;
assign addr[2185]= 2012691075;
assign addr[2186]= 2025707632;
assign addr[2187]= 2038081698;
assign addr[2188]= 2049809346;
assign addr[2189]= 2060886858;
assign addr[2190]= 2071310720;
assign addr[2191]= 2081077626;
assign addr[2192]= 2090184478;
assign addr[2193]= 2098628387;
assign addr[2194]= 2106406677;
assign addr[2195]= 2113516878;
assign addr[2196]= 2119956737;
assign addr[2197]= 2125724211;
assign addr[2198]= 2130817471;
assign addr[2199]= 2135234901;
assign addr[2200]= 2138975100;
assign addr[2201]= 2142036881;
assign addr[2202]= 2144419275;
assign addr[2203]= 2146121524;
assign addr[2204]= 2147143090;
assign addr[2205]= 2147483648;
assign addr[2206]= 2147143090;
assign addr[2207]= 2146121524;
assign addr[2208]= 2144419275;
assign addr[2209]= 2142036881;
assign addr[2210]= 2138975100;
assign addr[2211]= 2135234901;
assign addr[2212]= 2130817471;
assign addr[2213]= 2125724211;
assign addr[2214]= 2119956737;
assign addr[2215]= 2113516878;
assign addr[2216]= 2106406677;
assign addr[2217]= 2098628387;
assign addr[2218]= 2090184478;
assign addr[2219]= 2081077626;
assign addr[2220]= 2071310720;
assign addr[2221]= 2060886858;
assign addr[2222]= 2049809346;
assign addr[2223]= 2038081698;
assign addr[2224]= 2025707632;
assign addr[2225]= 2012691075;
assign addr[2226]= 1999036154;
assign addr[2227]= 1984747199;
assign addr[2228]= 1969828744;
assign addr[2229]= 1954285520;
assign addr[2230]= 1938122457;
assign addr[2231]= 1921344681;
assign addr[2232]= 1903957513;
assign addr[2233]= 1885966468;
assign addr[2234]= 1867377253;
assign addr[2235]= 1848195763;
assign addr[2236]= 1828428082;
assign addr[2237]= 1808080480;
assign addr[2238]= 1787159411;
assign addr[2239]= 1765671509;
assign addr[2240]= 1743623590;
assign addr[2241]= 1721022648;
assign addr[2242]= 1697875851;
assign addr[2243]= 1674190539;
assign addr[2244]= 1649974225;
assign addr[2245]= 1625234591;
assign addr[2246]= 1599979481;
assign addr[2247]= 1574216908;
assign addr[2248]= 1547955041;
assign addr[2249]= 1521202211;
assign addr[2250]= 1493966902;
assign addr[2251]= 1466257752;
assign addr[2252]= 1438083551;
assign addr[2253]= 1409453233;
assign addr[2254]= 1380375881;
assign addr[2255]= 1350860716;
assign addr[2256]= 1320917099;
assign addr[2257]= 1290554528;
assign addr[2258]= 1259782632;
assign addr[2259]= 1228611172;
assign addr[2260]= 1197050035;
assign addr[2261]= 1165109230;
assign addr[2262]= 1132798888;
assign addr[2263]= 1100129257;
assign addr[2264]= 1067110699;
assign addr[2265]= 1033753687;
assign addr[2266]= 1000068799;
assign addr[2267]= 966066720;
assign addr[2268]= 931758235;
assign addr[2269]= 897154224;
assign addr[2270]= 862265664;
assign addr[2271]= 827103620;
assign addr[2272]= 791679244;
assign addr[2273]= 756003771;
assign addr[2274]= 720088517;
assign addr[2275]= 683944874;
assign addr[2276]= 647584304;
assign addr[2277]= 611018340;
assign addr[2278]= 574258580;
assign addr[2279]= 537316682;
assign addr[2280]= 500204365;
assign addr[2281]= 462933398;
assign addr[2282]= 425515602;
assign addr[2283]= 387962847;
assign addr[2284]= 350287041;
assign addr[2285]= 312500135;
assign addr[2286]= 274614114;
assign addr[2287]= 236640993;
assign addr[2288]= 198592817;
assign addr[2289]= 160481654;
assign addr[2290]= 122319591;
assign addr[2291]= 84118732;
assign addr[2292]= 45891193;
assign addr[2293]= 7649098;
assign addr[2294]= -30595422;
assign addr[2295]= -68830239;
assign addr[2296]= -107043224;
assign addr[2297]= -145222259;
assign addr[2298]= -183355234;
assign addr[2299]= -221430054;
assign addr[2300]= -259434643;
assign addr[2301]= -297356948;
assign addr[2302]= -335184940;
assign addr[2303]= -372906622;
assign addr[2304]= -410510029;
assign addr[2305]= -447983235;
assign addr[2306]= -485314355;
assign addr[2307]= -522491548;
assign addr[2308]= -559503022;
assign addr[2309]= -596337040;
assign addr[2310]= -632981917;
assign addr[2311]= -669426032;
assign addr[2312]= -705657826;
assign addr[2313]= -741665807;
assign addr[2314]= -777438554;
assign addr[2315]= -812964722;
assign addr[2316]= -848233042;
assign addr[2317]= -883232329;
assign addr[2318]= -917951481;
assign addr[2319]= -952379488;
assign addr[2320]= -986505429;
assign addr[2321]= -1020318481;
assign addr[2322]= -1053807919;
assign addr[2323]= -1086963121;
assign addr[2324]= -1119773573;
assign addr[2325]= -1152228866;
assign addr[2326]= -1184318708;
assign addr[2327]= -1216032921;
assign addr[2328]= -1247361445;
assign addr[2329]= -1278294345;
assign addr[2330]= -1308821808;
assign addr[2331]= -1338934154;
assign addr[2332]= -1368621831;
assign addr[2333]= -1397875423;
assign addr[2334]= -1426685652;
assign addr[2335]= -1455043381;
assign addr[2336]= -1482939614;
assign addr[2337]= -1510365504;
assign addr[2338]= -1537312353;
assign addr[2339]= -1563771613;
assign addr[2340]= -1589734894;
assign addr[2341]= -1615193959;
assign addr[2342]= -1640140734;
assign addr[2343]= -1664567307;
assign addr[2344]= -1688465931;
assign addr[2345]= -1711829025;
assign addr[2346]= -1734649179;
assign addr[2347]= -1756919156;
assign addr[2348]= -1778631892;
assign addr[2349]= -1799780501;
assign addr[2350]= -1820358275;
assign addr[2351]= -1840358687;
assign addr[2352]= -1859775393;
assign addr[2353]= -1878602237;
assign addr[2354]= -1896833245;
assign addr[2355]= -1914462636;
assign addr[2356]= -1931484818;
assign addr[2357]= -1947894393;
assign addr[2358]= -1963686155;
assign addr[2359]= -1978855097;
assign addr[2360]= -1993396407;
assign addr[2361]= -2007305472;
assign addr[2362]= -2020577882;
assign addr[2363]= -2033209426;
assign addr[2364]= -2045196100;
assign addr[2365]= -2056534099;
assign addr[2366]= -2067219829;
assign addr[2367]= -2077249901;
assign addr[2368]= -2086621133;
assign addr[2369]= -2095330553;
assign addr[2370]= -2103375398;
assign addr[2371]= -2110753117;
assign addr[2372]= -2117461370;
assign addr[2373]= -2123498030;
assign addr[2374]= -2128861181;
assign addr[2375]= -2133549123;
assign addr[2376]= -2137560369;
assign addr[2377]= -2140893646;
assign addr[2378]= -2143547897;
assign addr[2379]= -2145522281;
assign addr[2380]= -2146816171;
assign addr[2381]= -2147429158;
assign addr[2382]= -2147361045;
assign addr[2383]= -2146611856;
assign addr[2384]= -2145181827;
assign addr[2385]= -2143071413;
assign addr[2386]= -2140281282;
assign addr[2387]= -2136812319;
assign addr[2388]= -2132665626;
assign addr[2389]= -2127842516;
assign addr[2390]= -2122344521;
assign addr[2391]= -2116173382;
assign addr[2392]= -2109331059;
assign addr[2393]= -2101819720;
assign addr[2394]= -2093641749;
assign addr[2395]= -2084799740;
assign addr[2396]= -2075296495;
assign addr[2397]= -2065135031;
assign addr[2398]= -2054318569;
assign addr[2399]= -2042850540;
assign addr[2400]= -2030734582;
assign addr[2401]= -2017974537;
assign addr[2402]= -2004574453;
assign addr[2403]= -1990538579;
assign addr[2404]= -1975871368;
assign addr[2405]= -1960577471;
assign addr[2406]= -1944661739;
assign addr[2407]= -1928129220;
assign addr[2408]= -1910985158;
assign addr[2409]= -1893234990;
assign addr[2410]= -1874884346;
assign addr[2411]= -1855939047;
assign addr[2412]= -1836405100;
assign addr[2413]= -1816288703;
assign addr[2414]= -1795596234;
assign addr[2415]= -1774334257;
assign addr[2416]= -1752509516;
assign addr[2417]= -1730128933;
assign addr[2418]= -1707199606;
assign addr[2419]= -1683728808;
assign addr[2420]= -1659723983;
assign addr[2421]= -1635192744;
assign addr[2422]= -1610142873;
assign addr[2423]= -1584582314;
assign addr[2424]= -1558519173;
assign addr[2425]= -1531961719;
assign addr[2426]= -1504918373;
assign addr[2427]= -1477397714;
assign addr[2428]= -1449408469;
assign addr[2429]= -1420959516;
assign addr[2430]= -1392059879;
assign addr[2431]= -1362718723;
assign addr[2432]= -1332945355;
assign addr[2433]= -1302749217;
assign addr[2434]= -1272139887;
assign addr[2435]= -1241127074;
assign addr[2436]= -1209720613;
assign addr[2437]= -1177930466;
assign addr[2438]= -1145766716;
assign addr[2439]= -1113239564;
assign addr[2440]= -1080359326;
assign addr[2441]= -1047136432;
assign addr[2442]= -1013581418;
assign addr[2443]= -979704927;
assign addr[2444]= -945517704;
assign addr[2445]= -911030591;
assign addr[2446]= -876254528;
assign addr[2447]= -841200544;
assign addr[2448]= -805879757;
assign addr[2449]= -770303369;
assign addr[2450]= -734482665;
assign addr[2451]= -698429006;
assign addr[2452]= -662153826;
assign addr[2453]= -625668632;
assign addr[2454]= -588984994;
assign addr[2455]= -552114549;
assign addr[2456]= -515068990;
assign addr[2457]= -477860067;
assign addr[2458]= -440499581;
assign addr[2459]= -402999383;
assign addr[2460]= -365371365;
assign addr[2461]= -327627463;
assign addr[2462]= -289779648;
assign addr[2463]= -251839923;
assign addr[2464]= -213820322;
assign addr[2465]= -175732905;
assign addr[2466]= -137589750;
assign addr[2467]= -99402956;
assign addr[2468]= -61184634;
assign addr[2469]= -22946906;
assign addr[2470]= 15298099;
assign addr[2471]= 53538253;
assign addr[2472]= 91761426;
assign addr[2473]= 129955495;
assign addr[2474]= 168108346;
assign addr[2475]= 206207878;
assign addr[2476]= 244242007;
assign addr[2477]= 282198671;
assign addr[2478]= 320065829;
assign addr[2479]= 357831473;
assign addr[2480]= 395483624;
assign addr[2481]= 433010339;
assign addr[2482]= 470399716;
assign addr[2483]= 507639898;
assign addr[2484]= 544719071;
assign addr[2485]= 581625477;
assign addr[2486]= 618347408;
assign addr[2487]= 654873219;
assign addr[2488]= 691191324;
assign addr[2489]= 727290205;
assign addr[2490]= 763158411;
assign addr[2491]= 798784567;
assign addr[2492]= 834157373;
assign addr[2493]= 869265610;
assign addr[2494]= 904098143;
assign addr[2495]= 938643924;
assign addr[2496]= 972891995;
assign addr[2497]= 1006831495;
assign addr[2498]= 1040451659;
assign addr[2499]= 1073741824;
assign addr[2500]= 1106691431;
assign addr[2501]= 1139290029;
assign addr[2502]= 1171527280;
assign addr[2503]= 1203392958;
assign addr[2504]= 1234876957;
assign addr[2505]= 1265969291;
assign addr[2506]= 1296660098;
assign addr[2507]= 1326939644;
assign addr[2508]= 1356798326;
assign addr[2509]= 1386226674;
assign addr[2510]= 1415215352;
assign addr[2511]= 1443755168;
assign addr[2512]= 1471837070;
assign addr[2513]= 1499452149;
assign addr[2514]= 1526591649;
assign addr[2515]= 1553246960;
assign addr[2516]= 1579409630;
assign addr[2517]= 1605071359;
assign addr[2518]= 1630224009;
assign addr[2519]= 1654859602;
assign addr[2520]= 1678970324;
assign addr[2521]= 1702548529;
assign addr[2522]= 1725586737;
assign addr[2523]= 1748077642;
assign addr[2524]= 1770014111;
assign addr[2525]= 1791389186;
assign addr[2526]= 1812196087;
assign addr[2527]= 1832428215;
assign addr[2528]= 1852079154;
assign addr[2529]= 1871142669;
assign addr[2530]= 1889612716;
assign addr[2531]= 1907483436;
assign addr[2532]= 1924749160;
assign addr[2533]= 1941404413;
assign addr[2534]= 1957443913;
assign addr[2535]= 1972862571;
assign addr[2536]= 1987655498;
assign addr[2537]= 2001818002;
assign addr[2538]= 2015345591;
assign addr[2539]= 2028233973;
assign addr[2540]= 2040479063;
assign addr[2541]= 2052076975;
assign addr[2542]= 2063024031;
assign addr[2543]= 2073316760;
assign addr[2544]= 2082951896;
assign addr[2545]= 2091926384;
assign addr[2546]= 2100237377;
assign addr[2547]= 2107882239;
assign addr[2548]= 2114858546;
assign addr[2549]= 2121164085;
assign addr[2550]= 2126796855;
assign addr[2551]= 2131755071;
assign addr[2552]= 2136037160;
assign addr[2553]= 2139641764;
assign addr[2554]= 2142567738;
assign addr[2555]= 2144814157;
assign addr[2556]= 2146380306;
assign addr[2557]= 2147265689;
assign addr[2558]= 2147470025;
assign addr[2559]= 2146993250;
assign addr[2560]= 2145835515;
assign addr[2561]= 2143997187;
assign addr[2562]= 2141478848;
assign addr[2563]= 2138281298;
assign addr[2564]= 2134405552;
assign addr[2565]= 2129852837;
assign addr[2566]= 2124624598;
assign addr[2567]= 2118722494;
assign addr[2568]= 2112148396;
assign addr[2569]= 2104904390;
assign addr[2570]= 2096992772;
assign addr[2571]= 2088416053;
assign addr[2572]= 2079176953;
assign addr[2573]= 2069278401;
assign addr[2574]= 2058723538;
assign addr[2575]= 2047515711;
assign addr[2576]= 2035658475;
assign addr[2577]= 2023155591;
assign addr[2578]= 2010011024;
assign addr[2579]= 1996228943;
assign addr[2580]= 1981813720;
assign addr[2581]= 1966769926;
assign addr[2582]= 1951102334;
assign addr[2583]= 1934815911;
assign addr[2584]= 1917915825;
assign addr[2585]= 1900407434;
assign addr[2586]= 1882296293;
assign addr[2587]= 1863588145;
assign addr[2588]= 1844288924;
assign addr[2589]= 1824404752;
assign addr[2590]= 1803941934;
assign addr[2591]= 1782906961;
assign addr[2592]= 1761306505;
assign addr[2593]= 1739147417;
assign addr[2594]= 1716436725;
assign addr[2595]= 1693181631;
assign addr[2596]= 1669389513;
assign addr[2597]= 1645067915;
assign addr[2598]= 1620224553;
assign addr[2599]= 1594867305;
assign addr[2600]= 1569004214;
assign addr[2601]= 1542643483;
assign addr[2602]= 1515793473;
assign addr[2603]= 1488462700;
assign addr[2604]= 1460659832;
assign addr[2605]= 1432393688;
assign addr[2606]= 1403673233;
assign addr[2607]= 1374507575;
assign addr[2608]= 1344905966;
assign addr[2609]= 1314877795;
assign addr[2610]= 1284432584;
assign addr[2611]= 1253579991;
assign addr[2612]= 1222329801;
assign addr[2613]= 1190691925;
assign addr[2614]= 1158676398;
assign addr[2615]= 1126293375;
assign addr[2616]= 1093553126;
assign addr[2617]= 1060466036;
assign addr[2618]= 1027042599;
assign addr[2619]= 993293415;
assign addr[2620]= 959229189;
assign addr[2621]= 924860725;
assign addr[2622]= 890198924;
assign addr[2623]= 855254778;
assign addr[2624]= 820039373;
assign addr[2625]= 784563876;
assign addr[2626]= 748839539;
assign addr[2627]= 712877694;
assign addr[2628]= 676689746;
assign addr[2629]= 640287172;
assign addr[2630]= 603681519;
assign addr[2631]= 566884397;
assign addr[2632]= 529907477;
assign addr[2633]= 492762486;
assign addr[2634]= 455461206;
assign addr[2635]= 418015468;
assign addr[2636]= 380437148;
assign addr[2637]= 342738165;
assign addr[2638]= 304930476;
assign addr[2639]= 267026072;
assign addr[2640]= 229036977;
assign addr[2641]= 190975237;
assign addr[2642]= 152852926;
assign addr[2643]= 114682135;
assign addr[2644]= 76474970;
assign addr[2645]= 38243550;
assign addr[2646]= 0;
assign addr[2647]= -38243550;
assign addr[2648]= -76474970;
assign addr[2649]= -114682135;
assign addr[2650]= -152852926;
assign addr[2651]= -190975237;
assign addr[2652]= -229036977;
assign addr[2653]= -267026072;
assign addr[2654]= -304930476;
assign addr[2655]= -342738165;
assign addr[2656]= -380437148;
assign addr[2657]= -418015468;
assign addr[2658]= -455461206;
assign addr[2659]= -492762486;
assign addr[2660]= -529907477;
assign addr[2661]= -566884397;
assign addr[2662]= -603681519;
assign addr[2663]= -640287172;
assign addr[2664]= -676689746;
assign addr[2665]= -712877694;
assign addr[2666]= -748839539;
assign addr[2667]= -784563876;
assign addr[2668]= -820039373;
assign addr[2669]= -855254778;
assign addr[2670]= -890198924;
assign addr[2671]= -924860725;
assign addr[2672]= -959229189;
assign addr[2673]= -993293415;
assign addr[2674]= -1027042599;
assign addr[2675]= -1060466036;
assign addr[2676]= -1093553126;
assign addr[2677]= -1126293375;
assign addr[2678]= -1158676398;
assign addr[2679]= -1190691925;
assign addr[2680]= -1222329801;
assign addr[2681]= -1253579991;
assign addr[2682]= -1284432584;
assign addr[2683]= -1314877795;
assign addr[2684]= -1344905966;
assign addr[2685]= -1374507575;
assign addr[2686]= -1403673233;
assign addr[2687]= -1432393688;
assign addr[2688]= -1460659832;
assign addr[2689]= -1488462700;
assign addr[2690]= -1515793473;
assign addr[2691]= -1542643483;
assign addr[2692]= -1569004214;
assign addr[2693]= -1594867305;
assign addr[2694]= -1620224553;
assign addr[2695]= -1645067915;
assign addr[2696]= -1669389513;
assign addr[2697]= -1693181631;
assign addr[2698]= -1716436725;
assign addr[2699]= -1739147417;
assign addr[2700]= -1761306505;
assign addr[2701]= -1782906961;
assign addr[2702]= -1803941934;
assign addr[2703]= -1824404752;
assign addr[2704]= -1844288924;
assign addr[2705]= -1863588145;
assign addr[2706]= -1882296293;
assign addr[2707]= -1900407434;
assign addr[2708]= -1917915825;
assign addr[2709]= -1934815911;
assign addr[2710]= -1951102334;
assign addr[2711]= -1966769926;
assign addr[2712]= -1981813720;
assign addr[2713]= -1996228943;
assign addr[2714]= -2010011024;
assign addr[2715]= -2023155591;
assign addr[2716]= -2035658475;
assign addr[2717]= -2047515711;
assign addr[2718]= -2058723538;
assign addr[2719]= -2069278401;
assign addr[2720]= -2079176953;
assign addr[2721]= -2088416053;
assign addr[2722]= -2096992772;
assign addr[2723]= -2104904390;
assign addr[2724]= -2112148396;
assign addr[2725]= -2118722494;
assign addr[2726]= -2124624598;
assign addr[2727]= -2129852837;
assign addr[2728]= -2134405552;
assign addr[2729]= -2138281298;
assign addr[2730]= -2141478848;
assign addr[2731]= -2143997187;
assign addr[2732]= -2145835515;
assign addr[2733]= -2146993250;
assign addr[2734]= -2147470025;
assign addr[2735]= -2147265689;
assign addr[2736]= -2146380306;
assign addr[2737]= -2144814157;
assign addr[2738]= -2142567738;
assign addr[2739]= -2139641764;
assign addr[2740]= -2136037160;
assign addr[2741]= -2131755071;
assign addr[2742]= -2126796855;
assign addr[2743]= -2121164085;
assign addr[2744]= -2114858546;
assign addr[2745]= -2107882239;
assign addr[2746]= -2100237377;
assign addr[2747]= -2091926384;
assign addr[2748]= -2082951896;
assign addr[2749]= -2073316760;
assign addr[2750]= -2063024031;
assign addr[2751]= -2052076975;
assign addr[2752]= -2040479063;
assign addr[2753]= -2028233973;
assign addr[2754]= -2015345591;
assign addr[2755]= -2001818002;
assign addr[2756]= -1987655498;
assign addr[2757]= -1972862571;
assign addr[2758]= -1957443913;
assign addr[2759]= -1941404413;
assign addr[2760]= -1924749160;
assign addr[2761]= -1907483436;
assign addr[2762]= -1889612716;
assign addr[2763]= -1871142669;
assign addr[2764]= -1852079154;
assign addr[2765]= -1832428215;
assign addr[2766]= -1812196087;
assign addr[2767]= -1791389186;
assign addr[2768]= -1770014111;
assign addr[2769]= -1748077642;
assign addr[2770]= -1725586737;
assign addr[2771]= -1702548529;
assign addr[2772]= -1678970324;
assign addr[2773]= -1654859602;
assign addr[2774]= -1630224009;
assign addr[2775]= -1605071359;
assign addr[2776]= -1579409630;
assign addr[2777]= -1553246960;
assign addr[2778]= -1526591649;
assign addr[2779]= -1499452149;
assign addr[2780]= -1471837070;
assign addr[2781]= -1443755168;
assign addr[2782]= -1415215352;
assign addr[2783]= -1386226674;
assign addr[2784]= -1356798326;
assign addr[2785]= -1326939644;
assign addr[2786]= -1296660098;
assign addr[2787]= -1265969291;
assign addr[2788]= -1234876957;
assign addr[2789]= -1203392958;
assign addr[2790]= -1171527280;
assign addr[2791]= -1139290029;
assign addr[2792]= -1106691431;
assign addr[2793]= -1073741824;
assign addr[2794]= -1040451659;
assign addr[2795]= -1006831495;
assign addr[2796]= -972891995;
assign addr[2797]= -938643924;
assign addr[2798]= -904098143;
assign addr[2799]= -869265610;
assign addr[2800]= -834157373;
assign addr[2801]= -798784567;
assign addr[2802]= -763158411;
assign addr[2803]= -727290205;
assign addr[2804]= -691191324;
assign addr[2805]= -654873219;
assign addr[2806]= -618347408;
assign addr[2807]= -581625477;
assign addr[2808]= -544719071;
assign addr[2809]= -507639898;
assign addr[2810]= -470399716;
assign addr[2811]= -433010339;
assign addr[2812]= -395483624;
assign addr[2813]= -357831473;
assign addr[2814]= -320065829;
assign addr[2815]= -282198671;
assign addr[2816]= -244242007;
assign addr[2817]= -206207878;
assign addr[2818]= -168108346;
assign addr[2819]= -129955495;
assign addr[2820]= -91761426;
assign addr[2821]= -53538253;
assign addr[2822]= -15298099;
assign addr[2823]= 22946906;
assign addr[2824]= 61184634;
assign addr[2825]= 99402956;
assign addr[2826]= 137589750;
assign addr[2827]= 175732905;
assign addr[2828]= 213820322;
assign addr[2829]= 251839923;
assign addr[2830]= 289779648;
assign addr[2831]= 327627463;
assign addr[2832]= 365371365;
assign addr[2833]= 402999383;
assign addr[2834]= 440499581;
assign addr[2835]= 477860067;
assign addr[2836]= 515068990;
assign addr[2837]= 552114549;
assign addr[2838]= 588984994;
assign addr[2839]= 625668632;
assign addr[2840]= 662153826;
assign addr[2841]= 698429006;
assign addr[2842]= 734482665;
assign addr[2843]= 770303369;
assign addr[2844]= 805879757;
assign addr[2845]= 841200544;
assign addr[2846]= 876254528;
assign addr[2847]= 911030591;
assign addr[2848]= 945517704;
assign addr[2849]= 979704927;
assign addr[2850]= 1013581418;
assign addr[2851]= 1047136432;
assign addr[2852]= 1080359326;
assign addr[2853]= 1113239564;
assign addr[2854]= 1145766716;
assign addr[2855]= 1177930466;
assign addr[2856]= 1209720613;
assign addr[2857]= 1241127074;
assign addr[2858]= 1272139887;
assign addr[2859]= 1302749217;
assign addr[2860]= 1332945355;
assign addr[2861]= 1362718723;
assign addr[2862]= 1392059879;
assign addr[2863]= 1420959516;
assign addr[2864]= 1449408469;
assign addr[2865]= 1477397714;
assign addr[2866]= 1504918373;
assign addr[2867]= 1531961719;
assign addr[2868]= 1558519173;
assign addr[2869]= 1584582314;
assign addr[2870]= 1610142873;
assign addr[2871]= 1635192744;
assign addr[2872]= 1659723983;
assign addr[2873]= 1683728808;
assign addr[2874]= 1707199606;
assign addr[2875]= 1730128933;
assign addr[2876]= 1752509516;
assign addr[2877]= 1774334257;
assign addr[2878]= 1795596234;
assign addr[2879]= 1816288703;
assign addr[2880]= 1836405100;
assign addr[2881]= 1855939047;
assign addr[2882]= 1874884346;
assign addr[2883]= 1893234990;
assign addr[2884]= 1910985158;
assign addr[2885]= 1928129220;
assign addr[2886]= 1944661739;
assign addr[2887]= 1960577471;
assign addr[2888]= 1975871368;
assign addr[2889]= 1990538579;
assign addr[2890]= 2004574453;
assign addr[2891]= 2017974537;
assign addr[2892]= 2030734582;
assign addr[2893]= 2042850540;
assign addr[2894]= 2054318569;
assign addr[2895]= 2065135031;
assign addr[2896]= 2075296495;
assign addr[2897]= 2084799740;
assign addr[2898]= 2093641749;
assign addr[2899]= 2101819720;
assign addr[2900]= 2109331059;
assign addr[2901]= 2116173382;
assign addr[2902]= 2122344521;
assign addr[2903]= 2127842516;
assign addr[2904]= 2132665626;
assign addr[2905]= 2136812319;
assign addr[2906]= 2140281282;
assign addr[2907]= 2143071413;
assign addr[2908]= 2145181827;
assign addr[2909]= 2146611856;
assign addr[2910]= 2147361045;
assign addr[2911]= 2147429158;
assign addr[2912]= 2146816171;
assign addr[2913]= 2145522281;
assign addr[2914]= 2143547897;
assign addr[2915]= 2140893646;
assign addr[2916]= 2137560369;
assign addr[2917]= 2133549123;
assign addr[2918]= 2128861181;
assign addr[2919]= 2123498030;
assign addr[2920]= 2117461370;
assign addr[2921]= 2110753117;
assign addr[2922]= 2103375398;
assign addr[2923]= 2095330553;
assign addr[2924]= 2086621133;
assign addr[2925]= 2077249901;
assign addr[2926]= 2067219829;
assign addr[2927]= 2056534099;
assign addr[2928]= 2045196100;
assign addr[2929]= 2033209426;
assign addr[2930]= 2020577882;
assign addr[2931]= 2007305472;
assign addr[2932]= 1993396407;
assign addr[2933]= 1978855097;
assign addr[2934]= 1963686155;
assign addr[2935]= 1947894393;
assign addr[2936]= 1931484818;
assign addr[2937]= 1914462636;
assign addr[2938]= 1896833245;
assign addr[2939]= 1878602237;
assign addr[2940]= 1859775393;
assign addr[2941]= 1840358687;
assign addr[2942]= 1820358275;
assign addr[2943]= 1799780501;
assign addr[2944]= 1778631892;
assign addr[2945]= 1756919156;
assign addr[2946]= 1734649179;
assign addr[2947]= 1711829025;
assign addr[2948]= 1688465931;
assign addr[2949]= 1664567307;
assign addr[2950]= 1640140734;
assign addr[2951]= 1615193959;
assign addr[2952]= 1589734894;
assign addr[2953]= 1563771613;
assign addr[2954]= 1537312353;
assign addr[2955]= 1510365504;
assign addr[2956]= 1482939614;
assign addr[2957]= 1455043381;
assign addr[2958]= 1426685652;
assign addr[2959]= 1397875423;
assign addr[2960]= 1368621831;
assign addr[2961]= 1338934154;
assign addr[2962]= 1308821808;
assign addr[2963]= 1278294345;
assign addr[2964]= 1247361445;
assign addr[2965]= 1216032921;
assign addr[2966]= 1184318708;
assign addr[2967]= 1152228866;
assign addr[2968]= 1119773573;
assign addr[2969]= 1086963121;
assign addr[2970]= 1053807919;
assign addr[2971]= 1020318481;
assign addr[2972]= 986505429;
assign addr[2973]= 952379488;
assign addr[2974]= 917951481;
assign addr[2975]= 883232329;
assign addr[2976]= 848233042;
assign addr[2977]= 812964722;
assign addr[2978]= 777438554;
assign addr[2979]= 741665807;
assign addr[2980]= 705657826;
assign addr[2981]= 669426032;
assign addr[2982]= 632981917;
assign addr[2983]= 596337040;
assign addr[2984]= 559503022;
assign addr[2985]= 522491548;
assign addr[2986]= 485314355;
assign addr[2987]= 447983235;
assign addr[2988]= 410510029;
assign addr[2989]= 372906622;
assign addr[2990]= 335184940;
assign addr[2991]= 297356948;
assign addr[2992]= 259434643;
assign addr[2993]= 221430054;
assign addr[2994]= 183355234;
assign addr[2995]= 145222259;
assign addr[2996]= 107043224;
assign addr[2997]= 68830239;
assign addr[2998]= 30595422;
assign addr[2999]= -7649098;
assign addr[3000]= -45891193;
assign addr[3001]= -84118732;
assign addr[3002]= -122319591;
assign addr[3003]= -160481654;
assign addr[3004]= -198592817;
assign addr[3005]= -236640993;
assign addr[3006]= -274614114;
assign addr[3007]= -312500135;
assign addr[3008]= -350287041;
assign addr[3009]= -387962847;
assign addr[3010]= -425515602;
assign addr[3011]= -462933398;
assign addr[3012]= -500204365;
assign addr[3013]= -537316682;
assign addr[3014]= -574258580;
assign addr[3015]= -611018340;
assign addr[3016]= -647584304;
assign addr[3017]= -683944874;
assign addr[3018]= -720088517;
assign addr[3019]= -756003771;
assign addr[3020]= -791679244;
assign addr[3021]= -827103620;
assign addr[3022]= -862265664;
assign addr[3023]= -897154224;
assign addr[3024]= -931758235;
assign addr[3025]= -966066720;
assign addr[3026]= -1000068799;
assign addr[3027]= -1033753687;
assign addr[3028]= -1067110699;
assign addr[3029]= -1100129257;
assign addr[3030]= -1132798888;
assign addr[3031]= -1165109230;
assign addr[3032]= -1197050035;
assign addr[3033]= -1228611172;
assign addr[3034]= -1259782632;
assign addr[3035]= -1290554528;
assign addr[3036]= -1320917099;
assign addr[3037]= -1350860716;
assign addr[3038]= -1380375881;
assign addr[3039]= -1409453233;
assign addr[3040]= -1438083551;
assign addr[3041]= -1466257752;
assign addr[3042]= -1493966902;
assign addr[3043]= -1521202211;
assign addr[3044]= -1547955041;
assign addr[3045]= -1574216908;
assign addr[3046]= -1599979481;
assign addr[3047]= -1625234591;
assign addr[3048]= -1649974225;
assign addr[3049]= -1674190539;
assign addr[3050]= -1697875851;
assign addr[3051]= -1721022648;
assign addr[3052]= -1743623590;
assign addr[3053]= -1765671509;
assign addr[3054]= -1787159411;
assign addr[3055]= -1808080480;
assign addr[3056]= -1828428082;
assign addr[3057]= -1848195763;
assign addr[3058]= -1867377253;
assign addr[3059]= -1885966468;
assign addr[3060]= -1903957513;
assign addr[3061]= -1921344681;
assign addr[3062]= -1938122457;
assign addr[3063]= -1954285520;
assign addr[3064]= -1969828744;
assign addr[3065]= -1984747199;
assign addr[3066]= -1999036154;
assign addr[3067]= -2012691075;
assign addr[3068]= -2025707632;
assign addr[3069]= -2038081698;
assign addr[3070]= -2049809346;
assign addr[3071]= -2060886858;
assign addr[3072]= -2071310720;
assign addr[3073]= -2081077626;
assign addr[3074]= -2090184478;
assign addr[3075]= -2098628387;
assign addr[3076]= -2106406677;
assign addr[3077]= -2113516878;
assign addr[3078]= -2119956737;
assign addr[3079]= -2125724211;
assign addr[3080]= -2130817471;
assign addr[3081]= -2135234901;
assign addr[3082]= -2138975100;
assign addr[3083]= -2142036881;
assign addr[3084]= -2144419275;
assign addr[3085]= -2146121524;
assign addr[3086]= -2147143090;
assign addr[3087]= -2147483648;
assign addr[3088]= -2147143090;
assign addr[3089]= -2146121524;
assign addr[3090]= -2144419275;
assign addr[3091]= -2142036881;
assign addr[3092]= -2138975100;
assign addr[3093]= -2135234901;
assign addr[3094]= -2130817471;
assign addr[3095]= -2125724211;
assign addr[3096]= -2119956737;
assign addr[3097]= -2113516878;
assign addr[3098]= -2106406677;
assign addr[3099]= -2098628387;
assign addr[3100]= -2090184478;
assign addr[3101]= -2081077626;
assign addr[3102]= -2071310720;
assign addr[3103]= -2060886858;
assign addr[3104]= -2049809346;
assign addr[3105]= -2038081698;
assign addr[3106]= -2025707632;
assign addr[3107]= -2012691075;
assign addr[3108]= -1999036154;
assign addr[3109]= -1984747199;
assign addr[3110]= -1969828744;
assign addr[3111]= -1954285520;
assign addr[3112]= -1938122457;
assign addr[3113]= -1921344681;
assign addr[3114]= -1903957513;
assign addr[3115]= -1885966468;
assign addr[3116]= -1867377253;
assign addr[3117]= -1848195763;
assign addr[3118]= -1828428082;
assign addr[3119]= -1808080480;
assign addr[3120]= -1787159411;
assign addr[3121]= -1765671509;
assign addr[3122]= -1743623590;
assign addr[3123]= -1721022648;
assign addr[3124]= -1697875851;
assign addr[3125]= -1674190539;
assign addr[3126]= -1649974225;
assign addr[3127]= -1625234591;
assign addr[3128]= -1599979481;
assign addr[3129]= -1574216908;
assign addr[3130]= -1547955041;
assign addr[3131]= -1521202211;
assign addr[3132]= -1493966902;
assign addr[3133]= -1466257752;
assign addr[3134]= -1438083551;
assign addr[3135]= -1409453233;
assign addr[3136]= -1380375881;
assign addr[3137]= -1350860716;
assign addr[3138]= -1320917099;
assign addr[3139]= -1290554528;
assign addr[3140]= -1259782632;
assign addr[3141]= -1228611172;
assign addr[3142]= -1197050035;
assign addr[3143]= -1165109230;
assign addr[3144]= -1132798888;
assign addr[3145]= -1100129257;
assign addr[3146]= -1067110699;
assign addr[3147]= -1033753687;
assign addr[3148]= -1000068799;
assign addr[3149]= -966066720;
assign addr[3150]= -931758235;
assign addr[3151]= -897154224;
assign addr[3152]= -862265664;
assign addr[3153]= -827103620;
assign addr[3154]= -791679244;
assign addr[3155]= -756003771;
assign addr[3156]= -720088517;
assign addr[3157]= -683944874;
assign addr[3158]= -647584304;
assign addr[3159]= -611018340;
assign addr[3160]= -574258580;
assign addr[3161]= -537316682;
assign addr[3162]= -500204365;
assign addr[3163]= -462933398;
assign addr[3164]= -425515602;
assign addr[3165]= -387962847;
assign addr[3166]= -350287041;
assign addr[3167]= -312500135;
assign addr[3168]= -274614114;
assign addr[3169]= -236640993;
assign addr[3170]= -198592817;
assign addr[3171]= -160481654;
assign addr[3172]= -122319591;
assign addr[3173]= -84118732;
assign addr[3174]= -45891193;
assign addr[3175]= -7649098;
assign addr[3176]= 30595422;
assign addr[3177]= 68830239;
assign addr[3178]= 107043224;
assign addr[3179]= 145222259;
assign addr[3180]= 183355234;
assign addr[3181]= 221430054;
assign addr[3182]= 259434643;
assign addr[3183]= 297356948;
assign addr[3184]= 335184940;
assign addr[3185]= 372906622;
assign addr[3186]= 410510029;
assign addr[3187]= 447983235;
assign addr[3188]= 485314355;
assign addr[3189]= 522491548;
assign addr[3190]= 559503022;
assign addr[3191]= 596337040;
assign addr[3192]= 632981917;
assign addr[3193]= 669426032;
assign addr[3194]= 705657826;
assign addr[3195]= 741665807;
assign addr[3196]= 777438554;
assign addr[3197]= 812964722;
assign addr[3198]= 848233042;
assign addr[3199]= 883232329;
assign addr[3200]= 917951481;
assign addr[3201]= 952379488;
assign addr[3202]= 986505429;
assign addr[3203]= 1020318481;
assign addr[3204]= 1053807919;
assign addr[3205]= 1086963121;
assign addr[3206]= 1119773573;
assign addr[3207]= 1152228866;
assign addr[3208]= 1184318708;
assign addr[3209]= 1216032921;
assign addr[3210]= 1247361445;
assign addr[3211]= 1278294345;
assign addr[3212]= 1308821808;
assign addr[3213]= 1338934154;
assign addr[3214]= 1368621831;
assign addr[3215]= 1397875423;
assign addr[3216]= 1426685652;
assign addr[3217]= 1455043381;
assign addr[3218]= 1482939614;
assign addr[3219]= 1510365504;
assign addr[3220]= 1537312353;
assign addr[3221]= 1563771613;
assign addr[3222]= 1589734894;
assign addr[3223]= 1615193959;
assign addr[3224]= 1640140734;
assign addr[3225]= 1664567307;
assign addr[3226]= 1688465931;
assign addr[3227]= 1711829025;
assign addr[3228]= 1734649179;
assign addr[3229]= 1756919156;
assign addr[3230]= 1778631892;
assign addr[3231]= 1799780501;
assign addr[3232]= 1820358275;
assign addr[3233]= 1840358687;
assign addr[3234]= 1859775393;
assign addr[3235]= 1878602237;
assign addr[3236]= 1896833245;
assign addr[3237]= 1914462636;
assign addr[3238]= 1931484818;
assign addr[3239]= 1947894393;
assign addr[3240]= 1963686155;
assign addr[3241]= 1978855097;
assign addr[3242]= 1993396407;
assign addr[3243]= 2007305472;
assign addr[3244]= 2020577882;
assign addr[3245]= 2033209426;
assign addr[3246]= 2045196100;
assign addr[3247]= 2056534099;
assign addr[3248]= 2067219829;
assign addr[3249]= 2077249901;
assign addr[3250]= 2086621133;
assign addr[3251]= 2095330553;
assign addr[3252]= 2103375398;
assign addr[3253]= 2110753117;
assign addr[3254]= 2117461370;
assign addr[3255]= 2123498030;
assign addr[3256]= 2128861181;
assign addr[3257]= 2133549123;
assign addr[3258]= 2137560369;
assign addr[3259]= 2140893646;
assign addr[3260]= 2143547897;
assign addr[3261]= 2145522281;
assign addr[3262]= 2146816171;
assign addr[3263]= 2147429158;
assign addr[3264]= 2147361045;
assign addr[3265]= 2146611856;
assign addr[3266]= 2145181827;
assign addr[3267]= 2143071413;
assign addr[3268]= 2140281282;
assign addr[3269]= 2136812319;
assign addr[3270]= 2132665626;
assign addr[3271]= 2127842516;
assign addr[3272]= 2122344521;
assign addr[3273]= 2116173382;
assign addr[3274]= 2109331059;
assign addr[3275]= 2101819720;
assign addr[3276]= 2093641749;
assign addr[3277]= 2084799740;
assign addr[3278]= 2075296495;
assign addr[3279]= 2065135031;
assign addr[3280]= 2054318569;
assign addr[3281]= 2042850540;
assign addr[3282]= 2030734582;
assign addr[3283]= 2017974537;
assign addr[3284]= 2004574453;
assign addr[3285]= 1990538579;
assign addr[3286]= 1975871368;
assign addr[3287]= 1960577471;
assign addr[3288]= 1944661739;
assign addr[3289]= 1928129220;
assign addr[3290]= 1910985158;
assign addr[3291]= 1893234990;
assign addr[3292]= 1874884346;
assign addr[3293]= 1855939047;
assign addr[3294]= 1836405100;
assign addr[3295]= 1816288703;
assign addr[3296]= 1795596234;
assign addr[3297]= 1774334257;
assign addr[3298]= 1752509516;
assign addr[3299]= 1730128933;
assign addr[3300]= 1707199606;
assign addr[3301]= 1683728808;
assign addr[3302]= 1659723983;
assign addr[3303]= 1635192744;
assign addr[3304]= 1610142873;
assign addr[3305]= 1584582314;
assign addr[3306]= 1558519173;
assign addr[3307]= 1531961719;
assign addr[3308]= 1504918373;
assign addr[3309]= 1477397714;
assign addr[3310]= 1449408469;
assign addr[3311]= 1420959516;
assign addr[3312]= 1392059879;
assign addr[3313]= 1362718723;
assign addr[3314]= 1332945355;
assign addr[3315]= 1302749217;
assign addr[3316]= 1272139887;
assign addr[3317]= 1241127074;
assign addr[3318]= 1209720613;
assign addr[3319]= 1177930466;
assign addr[3320]= 1145766716;
assign addr[3321]= 1113239564;
assign addr[3322]= 1080359326;
assign addr[3323]= 1047136432;
assign addr[3324]= 1013581418;
assign addr[3325]= 979704927;
assign addr[3326]= 945517704;
assign addr[3327]= 911030591;
assign addr[3328]= 876254528;
assign addr[3329]= 841200544;
assign addr[3330]= 805879757;
assign addr[3331]= 770303369;
assign addr[3332]= 734482665;
assign addr[3333]= 698429006;
assign addr[3334]= 662153826;
assign addr[3335]= 625668632;
assign addr[3336]= 588984994;
assign addr[3337]= 552114549;
assign addr[3338]= 515068990;
assign addr[3339]= 477860067;
assign addr[3340]= 440499581;
assign addr[3341]= 402999383;
assign addr[3342]= 365371365;
assign addr[3343]= 327627463;
assign addr[3344]= 289779648;
assign addr[3345]= 251839923;
assign addr[3346]= 213820322;
assign addr[3347]= 175732905;
assign addr[3348]= 137589750;
assign addr[3349]= 99402956;
assign addr[3350]= 61184634;
assign addr[3351]= 22946906;
assign addr[3352]= -15298099;
assign addr[3353]= -53538253;
assign addr[3354]= -91761426;
assign addr[3355]= -129955495;
assign addr[3356]= -168108346;
assign addr[3357]= -206207878;
assign addr[3358]= -244242007;
assign addr[3359]= -282198671;
assign addr[3360]= -320065829;
assign addr[3361]= -357831473;
assign addr[3362]= -395483624;
assign addr[3363]= -433010339;
assign addr[3364]= -470399716;
assign addr[3365]= -507639898;
assign addr[3366]= -544719071;
assign addr[3367]= -581625477;
assign addr[3368]= -618347408;
assign addr[3369]= -654873219;
assign addr[3370]= -691191324;
assign addr[3371]= -727290205;
assign addr[3372]= -763158411;
assign addr[3373]= -798784567;
assign addr[3374]= -834157373;
assign addr[3375]= -869265610;
assign addr[3376]= -904098143;
assign addr[3377]= -938643924;
assign addr[3378]= -972891995;
assign addr[3379]= -1006831495;
assign addr[3380]= -1040451659;
assign addr[3381]= -1073741824;
assign addr[3382]= -1106691431;
assign addr[3383]= -1139290029;
assign addr[3384]= -1171527280;
assign addr[3385]= -1203392958;
assign addr[3386]= -1234876957;
assign addr[3387]= -1265969291;
assign addr[3388]= -1296660098;
assign addr[3389]= -1326939644;
assign addr[3390]= -1356798326;
assign addr[3391]= -1386226674;
assign addr[3392]= -1415215352;
assign addr[3393]= -1443755168;
assign addr[3394]= -1471837070;
assign addr[3395]= -1499452149;
assign addr[3396]= -1526591649;
assign addr[3397]= -1553246960;
assign addr[3398]= -1579409630;
assign addr[3399]= -1605071359;
assign addr[3400]= -1630224009;
assign addr[3401]= -1654859602;
assign addr[3402]= -1678970324;
assign addr[3403]= -1702548529;
assign addr[3404]= -1725586737;
assign addr[3405]= -1748077642;
assign addr[3406]= -1770014111;
assign addr[3407]= -1791389186;
assign addr[3408]= -1812196087;
assign addr[3409]= -1832428215;
assign addr[3410]= -1852079154;
assign addr[3411]= -1871142669;
assign addr[3412]= -1889612716;
assign addr[3413]= -1907483436;
assign addr[3414]= -1924749160;
assign addr[3415]= -1941404413;
assign addr[3416]= -1957443913;
assign addr[3417]= -1972862571;
assign addr[3418]= -1987655498;
assign addr[3419]= -2001818002;
assign addr[3420]= -2015345591;
assign addr[3421]= -2028233973;
assign addr[3422]= -2040479063;
assign addr[3423]= -2052076975;
assign addr[3424]= -2063024031;
assign addr[3425]= -2073316760;
assign addr[3426]= -2082951896;
assign addr[3427]= -2091926384;
assign addr[3428]= -2100237377;
assign addr[3429]= -2107882239;
assign addr[3430]= -2114858546;
assign addr[3431]= -2121164085;
assign addr[3432]= -2126796855;
assign addr[3433]= -2131755071;
assign addr[3434]= -2136037160;
assign addr[3435]= -2139641764;
assign addr[3436]= -2142567738;
assign addr[3437]= -2144814157;
assign addr[3438]= -2146380306;
assign addr[3439]= -2147265689;
assign addr[3440]= -2147470025;
assign addr[3441]= -2146993250;
assign addr[3442]= -2145835515;
assign addr[3443]= -2143997187;
assign addr[3444]= -2141478848;
assign addr[3445]= -2138281298;
assign addr[3446]= -2134405552;
assign addr[3447]= -2129852837;
assign addr[3448]= -2124624598;
assign addr[3449]= -2118722494;
assign addr[3450]= -2112148396;
assign addr[3451]= -2104904390;
assign addr[3452]= -2096992772;
assign addr[3453]= -2088416053;
assign addr[3454]= -2079176953;
assign addr[3455]= -2069278401;
assign addr[3456]= -2058723538;
assign addr[3457]= -2047515711;
assign addr[3458]= -2035658475;
assign addr[3459]= -2023155591;
assign addr[3460]= -2010011024;
assign addr[3461]= -1996228943;
assign addr[3462]= -1981813720;
assign addr[3463]= -1966769926;
assign addr[3464]= -1951102334;
assign addr[3465]= -1934815911;
assign addr[3466]= -1917915825;
assign addr[3467]= -1900407434;
assign addr[3468]= -1882296293;
assign addr[3469]= -1863588145;
assign addr[3470]= -1844288924;
assign addr[3471]= -1824404752;
assign addr[3472]= -1803941934;
assign addr[3473]= -1782906961;
assign addr[3474]= -1761306505;
assign addr[3475]= -1739147417;
assign addr[3476]= -1716436725;
assign addr[3477]= -1693181631;
assign addr[3478]= -1669389513;
assign addr[3479]= -1645067915;
assign addr[3480]= -1620224553;
assign addr[3481]= -1594867305;
assign addr[3482]= -1569004214;
assign addr[3483]= -1542643483;
assign addr[3484]= -1515793473;
assign addr[3485]= -1488462700;
assign addr[3486]= -1460659832;
assign addr[3487]= -1432393688;
assign addr[3488]= -1403673233;
assign addr[3489]= -1374507575;
assign addr[3490]= -1344905966;
assign addr[3491]= -1314877795;
assign addr[3492]= -1284432584;
assign addr[3493]= -1253579991;
assign addr[3494]= -1222329801;
assign addr[3495]= -1190691925;
assign addr[3496]= -1158676398;
assign addr[3497]= -1126293375;
assign addr[3498]= -1093553126;
assign addr[3499]= -1060466036;
assign addr[3500]= -1027042599;
assign addr[3501]= -993293415;
assign addr[3502]= -959229189;
assign addr[3503]= -924860725;
assign addr[3504]= -890198924;
assign addr[3505]= -855254778;
assign addr[3506]= -820039373;
assign addr[3507]= -784563876;
assign addr[3508]= -748839539;
assign addr[3509]= -712877694;
assign addr[3510]= -676689746;
assign addr[3511]= -640287172;
assign addr[3512]= -603681519;
assign addr[3513]= -566884397;
assign addr[3514]= -529907477;
assign addr[3515]= -492762486;
assign addr[3516]= -455461206;
assign addr[3517]= -418015468;
assign addr[3518]= -380437148;
assign addr[3519]= -342738165;
assign addr[3520]= -304930476;
assign addr[3521]= -267026072;
assign addr[3522]= -229036977;
assign addr[3523]= -190975237;
assign addr[3524]= -152852926;
assign addr[3525]= -114682135;
assign addr[3526]= -76474970;
assign addr[3527]= -38243550;
assign addr[3528]= 0;
assign addr[3529]= 38243550;
assign addr[3530]= 76474970;
assign addr[3531]= 114682135;
assign addr[3532]= 152852926;
assign addr[3533]= 190975237;
assign addr[3534]= 229036977;
assign addr[3535]= 267026072;
assign addr[3536]= 304930476;
assign addr[3537]= 342738165;
assign addr[3538]= 380437148;
assign addr[3539]= 418015468;
assign addr[3540]= 455461206;
assign addr[3541]= 492762486;
assign addr[3542]= 529907477;
assign addr[3543]= 566884397;
assign addr[3544]= 603681519;
assign addr[3545]= 640287172;
assign addr[3546]= 676689746;
assign addr[3547]= 712877694;
assign addr[3548]= 748839539;
assign addr[3549]= 784563876;
assign addr[3550]= 820039373;
assign addr[3551]= 855254778;
assign addr[3552]= 890198924;
assign addr[3553]= 924860725;
assign addr[3554]= 959229189;
assign addr[3555]= 993293415;
assign addr[3556]= 1027042599;
assign addr[3557]= 1060466036;
assign addr[3558]= 1093553126;
assign addr[3559]= 1126293375;
assign addr[3560]= 1158676398;
assign addr[3561]= 1190691925;
assign addr[3562]= 1222329801;
assign addr[3563]= 1253579991;
assign addr[3564]= 1284432584;
assign addr[3565]= 1314877795;
assign addr[3566]= 1344905966;
assign addr[3567]= 1374507575;
assign addr[3568]= 1403673233;
assign addr[3569]= 1432393688;
assign addr[3570]= 1460659832;
assign addr[3571]= 1488462700;
assign addr[3572]= 1515793473;
assign addr[3573]= 1542643483;
assign addr[3574]= 1569004214;
assign addr[3575]= 1594867305;
assign addr[3576]= 1620224553;
assign addr[3577]= 1645067915;
assign addr[3578]= 1669389513;
assign addr[3579]= 1693181631;
assign addr[3580]= 1716436725;
assign addr[3581]= 1739147417;
assign addr[3582]= 1761306505;
assign addr[3583]= 1782906961;
assign addr[3584]= 1803941934;
assign addr[3585]= 1824404752;
assign addr[3586]= 1844288924;
assign addr[3587]= 1863588145;
assign addr[3588]= 1882296293;
assign addr[3589]= 1900407434;
assign addr[3590]= 1917915825;
assign addr[3591]= 1934815911;
assign addr[3592]= 1951102334;
assign addr[3593]= 1966769926;
assign addr[3594]= 1981813720;
assign addr[3595]= 1996228943;
assign addr[3596]= 2010011024;
assign addr[3597]= 2023155591;
assign addr[3598]= 2035658475;
assign addr[3599]= 2047515711;
assign addr[3600]= 2058723538;
assign addr[3601]= 2069278401;
assign addr[3602]= 2079176953;
assign addr[3603]= 2088416053;
assign addr[3604]= 2096992772;
assign addr[3605]= 2104904390;
assign addr[3606]= 2112148396;
assign addr[3607]= 2118722494;
assign addr[3608]= 2124624598;
assign addr[3609]= 2129852837;
assign addr[3610]= 2134405552;
assign addr[3611]= 2138281298;
assign addr[3612]= 2141478848;
assign addr[3613]= 2143997187;
assign addr[3614]= 2145835515;
assign addr[3615]= 2146993250;
assign addr[3616]= 2147470025;
assign addr[3617]= 2147265689;
assign addr[3618]= 2146380306;
assign addr[3619]= 2144814157;
assign addr[3620]= 2142567738;
assign addr[3621]= 2139641764;
assign addr[3622]= 2136037160;
assign addr[3623]= 2131755071;
assign addr[3624]= 2126796855;
assign addr[3625]= 2121164085;
assign addr[3626]= 2114858546;
assign addr[3627]= 2107882239;
assign addr[3628]= 2100237377;
assign addr[3629]= 2091926384;
assign addr[3630]= 2082951896;
assign addr[3631]= 2073316760;
assign addr[3632]= 2063024031;
assign addr[3633]= 2052076975;
assign addr[3634]= 2040479063;
assign addr[3635]= 2028233973;
assign addr[3636]= 2015345591;
assign addr[3637]= 2001818002;
assign addr[3638]= 1987655498;
assign addr[3639]= 1972862571;
assign addr[3640]= 1957443913;
assign addr[3641]= 1941404413;
assign addr[3642]= 1924749160;
assign addr[3643]= 1907483436;
assign addr[3644]= 1889612716;
assign addr[3645]= 1871142669;
assign addr[3646]= 1852079154;
assign addr[3647]= 1832428215;
assign addr[3648]= 1812196087;
assign addr[3649]= 1791389186;
assign addr[3650]= 1770014111;
assign addr[3651]= 1748077642;
assign addr[3652]= 1725586737;
assign addr[3653]= 1702548529;
assign addr[3654]= 1678970324;
assign addr[3655]= 1654859602;
assign addr[3656]= 1630224009;
assign addr[3657]= 1605071359;
assign addr[3658]= 1579409630;
assign addr[3659]= 1553246960;
assign addr[3660]= 1526591649;
assign addr[3661]= 1499452149;
assign addr[3662]= 1471837070;
assign addr[3663]= 1443755168;
assign addr[3664]= 1415215352;
assign addr[3665]= 1386226674;
assign addr[3666]= 1356798326;
assign addr[3667]= 1326939644;
assign addr[3668]= 1296660098;
assign addr[3669]= 1265969291;
assign addr[3670]= 1234876957;
assign addr[3671]= 1203392958;
assign addr[3672]= 1171527280;
assign addr[3673]= 1139290029;
assign addr[3674]= 1106691431;
assign addr[3675]= 1073741824;
assign addr[3676]= 1040451659;
assign addr[3677]= 1006831495;
assign addr[3678]= 972891995;
assign addr[3679]= 938643924;
assign addr[3680]= 904098143;
assign addr[3681]= 869265610;
assign addr[3682]= 834157373;
assign addr[3683]= 798784567;
assign addr[3684]= 763158411;
assign addr[3685]= 727290205;
assign addr[3686]= 691191324;
assign addr[3687]= 654873219;
assign addr[3688]= 618347408;
assign addr[3689]= 581625477;
assign addr[3690]= 544719071;
assign addr[3691]= 507639898;
assign addr[3692]= 470399716;
assign addr[3693]= 433010339;
assign addr[3694]= 395483624;
assign addr[3695]= 357831473;
assign addr[3696]= 320065829;
assign addr[3697]= 282198671;
assign addr[3698]= 244242007;
assign addr[3699]= 206207878;
assign addr[3700]= 168108346;
assign addr[3701]= 129955495;
assign addr[3702]= 91761426;
assign addr[3703]= 53538253;
assign addr[3704]= 15298099;
assign addr[3705]= -22946906;
assign addr[3706]= -61184634;
assign addr[3707]= -99402956;
assign addr[3708]= -137589750;
assign addr[3709]= -175732905;
assign addr[3710]= -213820322;
assign addr[3711]= -251839923;
assign addr[3712]= -289779648;
assign addr[3713]= -327627463;
assign addr[3714]= -365371365;
assign addr[3715]= -402999383;
assign addr[3716]= -440499581;
assign addr[3717]= -477860067;
assign addr[3718]= -515068990;
assign addr[3719]= -552114549;
assign addr[3720]= -588984994;
assign addr[3721]= -625668632;
assign addr[3722]= -662153826;
assign addr[3723]= -698429006;
assign addr[3724]= -734482665;
assign addr[3725]= -770303369;
assign addr[3726]= -805879757;
assign addr[3727]= -841200544;
assign addr[3728]= -876254528;
assign addr[3729]= -911030591;
assign addr[3730]= -945517704;
assign addr[3731]= -979704927;
assign addr[3732]= -1013581418;
assign addr[3733]= -1047136432;
assign addr[3734]= -1080359326;
assign addr[3735]= -1113239564;
assign addr[3736]= -1145766716;
assign addr[3737]= -1177930466;
assign addr[3738]= -1209720613;
assign addr[3739]= -1241127074;
assign addr[3740]= -1272139887;
assign addr[3741]= -1302749217;
assign addr[3742]= -1332945355;
assign addr[3743]= -1362718723;
assign addr[3744]= -1392059879;
assign addr[3745]= -1420959516;
assign addr[3746]= -1449408469;
assign addr[3747]= -1477397714;
assign addr[3748]= -1504918373;
assign addr[3749]= -1531961719;
assign addr[3750]= -1558519173;
assign addr[3751]= -1584582314;
assign addr[3752]= -1610142873;
assign addr[3753]= -1635192744;
assign addr[3754]= -1659723983;
assign addr[3755]= -1683728808;
assign addr[3756]= -1707199606;
assign addr[3757]= -1730128933;
assign addr[3758]= -1752509516;
assign addr[3759]= -1774334257;
assign addr[3760]= -1795596234;
assign addr[3761]= -1816288703;
assign addr[3762]= -1836405100;
assign addr[3763]= -1855939047;
assign addr[3764]= -1874884346;
assign addr[3765]= -1893234990;
assign addr[3766]= -1910985158;
assign addr[3767]= -1928129220;
assign addr[3768]= -1944661739;
assign addr[3769]= -1960577471;
assign addr[3770]= -1975871368;
assign addr[3771]= -1990538579;
assign addr[3772]= -2004574453;
assign addr[3773]= -2017974537;
assign addr[3774]= -2030734582;
assign addr[3775]= -2042850540;
assign addr[3776]= -2054318569;
assign addr[3777]= -2065135031;
assign addr[3778]= -2075296495;
assign addr[3779]= -2084799740;
assign addr[3780]= -2093641749;
assign addr[3781]= -2101819720;
assign addr[3782]= -2109331059;
assign addr[3783]= -2116173382;
assign addr[3784]= -2122344521;
assign addr[3785]= -2127842516;
assign addr[3786]= -2132665626;
assign addr[3787]= -2136812319;
assign addr[3788]= -2140281282;
assign addr[3789]= -2143071413;
assign addr[3790]= -2145181827;
assign addr[3791]= -2146611856;
assign addr[3792]= -2147361045;
assign addr[3793]= -2147429158;
assign addr[3794]= -2146816171;
assign addr[3795]= -2145522281;
assign addr[3796]= -2143547897;
assign addr[3797]= -2140893646;
assign addr[3798]= -2137560369;
assign addr[3799]= -2133549123;
assign addr[3800]= -2128861181;
assign addr[3801]= -2123498030;
assign addr[3802]= -2117461370;
assign addr[3803]= -2110753117;
assign addr[3804]= -2103375398;
assign addr[3805]= -2095330553;
assign addr[3806]= -2086621133;
assign addr[3807]= -2077249901;
assign addr[3808]= -2067219829;
assign addr[3809]= -2056534099;
assign addr[3810]= -2045196100;
assign addr[3811]= -2033209426;
assign addr[3812]= -2020577882;
assign addr[3813]= -2007305472;
assign addr[3814]= -1993396407;
assign addr[3815]= -1978855097;
assign addr[3816]= -1963686155;
assign addr[3817]= -1947894393;
assign addr[3818]= -1931484818;
assign addr[3819]= -1914462636;
assign addr[3820]= -1896833245;
assign addr[3821]= -1878602237;
assign addr[3822]= -1859775393;
assign addr[3823]= -1840358687;
assign addr[3824]= -1820358275;
assign addr[3825]= -1799780501;
assign addr[3826]= -1778631892;
assign addr[3827]= -1756919156;
assign addr[3828]= -1734649179;
assign addr[3829]= -1711829025;
assign addr[3830]= -1688465931;
assign addr[3831]= -1664567307;
assign addr[3832]= -1640140734;
assign addr[3833]= -1615193959;
assign addr[3834]= -1589734894;
assign addr[3835]= -1563771613;
assign addr[3836]= -1537312353;
assign addr[3837]= -1510365504;
assign addr[3838]= -1482939614;
assign addr[3839]= -1455043381;
assign addr[3840]= -1426685652;
assign addr[3841]= -1397875423;
assign addr[3842]= -1368621831;
assign addr[3843]= -1338934154;
assign addr[3844]= -1308821808;
assign addr[3845]= -1278294345;
assign addr[3846]= -1247361445;
assign addr[3847]= -1216032921;
assign addr[3848]= -1184318708;
assign addr[3849]= -1152228866;
assign addr[3850]= -1119773573;
assign addr[3851]= -1086963121;
assign addr[3852]= -1053807919;
assign addr[3853]= -1020318481;
assign addr[3854]= -986505429;
assign addr[3855]= -952379488;
assign addr[3856]= -917951481;
assign addr[3857]= -883232329;
assign addr[3858]= -848233042;
assign addr[3859]= -812964722;
assign addr[3860]= -777438554;
assign addr[3861]= -741665807;
assign addr[3862]= -705657826;
assign addr[3863]= -669426032;
assign addr[3864]= -632981917;
assign addr[3865]= -596337040;
assign addr[3866]= -559503022;
assign addr[3867]= -522491548;
assign addr[3868]= -485314355;
assign addr[3869]= -447983235;
assign addr[3870]= -410510029;
assign addr[3871]= -372906622;
assign addr[3872]= -335184940;
assign addr[3873]= -297356948;
assign addr[3874]= -259434643;
assign addr[3875]= -221430054;
assign addr[3876]= -183355234;
assign addr[3877]= -145222259;
assign addr[3878]= -107043224;
assign addr[3879]= -68830239;
assign addr[3880]= -30595422;
assign addr[3881]= 7649098;
assign addr[3882]= 45891193;
assign addr[3883]= 84118732;
assign addr[3884]= 122319591;
assign addr[3885]= 160481654;
assign addr[3886]= 198592817;
assign addr[3887]= 236640993;
assign addr[3888]= 274614114;
assign addr[3889]= 312500135;
assign addr[3890]= 350287041;
assign addr[3891]= 387962847;
assign addr[3892]= 425515602;
assign addr[3893]= 462933398;
assign addr[3894]= 500204365;
assign addr[3895]= 537316682;
assign addr[3896]= 574258580;
assign addr[3897]= 611018340;
assign addr[3898]= 647584304;
assign addr[3899]= 683944874;
assign addr[3900]= 720088517;
assign addr[3901]= 756003771;
assign addr[3902]= 791679244;
assign addr[3903]= 827103620;
assign addr[3904]= 862265664;
assign addr[3905]= 897154224;
assign addr[3906]= 931758235;
assign addr[3907]= 966066720;
assign addr[3908]= 1000068799;
assign addr[3909]= 1033753687;
assign addr[3910]= 1067110699;
assign addr[3911]= 1100129257;
assign addr[3912]= 1132798888;
assign addr[3913]= 1165109230;
assign addr[3914]= 1197050035;
assign addr[3915]= 1228611172;
assign addr[3916]= 1259782632;
assign addr[3917]= 1290554528;
assign addr[3918]= 1320917099;
assign addr[3919]= 1350860716;
assign addr[3920]= 1380375881;
assign addr[3921]= 1409453233;
assign addr[3922]= 1438083551;
assign addr[3923]= 1466257752;
assign addr[3924]= 1493966902;
assign addr[3925]= 1521202211;
assign addr[3926]= 1547955041;
assign addr[3927]= 1574216908;
assign addr[3928]= 1599979481;
assign addr[3929]= 1625234591;
assign addr[3930]= 1649974225;
assign addr[3931]= 1674190539;
assign addr[3932]= 1697875851;
assign addr[3933]= 1721022648;
assign addr[3934]= 1743623590;
assign addr[3935]= 1765671509;
assign addr[3936]= 1787159411;
assign addr[3937]= 1808080480;
assign addr[3938]= 1828428082;
assign addr[3939]= 1848195763;
assign addr[3940]= 1867377253;
assign addr[3941]= 1885966468;
assign addr[3942]= 1903957513;
assign addr[3943]= 1921344681;
assign addr[3944]= 1938122457;
assign addr[3945]= 1954285520;
assign addr[3946]= 1969828744;
assign addr[3947]= 1984747199;
assign addr[3948]= 1999036154;
assign addr[3949]= 2012691075;
assign addr[3950]= 2025707632;
assign addr[3951]= 2038081698;
assign addr[3952]= 2049809346;
assign addr[3953]= 2060886858;
assign addr[3954]= 2071310720;
assign addr[3955]= 2081077626;
assign addr[3956]= 2090184478;
assign addr[3957]= 2098628387;
assign addr[3958]= 2106406677;
assign addr[3959]= 2113516878;
assign addr[3960]= 2119956737;
assign addr[3961]= 2125724211;
assign addr[3962]= 2130817471;
assign addr[3963]= 2135234901;
assign addr[3964]= 2138975100;
assign addr[3965]= 2142036881;
assign addr[3966]= 2144419275;
assign addr[3967]= 2146121524;
assign addr[3968]= 2147143090;
assign addr[3969]= 2147483648;
assign addr[3970]= 2147143090;
assign addr[3971]= 2146121524;
assign addr[3972]= 2144419275;
assign addr[3973]= 2142036881;
assign addr[3974]= 2138975100;
assign addr[3975]= 2135234901;
assign addr[3976]= 2130817471;
assign addr[3977]= 2125724211;
assign addr[3978]= 2119956737;
assign addr[3979]= 2113516878;
assign addr[3980]= 2106406677;
assign addr[3981]= 2098628387;
assign addr[3982]= 2090184478;
assign addr[3983]= 2081077626;
assign addr[3984]= 2071310720;
assign addr[3985]= 2060886858;
assign addr[3986]= 2049809346;
assign addr[3987]= 2038081698;
assign addr[3988]= 2025707632;
assign addr[3989]= 2012691075;
assign addr[3990]= 1999036154;
assign addr[3991]= 1984747199;
assign addr[3992]= 1969828744;
assign addr[3993]= 1954285520;
assign addr[3994]= 1938122457;
assign addr[3995]= 1921344681;
assign addr[3996]= 1903957513;
assign addr[3997]= 1885966468;
assign addr[3998]= 1867377253;
assign addr[3999]= 1848195763;
assign addr[4000]= 1828428082;
assign addr[4001]= 1808080480;
assign addr[4002]= 1787159411;
assign addr[4003]= 1765671509;
assign addr[4004]= 1743623590;
assign addr[4005]= 1721022648;
assign addr[4006]= 1697875851;
assign addr[4007]= 1674190539;
assign addr[4008]= 1649974225;
assign addr[4009]= 1625234591;
assign addr[4010]= 1599979481;
assign addr[4011]= 1574216908;
assign addr[4012]= 1547955041;
assign addr[4013]= 1521202211;
assign addr[4014]= 1493966902;
assign addr[4015]= 1466257752;
assign addr[4016]= 1438083551;
assign addr[4017]= 1409453233;
assign addr[4018]= 1380375881;
assign addr[4019]= 1350860716;
assign addr[4020]= 1320917099;
assign addr[4021]= 1290554528;
assign addr[4022]= 1259782632;
assign addr[4023]= 1228611172;
assign addr[4024]= 1197050035;
assign addr[4025]= 1165109230;
assign addr[4026]= 1132798888;
assign addr[4027]= 1100129257;
assign addr[4028]= 1067110699;
assign addr[4029]= 1033753687;
assign addr[4030]= 1000068799;
assign addr[4031]= 966066720;
assign addr[4032]= 931758235;
assign addr[4033]= 897154224;
assign addr[4034]= 862265664;
assign addr[4035]= 827103620;
assign addr[4036]= 791679244;
assign addr[4037]= 756003771;
assign addr[4038]= 720088517;
assign addr[4039]= 683944874;
assign addr[4040]= 647584304;
assign addr[4041]= 611018340;
assign addr[4042]= 574258580;
assign addr[4043]= 537316682;
assign addr[4044]= 500204365;
assign addr[4045]= 462933398;
assign addr[4046]= 425515602;
assign addr[4047]= 387962847;
assign addr[4048]= 350287041;
assign addr[4049]= 312500135;
assign addr[4050]= 274614114;
assign addr[4051]= 236640993;
assign addr[4052]= 198592817;
assign addr[4053]= 160481654;
assign addr[4054]= 122319591;
assign addr[4055]= 84118732;
assign addr[4056]= 45891193;
assign addr[4057]= 7649098;
assign addr[4058]= -30595422;
assign addr[4059]= -68830239;
assign addr[4060]= -107043224;
assign addr[4061]= -145222259;
assign addr[4062]= -183355234;
assign addr[4063]= -221430054;
assign addr[4064]= -259434643;
assign addr[4065]= -297356948;
assign addr[4066]= -335184940;
assign addr[4067]= -372906622;
assign addr[4068]= -410510029;
assign addr[4069]= -447983235;
assign addr[4070]= -485314355;
assign addr[4071]= -522491548;
assign addr[4072]= -559503022;
assign addr[4073]= -596337040;
assign addr[4074]= -632981917;
assign addr[4075]= -669426032;
assign addr[4076]= -705657826;
assign addr[4077]= -741665807;
assign addr[4078]= -777438554;
assign addr[4079]= -812964722;
assign addr[4080]= -848233042;
assign addr[4081]= -883232329;
assign addr[4082]= -917951481;
assign addr[4083]= -952379488;
assign addr[4084]= -986505429;
assign addr[4085]= -1020318481;
assign addr[4086]= -1053807919;
assign addr[4087]= -1086963121;
assign addr[4088]= -1119773573;
assign addr[4089]= -1152228866;
assign addr[4090]= -1184318708;
assign addr[4091]= -1216032921;
assign addr[4092]= -1247361445;
assign addr[4093]= -1278294345;
assign addr[4094]= -1308821808;
assign addr[4095]= -1338934154;
assign addr[4096]= -1368621831;
assign addr[4097]= -1397875423;
assign addr[4098]= -1426685652;
assign addr[4099]= -1455043381;
assign addr[4100]= -1482939614;
assign addr[4101]= -1510365504;
assign addr[4102]= -1537312353;
assign addr[4103]= -1563771613;
assign addr[4104]= -1589734894;
assign addr[4105]= -1615193959;
assign addr[4106]= -1640140734;
assign addr[4107]= -1664567307;
assign addr[4108]= -1688465931;
assign addr[4109]= -1711829025;
assign addr[4110]= -1734649179;
assign addr[4111]= -1756919156;
assign addr[4112]= -1778631892;
assign addr[4113]= -1799780501;
assign addr[4114]= -1820358275;
assign addr[4115]= -1840358687;
assign addr[4116]= -1859775393;
assign addr[4117]= -1878602237;
assign addr[4118]= -1896833245;
assign addr[4119]= -1914462636;
assign addr[4120]= -1931484818;
assign addr[4121]= -1947894393;
assign addr[4122]= -1963686155;
assign addr[4123]= -1978855097;
assign addr[4124]= -1993396407;
assign addr[4125]= -2007305472;
assign addr[4126]= -2020577882;
assign addr[4127]= -2033209426;
assign addr[4128]= -2045196100;
assign addr[4129]= -2056534099;
assign addr[4130]= -2067219829;
assign addr[4131]= -2077249901;
assign addr[4132]= -2086621133;
assign addr[4133]= -2095330553;
assign addr[4134]= -2103375398;
assign addr[4135]= -2110753117;
assign addr[4136]= -2117461370;
assign addr[4137]= -2123498030;
assign addr[4138]= -2128861181;
assign addr[4139]= -2133549123;
assign addr[4140]= -2137560369;
assign addr[4141]= -2140893646;
assign addr[4142]= -2143547897;
assign addr[4143]= -2145522281;
assign addr[4144]= -2146816171;
assign addr[4145]= -2147429158;
assign addr[4146]= -2147361045;
assign addr[4147]= -2146611856;
assign addr[4148]= -2145181827;
assign addr[4149]= -2143071413;
assign addr[4150]= -2140281282;
assign addr[4151]= -2136812319;
assign addr[4152]= -2132665626;
assign addr[4153]= -2127842516;
assign addr[4154]= -2122344521;
assign addr[4155]= -2116173382;
assign addr[4156]= -2109331059;
assign addr[4157]= -2101819720;
assign addr[4158]= -2093641749;
assign addr[4159]= -2084799740;
assign addr[4160]= -2075296495;
assign addr[4161]= -2065135031;
assign addr[4162]= -2054318569;
assign addr[4163]= -2042850540;
assign addr[4164]= -2030734582;
assign addr[4165]= -2017974537;
assign addr[4166]= -2004574453;
assign addr[4167]= -1990538579;
assign addr[4168]= -1975871368;
assign addr[4169]= -1960577471;
assign addr[4170]= -1944661739;
assign addr[4171]= -1928129220;
assign addr[4172]= -1910985158;
assign addr[4173]= -1893234990;
assign addr[4174]= -1874884346;
assign addr[4175]= -1855939047;
assign addr[4176]= -1836405100;
assign addr[4177]= -1816288703;
assign addr[4178]= -1795596234;
assign addr[4179]= -1774334257;
assign addr[4180]= -1752509516;
assign addr[4181]= -1730128933;
assign addr[4182]= -1707199606;
assign addr[4183]= -1683728808;
assign addr[4184]= -1659723983;
assign addr[4185]= -1635192744;
assign addr[4186]= -1610142873;
assign addr[4187]= -1584582314;
assign addr[4188]= -1558519173;
assign addr[4189]= -1531961719;
assign addr[4190]= -1504918373;
assign addr[4191]= -1477397714;
assign addr[4192]= -1449408469;
assign addr[4193]= -1420959516;
assign addr[4194]= -1392059879;
assign addr[4195]= -1362718723;
assign addr[4196]= -1332945355;
assign addr[4197]= -1302749217;
assign addr[4198]= -1272139887;
assign addr[4199]= -1241127074;
assign addr[4200]= -1209720613;
assign addr[4201]= -1177930466;
assign addr[4202]= -1145766716;
assign addr[4203]= -1113239564;
assign addr[4204]= -1080359326;
assign addr[4205]= -1047136432;
assign addr[4206]= -1013581418;
assign addr[4207]= -979704927;
assign addr[4208]= -945517704;
assign addr[4209]= -911030591;
assign addr[4210]= -876254528;
assign addr[4211]= -841200544;
assign addr[4212]= -805879757;
assign addr[4213]= -770303369;
assign addr[4214]= -734482665;
assign addr[4215]= -698429006;
assign addr[4216]= -662153826;
assign addr[4217]= -625668632;
assign addr[4218]= -588984994;
assign addr[4219]= -552114549;
assign addr[4220]= -515068990;
assign addr[4221]= -477860067;
assign addr[4222]= -440499581;
assign addr[4223]= -402999383;
assign addr[4224]= -365371365;
assign addr[4225]= -327627463;
assign addr[4226]= -289779648;
assign addr[4227]= -251839923;
assign addr[4228]= -213820322;
assign addr[4229]= -175732905;
assign addr[4230]= -137589750;
assign addr[4231]= -99402956;
assign addr[4232]= -61184634;
assign addr[4233]= -22946906;
assign addr[4234]= 15298099;
assign addr[4235]= 53538253;
assign addr[4236]= 91761426;
assign addr[4237]= 129955495;
assign addr[4238]= 168108346;
assign addr[4239]= 206207878;
assign addr[4240]= 244242007;
assign addr[4241]= 282198671;
assign addr[4242]= 320065829;
assign addr[4243]= 357831473;
assign addr[4244]= 395483624;
assign addr[4245]= 433010339;
assign addr[4246]= 470399716;
assign addr[4247]= 507639898;
assign addr[4248]= 544719071;
assign addr[4249]= 581625477;
assign addr[4250]= 618347408;
assign addr[4251]= 654873219;
assign addr[4252]= 691191324;
assign addr[4253]= 727290205;
assign addr[4254]= 763158411;
assign addr[4255]= 798784567;
assign addr[4256]= 834157373;
assign addr[4257]= 869265610;
assign addr[4258]= 904098143;
assign addr[4259]= 938643924;
assign addr[4260]= 972891995;
assign addr[4261]= 1006831495;
assign addr[4262]= 1040451659;
assign addr[4263]= 1073741824;
assign addr[4264]= 1106691431;
assign addr[4265]= 1139290029;
assign addr[4266]= 1171527280;
assign addr[4267]= 1203392958;
assign addr[4268]= 1234876957;
assign addr[4269]= 1265969291;
assign addr[4270]= 1296660098;
assign addr[4271]= 1326939644;
assign addr[4272]= 1356798326;
assign addr[4273]= 1386226674;
assign addr[4274]= 1415215352;
assign addr[4275]= 1443755168;
assign addr[4276]= 1471837070;
assign addr[4277]= 1499452149;
assign addr[4278]= 1526591649;
assign addr[4279]= 1553246960;
assign addr[4280]= 1579409630;
assign addr[4281]= 1605071359;
assign addr[4282]= 1630224009;
assign addr[4283]= 1654859602;
assign addr[4284]= 1678970324;
assign addr[4285]= 1702548529;
assign addr[4286]= 1725586737;
assign addr[4287]= 1748077642;
assign addr[4288]= 1770014111;
assign addr[4289]= 1791389186;
assign addr[4290]= 1812196087;
assign addr[4291]= 1832428215;
assign addr[4292]= 1852079154;
assign addr[4293]= 1871142669;
assign addr[4294]= 1889612716;
assign addr[4295]= 1907483436;
assign addr[4296]= 1924749160;
assign addr[4297]= 1941404413;
assign addr[4298]= 1957443913;
assign addr[4299]= 1972862571;
assign addr[4300]= 1987655498;
assign addr[4301]= 2001818002;
assign addr[4302]= 2015345591;
assign addr[4303]= 2028233973;
assign addr[4304]= 2040479063;
assign addr[4305]= 2052076975;
assign addr[4306]= 2063024031;
assign addr[4307]= 2073316760;
assign addr[4308]= 2082951896;
assign addr[4309]= 2091926384;
assign addr[4310]= 2100237377;
assign addr[4311]= 2107882239;
assign addr[4312]= 2114858546;
assign addr[4313]= 2121164085;
assign addr[4314]= 2126796855;
assign addr[4315]= 2131755071;
assign addr[4316]= 2136037160;
assign addr[4317]= 2139641764;
assign addr[4318]= 2142567738;
assign addr[4319]= 2144814157;
assign addr[4320]= 2146380306;
assign addr[4321]= 2147265689;
assign addr[4322]= 2147470025;
assign addr[4323]= 2146993250;
assign addr[4324]= 2145835515;
assign addr[4325]= 2143997187;
assign addr[4326]= 2141478848;
assign addr[4327]= 2138281298;
assign addr[4328]= 2134405552;
assign addr[4329]= 2129852837;
assign addr[4330]= 2124624598;
assign addr[4331]= 2118722494;
assign addr[4332]= 2112148396;
assign addr[4333]= 2104904390;
assign addr[4334]= 2096992772;
assign addr[4335]= 2088416053;
assign addr[4336]= 2079176953;
assign addr[4337]= 2069278401;
assign addr[4338]= 2058723538;
assign addr[4339]= 2047515711;
assign addr[4340]= 2035658475;
assign addr[4341]= 2023155591;
assign addr[4342]= 2010011024;
assign addr[4343]= 1996228943;
assign addr[4344]= 1981813720;
assign addr[4345]= 1966769926;
assign addr[4346]= 1951102334;
assign addr[4347]= 1934815911;
assign addr[4348]= 1917915825;
assign addr[4349]= 1900407434;
assign addr[4350]= 1882296293;
assign addr[4351]= 1863588145;
assign addr[4352]= 1844288924;
assign addr[4353]= 1824404752;
assign addr[4354]= 1803941934;
assign addr[4355]= 1782906961;
assign addr[4356]= 1761306505;
assign addr[4357]= 1739147417;
assign addr[4358]= 1716436725;
assign addr[4359]= 1693181631;
assign addr[4360]= 1669389513;
assign addr[4361]= 1645067915;
assign addr[4362]= 1620224553;
assign addr[4363]= 1594867305;
assign addr[4364]= 1569004214;
assign addr[4365]= 1542643483;
assign addr[4366]= 1515793473;
assign addr[4367]= 1488462700;
assign addr[4368]= 1460659832;
assign addr[4369]= 1432393688;
assign addr[4370]= 1403673233;
assign addr[4371]= 1374507575;
assign addr[4372]= 1344905966;
assign addr[4373]= 1314877795;
assign addr[4374]= 1284432584;
assign addr[4375]= 1253579991;
assign addr[4376]= 1222329801;
assign addr[4377]= 1190691925;
assign addr[4378]= 1158676398;
assign addr[4379]= 1126293375;
assign addr[4380]= 1093553126;
assign addr[4381]= 1060466036;
assign addr[4382]= 1027042599;
assign addr[4383]= 993293415;
assign addr[4384]= 959229189;
assign addr[4385]= 924860725;
assign addr[4386]= 890198924;
assign addr[4387]= 855254778;
assign addr[4388]= 820039373;
assign addr[4389]= 784563876;
assign addr[4390]= 748839539;
assign addr[4391]= 712877694;
assign addr[4392]= 676689746;
assign addr[4393]= 640287172;
assign addr[4394]= 603681519;
assign addr[4395]= 566884397;
assign addr[4396]= 529907477;
assign addr[4397]= 492762486;
assign addr[4398]= 455461206;
assign addr[4399]= 418015468;
assign addr[4400]= 380437148;
assign addr[4401]= 342738165;
assign addr[4402]= 304930476;
assign addr[4403]= 267026072;
assign addr[4404]= 229036977;
assign addr[4405]= 190975237;
assign addr[4406]= 152852926;
assign addr[4407]= 114682135;
assign addr[4408]= 76474970;
assign addr[4409]= 38243550;
assign addr[4410]= 0;
assign addr[4411]= -38243550;
assign addr[4412]= -76474970;
assign addr[4413]= -114682135;
assign addr[4414]= -152852926;
assign addr[4415]= -190975237;
assign addr[4416]= -229036977;
assign addr[4417]= -267026072;
assign addr[4418]= -304930476;
assign addr[4419]= -342738165;
assign addr[4420]= -380437148;
assign addr[4421]= -418015468;
assign addr[4422]= -455461206;
assign addr[4423]= -492762486;
assign addr[4424]= -529907477;
assign addr[4425]= -566884397;
assign addr[4426]= -603681519;
assign addr[4427]= -640287172;
assign addr[4428]= -676689746;
assign addr[4429]= -712877694;
assign addr[4430]= -748839539;
assign addr[4431]= -784563876;
assign addr[4432]= -820039373;
assign addr[4433]= -855254778;
assign addr[4434]= -890198924;
assign addr[4435]= -924860725;
assign addr[4436]= -959229189;
assign addr[4437]= -993293415;
assign addr[4438]= -1027042599;
assign addr[4439]= -1060466036;
assign addr[4440]= -1093553126;
assign addr[4441]= -1126293375;
assign addr[4442]= -1158676398;
assign addr[4443]= -1190691925;
assign addr[4444]= -1222329801;
assign addr[4445]= -1253579991;
assign addr[4446]= -1284432584;
assign addr[4447]= -1314877795;
assign addr[4448]= -1344905966;
assign addr[4449]= -1374507575;
assign addr[4450]= -1403673233;
assign addr[4451]= -1432393688;
assign addr[4452]= -1460659832;
assign addr[4453]= -1488462700;
assign addr[4454]= -1515793473;
assign addr[4455]= -1542643483;
assign addr[4456]= -1569004214;
assign addr[4457]= -1594867305;
assign addr[4458]= -1620224553;
assign addr[4459]= -1645067915;
assign addr[4460]= -1669389513;
assign addr[4461]= -1693181631;
assign addr[4462]= -1716436725;
assign addr[4463]= -1739147417;
assign addr[4464]= -1761306505;
assign addr[4465]= -1782906961;
assign addr[4466]= -1803941934;
assign addr[4467]= -1824404752;
assign addr[4468]= -1844288924;
assign addr[4469]= -1863588145;
assign addr[4470]= -1882296293;
assign addr[4471]= -1900407434;
assign addr[4472]= -1917915825;
assign addr[4473]= -1934815911;
assign addr[4474]= -1951102334;
assign addr[4475]= -1966769926;
assign addr[4476]= -1981813720;
assign addr[4477]= -1996228943;
assign addr[4478]= -2010011024;
assign addr[4479]= -2023155591;
assign addr[4480]= -2035658475;
assign addr[4481]= -2047515711;
assign addr[4482]= -2058723538;
assign addr[4483]= -2069278401;
assign addr[4484]= -2079176953;
assign addr[4485]= -2088416053;
assign addr[4486]= -2096992772;
assign addr[4487]= -2104904390;
assign addr[4488]= -2112148396;
assign addr[4489]= -2118722494;
assign addr[4490]= -2124624598;
assign addr[4491]= -2129852837;
assign addr[4492]= -2134405552;
assign addr[4493]= -2138281298;
assign addr[4494]= -2141478848;
assign addr[4495]= -2143997187;
assign addr[4496]= -2145835515;
assign addr[4497]= -2146993250;
assign addr[4498]= -2147470025;
assign addr[4499]= -2147265689;
assign addr[4500]= -2146380306;
assign addr[4501]= -2144814157;
assign addr[4502]= -2142567738;
assign addr[4503]= -2139641764;
assign addr[4504]= -2136037160;
assign addr[4505]= -2131755071;
assign addr[4506]= -2126796855;
assign addr[4507]= -2121164085;
assign addr[4508]= -2114858546;
assign addr[4509]= -2107882239;
assign addr[4510]= -2100237377;
assign addr[4511]= -2091926384;
assign addr[4512]= -2082951896;
assign addr[4513]= -2073316760;
assign addr[4514]= -2063024031;
assign addr[4515]= -2052076975;
assign addr[4516]= -2040479063;
assign addr[4517]= -2028233973;
assign addr[4518]= -2015345591;
assign addr[4519]= -2001818002;
assign addr[4520]= -1987655498;
assign addr[4521]= -1972862571;
assign addr[4522]= -1957443913;
assign addr[4523]= -1941404413;
assign addr[4524]= -1924749160;
assign addr[4525]= -1907483436;
assign addr[4526]= -1889612716;
assign addr[4527]= -1871142669;
assign addr[4528]= -1852079154;
assign addr[4529]= -1832428215;
assign addr[4530]= -1812196087;
assign addr[4531]= -1791389186;
assign addr[4532]= -1770014111;
assign addr[4533]= -1748077642;
assign addr[4534]= -1725586737;
assign addr[4535]= -1702548529;
assign addr[4536]= -1678970324;
assign addr[4537]= -1654859602;
assign addr[4538]= -1630224009;
assign addr[4539]= -1605071359;
assign addr[4540]= -1579409630;
assign addr[4541]= -1553246960;
assign addr[4542]= -1526591649;
assign addr[4543]= -1499452149;
assign addr[4544]= -1471837070;
assign addr[4545]= -1443755168;
assign addr[4546]= -1415215352;
assign addr[4547]= -1386226674;
assign addr[4548]= -1356798326;
assign addr[4549]= -1326939644;
assign addr[4550]= -1296660098;
assign addr[4551]= -1265969291;
assign addr[4552]= -1234876957;
assign addr[4553]= -1203392958;
assign addr[4554]= -1171527280;
assign addr[4555]= -1139290029;
assign addr[4556]= -1106691431;
assign addr[4557]= -1073741824;
assign addr[4558]= -1040451659;
assign addr[4559]= -1006831495;
assign addr[4560]= -972891995;
assign addr[4561]= -938643924;
assign addr[4562]= -904098143;
assign addr[4563]= -869265610;
assign addr[4564]= -834157373;
assign addr[4565]= -798784567;
assign addr[4566]= -763158411;
assign addr[4567]= -727290205;
assign addr[4568]= -691191324;
assign addr[4569]= -654873219;
assign addr[4570]= -618347408;
assign addr[4571]= -581625477;
assign addr[4572]= -544719071;
assign addr[4573]= -507639898;
assign addr[4574]= -470399716;
assign addr[4575]= -433010339;
assign addr[4576]= -395483624;
assign addr[4577]= -357831473;
assign addr[4578]= -320065829;
assign addr[4579]= -282198671;
assign addr[4580]= -244242007;
assign addr[4581]= -206207878;
assign addr[4582]= -168108346;
assign addr[4583]= -129955495;
assign addr[4584]= -91761426;
assign addr[4585]= -53538253;
assign addr[4586]= -15298099;
assign addr[4587]= 22946906;
assign addr[4588]= 61184634;
assign addr[4589]= 99402956;
assign addr[4590]= 137589750;
assign addr[4591]= 175732905;
assign addr[4592]= 213820322;
assign addr[4593]= 251839923;
assign addr[4594]= 289779648;
assign addr[4595]= 327627463;
assign addr[4596]= 365371365;
assign addr[4597]= 402999383;
assign addr[4598]= 440499581;
assign addr[4599]= 477860067;
assign addr[4600]= 515068990;
assign addr[4601]= 552114549;
assign addr[4602]= 588984994;
assign addr[4603]= 625668632;
assign addr[4604]= 662153826;
assign addr[4605]= 698429006;
assign addr[4606]= 734482665;
assign addr[4607]= 770303369;
assign addr[4608]= 805879757;
assign addr[4609]= 841200544;
assign addr[4610]= 876254528;
assign addr[4611]= 911030591;
assign addr[4612]= 945517704;
assign addr[4613]= 979704927;
assign addr[4614]= 1013581418;
assign addr[4615]= 1047136432;
assign addr[4616]= 1080359326;
assign addr[4617]= 1113239564;
assign addr[4618]= 1145766716;
assign addr[4619]= 1177930466;
assign addr[4620]= 1209720613;
assign addr[4621]= 1241127074;
assign addr[4622]= 1272139887;
assign addr[4623]= 1302749217;
assign addr[4624]= 1332945355;
assign addr[4625]= 1362718723;
assign addr[4626]= 1392059879;
assign addr[4627]= 1420959516;
assign addr[4628]= 1449408469;
assign addr[4629]= 1477397714;
assign addr[4630]= 1504918373;
assign addr[4631]= 1531961719;
assign addr[4632]= 1558519173;
assign addr[4633]= 1584582314;
assign addr[4634]= 1610142873;
assign addr[4635]= 1635192744;
assign addr[4636]= 1659723983;
assign addr[4637]= 1683728808;
assign addr[4638]= 1707199606;
assign addr[4639]= 1730128933;
assign addr[4640]= 1752509516;
assign addr[4641]= 1774334257;
assign addr[4642]= 1795596234;
assign addr[4643]= 1816288703;
assign addr[4644]= 1836405100;
assign addr[4645]= 1855939047;
assign addr[4646]= 1874884346;
assign addr[4647]= 1893234990;
assign addr[4648]= 1910985158;
assign addr[4649]= 1928129220;
assign addr[4650]= 1944661739;
assign addr[4651]= 1960577471;
assign addr[4652]= 1975871368;
assign addr[4653]= 1990538579;
assign addr[4654]= 2004574453;
assign addr[4655]= 2017974537;
assign addr[4656]= 2030734582;
assign addr[4657]= 2042850540;
assign addr[4658]= 2054318569;
assign addr[4659]= 2065135031;
assign addr[4660]= 2075296495;
assign addr[4661]= 2084799740;
assign addr[4662]= 2093641749;
assign addr[4663]= 2101819720;
assign addr[4664]= 2109331059;
assign addr[4665]= 2116173382;
assign addr[4666]= 2122344521;
assign addr[4667]= 2127842516;
assign addr[4668]= 2132665626;
assign addr[4669]= 2136812319;
assign addr[4670]= 2140281282;
assign addr[4671]= 2143071413;
assign addr[4672]= 2145181827;
assign addr[4673]= 2146611856;
assign addr[4674]= 2147361045;
assign addr[4675]= 2147429158;
assign addr[4676]= 2146816171;
assign addr[4677]= 2145522281;
assign addr[4678]= 2143547897;
assign addr[4679]= 2140893646;
assign addr[4680]= 2137560369;
assign addr[4681]= 2133549123;
assign addr[4682]= 2128861181;
assign addr[4683]= 2123498030;
assign addr[4684]= 2117461370;
assign addr[4685]= 2110753117;
assign addr[4686]= 2103375398;
assign addr[4687]= 2095330553;
assign addr[4688]= 2086621133;
assign addr[4689]= 2077249901;
assign addr[4690]= 2067219829;
assign addr[4691]= 2056534099;
assign addr[4692]= 2045196100;
assign addr[4693]= 2033209426;
assign addr[4694]= 2020577882;
assign addr[4695]= 2007305472;
assign addr[4696]= 1993396407;
assign addr[4697]= 1978855097;
assign addr[4698]= 1963686155;
assign addr[4699]= 1947894393;
assign addr[4700]= 1931484818;
assign addr[4701]= 1914462636;
assign addr[4702]= 1896833245;
assign addr[4703]= 1878602237;
assign addr[4704]= 1859775393;
assign addr[4705]= 1840358687;
assign addr[4706]= 1820358275;
assign addr[4707]= 1799780501;
assign addr[4708]= 1778631892;
assign addr[4709]= 1756919156;
assign addr[4710]= 1734649179;
assign addr[4711]= 1711829025;
assign addr[4712]= 1688465931;
assign addr[4713]= 1664567307;
assign addr[4714]= 1640140734;
assign addr[4715]= 1615193959;
assign addr[4716]= 1589734894;
assign addr[4717]= 1563771613;
assign addr[4718]= 1537312353;
assign addr[4719]= 1510365504;
assign addr[4720]= 1482939614;
assign addr[4721]= 1455043381;
assign addr[4722]= 1426685652;
assign addr[4723]= 1397875423;
assign addr[4724]= 1368621831;
assign addr[4725]= 1338934154;
assign addr[4726]= 1308821808;
assign addr[4727]= 1278294345;
assign addr[4728]= 1247361445;
assign addr[4729]= 1216032921;
assign addr[4730]= 1184318708;
assign addr[4731]= 1152228866;
assign addr[4732]= 1119773573;
assign addr[4733]= 1086963121;
assign addr[4734]= 1053807919;
assign addr[4735]= 1020318481;
assign addr[4736]= 986505429;
assign addr[4737]= 952379488;
assign addr[4738]= 917951481;
assign addr[4739]= 883232329;
assign addr[4740]= 848233042;
assign addr[4741]= 812964722;
assign addr[4742]= 777438554;
assign addr[4743]= 741665807;
assign addr[4744]= 705657826;
assign addr[4745]= 669426032;
assign addr[4746]= 632981917;
assign addr[4747]= 596337040;
assign addr[4748]= 559503022;
assign addr[4749]= 522491548;
assign addr[4750]= 485314355;
assign addr[4751]= 447983235;
assign addr[4752]= 410510029;
assign addr[4753]= 372906622;
assign addr[4754]= 335184940;
assign addr[4755]= 297356948;
assign addr[4756]= 259434643;
assign addr[4757]= 221430054;
assign addr[4758]= 183355234;
assign addr[4759]= 145222259;
assign addr[4760]= 107043224;
assign addr[4761]= 68830239;
assign addr[4762]= 30595422;
assign addr[4763]= -7649098;
assign addr[4764]= -45891193;
assign addr[4765]= -84118732;
assign addr[4766]= -122319591;
assign addr[4767]= -160481654;
assign addr[4768]= -198592817;
assign addr[4769]= -236640993;
assign addr[4770]= -274614114;
assign addr[4771]= -312500135;
assign addr[4772]= -350287041;
assign addr[4773]= -387962847;
assign addr[4774]= -425515602;
assign addr[4775]= -462933398;
assign addr[4776]= -500204365;
assign addr[4777]= -537316682;
assign addr[4778]= -574258580;
assign addr[4779]= -611018340;
assign addr[4780]= -647584304;
assign addr[4781]= -683944874;
assign addr[4782]= -720088517;
assign addr[4783]= -756003771;
assign addr[4784]= -791679244;
assign addr[4785]= -827103620;
assign addr[4786]= -862265664;
assign addr[4787]= -897154224;
assign addr[4788]= -931758235;
assign addr[4789]= -966066720;
assign addr[4790]= -1000068799;
assign addr[4791]= -1033753687;
assign addr[4792]= -1067110699;
assign addr[4793]= -1100129257;
assign addr[4794]= -1132798888;
assign addr[4795]= -1165109230;
assign addr[4796]= -1197050035;
assign addr[4797]= -1228611172;
assign addr[4798]= -1259782632;
assign addr[4799]= -1290554528;
assign addr[4800]= -1320917099;
assign addr[4801]= -1350860716;
assign addr[4802]= -1380375881;
assign addr[4803]= -1409453233;
assign addr[4804]= -1438083551;
assign addr[4805]= -1466257752;
assign addr[4806]= -1493966902;
assign addr[4807]= -1521202211;
assign addr[4808]= -1547955041;
assign addr[4809]= -1574216908;
assign addr[4810]= -1599979481;
assign addr[4811]= -1625234591;
assign addr[4812]= -1649974225;
assign addr[4813]= -1674190539;
assign addr[4814]= -1697875851;
assign addr[4815]= -1721022648;
assign addr[4816]= -1743623590;
assign addr[4817]= -1765671509;
assign addr[4818]= -1787159411;
assign addr[4819]= -1808080480;
assign addr[4820]= -1828428082;
assign addr[4821]= -1848195763;
assign addr[4822]= -1867377253;
assign addr[4823]= -1885966468;
assign addr[4824]= -1903957513;
assign addr[4825]= -1921344681;
assign addr[4826]= -1938122457;
assign addr[4827]= -1954285520;
assign addr[4828]= -1969828744;
assign addr[4829]= -1984747199;
assign addr[4830]= -1999036154;
assign addr[4831]= -2012691075;
assign addr[4832]= -2025707632;
assign addr[4833]= -2038081698;
assign addr[4834]= -2049809346;
assign addr[4835]= -2060886858;
assign addr[4836]= -2071310720;
assign addr[4837]= -2081077626;
assign addr[4838]= -2090184478;
assign addr[4839]= -2098628387;
assign addr[4840]= -2106406677;
assign addr[4841]= -2113516878;
assign addr[4842]= -2119956737;
assign addr[4843]= -2125724211;
assign addr[4844]= -2130817471;
assign addr[4845]= -2135234901;
assign addr[4846]= -2138975100;
assign addr[4847]= -2142036881;
assign addr[4848]= -2144419275;
assign addr[4849]= -2146121524;
assign addr[4850]= -2147143090;
assign addr[4851]= -2147483648;
assign addr[4852]= -2147143090;
assign addr[4853]= -2146121524;
assign addr[4854]= -2144419275;
assign addr[4855]= -2142036881;
assign addr[4856]= -2138975100;
assign addr[4857]= -2135234901;
assign addr[4858]= -2130817471;
assign addr[4859]= -2125724211;
assign addr[4860]= -2119956737;
assign addr[4861]= -2113516878;
assign addr[4862]= -2106406677;
assign addr[4863]= -2098628387;
assign addr[4864]= -2090184478;
assign addr[4865]= -2081077626;
assign addr[4866]= -2071310720;
assign addr[4867]= -2060886858;
assign addr[4868]= -2049809346;
assign addr[4869]= -2038081698;
assign addr[4870]= -2025707632;
assign addr[4871]= -2012691075;
assign addr[4872]= -1999036154;
assign addr[4873]= -1984747199;
assign addr[4874]= -1969828744;
assign addr[4875]= -1954285520;
assign addr[4876]= -1938122457;
assign addr[4877]= -1921344681;
assign addr[4878]= -1903957513;
assign addr[4879]= -1885966468;
assign addr[4880]= -1867377253;
assign addr[4881]= -1848195763;
assign addr[4882]= -1828428082;
assign addr[4883]= -1808080480;
assign addr[4884]= -1787159411;
assign addr[4885]= -1765671509;
assign addr[4886]= -1743623590;
assign addr[4887]= -1721022648;
assign addr[4888]= -1697875851;
assign addr[4889]= -1674190539;
assign addr[4890]= -1649974225;
assign addr[4891]= -1625234591;
assign addr[4892]= -1599979481;
assign addr[4893]= -1574216908;
assign addr[4894]= -1547955041;
assign addr[4895]= -1521202211;
assign addr[4896]= -1493966902;
assign addr[4897]= -1466257752;
assign addr[4898]= -1438083551;
assign addr[4899]= -1409453233;
assign addr[4900]= -1380375881;
assign addr[4901]= -1350860716;
assign addr[4902]= -1320917099;
assign addr[4903]= -1290554528;
assign addr[4904]= -1259782632;
assign addr[4905]= -1228611172;
assign addr[4906]= -1197050035;
assign addr[4907]= -1165109230;
assign addr[4908]= -1132798888;
assign addr[4909]= -1100129257;
assign addr[4910]= -1067110699;
assign addr[4911]= -1033753687;
assign addr[4912]= -1000068799;
assign addr[4913]= -966066720;
assign addr[4914]= -931758235;
assign addr[4915]= -897154224;
assign addr[4916]= -862265664;
assign addr[4917]= -827103620;
assign addr[4918]= -791679244;
assign addr[4919]= -756003771;
assign addr[4920]= -720088517;
assign addr[4921]= -683944874;
assign addr[4922]= -647584304;
assign addr[4923]= -611018340;
assign addr[4924]= -574258580;
assign addr[4925]= -537316682;
assign addr[4926]= -500204365;
assign addr[4927]= -462933398;
assign addr[4928]= -425515602;
assign addr[4929]= -387962847;
assign addr[4930]= -350287041;
assign addr[4931]= -312500135;
assign addr[4932]= -274614114;
assign addr[4933]= -236640993;
assign addr[4934]= -198592817;
assign addr[4935]= -160481654;
assign addr[4936]= -122319591;
assign addr[4937]= -84118732;
assign addr[4938]= -45891193;
assign addr[4939]= -7649098;
assign addr[4940]= 30595422;
assign addr[4941]= 68830239;
assign addr[4942]= 107043224;
assign addr[4943]= 145222259;
assign addr[4944]= 183355234;
assign addr[4945]= 221430054;
assign addr[4946]= 259434643;
assign addr[4947]= 297356948;
assign addr[4948]= 335184940;
assign addr[4949]= 372906622;
assign addr[4950]= 410510029;
assign addr[4951]= 447983235;
assign addr[4952]= 485314355;
assign addr[4953]= 522491548;
assign addr[4954]= 559503022;
assign addr[4955]= 596337040;
assign addr[4956]= 632981917;
assign addr[4957]= 669426032;
assign addr[4958]= 705657826;
assign addr[4959]= 741665807;
assign addr[4960]= 777438554;
assign addr[4961]= 812964722;
assign addr[4962]= 848233042;
assign addr[4963]= 883232329;
assign addr[4964]= 917951481;
assign addr[4965]= 952379488;
assign addr[4966]= 986505429;
assign addr[4967]= 1020318481;
assign addr[4968]= 1053807919;
assign addr[4969]= 1086963121;
assign addr[4970]= 1119773573;
assign addr[4971]= 1152228866;
assign addr[4972]= 1184318708;
assign addr[4973]= 1216032921;
assign addr[4974]= 1247361445;
assign addr[4975]= 1278294345;
assign addr[4976]= 1308821808;
assign addr[4977]= 1338934154;
assign addr[4978]= 1368621831;
assign addr[4979]= 1397875423;
assign addr[4980]= 1426685652;
assign addr[4981]= 1455043381;
assign addr[4982]= 1482939614;
assign addr[4983]= 1510365504;
assign addr[4984]= 1537312353;
assign addr[4985]= 1563771613;
assign addr[4986]= 1589734894;
assign addr[4987]= 1615193959;
assign addr[4988]= 1640140734;
assign addr[4989]= 1664567307;
assign addr[4990]= 1688465931;
assign addr[4991]= 1711829025;
assign addr[4992]= 1734649179;
assign addr[4993]= 1756919156;
assign addr[4994]= 1778631892;
assign addr[4995]= 1799780501;
assign addr[4996]= 1820358275;
assign addr[4997]= 1840358687;
assign addr[4998]= 1859775393;
assign addr[4999]= 1878602237;
assign addr[5000]= 1896833245;
assign addr[5001]= 1914462636;
assign addr[5002]= 1931484818;
assign addr[5003]= 1947894393;
assign addr[5004]= 1963686155;
assign addr[5005]= 1978855097;
assign addr[5006]= 1993396407;
assign addr[5007]= 2007305472;
assign addr[5008]= 2020577882;
assign addr[5009]= 2033209426;
assign addr[5010]= 2045196100;
assign addr[5011]= 2056534099;
assign addr[5012]= 2067219829;
assign addr[5013]= 2077249901;
assign addr[5014]= 2086621133;
assign addr[5015]= 2095330553;
assign addr[5016]= 2103375398;
assign addr[5017]= 2110753117;
assign addr[5018]= 2117461370;
assign addr[5019]= 2123498030;
assign addr[5020]= 2128861181;
assign addr[5021]= 2133549123;
assign addr[5022]= 2137560369;
assign addr[5023]= 2140893646;
assign addr[5024]= 2143547897;
assign addr[5025]= 2145522281;
assign addr[5026]= 2146816171;
assign addr[5027]= 2147429158;
assign addr[5028]= 2147361045;
assign addr[5029]= 2146611856;
assign addr[5030]= 2145181827;
assign addr[5031]= 2143071413;
assign addr[5032]= 2140281282;
assign addr[5033]= 2136812319;
assign addr[5034]= 2132665626;
assign addr[5035]= 2127842516;
assign addr[5036]= 2122344521;
assign addr[5037]= 2116173382;
assign addr[5038]= 2109331059;
assign addr[5039]= 2101819720;
assign addr[5040]= 2093641749;
assign addr[5041]= 2084799740;
assign addr[5042]= 2075296495;
assign addr[5043]= 2065135031;
assign addr[5044]= 2054318569;
assign addr[5045]= 2042850540;
assign addr[5046]= 2030734582;
assign addr[5047]= 2017974537;
assign addr[5048]= 2004574453;
assign addr[5049]= 1990538579;
assign addr[5050]= 1975871368;
assign addr[5051]= 1960577471;
assign addr[5052]= 1944661739;
assign addr[5053]= 1928129220;
assign addr[5054]= 1910985158;
assign addr[5055]= 1893234990;
assign addr[5056]= 1874884346;
assign addr[5057]= 1855939047;
assign addr[5058]= 1836405100;
assign addr[5059]= 1816288703;
assign addr[5060]= 1795596234;
assign addr[5061]= 1774334257;
assign addr[5062]= 1752509516;
assign addr[5063]= 1730128933;
assign addr[5064]= 1707199606;
assign addr[5065]= 1683728808;
assign addr[5066]= 1659723983;
assign addr[5067]= 1635192744;
assign addr[5068]= 1610142873;
assign addr[5069]= 1584582314;
assign addr[5070]= 1558519173;
assign addr[5071]= 1531961719;
assign addr[5072]= 1504918373;
assign addr[5073]= 1477397714;
assign addr[5074]= 1449408469;
assign addr[5075]= 1420959516;
assign addr[5076]= 1392059879;
assign addr[5077]= 1362718723;
assign addr[5078]= 1332945355;
assign addr[5079]= 1302749217;
assign addr[5080]= 1272139887;
assign addr[5081]= 1241127074;
assign addr[5082]= 1209720613;
assign addr[5083]= 1177930466;
assign addr[5084]= 1145766716;
assign addr[5085]= 1113239564;
assign addr[5086]= 1080359326;
assign addr[5087]= 1047136432;
assign addr[5088]= 1013581418;
assign addr[5089]= 979704927;
assign addr[5090]= 945517704;
assign addr[5091]= 911030591;
assign addr[5092]= 876254528;
assign addr[5093]= 841200544;
assign addr[5094]= 805879757;
assign addr[5095]= 770303369;
assign addr[5096]= 734482665;
assign addr[5097]= 698429006;
assign addr[5098]= 662153826;
assign addr[5099]= 625668632;
assign addr[5100]= 588984994;
assign addr[5101]= 552114549;
assign addr[5102]= 515068990;
assign addr[5103]= 477860067;
assign addr[5104]= 440499581;
assign addr[5105]= 402999383;
assign addr[5106]= 365371365;
assign addr[5107]= 327627463;
assign addr[5108]= 289779648;
assign addr[5109]= 251839923;
assign addr[5110]= 213820322;
assign addr[5111]= 175732905;
assign addr[5112]= 137589750;
assign addr[5113]= 99402956;
assign addr[5114]= 61184634;
assign addr[5115]= 22946906;
assign addr[5116]= -15298099;
assign addr[5117]= -53538253;
assign addr[5118]= -91761426;
assign addr[5119]= -129955495;
assign addr[5120]= -168108346;
assign addr[5121]= -206207878;
assign addr[5122]= -244242007;
assign addr[5123]= -282198671;
assign addr[5124]= -320065829;
assign addr[5125]= -357831473;
assign addr[5126]= -395483624;
assign addr[5127]= -433010339;
assign addr[5128]= -470399716;
assign addr[5129]= -507639898;
assign addr[5130]= -544719071;
assign addr[5131]= -581625477;
assign addr[5132]= -618347408;
assign addr[5133]= -654873219;
assign addr[5134]= -691191324;
assign addr[5135]= -727290205;
assign addr[5136]= -763158411;
assign addr[5137]= -798784567;
assign addr[5138]= -834157373;
assign addr[5139]= -869265610;
assign addr[5140]= -904098143;
assign addr[5141]= -938643924;
assign addr[5142]= -972891995;
assign addr[5143]= -1006831495;
assign addr[5144]= -1040451659;
assign addr[5145]= -1073741824;
assign addr[5146]= -1106691431;
assign addr[5147]= -1139290029;
assign addr[5148]= -1171527280;
assign addr[5149]= -1203392958;
assign addr[5150]= -1234876957;
assign addr[5151]= -1265969291;
assign addr[5152]= -1296660098;
assign addr[5153]= -1326939644;
assign addr[5154]= -1356798326;
assign addr[5155]= -1386226674;
assign addr[5156]= -1415215352;
assign addr[5157]= -1443755168;
assign addr[5158]= -1471837070;
assign addr[5159]= -1499452149;
assign addr[5160]= -1526591649;
assign addr[5161]= -1553246960;
assign addr[5162]= -1579409630;
assign addr[5163]= -1605071359;
assign addr[5164]= -1630224009;
assign addr[5165]= -1654859602;
assign addr[5166]= -1678970324;
assign addr[5167]= -1702548529;
assign addr[5168]= -1725586737;
assign addr[5169]= -1748077642;
assign addr[5170]= -1770014111;
assign addr[5171]= -1791389186;
assign addr[5172]= -1812196087;
assign addr[5173]= -1832428215;
assign addr[5174]= -1852079154;
assign addr[5175]= -1871142669;
assign addr[5176]= -1889612716;
assign addr[5177]= -1907483436;
assign addr[5178]= -1924749160;
assign addr[5179]= -1941404413;
assign addr[5180]= -1957443913;
assign addr[5181]= -1972862571;
assign addr[5182]= -1987655498;
assign addr[5183]= -2001818002;
assign addr[5184]= -2015345591;
assign addr[5185]= -2028233973;
assign addr[5186]= -2040479063;
assign addr[5187]= -2052076975;
assign addr[5188]= -2063024031;
assign addr[5189]= -2073316760;
assign addr[5190]= -2082951896;
assign addr[5191]= -2091926384;
assign addr[5192]= -2100237377;
assign addr[5193]= -2107882239;
assign addr[5194]= -2114858546;
assign addr[5195]= -2121164085;
assign addr[5196]= -2126796855;
assign addr[5197]= -2131755071;
assign addr[5198]= -2136037160;
assign addr[5199]= -2139641764;
assign addr[5200]= -2142567738;
assign addr[5201]= -2144814157;
assign addr[5202]= -2146380306;
assign addr[5203]= -2147265689;
assign addr[5204]= -2147470025;
assign addr[5205]= -2146993250;
assign addr[5206]= -2145835515;
assign addr[5207]= -2143997187;
assign addr[5208]= -2141478848;
assign addr[5209]= -2138281298;
assign addr[5210]= -2134405552;
assign addr[5211]= -2129852837;
assign addr[5212]= -2124624598;
assign addr[5213]= -2118722494;
assign addr[5214]= -2112148396;
assign addr[5215]= -2104904390;
assign addr[5216]= -2096992772;
assign addr[5217]= -2088416053;
assign addr[5218]= -2079176953;
assign addr[5219]= -2069278401;
assign addr[5220]= -2058723538;
assign addr[5221]= -2047515711;
assign addr[5222]= -2035658475;
assign addr[5223]= -2023155591;
assign addr[5224]= -2010011024;
assign addr[5225]= -1996228943;
assign addr[5226]= -1981813720;
assign addr[5227]= -1966769926;
assign addr[5228]= -1951102334;
assign addr[5229]= -1934815911;
assign addr[5230]= -1917915825;
assign addr[5231]= -1900407434;
assign addr[5232]= -1882296293;
assign addr[5233]= -1863588145;
assign addr[5234]= -1844288924;
assign addr[5235]= -1824404752;
assign addr[5236]= -1803941934;
assign addr[5237]= -1782906961;
assign addr[5238]= -1761306505;
assign addr[5239]= -1739147417;
assign addr[5240]= -1716436725;
assign addr[5241]= -1693181631;
assign addr[5242]= -1669389513;
assign addr[5243]= -1645067915;
assign addr[5244]= -1620224553;
assign addr[5245]= -1594867305;
assign addr[5246]= -1569004214;
assign addr[5247]= -1542643483;
assign addr[5248]= -1515793473;
assign addr[5249]= -1488462700;
assign addr[5250]= -1460659832;
assign addr[5251]= -1432393688;
assign addr[5252]= -1403673233;
assign addr[5253]= -1374507575;
assign addr[5254]= -1344905966;
assign addr[5255]= -1314877795;
assign addr[5256]= -1284432584;
assign addr[5257]= -1253579991;
assign addr[5258]= -1222329801;
assign addr[5259]= -1190691925;
assign addr[5260]= -1158676398;
assign addr[5261]= -1126293375;
assign addr[5262]= -1093553126;
assign addr[5263]= -1060466036;
assign addr[5264]= -1027042599;
assign addr[5265]= -993293415;
assign addr[5266]= -959229189;
assign addr[5267]= -924860725;
assign addr[5268]= -890198924;
assign addr[5269]= -855254778;
assign addr[5270]= -820039373;
assign addr[5271]= -784563876;
assign addr[5272]= -748839539;
assign addr[5273]= -712877694;
assign addr[5274]= -676689746;
assign addr[5275]= -640287172;
assign addr[5276]= -603681519;
assign addr[5277]= -566884397;
assign addr[5278]= -529907477;
assign addr[5279]= -492762486;
assign addr[5280]= -455461206;
assign addr[5281]= -418015468;
assign addr[5282]= -380437148;
assign addr[5283]= -342738165;
assign addr[5284]= -304930476;
assign addr[5285]= -267026072;
assign addr[5286]= -229036977;
assign addr[5287]= -190975237;
assign addr[5288]= -152852926;
assign addr[5289]= -114682135;
assign addr[5290]= -76474970;
assign addr[5291]= -38243550;
assign addr[5292]= 0;
assign addr[5293]= 38243550;
assign addr[5294]= 76474970;
assign addr[5295]= 114682135;
assign addr[5296]= 152852926;
assign addr[5297]= 190975237;
assign addr[5298]= 229036977;
assign addr[5299]= 267026072;
assign addr[5300]= 304930476;
assign addr[5301]= 342738165;
assign addr[5302]= 380437148;
assign addr[5303]= 418015468;
assign addr[5304]= 455461206;
assign addr[5305]= 492762486;
assign addr[5306]= 529907477;
assign addr[5307]= 566884397;
assign addr[5308]= 603681519;
assign addr[5309]= 640287172;
assign addr[5310]= 676689746;
assign addr[5311]= 712877694;
assign addr[5312]= 748839539;
assign addr[5313]= 784563876;
assign addr[5314]= 820039373;
assign addr[5315]= 855254778;
assign addr[5316]= 890198924;
assign addr[5317]= 924860725;
assign addr[5318]= 959229189;
assign addr[5319]= 993293415;
assign addr[5320]= 1027042599;
assign addr[5321]= 1060466036;
assign addr[5322]= 1093553126;
assign addr[5323]= 1126293375;
assign addr[5324]= 1158676398;
assign addr[5325]= 1190691925;
assign addr[5326]= 1222329801;
assign addr[5327]= 1253579991;
assign addr[5328]= 1284432584;
assign addr[5329]= 1314877795;
assign addr[5330]= 1344905966;
assign addr[5331]= 1374507575;
assign addr[5332]= 1403673233;
assign addr[5333]= 1432393688;
assign addr[5334]= 1460659832;
assign addr[5335]= 1488462700;
assign addr[5336]= 1515793473;
assign addr[5337]= 1542643483;
assign addr[5338]= 1569004214;
assign addr[5339]= 1594867305;
assign addr[5340]= 1620224553;
assign addr[5341]= 1645067915;
assign addr[5342]= 1669389513;
assign addr[5343]= 1693181631;
assign addr[5344]= 1716436725;
assign addr[5345]= 1739147417;
assign addr[5346]= 1761306505;
assign addr[5347]= 1782906961;
assign addr[5348]= 1803941934;
assign addr[5349]= 1824404752;
assign addr[5350]= 1844288924;
assign addr[5351]= 1863588145;
assign addr[5352]= 1882296293;
assign addr[5353]= 1900407434;
assign addr[5354]= 1917915825;
assign addr[5355]= 1934815911;
assign addr[5356]= 1951102334;
assign addr[5357]= 1966769926;
assign addr[5358]= 1981813720;
assign addr[5359]= 1996228943;
assign addr[5360]= 2010011024;
assign addr[5361]= 2023155591;
assign addr[5362]= 2035658475;
assign addr[5363]= 2047515711;
assign addr[5364]= 2058723538;
assign addr[5365]= 2069278401;
assign addr[5366]= 2079176953;
assign addr[5367]= 2088416053;
assign addr[5368]= 2096992772;
assign addr[5369]= 2104904390;
assign addr[5370]= 2112148396;
assign addr[5371]= 2118722494;
assign addr[5372]= 2124624598;
assign addr[5373]= 2129852837;
assign addr[5374]= 2134405552;
assign addr[5375]= 2138281298;
assign addr[5376]= 2141478848;
assign addr[5377]= 2143997187;
assign addr[5378]= 2145835515;
assign addr[5379]= 2146993250;
assign addr[5380]= 2147470025;
assign addr[5381]= 2147265689;
assign addr[5382]= 2146380306;
assign addr[5383]= 2144814157;
assign addr[5384]= 2142567738;
assign addr[5385]= 2139641764;
assign addr[5386]= 2136037160;
assign addr[5387]= 2131755071;
assign addr[5388]= 2126796855;
assign addr[5389]= 2121164085;
assign addr[5390]= 2114858546;
assign addr[5391]= 2107882239;
assign addr[5392]= 2100237377;
assign addr[5393]= 2091926384;
assign addr[5394]= 2082951896;
assign addr[5395]= 2073316760;
assign addr[5396]= 2063024031;
assign addr[5397]= 2052076975;
assign addr[5398]= 2040479063;
assign addr[5399]= 2028233973;
assign addr[5400]= 2015345591;
assign addr[5401]= 2001818002;
assign addr[5402]= 1987655498;
assign addr[5403]= 1972862571;
assign addr[5404]= 1957443913;
assign addr[5405]= 1941404413;
assign addr[5406]= 1924749160;
assign addr[5407]= 1907483436;
assign addr[5408]= 1889612716;
assign addr[5409]= 1871142669;
assign addr[5410]= 1852079154;
assign addr[5411]= 1832428215;
assign addr[5412]= 1812196087;
assign addr[5413]= 1791389186;
assign addr[5414]= 1770014111;
assign addr[5415]= 1748077642;
assign addr[5416]= 1725586737;
assign addr[5417]= 1702548529;
assign addr[5418]= 1678970324;
assign addr[5419]= 1654859602;
assign addr[5420]= 1630224009;
assign addr[5421]= 1605071359;
assign addr[5422]= 1579409630;
assign addr[5423]= 1553246960;
assign addr[5424]= 1526591649;
assign addr[5425]= 1499452149;
assign addr[5426]= 1471837070;
assign addr[5427]= 1443755168;
assign addr[5428]= 1415215352;
assign addr[5429]= 1386226674;
assign addr[5430]= 1356798326;
assign addr[5431]= 1326939644;
assign addr[5432]= 1296660098;
assign addr[5433]= 1265969291;
assign addr[5434]= 1234876957;
assign addr[5435]= 1203392958;
assign addr[5436]= 1171527280;
assign addr[5437]= 1139290029;
assign addr[5438]= 1106691431;
assign addr[5439]= 1073741824;
assign addr[5440]= 1040451659;
assign addr[5441]= 1006831495;
assign addr[5442]= 972891995;
assign addr[5443]= 938643924;
assign addr[5444]= 904098143;
assign addr[5445]= 869265610;
assign addr[5446]= 834157373;
assign addr[5447]= 798784567;
assign addr[5448]= 763158411;
assign addr[5449]= 727290205;
assign addr[5450]= 691191324;
assign addr[5451]= 654873219;
assign addr[5452]= 618347408;
assign addr[5453]= 581625477;
assign addr[5454]= 544719071;
assign addr[5455]= 507639898;
assign addr[5456]= 470399716;
assign addr[5457]= 433010339;
assign addr[5458]= 395483624;
assign addr[5459]= 357831473;
assign addr[5460]= 320065829;
assign addr[5461]= 282198671;
assign addr[5462]= 244242007;
assign addr[5463]= 206207878;
assign addr[5464]= 168108346;
assign addr[5465]= 129955495;
assign addr[5466]= 91761426;
assign addr[5467]= 53538253;
assign addr[5468]= 15298099;
assign addr[5469]= -22946906;
assign addr[5470]= -61184634;
assign addr[5471]= -99402956;
assign addr[5472]= -137589750;
assign addr[5473]= -175732905;
assign addr[5474]= -213820322;
assign addr[5475]= -251839923;
assign addr[5476]= -289779648;
assign addr[5477]= -327627463;
assign addr[5478]= -365371365;
assign addr[5479]= -402999383;
assign addr[5480]= -440499581;
assign addr[5481]= -477860067;
assign addr[5482]= -515068990;
assign addr[5483]= -552114549;
assign addr[5484]= -588984994;
assign addr[5485]= -625668632;
assign addr[5486]= -662153826;
assign addr[5487]= -698429006;
assign addr[5488]= -734482665;
assign addr[5489]= -770303369;
assign addr[5490]= -805879757;
assign addr[5491]= -841200544;
assign addr[5492]= -876254528;
assign addr[5493]= -911030591;
assign addr[5494]= -945517704;
assign addr[5495]= -979704927;
assign addr[5496]= -1013581418;
assign addr[5497]= -1047136432;
assign addr[5498]= -1080359326;
assign addr[5499]= -1113239564;
assign addr[5500]= -1145766716;
assign addr[5501]= -1177930466;
assign addr[5502]= -1209720613;
assign addr[5503]= -1241127074;
assign addr[5504]= -1272139887;
assign addr[5505]= -1302749217;
assign addr[5506]= -1332945355;
assign addr[5507]= -1362718723;
assign addr[5508]= -1392059879;
assign addr[5509]= -1420959516;
assign addr[5510]= -1449408469;
assign addr[5511]= -1477397714;
assign addr[5512]= -1504918373;
assign addr[5513]= -1531961719;
assign addr[5514]= -1558519173;
assign addr[5515]= -1584582314;
assign addr[5516]= -1610142873;
assign addr[5517]= -1635192744;
assign addr[5518]= -1659723983;
assign addr[5519]= -1683728808;
assign addr[5520]= -1707199606;
assign addr[5521]= -1730128933;
assign addr[5522]= -1752509516;
assign addr[5523]= -1774334257;
assign addr[5524]= -1795596234;
assign addr[5525]= -1816288703;
assign addr[5526]= -1836405100;
assign addr[5527]= -1855939047;
assign addr[5528]= -1874884346;
assign addr[5529]= -1893234990;
assign addr[5530]= -1910985158;
assign addr[5531]= -1928129220;
assign addr[5532]= -1944661739;
assign addr[5533]= -1960577471;
assign addr[5534]= -1975871368;
assign addr[5535]= -1990538579;
assign addr[5536]= -2004574453;
assign addr[5537]= -2017974537;
assign addr[5538]= -2030734582;
assign addr[5539]= -2042850540;
assign addr[5540]= -2054318569;
assign addr[5541]= -2065135031;
assign addr[5542]= -2075296495;
assign addr[5543]= -2084799740;
assign addr[5544]= -2093641749;
assign addr[5545]= -2101819720;
assign addr[5546]= -2109331059;
assign addr[5547]= -2116173382;
assign addr[5548]= -2122344521;
assign addr[5549]= -2127842516;
assign addr[5550]= -2132665626;
assign addr[5551]= -2136812319;
assign addr[5552]= -2140281282;
assign addr[5553]= -2143071413;
assign addr[5554]= -2145181827;
assign addr[5555]= -2146611856;
assign addr[5556]= -2147361045;
assign addr[5557]= -2147429158;
assign addr[5558]= -2146816171;
assign addr[5559]= -2145522281;
assign addr[5560]= -2143547897;
assign addr[5561]= -2140893646;
assign addr[5562]= -2137560369;
assign addr[5563]= -2133549123;
assign addr[5564]= -2128861181;
assign addr[5565]= -2123498030;
assign addr[5566]= -2117461370;
assign addr[5567]= -2110753117;
assign addr[5568]= -2103375398;
assign addr[5569]= -2095330553;
assign addr[5570]= -2086621133;
assign addr[5571]= -2077249901;
assign addr[5572]= -2067219829;
assign addr[5573]= -2056534099;
assign addr[5574]= -2045196100;
assign addr[5575]= -2033209426;
assign addr[5576]= -2020577882;
assign addr[5577]= -2007305472;
assign addr[5578]= -1993396407;
assign addr[5579]= -1978855097;
assign addr[5580]= -1963686155;
assign addr[5581]= -1947894393;
assign addr[5582]= -1931484818;
assign addr[5583]= -1914462636;
assign addr[5584]= -1896833245;
assign addr[5585]= -1878602237;
assign addr[5586]= -1859775393;
assign addr[5587]= -1840358687;
assign addr[5588]= -1820358275;
assign addr[5589]= -1799780501;
assign addr[5590]= -1778631892;
assign addr[5591]= -1756919156;
assign addr[5592]= -1734649179;
assign addr[5593]= -1711829025;
assign addr[5594]= -1688465931;
assign addr[5595]= -1664567307;
assign addr[5596]= -1640140734;
assign addr[5597]= -1615193959;
assign addr[5598]= -1589734894;
assign addr[5599]= -1563771613;
assign addr[5600]= -1537312353;
assign addr[5601]= -1510365504;
assign addr[5602]= -1482939614;
assign addr[5603]= -1455043381;
assign addr[5604]= -1426685652;
assign addr[5605]= -1397875423;
assign addr[5606]= -1368621831;
assign addr[5607]= -1338934154;
assign addr[5608]= -1308821808;
assign addr[5609]= -1278294345;
assign addr[5610]= -1247361445;
assign addr[5611]= -1216032921;
assign addr[5612]= -1184318708;
assign addr[5613]= -1152228866;
assign addr[5614]= -1119773573;
assign addr[5615]= -1086963121;
assign addr[5616]= -1053807919;
assign addr[5617]= -1020318481;
assign addr[5618]= -986505429;
assign addr[5619]= -952379488;
assign addr[5620]= -917951481;
assign addr[5621]= -883232329;
assign addr[5622]= -848233042;
assign addr[5623]= -812964722;
assign addr[5624]= -777438554;
assign addr[5625]= -741665807;
assign addr[5626]= -705657826;
assign addr[5627]= -669426032;
assign addr[5628]= -632981917;
assign addr[5629]= -596337040;
assign addr[5630]= -559503022;
assign addr[5631]= -522491548;
assign addr[5632]= -485314355;
assign addr[5633]= -447983235;
assign addr[5634]= -410510029;
assign addr[5635]= -372906622;
assign addr[5636]= -335184940;
assign addr[5637]= -297356948;
assign addr[5638]= -259434643;
assign addr[5639]= -221430054;
assign addr[5640]= -183355234;
assign addr[5641]= -145222259;
assign addr[5642]= -107043224;
assign addr[5643]= -68830239;
assign addr[5644]= -30595422;
assign addr[5645]= 7649098;
assign addr[5646]= 45891193;
assign addr[5647]= 84118732;
assign addr[5648]= 122319591;
assign addr[5649]= 160481654;
assign addr[5650]= 198592817;
assign addr[5651]= 236640993;
assign addr[5652]= 274614114;
assign addr[5653]= 312500135;
assign addr[5654]= 350287041;
assign addr[5655]= 387962847;
assign addr[5656]= 425515602;
assign addr[5657]= 462933398;
assign addr[5658]= 500204365;
assign addr[5659]= 537316682;
assign addr[5660]= 574258580;
assign addr[5661]= 611018340;
assign addr[5662]= 647584304;
assign addr[5663]= 683944874;
assign addr[5664]= 720088517;
assign addr[5665]= 756003771;
assign addr[5666]= 791679244;
assign addr[5667]= 827103620;
assign addr[5668]= 862265664;
assign addr[5669]= 897154224;
assign addr[5670]= 931758235;
assign addr[5671]= 966066720;
assign addr[5672]= 1000068799;
assign addr[5673]= 1033753687;
assign addr[5674]= 1067110699;
assign addr[5675]= 1100129257;
assign addr[5676]= 1132798888;
assign addr[5677]= 1165109230;
assign addr[5678]= 1197050035;
assign addr[5679]= 1228611172;
assign addr[5680]= 1259782632;
assign addr[5681]= 1290554528;
assign addr[5682]= 1320917099;
assign addr[5683]= 1350860716;
assign addr[5684]= 1380375881;
assign addr[5685]= 1409453233;
assign addr[5686]= 1438083551;
assign addr[5687]= 1466257752;
assign addr[5688]= 1493966902;
assign addr[5689]= 1521202211;
assign addr[5690]= 1547955041;
assign addr[5691]= 1574216908;
assign addr[5692]= 1599979481;
assign addr[5693]= 1625234591;
assign addr[5694]= 1649974225;
assign addr[5695]= 1674190539;
assign addr[5696]= 1697875851;
assign addr[5697]= 1721022648;
assign addr[5698]= 1743623590;
assign addr[5699]= 1765671509;
assign addr[5700]= 1787159411;
assign addr[5701]= 1808080480;
assign addr[5702]= 1828428082;
assign addr[5703]= 1848195763;
assign addr[5704]= 1867377253;
assign addr[5705]= 1885966468;
assign addr[5706]= 1903957513;
assign addr[5707]= 1921344681;
assign addr[5708]= 1938122457;
assign addr[5709]= 1954285520;
assign addr[5710]= 1969828744;
assign addr[5711]= 1984747199;
assign addr[5712]= 1999036154;
assign addr[5713]= 2012691075;
assign addr[5714]= 2025707632;
assign addr[5715]= 2038081698;
assign addr[5716]= 2049809346;
assign addr[5717]= 2060886858;
assign addr[5718]= 2071310720;
assign addr[5719]= 2081077626;
assign addr[5720]= 2090184478;
assign addr[5721]= 2098628387;
assign addr[5722]= 2106406677;
assign addr[5723]= 2113516878;
assign addr[5724]= 2119956737;
assign addr[5725]= 2125724211;
assign addr[5726]= 2130817471;
assign addr[5727]= 2135234901;
assign addr[5728]= 2138975100;
assign addr[5729]= 2142036881;
assign addr[5730]= 2144419275;
assign addr[5731]= 2146121524;
assign addr[5732]= 2147143090;
assign addr[5733]= 2147483648;
assign addr[5734]= 2147143090;
assign addr[5735]= 2146121524;
assign addr[5736]= 2144419275;
assign addr[5737]= 2142036881;
assign addr[5738]= 2138975100;
assign addr[5739]= 2135234901;
assign addr[5740]= 2130817471;
assign addr[5741]= 2125724211;
assign addr[5742]= 2119956737;
assign addr[5743]= 2113516878;
assign addr[5744]= 2106406677;
assign addr[5745]= 2098628387;
assign addr[5746]= 2090184478;
assign addr[5747]= 2081077626;
assign addr[5748]= 2071310720;
assign addr[5749]= 2060886858;
assign addr[5750]= 2049809346;
assign addr[5751]= 2038081698;
assign addr[5752]= 2025707632;
assign addr[5753]= 2012691075;
assign addr[5754]= 1999036154;
assign addr[5755]= 1984747199;
assign addr[5756]= 1969828744;
assign addr[5757]= 1954285520;
assign addr[5758]= 1938122457;
assign addr[5759]= 1921344681;
assign addr[5760]= 1903957513;
assign addr[5761]= 1885966468;
assign addr[5762]= 1867377253;
assign addr[5763]= 1848195763;
assign addr[5764]= 1828428082;
assign addr[5765]= 1808080480;
assign addr[5766]= 1787159411;
assign addr[5767]= 1765671509;
assign addr[5768]= 1743623590;
assign addr[5769]= 1721022648;
assign addr[5770]= 1697875851;
assign addr[5771]= 1674190539;
assign addr[5772]= 1649974225;
assign addr[5773]= 1625234591;
assign addr[5774]= 1599979481;
assign addr[5775]= 1574216908;
assign addr[5776]= 1547955041;
assign addr[5777]= 1521202211;
assign addr[5778]= 1493966902;
assign addr[5779]= 1466257752;
assign addr[5780]= 1438083551;
assign addr[5781]= 1409453233;
assign addr[5782]= 1380375881;
assign addr[5783]= 1350860716;
assign addr[5784]= 1320917099;
assign addr[5785]= 1290554528;
assign addr[5786]= 1259782632;
assign addr[5787]= 1228611172;
assign addr[5788]= 1197050035;
assign addr[5789]= 1165109230;
assign addr[5790]= 1132798888;
assign addr[5791]= 1100129257;
assign addr[5792]= 1067110699;
assign addr[5793]= 1033753687;
assign addr[5794]= 1000068799;
assign addr[5795]= 966066720;
assign addr[5796]= 931758235;
assign addr[5797]= 897154224;
assign addr[5798]= 862265664;
assign addr[5799]= 827103620;
assign addr[5800]= 791679244;
assign addr[5801]= 756003771;
assign addr[5802]= 720088517;
assign addr[5803]= 683944874;
assign addr[5804]= 647584304;
assign addr[5805]= 611018340;
assign addr[5806]= 574258580;
assign addr[5807]= 537316682;
assign addr[5808]= 500204365;
assign addr[5809]= 462933398;
assign addr[5810]= 425515602;
assign addr[5811]= 387962847;
assign addr[5812]= 350287041;
assign addr[5813]= 312500135;
assign addr[5814]= 274614114;
assign addr[5815]= 236640993;
assign addr[5816]= 198592817;
assign addr[5817]= 160481654;
assign addr[5818]= 122319591;
assign addr[5819]= 84118732;
assign addr[5820]= 45891193;
assign addr[5821]= 7649098;
assign addr[5822]= -30595422;
assign addr[5823]= -68830239;
assign addr[5824]= -107043224;
assign addr[5825]= -145222259;
assign addr[5826]= -183355234;
assign addr[5827]= -221430054;
assign addr[5828]= -259434643;
assign addr[5829]= -297356948;
assign addr[5830]= -335184940;
assign addr[5831]= -372906622;
assign addr[5832]= -410510029;
assign addr[5833]= -447983235;
assign addr[5834]= -485314355;
assign addr[5835]= -522491548;
assign addr[5836]= -559503022;
assign addr[5837]= -596337040;
assign addr[5838]= -632981917;
assign addr[5839]= -669426032;
assign addr[5840]= -705657826;
assign addr[5841]= -741665807;
assign addr[5842]= -777438554;
assign addr[5843]= -812964722;
assign addr[5844]= -848233042;
assign addr[5845]= -883232329;
assign addr[5846]= -917951481;
assign addr[5847]= -952379488;
assign addr[5848]= -986505429;
assign addr[5849]= -1020318481;
assign addr[5850]= -1053807919;
assign addr[5851]= -1086963121;
assign addr[5852]= -1119773573;
assign addr[5853]= -1152228866;
assign addr[5854]= -1184318708;
assign addr[5855]= -1216032921;
assign addr[5856]= -1247361445;
assign addr[5857]= -1278294345;
assign addr[5858]= -1308821808;
assign addr[5859]= -1338934154;
assign addr[5860]= -1368621831;
assign addr[5861]= -1397875423;
assign addr[5862]= -1426685652;
assign addr[5863]= -1455043381;
assign addr[5864]= -1482939614;
assign addr[5865]= -1510365504;
assign addr[5866]= -1537312353;
assign addr[5867]= -1563771613;
assign addr[5868]= -1589734894;
assign addr[5869]= -1615193959;
assign addr[5870]= -1640140734;
assign addr[5871]= -1664567307;
assign addr[5872]= -1688465931;
assign addr[5873]= -1711829025;
assign addr[5874]= -1734649179;
assign addr[5875]= -1756919156;
assign addr[5876]= -1778631892;
assign addr[5877]= -1799780501;
assign addr[5878]= -1820358275;
assign addr[5879]= -1840358687;
assign addr[5880]= -1859775393;
assign addr[5881]= -1878602237;
assign addr[5882]= -1896833245;
assign addr[5883]= -1914462636;
assign addr[5884]= -1931484818;
assign addr[5885]= -1947894393;
assign addr[5886]= -1963686155;
assign addr[5887]= -1978855097;
assign addr[5888]= -1993396407;
assign addr[5889]= -2007305472;
assign addr[5890]= -2020577882;
assign addr[5891]= -2033209426;
assign addr[5892]= -2045196100;
assign addr[5893]= -2056534099;
assign addr[5894]= -2067219829;
assign addr[5895]= -2077249901;
assign addr[5896]= -2086621133;
assign addr[5897]= -2095330553;
assign addr[5898]= -2103375398;
assign addr[5899]= -2110753117;
assign addr[5900]= -2117461370;
assign addr[5901]= -2123498030;
assign addr[5902]= -2128861181;
assign addr[5903]= -2133549123;
assign addr[5904]= -2137560369;
assign addr[5905]= -2140893646;
assign addr[5906]= -2143547897;
assign addr[5907]= -2145522281;
assign addr[5908]= -2146816171;
assign addr[5909]= -2147429158;
assign addr[5910]= -2147361045;
assign addr[5911]= -2146611856;
assign addr[5912]= -2145181827;
assign addr[5913]= -2143071413;
assign addr[5914]= -2140281282;
assign addr[5915]= -2136812319;
assign addr[5916]= -2132665626;
assign addr[5917]= -2127842516;
assign addr[5918]= -2122344521;
assign addr[5919]= -2116173382;
assign addr[5920]= -2109331059;
assign addr[5921]= -2101819720;
assign addr[5922]= -2093641749;
assign addr[5923]= -2084799740;
assign addr[5924]= -2075296495;
assign addr[5925]= -2065135031;
assign addr[5926]= -2054318569;
assign addr[5927]= -2042850540;
assign addr[5928]= -2030734582;
assign addr[5929]= -2017974537;
assign addr[5930]= -2004574453;
assign addr[5931]= -1990538579;
assign addr[5932]= -1975871368;
assign addr[5933]= -1960577471;
assign addr[5934]= -1944661739;
assign addr[5935]= -1928129220;
assign addr[5936]= -1910985158;
assign addr[5937]= -1893234990;
assign addr[5938]= -1874884346;
assign addr[5939]= -1855939047;
assign addr[5940]= -1836405100;
assign addr[5941]= -1816288703;
assign addr[5942]= -1795596234;
assign addr[5943]= -1774334257;
assign addr[5944]= -1752509516;
assign addr[5945]= -1730128933;
assign addr[5946]= -1707199606;
assign addr[5947]= -1683728808;
assign addr[5948]= -1659723983;
assign addr[5949]= -1635192744;
assign addr[5950]= -1610142873;
assign addr[5951]= -1584582314;
assign addr[5952]= -1558519173;
assign addr[5953]= -1531961719;
assign addr[5954]= -1504918373;
assign addr[5955]= -1477397714;
assign addr[5956]= -1449408469;
assign addr[5957]= -1420959516;
assign addr[5958]= -1392059879;
assign addr[5959]= -1362718723;
assign addr[5960]= -1332945355;
assign addr[5961]= -1302749217;
assign addr[5962]= -1272139887;
assign addr[5963]= -1241127074;
assign addr[5964]= -1209720613;
assign addr[5965]= -1177930466;
assign addr[5966]= -1145766716;
assign addr[5967]= -1113239564;
assign addr[5968]= -1080359326;
assign addr[5969]= -1047136432;
assign addr[5970]= -1013581418;
assign addr[5971]= -979704927;
assign addr[5972]= -945517704;
assign addr[5973]= -911030591;
assign addr[5974]= -876254528;
assign addr[5975]= -841200544;
assign addr[5976]= -805879757;
assign addr[5977]= -770303369;
assign addr[5978]= -734482665;
assign addr[5979]= -698429006;
assign addr[5980]= -662153826;
assign addr[5981]= -625668632;
assign addr[5982]= -588984994;
assign addr[5983]= -552114549;
assign addr[5984]= -515068990;
assign addr[5985]= -477860067;
assign addr[5986]= -440499581;
assign addr[5987]= -402999383;
assign addr[5988]= -365371365;
assign addr[5989]= -327627463;
assign addr[5990]= -289779648;
assign addr[5991]= -251839923;
assign addr[5992]= -213820322;
assign addr[5993]= -175732905;
assign addr[5994]= -137589750;
assign addr[5995]= -99402956;
assign addr[5996]= -61184634;
assign addr[5997]= -22946906;
assign addr[5998]= 15298099;
assign addr[5999]= 53538253;
assign addr[6000]= 91761426;
assign addr[6001]= 129955495;
assign addr[6002]= 168108346;
assign addr[6003]= 206207878;
assign addr[6004]= 244242007;
assign addr[6005]= 282198671;
assign addr[6006]= 320065829;
assign addr[6007]= 357831473;
assign addr[6008]= 395483624;
assign addr[6009]= 433010339;
assign addr[6010]= 470399716;
assign addr[6011]= 507639898;
assign addr[6012]= 544719071;
assign addr[6013]= 581625477;
assign addr[6014]= 618347408;
assign addr[6015]= 654873219;
assign addr[6016]= 691191324;
assign addr[6017]= 727290205;
assign addr[6018]= 763158411;
assign addr[6019]= 798784567;
assign addr[6020]= 834157373;
assign addr[6021]= 869265610;
assign addr[6022]= 904098143;
assign addr[6023]= 938643924;
assign addr[6024]= 972891995;
assign addr[6025]= 1006831495;
assign addr[6026]= 1040451659;
assign addr[6027]= 1073741824;
assign addr[6028]= 1106691431;
assign addr[6029]= 1139290029;
assign addr[6030]= 1171527280;
assign addr[6031]= 1203392958;
assign addr[6032]= 1234876957;
assign addr[6033]= 1265969291;
assign addr[6034]= 1296660098;
assign addr[6035]= 1326939644;
assign addr[6036]= 1356798326;
assign addr[6037]= 1386226674;
assign addr[6038]= 1415215352;
assign addr[6039]= 1443755168;
assign addr[6040]= 1471837070;
assign addr[6041]= 1499452149;
assign addr[6042]= 1526591649;
assign addr[6043]= 1553246960;
assign addr[6044]= 1579409630;
assign addr[6045]= 1605071359;
assign addr[6046]= 1630224009;
assign addr[6047]= 1654859602;
assign addr[6048]= 1678970324;
assign addr[6049]= 1702548529;
assign addr[6050]= 1725586737;
assign addr[6051]= 1748077642;
assign addr[6052]= 1770014111;
assign addr[6053]= 1791389186;
assign addr[6054]= 1812196087;
assign addr[6055]= 1832428215;
assign addr[6056]= 1852079154;
assign addr[6057]= 1871142669;
assign addr[6058]= 1889612716;
assign addr[6059]= 1907483436;
assign addr[6060]= 1924749160;
assign addr[6061]= 1941404413;
assign addr[6062]= 1957443913;
assign addr[6063]= 1972862571;
assign addr[6064]= 1987655498;
assign addr[6065]= 2001818002;
assign addr[6066]= 2015345591;
assign addr[6067]= 2028233973;
assign addr[6068]= 2040479063;
assign addr[6069]= 2052076975;
assign addr[6070]= 2063024031;
assign addr[6071]= 2073316760;
assign addr[6072]= 2082951896;
assign addr[6073]= 2091926384;
assign addr[6074]= 2100237377;
assign addr[6075]= 2107882239;
assign addr[6076]= 2114858546;
assign addr[6077]= 2121164085;
assign addr[6078]= 2126796855;
assign addr[6079]= 2131755071;
assign addr[6080]= 2136037160;
assign addr[6081]= 2139641764;
assign addr[6082]= 2142567738;
assign addr[6083]= 2144814157;
assign addr[6084]= 2146380306;
assign addr[6085]= 2147265689;
assign addr[6086]= 2147470025;
assign addr[6087]= 2146993250;
assign addr[6088]= 2145835515;
assign addr[6089]= 2143997187;
assign addr[6090]= 2141478848;
assign addr[6091]= 2138281298;
assign addr[6092]= 2134405552;
assign addr[6093]= 2129852837;
assign addr[6094]= 2124624598;
assign addr[6095]= 2118722494;
assign addr[6096]= 2112148396;
assign addr[6097]= 2104904390;
assign addr[6098]= 2096992772;
assign addr[6099]= 2088416053;
assign addr[6100]= 2079176953;
assign addr[6101]= 2069278401;
assign addr[6102]= 2058723538;
assign addr[6103]= 2047515711;
assign addr[6104]= 2035658475;
assign addr[6105]= 2023155591;
assign addr[6106]= 2010011024;
assign addr[6107]= 1996228943;
assign addr[6108]= 1981813720;
assign addr[6109]= 1966769926;
assign addr[6110]= 1951102334;
assign addr[6111]= 1934815911;
assign addr[6112]= 1917915825;
assign addr[6113]= 1900407434;
assign addr[6114]= 1882296293;
assign addr[6115]= 1863588145;
assign addr[6116]= 1844288924;
assign addr[6117]= 1824404752;
assign addr[6118]= 1803941934;
assign addr[6119]= 1782906961;
assign addr[6120]= 1761306505;
assign addr[6121]= 1739147417;
assign addr[6122]= 1716436725;
assign addr[6123]= 1693181631;
assign addr[6124]= 1669389513;
assign addr[6125]= 1645067915;
assign addr[6126]= 1620224553;
assign addr[6127]= 1594867305;
assign addr[6128]= 1569004214;
assign addr[6129]= 1542643483;
assign addr[6130]= 1515793473;
assign addr[6131]= 1488462700;
assign addr[6132]= 1460659832;
assign addr[6133]= 1432393688;
assign addr[6134]= 1403673233;
assign addr[6135]= 1374507575;
assign addr[6136]= 1344905966;
assign addr[6137]= 1314877795;
assign addr[6138]= 1284432584;
assign addr[6139]= 1253579991;
assign addr[6140]= 1222329801;
assign addr[6141]= 1190691925;
assign addr[6142]= 1158676398;
assign addr[6143]= 1126293375;
assign addr[6144]= 1093553126;
assign addr[6145]= 1060466036;
assign addr[6146]= 1027042599;
assign addr[6147]= 993293415;
assign addr[6148]= 959229189;
assign addr[6149]= 924860725;
assign addr[6150]= 890198924;
assign addr[6151]= 855254778;
assign addr[6152]= 820039373;
assign addr[6153]= 784563876;
assign addr[6154]= 748839539;
assign addr[6155]= 712877694;
assign addr[6156]= 676689746;
assign addr[6157]= 640287172;
assign addr[6158]= 603681519;
assign addr[6159]= 566884397;
assign addr[6160]= 529907477;
assign addr[6161]= 492762486;
assign addr[6162]= 455461206;
assign addr[6163]= 418015468;
assign addr[6164]= 380437148;
assign addr[6165]= 342738165;
assign addr[6166]= 304930476;
assign addr[6167]= 267026072;
assign addr[6168]= 229036977;
assign addr[6169]= 190975237;
assign addr[6170]= 152852926;
assign addr[6171]= 114682135;
assign addr[6172]= 76474970;
assign addr[6173]= 38243550;
assign addr[6174]= 0;
assign addr[6175]= -38243550;
assign addr[6176]= -76474970;
assign addr[6177]= -114682135;
assign addr[6178]= -152852926;
assign addr[6179]= -190975237;
assign addr[6180]= -229036977;
assign addr[6181]= -267026072;
assign addr[6182]= -304930476;
assign addr[6183]= -342738165;
assign addr[6184]= -380437148;
assign addr[6185]= -418015468;
assign addr[6186]= -455461206;
assign addr[6187]= -492762486;
assign addr[6188]= -529907477;
assign addr[6189]= -566884397;
assign addr[6190]= -603681519;
assign addr[6191]= -640287172;
assign addr[6192]= -676689746;
assign addr[6193]= -712877694;
assign addr[6194]= -748839539;
assign addr[6195]= -784563876;
assign addr[6196]= -820039373;
assign addr[6197]= -855254778;
assign addr[6198]= -890198924;
assign addr[6199]= -924860725;
assign addr[6200]= -959229189;
assign addr[6201]= -993293415;
assign addr[6202]= -1027042599;
assign addr[6203]= -1060466036;
assign addr[6204]= -1093553126;
assign addr[6205]= -1126293375;
assign addr[6206]= -1158676398;
assign addr[6207]= -1190691925;
assign addr[6208]= -1222329801;
assign addr[6209]= -1253579991;
assign addr[6210]= -1284432584;
assign addr[6211]= -1314877795;
assign addr[6212]= -1344905966;
assign addr[6213]= -1374507575;
assign addr[6214]= -1403673233;
assign addr[6215]= -1432393688;
assign addr[6216]= -1460659832;
assign addr[6217]= -1488462700;
assign addr[6218]= -1515793473;
assign addr[6219]= -1542643483;
assign addr[6220]= -1569004214;
assign addr[6221]= -1594867305;
assign addr[6222]= -1620224553;
assign addr[6223]= -1645067915;
assign addr[6224]= -1669389513;
assign addr[6225]= -1693181631;
assign addr[6226]= -1716436725;
assign addr[6227]= -1739147417;
assign addr[6228]= -1761306505;
assign addr[6229]= -1782906961;
assign addr[6230]= -1803941934;
assign addr[6231]= -1824404752;
assign addr[6232]= -1844288924;
assign addr[6233]= -1863588145;
assign addr[6234]= -1882296293;
assign addr[6235]= -1900407434;
assign addr[6236]= -1917915825;
assign addr[6237]= -1934815911;
assign addr[6238]= -1951102334;
assign addr[6239]= -1966769926;
assign addr[6240]= -1981813720;
assign addr[6241]= -1996228943;
assign addr[6242]= -2010011024;
assign addr[6243]= -2023155591;
assign addr[6244]= -2035658475;
assign addr[6245]= -2047515711;
assign addr[6246]= -2058723538;
assign addr[6247]= -2069278401;
assign addr[6248]= -2079176953;
assign addr[6249]= -2088416053;
assign addr[6250]= -2096992772;
assign addr[6251]= -2104904390;
assign addr[6252]= -2112148396;
assign addr[6253]= -2118722494;
assign addr[6254]= -2124624598;
assign addr[6255]= -2129852837;
assign addr[6256]= -2134405552;
assign addr[6257]= -2138281298;
assign addr[6258]= -2141478848;
assign addr[6259]= -2143997187;
assign addr[6260]= -2145835515;
assign addr[6261]= -2146993250;
assign addr[6262]= -2147470025;
assign addr[6263]= -2147265689;
assign addr[6264]= -2146380306;
assign addr[6265]= -2144814157;
assign addr[6266]= -2142567738;
assign addr[6267]= -2139641764;
assign addr[6268]= -2136037160;
assign addr[6269]= -2131755071;
assign addr[6270]= -2126796855;
assign addr[6271]= -2121164085;
assign addr[6272]= -2114858546;
assign addr[6273]= -2107882239;
assign addr[6274]= -2100237377;
assign addr[6275]= -2091926384;
assign addr[6276]= -2082951896;
assign addr[6277]= -2073316760;
assign addr[6278]= -2063024031;
assign addr[6279]= -2052076975;
assign addr[6280]= -2040479063;
assign addr[6281]= -2028233973;
assign addr[6282]= -2015345591;
assign addr[6283]= -2001818002;
assign addr[6284]= -1987655498;
assign addr[6285]= -1972862571;
assign addr[6286]= -1957443913;
assign addr[6287]= -1941404413;
assign addr[6288]= -1924749160;
assign addr[6289]= -1907483436;
assign addr[6290]= -1889612716;
assign addr[6291]= -1871142669;
assign addr[6292]= -1852079154;
assign addr[6293]= -1832428215;
assign addr[6294]= -1812196087;
assign addr[6295]= -1791389186;
assign addr[6296]= -1770014111;
assign addr[6297]= -1748077642;
assign addr[6298]= -1725586737;
assign addr[6299]= -1702548529;
assign addr[6300]= -1678970324;
assign addr[6301]= -1654859602;
assign addr[6302]= -1630224009;
assign addr[6303]= -1605071359;
assign addr[6304]= -1579409630;
assign addr[6305]= -1553246960;
assign addr[6306]= -1526591649;
assign addr[6307]= -1499452149;
assign addr[6308]= -1471837070;
assign addr[6309]= -1443755168;
assign addr[6310]= -1415215352;
assign addr[6311]= -1386226674;
assign addr[6312]= -1356798326;
assign addr[6313]= -1326939644;
assign addr[6314]= -1296660098;
assign addr[6315]= -1265969291;
assign addr[6316]= -1234876957;
assign addr[6317]= -1203392958;
assign addr[6318]= -1171527280;
assign addr[6319]= -1139290029;
assign addr[6320]= -1106691431;
assign addr[6321]= -1073741824;
assign addr[6322]= -1040451659;
assign addr[6323]= -1006831495;
assign addr[6324]= -972891995;
assign addr[6325]= -938643924;
assign addr[6326]= -904098143;
assign addr[6327]= -869265610;
assign addr[6328]= -834157373;
assign addr[6329]= -798784567;
assign addr[6330]= -763158411;
assign addr[6331]= -727290205;
assign addr[6332]= -691191324;
assign addr[6333]= -654873219;
assign addr[6334]= -618347408;
assign addr[6335]= -581625477;
assign addr[6336]= -544719071;
assign addr[6337]= -507639898;
assign addr[6338]= -470399716;
assign addr[6339]= -433010339;
assign addr[6340]= -395483624;
assign addr[6341]= -357831473;
assign addr[6342]= -320065829;
assign addr[6343]= -282198671;
assign addr[6344]= -244242007;
assign addr[6345]= -206207878;
assign addr[6346]= -168108346;
assign addr[6347]= -129955495;
assign addr[6348]= -91761426;
assign addr[6349]= -53538253;
assign addr[6350]= -15298099;
assign addr[6351]= 22946906;
assign addr[6352]= 61184634;
assign addr[6353]= 99402956;
assign addr[6354]= 137589750;
assign addr[6355]= 175732905;
assign addr[6356]= 213820322;
assign addr[6357]= 251839923;
assign addr[6358]= 289779648;
assign addr[6359]= 327627463;
assign addr[6360]= 365371365;
assign addr[6361]= 402999383;
assign addr[6362]= 440499581;
assign addr[6363]= 477860067;
assign addr[6364]= 515068990;
assign addr[6365]= 552114549;
assign addr[6366]= 588984994;
assign addr[6367]= 625668632;
assign addr[6368]= 662153826;
assign addr[6369]= 698429006;
assign addr[6370]= 734482665;
assign addr[6371]= 770303369;
assign addr[6372]= 805879757;
assign addr[6373]= 841200544;
assign addr[6374]= 876254528;
assign addr[6375]= 911030591;
assign addr[6376]= 945517704;
assign addr[6377]= 979704927;
assign addr[6378]= 1013581418;
assign addr[6379]= 1047136432;
assign addr[6380]= 1080359326;
assign addr[6381]= 1113239564;
assign addr[6382]= 1145766716;
assign addr[6383]= 1177930466;
assign addr[6384]= 1209720613;
assign addr[6385]= 1241127074;
assign addr[6386]= 1272139887;
assign addr[6387]= 1302749217;
assign addr[6388]= 1332945355;
assign addr[6389]= 1362718723;
assign addr[6390]= 1392059879;
assign addr[6391]= 1420959516;
assign addr[6392]= 1449408469;
assign addr[6393]= 1477397714;
assign addr[6394]= 1504918373;
assign addr[6395]= 1531961719;
assign addr[6396]= 1558519173;
assign addr[6397]= 1584582314;
assign addr[6398]= 1610142873;
assign addr[6399]= 1635192744;
assign addr[6400]= 1659723983;
assign addr[6401]= 1683728808;
assign addr[6402]= 1707199606;
assign addr[6403]= 1730128933;
assign addr[6404]= 1752509516;
assign addr[6405]= 1774334257;
assign addr[6406]= 1795596234;
assign addr[6407]= 1816288703;
assign addr[6408]= 1836405100;
assign addr[6409]= 1855939047;
assign addr[6410]= 1874884346;
assign addr[6411]= 1893234990;
assign addr[6412]= 1910985158;
assign addr[6413]= 1928129220;
assign addr[6414]= 1944661739;
assign addr[6415]= 1960577471;
assign addr[6416]= 1975871368;
assign addr[6417]= 1990538579;
assign addr[6418]= 2004574453;
assign addr[6419]= 2017974537;
assign addr[6420]= 2030734582;
assign addr[6421]= 2042850540;
assign addr[6422]= 2054318569;
assign addr[6423]= 2065135031;
assign addr[6424]= 2075296495;
assign addr[6425]= 2084799740;
assign addr[6426]= 2093641749;
assign addr[6427]= 2101819720;
assign addr[6428]= 2109331059;
assign addr[6429]= 2116173382;
assign addr[6430]= 2122344521;
assign addr[6431]= 2127842516;
assign addr[6432]= 2132665626;
assign addr[6433]= 2136812319;
assign addr[6434]= 2140281282;
assign addr[6435]= 2143071413;
assign addr[6436]= 2145181827;
assign addr[6437]= 2146611856;
assign addr[6438]= 2147361045;
assign addr[6439]= 2147429158;
assign addr[6440]= 2146816171;
assign addr[6441]= 2145522281;
assign addr[6442]= 2143547897;
assign addr[6443]= 2140893646;
assign addr[6444]= 2137560369;
assign addr[6445]= 2133549123;
assign addr[6446]= 2128861181;
assign addr[6447]= 2123498030;
assign addr[6448]= 2117461370;
assign addr[6449]= 2110753117;
assign addr[6450]= 2103375398;
assign addr[6451]= 2095330553;
assign addr[6452]= 2086621133;
assign addr[6453]= 2077249901;
assign addr[6454]= 2067219829;
assign addr[6455]= 2056534099;
assign addr[6456]= 2045196100;
assign addr[6457]= 2033209426;
assign addr[6458]= 2020577882;
assign addr[6459]= 2007305472;
assign addr[6460]= 1993396407;
assign addr[6461]= 1978855097;
assign addr[6462]= 1963686155;
assign addr[6463]= 1947894393;
assign addr[6464]= 1931484818;
assign addr[6465]= 1914462636;
assign addr[6466]= 1896833245;
assign addr[6467]= 1878602237;
assign addr[6468]= 1859775393;
assign addr[6469]= 1840358687;
assign addr[6470]= 1820358275;
assign addr[6471]= 1799780501;
assign addr[6472]= 1778631892;
assign addr[6473]= 1756919156;
assign addr[6474]= 1734649179;
assign addr[6475]= 1711829025;
assign addr[6476]= 1688465931;
assign addr[6477]= 1664567307;
assign addr[6478]= 1640140734;
assign addr[6479]= 1615193959;
assign addr[6480]= 1589734894;
assign addr[6481]= 1563771613;
assign addr[6482]= 1537312353;
assign addr[6483]= 1510365504;
assign addr[6484]= 1482939614;
assign addr[6485]= 1455043381;
assign addr[6486]= 1426685652;
assign addr[6487]= 1397875423;
assign addr[6488]= 1368621831;
assign addr[6489]= 1338934154;
assign addr[6490]= 1308821808;
assign addr[6491]= 1278294345;
assign addr[6492]= 1247361445;
assign addr[6493]= 1216032921;
assign addr[6494]= 1184318708;
assign addr[6495]= 1152228866;
assign addr[6496]= 1119773573;
assign addr[6497]= 1086963121;
assign addr[6498]= 1053807919;
assign addr[6499]= 1020318481;
assign addr[6500]= 986505429;
assign addr[6501]= 952379488;
assign addr[6502]= 917951481;
assign addr[6503]= 883232329;
assign addr[6504]= 848233042;
assign addr[6505]= 812964722;
assign addr[6506]= 777438554;
assign addr[6507]= 741665807;
assign addr[6508]= 705657826;
assign addr[6509]= 669426032;
assign addr[6510]= 632981917;
assign addr[6511]= 596337040;
assign addr[6512]= 559503022;
assign addr[6513]= 522491548;
assign addr[6514]= 485314355;
assign addr[6515]= 447983235;
assign addr[6516]= 410510029;
assign addr[6517]= 372906622;
assign addr[6518]= 335184940;
assign addr[6519]= 297356948;
assign addr[6520]= 259434643;
assign addr[6521]= 221430054;
assign addr[6522]= 183355234;
assign addr[6523]= 145222259;
assign addr[6524]= 107043224;
assign addr[6525]= 68830239;
assign addr[6526]= 30595422;
assign addr[6527]= -7649098;
assign addr[6528]= -45891193;
assign addr[6529]= -84118732;
assign addr[6530]= -122319591;
assign addr[6531]= -160481654;
assign addr[6532]= -198592817;
assign addr[6533]= -236640993;
assign addr[6534]= -274614114;
assign addr[6535]= -312500135;
assign addr[6536]= -350287041;
assign addr[6537]= -387962847;
assign addr[6538]= -425515602;
assign addr[6539]= -462933398;
assign addr[6540]= -500204365;
assign addr[6541]= -537316682;
assign addr[6542]= -574258580;
assign addr[6543]= -611018340;
assign addr[6544]= -647584304;
assign addr[6545]= -683944874;
assign addr[6546]= -720088517;
assign addr[6547]= -756003771;
assign addr[6548]= -791679244;
assign addr[6549]= -827103620;
assign addr[6550]= -862265664;
assign addr[6551]= -897154224;
assign addr[6552]= -931758235;
assign addr[6553]= -966066720;
assign addr[6554]= -1000068799;
assign addr[6555]= -1033753687;
assign addr[6556]= -1067110699;
assign addr[6557]= -1100129257;
assign addr[6558]= -1132798888;
assign addr[6559]= -1165109230;
assign addr[6560]= -1197050035;
assign addr[6561]= -1228611172;
assign addr[6562]= -1259782632;
assign addr[6563]= -1290554528;
assign addr[6564]= -1320917099;
assign addr[6565]= -1350860716;
assign addr[6566]= -1380375881;
assign addr[6567]= -1409453233;
assign addr[6568]= -1438083551;
assign addr[6569]= -1466257752;
assign addr[6570]= -1493966902;
assign addr[6571]= -1521202211;
assign addr[6572]= -1547955041;
assign addr[6573]= -1574216908;
assign addr[6574]= -1599979481;
assign addr[6575]= -1625234591;
assign addr[6576]= -1649974225;
assign addr[6577]= -1674190539;
assign addr[6578]= -1697875851;
assign addr[6579]= -1721022648;
assign addr[6580]= -1743623590;
assign addr[6581]= -1765671509;
assign addr[6582]= -1787159411;
assign addr[6583]= -1808080480;
assign addr[6584]= -1828428082;
assign addr[6585]= -1848195763;
assign addr[6586]= -1867377253;
assign addr[6587]= -1885966468;
assign addr[6588]= -1903957513;
assign addr[6589]= -1921344681;
assign addr[6590]= -1938122457;
assign addr[6591]= -1954285520;
assign addr[6592]= -1969828744;
assign addr[6593]= -1984747199;
assign addr[6594]= -1999036154;
assign addr[6595]= -2012691075;
assign addr[6596]= -2025707632;
assign addr[6597]= -2038081698;
assign addr[6598]= -2049809346;
assign addr[6599]= -2060886858;
assign addr[6600]= -2071310720;
assign addr[6601]= -2081077626;
assign addr[6602]= -2090184478;
assign addr[6603]= -2098628387;
assign addr[6604]= -2106406677;
assign addr[6605]= -2113516878;
assign addr[6606]= -2119956737;
assign addr[6607]= -2125724211;
assign addr[6608]= -2130817471;
assign addr[6609]= -2135234901;
assign addr[6610]= -2138975100;
assign addr[6611]= -2142036881;
assign addr[6612]= -2144419275;
assign addr[6613]= -2146121524;
assign addr[6614]= -2147143090;
assign addr[6615]= -2147483648;
assign addr[6616]= -2147143090;
assign addr[6617]= -2146121524;
assign addr[6618]= -2144419275;
assign addr[6619]= -2142036881;
assign addr[6620]= -2138975100;
assign addr[6621]= -2135234901;
assign addr[6622]= -2130817471;
assign addr[6623]= -2125724211;
assign addr[6624]= -2119956737;
assign addr[6625]= -2113516878;
assign addr[6626]= -2106406677;
assign addr[6627]= -2098628387;
assign addr[6628]= -2090184478;
assign addr[6629]= -2081077626;
assign addr[6630]= -2071310720;
assign addr[6631]= -2060886858;
assign addr[6632]= -2049809346;
assign addr[6633]= -2038081698;
assign addr[6634]= -2025707632;
assign addr[6635]= -2012691075;
assign addr[6636]= -1999036154;
assign addr[6637]= -1984747199;
assign addr[6638]= -1969828744;
assign addr[6639]= -1954285520;
assign addr[6640]= -1938122457;
assign addr[6641]= -1921344681;
assign addr[6642]= -1903957513;
assign addr[6643]= -1885966468;
assign addr[6644]= -1867377253;
assign addr[6645]= -1848195763;
assign addr[6646]= -1828428082;
assign addr[6647]= -1808080480;
assign addr[6648]= -1787159411;
assign addr[6649]= -1765671509;
assign addr[6650]= -1743623590;
assign addr[6651]= -1721022648;
assign addr[6652]= -1697875851;
assign addr[6653]= -1674190539;
assign addr[6654]= -1649974225;
assign addr[6655]= -1625234591;
assign addr[6656]= -1599979481;
assign addr[6657]= -1574216908;
assign addr[6658]= -1547955041;
assign addr[6659]= -1521202211;
assign addr[6660]= -1493966902;
assign addr[6661]= -1466257752;
assign addr[6662]= -1438083551;
assign addr[6663]= -1409453233;
assign addr[6664]= -1380375881;
assign addr[6665]= -1350860716;
assign addr[6666]= -1320917099;
assign addr[6667]= -1290554528;
assign addr[6668]= -1259782632;
assign addr[6669]= -1228611172;
assign addr[6670]= -1197050035;
assign addr[6671]= -1165109230;
assign addr[6672]= -1132798888;
assign addr[6673]= -1100129257;
assign addr[6674]= -1067110699;
assign addr[6675]= -1033753687;
assign addr[6676]= -1000068799;
assign addr[6677]= -966066720;
assign addr[6678]= -931758235;
assign addr[6679]= -897154224;
assign addr[6680]= -862265664;
assign addr[6681]= -827103620;
assign addr[6682]= -791679244;
assign addr[6683]= -756003771;
assign addr[6684]= -720088517;
assign addr[6685]= -683944874;
assign addr[6686]= -647584304;
assign addr[6687]= -611018340;
assign addr[6688]= -574258580;
assign addr[6689]= -537316682;
assign addr[6690]= -500204365;
assign addr[6691]= -462933398;
assign addr[6692]= -425515602;
assign addr[6693]= -387962847;
assign addr[6694]= -350287041;
assign addr[6695]= -312500135;
assign addr[6696]= -274614114;
assign addr[6697]= -236640993;
assign addr[6698]= -198592817;
assign addr[6699]= -160481654;
assign addr[6700]= -122319591;
assign addr[6701]= -84118732;
assign addr[6702]= -45891193;
assign addr[6703]= -7649098;
assign addr[6704]= 30595422;
assign addr[6705]= 68830239;
assign addr[6706]= 107043224;
assign addr[6707]= 145222259;
assign addr[6708]= 183355234;
assign addr[6709]= 221430054;
assign addr[6710]= 259434643;
assign addr[6711]= 297356948;
assign addr[6712]= 335184940;
assign addr[6713]= 372906622;
assign addr[6714]= 410510029;
assign addr[6715]= 447983235;
assign addr[6716]= 485314355;
assign addr[6717]= 522491548;
assign addr[6718]= 559503022;
assign addr[6719]= 596337040;
assign addr[6720]= 632981917;
assign addr[6721]= 669426032;
assign addr[6722]= 705657826;
assign addr[6723]= 741665807;
assign addr[6724]= 777438554;
assign addr[6725]= 812964722;
assign addr[6726]= 848233042;
assign addr[6727]= 883232329;
assign addr[6728]= 917951481;
assign addr[6729]= 952379488;
assign addr[6730]= 986505429;
assign addr[6731]= 1020318481;
assign addr[6732]= 1053807919;
assign addr[6733]= 1086963121;
assign addr[6734]= 1119773573;
assign addr[6735]= 1152228866;
assign addr[6736]= 1184318708;
assign addr[6737]= 1216032921;
assign addr[6738]= 1247361445;
assign addr[6739]= 1278294345;
assign addr[6740]= 1308821808;
assign addr[6741]= 1338934154;
assign addr[6742]= 1368621831;
assign addr[6743]= 1397875423;
assign addr[6744]= 1426685652;
assign addr[6745]= 1455043381;
assign addr[6746]= 1482939614;
assign addr[6747]= 1510365504;
assign addr[6748]= 1537312353;
assign addr[6749]= 1563771613;
assign addr[6750]= 1589734894;
assign addr[6751]= 1615193959;
assign addr[6752]= 1640140734;
assign addr[6753]= 1664567307;
assign addr[6754]= 1688465931;
assign addr[6755]= 1711829025;
assign addr[6756]= 1734649179;
assign addr[6757]= 1756919156;
assign addr[6758]= 1778631892;
assign addr[6759]= 1799780501;
assign addr[6760]= 1820358275;
assign addr[6761]= 1840358687;
assign addr[6762]= 1859775393;
assign addr[6763]= 1878602237;
assign addr[6764]= 1896833245;
assign addr[6765]= 1914462636;
assign addr[6766]= 1931484818;
assign addr[6767]= 1947894393;
assign addr[6768]= 1963686155;
assign addr[6769]= 1978855097;
assign addr[6770]= 1993396407;
assign addr[6771]= 2007305472;
assign addr[6772]= 2020577882;
assign addr[6773]= 2033209426;
assign addr[6774]= 2045196100;
assign addr[6775]= 2056534099;
assign addr[6776]= 2067219829;
assign addr[6777]= 2077249901;
assign addr[6778]= 2086621133;
assign addr[6779]= 2095330553;
assign addr[6780]= 2103375398;
assign addr[6781]= 2110753117;
assign addr[6782]= 2117461370;
assign addr[6783]= 2123498030;
assign addr[6784]= 2128861181;
assign addr[6785]= 2133549123;
assign addr[6786]= 2137560369;
assign addr[6787]= 2140893646;
assign addr[6788]= 2143547897;
assign addr[6789]= 2145522281;
assign addr[6790]= 2146816171;
assign addr[6791]= 2147429158;
assign addr[6792]= 2147361045;
assign addr[6793]= 2146611856;
assign addr[6794]= 2145181827;
assign addr[6795]= 2143071413;
assign addr[6796]= 2140281282;
assign addr[6797]= 2136812319;
assign addr[6798]= 2132665626;
assign addr[6799]= 2127842516;
assign addr[6800]= 2122344521;
assign addr[6801]= 2116173382;
assign addr[6802]= 2109331059;
assign addr[6803]= 2101819720;
assign addr[6804]= 2093641749;
assign addr[6805]= 2084799740;
assign addr[6806]= 2075296495;
assign addr[6807]= 2065135031;
assign addr[6808]= 2054318569;
assign addr[6809]= 2042850540;
assign addr[6810]= 2030734582;
assign addr[6811]= 2017974537;
assign addr[6812]= 2004574453;
assign addr[6813]= 1990538579;
assign addr[6814]= 1975871368;
assign addr[6815]= 1960577471;
assign addr[6816]= 1944661739;
assign addr[6817]= 1928129220;
assign addr[6818]= 1910985158;
assign addr[6819]= 1893234990;
assign addr[6820]= 1874884346;
assign addr[6821]= 1855939047;
assign addr[6822]= 1836405100;
assign addr[6823]= 1816288703;
assign addr[6824]= 1795596234;
assign addr[6825]= 1774334257;
assign addr[6826]= 1752509516;
assign addr[6827]= 1730128933;
assign addr[6828]= 1707199606;
assign addr[6829]= 1683728808;
assign addr[6830]= 1659723983;
assign addr[6831]= 1635192744;
assign addr[6832]= 1610142873;
assign addr[6833]= 1584582314;
assign addr[6834]= 1558519173;
assign addr[6835]= 1531961719;
assign addr[6836]= 1504918373;
assign addr[6837]= 1477397714;
assign addr[6838]= 1449408469;
assign addr[6839]= 1420959516;
assign addr[6840]= 1392059879;
assign addr[6841]= 1362718723;
assign addr[6842]= 1332945355;
assign addr[6843]= 1302749217;
assign addr[6844]= 1272139887;
assign addr[6845]= 1241127074;
assign addr[6846]= 1209720613;
assign addr[6847]= 1177930466;
assign addr[6848]= 1145766716;
assign addr[6849]= 1113239564;
assign addr[6850]= 1080359326;
assign addr[6851]= 1047136432;
assign addr[6852]= 1013581418;
assign addr[6853]= 979704927;
assign addr[6854]= 945517704;
assign addr[6855]= 911030591;
assign addr[6856]= 876254528;
assign addr[6857]= 841200544;
assign addr[6858]= 805879757;
assign addr[6859]= 770303369;
assign addr[6860]= 734482665;
assign addr[6861]= 698429006;
assign addr[6862]= 662153826;
assign addr[6863]= 625668632;
assign addr[6864]= 588984994;
assign addr[6865]= 552114549;
assign addr[6866]= 515068990;
assign addr[6867]= 477860067;
assign addr[6868]= 440499581;
assign addr[6869]= 402999383;
assign addr[6870]= 365371365;
assign addr[6871]= 327627463;
assign addr[6872]= 289779648;
assign addr[6873]= 251839923;
assign addr[6874]= 213820322;
assign addr[6875]= 175732905;
assign addr[6876]= 137589750;
assign addr[6877]= 99402956;
assign addr[6878]= 61184634;
assign addr[6879]= 22946906;
assign addr[6880]= -15298099;
assign addr[6881]= -53538253;
assign addr[6882]= -91761426;
assign addr[6883]= -129955495;
assign addr[6884]= -168108346;
assign addr[6885]= -206207878;
assign addr[6886]= -244242007;
assign addr[6887]= -282198671;
assign addr[6888]= -320065829;
assign addr[6889]= -357831473;
assign addr[6890]= -395483624;
assign addr[6891]= -433010339;
assign addr[6892]= -470399716;
assign addr[6893]= -507639898;
assign addr[6894]= -544719071;
assign addr[6895]= -581625477;
assign addr[6896]= -618347408;
assign addr[6897]= -654873219;
assign addr[6898]= -691191324;
assign addr[6899]= -727290205;
assign addr[6900]= -763158411;
assign addr[6901]= -798784567;
assign addr[6902]= -834157373;
assign addr[6903]= -869265610;
assign addr[6904]= -904098143;
assign addr[6905]= -938643924;
assign addr[6906]= -972891995;
assign addr[6907]= -1006831495;
assign addr[6908]= -1040451659;
assign addr[6909]= -1073741824;
assign addr[6910]= -1106691431;
assign addr[6911]= -1139290029;
assign addr[6912]= -1171527280;
assign addr[6913]= -1203392958;
assign addr[6914]= -1234876957;
assign addr[6915]= -1265969291;
assign addr[6916]= -1296660098;
assign addr[6917]= -1326939644;
assign addr[6918]= -1356798326;
assign addr[6919]= -1386226674;
assign addr[6920]= -1415215352;
assign addr[6921]= -1443755168;
assign addr[6922]= -1471837070;
assign addr[6923]= -1499452149;
assign addr[6924]= -1526591649;
assign addr[6925]= -1553246960;
assign addr[6926]= -1579409630;
assign addr[6927]= -1605071359;
assign addr[6928]= -1630224009;
assign addr[6929]= -1654859602;
assign addr[6930]= -1678970324;
assign addr[6931]= -1702548529;
assign addr[6932]= -1725586737;
assign addr[6933]= -1748077642;
assign addr[6934]= -1770014111;
assign addr[6935]= -1791389186;
assign addr[6936]= -1812196087;
assign addr[6937]= -1832428215;
assign addr[6938]= -1852079154;
assign addr[6939]= -1871142669;
assign addr[6940]= -1889612716;
assign addr[6941]= -1907483436;
assign addr[6942]= -1924749160;
assign addr[6943]= -1941404413;
assign addr[6944]= -1957443913;
assign addr[6945]= -1972862571;
assign addr[6946]= -1987655498;
assign addr[6947]= -2001818002;
assign addr[6948]= -2015345591;
assign addr[6949]= -2028233973;
assign addr[6950]= -2040479063;
assign addr[6951]= -2052076975;
assign addr[6952]= -2063024031;
assign addr[6953]= -2073316760;
assign addr[6954]= -2082951896;
assign addr[6955]= -2091926384;
assign addr[6956]= -2100237377;
assign addr[6957]= -2107882239;
assign addr[6958]= -2114858546;
assign addr[6959]= -2121164085;
assign addr[6960]= -2126796855;
assign addr[6961]= -2131755071;
assign addr[6962]= -2136037160;
assign addr[6963]= -2139641764;
assign addr[6964]= -2142567738;
assign addr[6965]= -2144814157;
assign addr[6966]= -2146380306;
assign addr[6967]= -2147265689;
assign addr[6968]= -2147470025;
assign addr[6969]= -2146993250;
assign addr[6970]= -2145835515;
assign addr[6971]= -2143997187;
assign addr[6972]= -2141478848;
assign addr[6973]= -2138281298;
assign addr[6974]= -2134405552;
assign addr[6975]= -2129852837;
assign addr[6976]= -2124624598;
assign addr[6977]= -2118722494;
assign addr[6978]= -2112148396;
assign addr[6979]= -2104904390;
assign addr[6980]= -2096992772;
assign addr[6981]= -2088416053;
assign addr[6982]= -2079176953;
assign addr[6983]= -2069278401;
assign addr[6984]= -2058723538;
assign addr[6985]= -2047515711;
assign addr[6986]= -2035658475;
assign addr[6987]= -2023155591;
assign addr[6988]= -2010011024;
assign addr[6989]= -1996228943;
assign addr[6990]= -1981813720;
assign addr[6991]= -1966769926;
assign addr[6992]= -1951102334;
assign addr[6993]= -1934815911;
assign addr[6994]= -1917915825;
assign addr[6995]= -1900407434;
assign addr[6996]= -1882296293;
assign addr[6997]= -1863588145;
assign addr[6998]= -1844288924;
assign addr[6999]= -1824404752;
assign addr[7000]= -1803941934;
assign addr[7001]= -1782906961;
assign addr[7002]= -1761306505;
assign addr[7003]= -1739147417;
assign addr[7004]= -1716436725;
assign addr[7005]= -1693181631;
assign addr[7006]= -1669389513;
assign addr[7007]= -1645067915;
assign addr[7008]= -1620224553;
assign addr[7009]= -1594867305;
assign addr[7010]= -1569004214;
assign addr[7011]= -1542643483;
assign addr[7012]= -1515793473;
assign addr[7013]= -1488462700;
assign addr[7014]= -1460659832;
assign addr[7015]= -1432393688;
assign addr[7016]= -1403673233;
assign addr[7017]= -1374507575;
assign addr[7018]= -1344905966;
assign addr[7019]= -1314877795;
assign addr[7020]= -1284432584;
assign addr[7021]= -1253579991;
assign addr[7022]= -1222329801;
assign addr[7023]= -1190691925;
assign addr[7024]= -1158676398;
assign addr[7025]= -1126293375;
assign addr[7026]= -1093553126;
assign addr[7027]= -1060466036;
assign addr[7028]= -1027042599;
assign addr[7029]= -993293415;
assign addr[7030]= -959229189;
assign addr[7031]= -924860725;
assign addr[7032]= -890198924;
assign addr[7033]= -855254778;
assign addr[7034]= -820039373;
assign addr[7035]= -784563876;
assign addr[7036]= -748839539;
assign addr[7037]= -712877694;
assign addr[7038]= -676689746;
assign addr[7039]= -640287172;
assign addr[7040]= -603681519;
assign addr[7041]= -566884397;
assign addr[7042]= -529907477;
assign addr[7043]= -492762486;
assign addr[7044]= -455461206;
assign addr[7045]= -418015468;
assign addr[7046]= -380437148;
assign addr[7047]= -342738165;
assign addr[7048]= -304930476;
assign addr[7049]= -267026072;
assign addr[7050]= -229036977;
assign addr[7051]= -190975237;
assign addr[7052]= -152852926;
assign addr[7053]= -114682135;
assign addr[7054]= -76474970;
assign addr[7055]= -38243550;
assign addr[7056]= 0;
assign addr[7057]= 38243550;
assign addr[7058]= 76474970;
assign addr[7059]= 114682135;
assign addr[7060]= 152852926;
assign addr[7061]= 190975237;
assign addr[7062]= 229036977;
assign addr[7063]= 267026072;
assign addr[7064]= 304930476;
assign addr[7065]= 342738165;
assign addr[7066]= 380437148;
assign addr[7067]= 418015468;
assign addr[7068]= 455461206;
assign addr[7069]= 492762486;
assign addr[7070]= 529907477;
assign addr[7071]= 566884397;
assign addr[7072]= 603681519;
assign addr[7073]= 640287172;
assign addr[7074]= 676689746;
assign addr[7075]= 712877694;
assign addr[7076]= 748839539;
assign addr[7077]= 784563876;
assign addr[7078]= 820039373;
assign addr[7079]= 855254778;
assign addr[7080]= 890198924;
assign addr[7081]= 924860725;
assign addr[7082]= 959229189;
assign addr[7083]= 993293415;
assign addr[7084]= 1027042599;
assign addr[7085]= 1060466036;
assign addr[7086]= 1093553126;
assign addr[7087]= 1126293375;
assign addr[7088]= 1158676398;
assign addr[7089]= 1190691925;
assign addr[7090]= 1222329801;
assign addr[7091]= 1253579991;
assign addr[7092]= 1284432584;
assign addr[7093]= 1314877795;
assign addr[7094]= 1344905966;
assign addr[7095]= 1374507575;
assign addr[7096]= 1403673233;
assign addr[7097]= 1432393688;
assign addr[7098]= 1460659832;
assign addr[7099]= 1488462700;
assign addr[7100]= 1515793473;
assign addr[7101]= 1542643483;
assign addr[7102]= 1569004214;
assign addr[7103]= 1594867305;
assign addr[7104]= 1620224553;
assign addr[7105]= 1645067915;
assign addr[7106]= 1669389513;
assign addr[7107]= 1693181631;
assign addr[7108]= 1716436725;
assign addr[7109]= 1739147417;
assign addr[7110]= 1761306505;
assign addr[7111]= 1782906961;
assign addr[7112]= 1803941934;
assign addr[7113]= 1824404752;
assign addr[7114]= 1844288924;
assign addr[7115]= 1863588145;
assign addr[7116]= 1882296293;
assign addr[7117]= 1900407434;
assign addr[7118]= 1917915825;
assign addr[7119]= 1934815911;
assign addr[7120]= 1951102334;
assign addr[7121]= 1966769926;
assign addr[7122]= 1981813720;
assign addr[7123]= 1996228943;
assign addr[7124]= 2010011024;
assign addr[7125]= 2023155591;
assign addr[7126]= 2035658475;
assign addr[7127]= 2047515711;
assign addr[7128]= 2058723538;
assign addr[7129]= 2069278401;
assign addr[7130]= 2079176953;
assign addr[7131]= 2088416053;
assign addr[7132]= 2096992772;
assign addr[7133]= 2104904390;
assign addr[7134]= 2112148396;
assign addr[7135]= 2118722494;
assign addr[7136]= 2124624598;
assign addr[7137]= 2129852837;
assign addr[7138]= 2134405552;
assign addr[7139]= 2138281298;
assign addr[7140]= 2141478848;
assign addr[7141]= 2143997187;
assign addr[7142]= 2145835515;
assign addr[7143]= 2146993250;
assign addr[7144]= 2147470025;
assign addr[7145]= 2147265689;
assign addr[7146]= 2146380306;
assign addr[7147]= 2144814157;
assign addr[7148]= 2142567738;
assign addr[7149]= 2139641764;
assign addr[7150]= 2136037160;
assign addr[7151]= 2131755071;
assign addr[7152]= 2126796855;
assign addr[7153]= 2121164085;
assign addr[7154]= 2114858546;
assign addr[7155]= 2107882239;
assign addr[7156]= 2100237377;
assign addr[7157]= 2091926384;
assign addr[7158]= 2082951896;
assign addr[7159]= 2073316760;
assign addr[7160]= 2063024031;
assign addr[7161]= 2052076975;
assign addr[7162]= 2040479063;
assign addr[7163]= 2028233973;
assign addr[7164]= 2015345591;
assign addr[7165]= 2001818002;
assign addr[7166]= 1987655498;
assign addr[7167]= 1972862571;
assign addr[7168]= 1957443913;
assign addr[7169]= 1941404413;
assign addr[7170]= 1924749160;
assign addr[7171]= 1907483436;
assign addr[7172]= 1889612716;
assign addr[7173]= 1871142669;
assign addr[7174]= 1852079154;
assign addr[7175]= 1832428215;
assign addr[7176]= 1812196087;
assign addr[7177]= 1791389186;
assign addr[7178]= 1770014111;
assign addr[7179]= 1748077642;
assign addr[7180]= 1725586737;
assign addr[7181]= 1702548529;
assign addr[7182]= 1678970324;
assign addr[7183]= 1654859602;
assign addr[7184]= 1630224009;
assign addr[7185]= 1605071359;
assign addr[7186]= 1579409630;
assign addr[7187]= 1553246960;
assign addr[7188]= 1526591649;
assign addr[7189]= 1499452149;
assign addr[7190]= 1471837070;
assign addr[7191]= 1443755168;
assign addr[7192]= 1415215352;
assign addr[7193]= 1386226674;
assign addr[7194]= 1356798326;
assign addr[7195]= 1326939644;
assign addr[7196]= 1296660098;
assign addr[7197]= 1265969291;
assign addr[7198]= 1234876957;
assign addr[7199]= 1203392958;
assign addr[7200]= 1171527280;
assign addr[7201]= 1139290029;
assign addr[7202]= 1106691431;
assign addr[7203]= 1073741824;
assign addr[7204]= 1040451659;
assign addr[7205]= 1006831495;
assign addr[7206]= 972891995;
assign addr[7207]= 938643924;
assign addr[7208]= 904098143;
assign addr[7209]= 869265610;
assign addr[7210]= 834157373;
assign addr[7211]= 798784567;
assign addr[7212]= 763158411;
assign addr[7213]= 727290205;
assign addr[7214]= 691191324;
assign addr[7215]= 654873219;
assign addr[7216]= 618347408;
assign addr[7217]= 581625477;
assign addr[7218]= 544719071;
assign addr[7219]= 507639898;
assign addr[7220]= 470399716;
assign addr[7221]= 433010339;
assign addr[7222]= 395483624;
assign addr[7223]= 357831473;
assign addr[7224]= 320065829;
assign addr[7225]= 282198671;
assign addr[7226]= 244242007;
assign addr[7227]= 206207878;
assign addr[7228]= 168108346;
assign addr[7229]= 129955495;
assign addr[7230]= 91761426;
assign addr[7231]= 53538253;
assign addr[7232]= 15298099;
assign addr[7233]= -22946906;
assign addr[7234]= -61184634;
assign addr[7235]= -99402956;
assign addr[7236]= -137589750;
assign addr[7237]= -175732905;
assign addr[7238]= -213820322;
assign addr[7239]= -251839923;
assign addr[7240]= -289779648;
assign addr[7241]= -327627463;
assign addr[7242]= -365371365;
assign addr[7243]= -402999383;
assign addr[7244]= -440499581;
assign addr[7245]= -477860067;
assign addr[7246]= -515068990;
assign addr[7247]= -552114549;
assign addr[7248]= -588984994;
assign addr[7249]= -625668632;
assign addr[7250]= -662153826;
assign addr[7251]= -698429006;
assign addr[7252]= -734482665;
assign addr[7253]= -770303369;
assign addr[7254]= -805879757;
assign addr[7255]= -841200544;
assign addr[7256]= -876254528;
assign addr[7257]= -911030591;
assign addr[7258]= -945517704;
assign addr[7259]= -979704927;
assign addr[7260]= -1013581418;
assign addr[7261]= -1047136432;
assign addr[7262]= -1080359326;
assign addr[7263]= -1113239564;
assign addr[7264]= -1145766716;
assign addr[7265]= -1177930466;
assign addr[7266]= -1209720613;
assign addr[7267]= -1241127074;
assign addr[7268]= -1272139887;
assign addr[7269]= -1302749217;
assign addr[7270]= -1332945355;
assign addr[7271]= -1362718723;
assign addr[7272]= -1392059879;
assign addr[7273]= -1420959516;
assign addr[7274]= -1449408469;
assign addr[7275]= -1477397714;
assign addr[7276]= -1504918373;
assign addr[7277]= -1531961719;
assign addr[7278]= -1558519173;
assign addr[7279]= -1584582314;
assign addr[7280]= -1610142873;
assign addr[7281]= -1635192744;
assign addr[7282]= -1659723983;
assign addr[7283]= -1683728808;
assign addr[7284]= -1707199606;
assign addr[7285]= -1730128933;
assign addr[7286]= -1752509516;
assign addr[7287]= -1774334257;
assign addr[7288]= -1795596234;
assign addr[7289]= -1816288703;
assign addr[7290]= -1836405100;
assign addr[7291]= -1855939047;
assign addr[7292]= -1874884346;
assign addr[7293]= -1893234990;
assign addr[7294]= -1910985158;
assign addr[7295]= -1928129220;
assign addr[7296]= -1944661739;
assign addr[7297]= -1960577471;
assign addr[7298]= -1975871368;
assign addr[7299]= -1990538579;
assign addr[7300]= -2004574453;
assign addr[7301]= -2017974537;
assign addr[7302]= -2030734582;
assign addr[7303]= -2042850540;
assign addr[7304]= -2054318569;
assign addr[7305]= -2065135031;
assign addr[7306]= -2075296495;
assign addr[7307]= -2084799740;
assign addr[7308]= -2093641749;
assign addr[7309]= -2101819720;
assign addr[7310]= -2109331059;
assign addr[7311]= -2116173382;
assign addr[7312]= -2122344521;
assign addr[7313]= -2127842516;
assign addr[7314]= -2132665626;
assign addr[7315]= -2136812319;
assign addr[7316]= -2140281282;
assign addr[7317]= -2143071413;
assign addr[7318]= -2145181827;
assign addr[7319]= -2146611856;
assign addr[7320]= -2147361045;
assign addr[7321]= -2147429158;
assign addr[7322]= -2146816171;
assign addr[7323]= -2145522281;
assign addr[7324]= -2143547897;
assign addr[7325]= -2140893646;
assign addr[7326]= -2137560369;
assign addr[7327]= -2133549123;
assign addr[7328]= -2128861181;
assign addr[7329]= -2123498030;
assign addr[7330]= -2117461370;
assign addr[7331]= -2110753117;
assign addr[7332]= -2103375398;
assign addr[7333]= -2095330553;
assign addr[7334]= -2086621133;
assign addr[7335]= -2077249901;
assign addr[7336]= -2067219829;
assign addr[7337]= -2056534099;
assign addr[7338]= -2045196100;
assign addr[7339]= -2033209426;
assign addr[7340]= -2020577882;
assign addr[7341]= -2007305472;
assign addr[7342]= -1993396407;
assign addr[7343]= -1978855097;
assign addr[7344]= -1963686155;
assign addr[7345]= -1947894393;
assign addr[7346]= -1931484818;
assign addr[7347]= -1914462636;
assign addr[7348]= -1896833245;
assign addr[7349]= -1878602237;
assign addr[7350]= -1859775393;
assign addr[7351]= -1840358687;
assign addr[7352]= -1820358275;
assign addr[7353]= -1799780501;
assign addr[7354]= -1778631892;
assign addr[7355]= -1756919156;
assign addr[7356]= -1734649179;
assign addr[7357]= -1711829025;
assign addr[7358]= -1688465931;
assign addr[7359]= -1664567307;
assign addr[7360]= -1640140734;
assign addr[7361]= -1615193959;
assign addr[7362]= -1589734894;
assign addr[7363]= -1563771613;
assign addr[7364]= -1537312353;
assign addr[7365]= -1510365504;
assign addr[7366]= -1482939614;
assign addr[7367]= -1455043381;
assign addr[7368]= -1426685652;
assign addr[7369]= -1397875423;
assign addr[7370]= -1368621831;
assign addr[7371]= -1338934154;
assign addr[7372]= -1308821808;
assign addr[7373]= -1278294345;
assign addr[7374]= -1247361445;
assign addr[7375]= -1216032921;
assign addr[7376]= -1184318708;
assign addr[7377]= -1152228866;
assign addr[7378]= -1119773573;
assign addr[7379]= -1086963121;
assign addr[7380]= -1053807919;
assign addr[7381]= -1020318481;
assign addr[7382]= -986505429;
assign addr[7383]= -952379488;
assign addr[7384]= -917951481;
assign addr[7385]= -883232329;
assign addr[7386]= -848233042;
assign addr[7387]= -812964722;
assign addr[7388]= -777438554;
assign addr[7389]= -741665807;
assign addr[7390]= -705657826;
assign addr[7391]= -669426032;
assign addr[7392]= -632981917;
assign addr[7393]= -596337040;
assign addr[7394]= -559503022;
assign addr[7395]= -522491548;
assign addr[7396]= -485314355;
assign addr[7397]= -447983235;
assign addr[7398]= -410510029;
assign addr[7399]= -372906622;
assign addr[7400]= -335184940;
assign addr[7401]= -297356948;
assign addr[7402]= -259434643;
assign addr[7403]= -221430054;
assign addr[7404]= -183355234;
assign addr[7405]= -145222259;
assign addr[7406]= -107043224;
assign addr[7407]= -68830239;
assign addr[7408]= -30595422;
assign addr[7409]= 7649098;
assign addr[7410]= 45891193;
assign addr[7411]= 84118732;
assign addr[7412]= 122319591;
assign addr[7413]= 160481654;
assign addr[7414]= 198592817;
assign addr[7415]= 236640993;
assign addr[7416]= 274614114;
assign addr[7417]= 312500135;
assign addr[7418]= 350287041;
assign addr[7419]= 387962847;
assign addr[7420]= 425515602;
assign addr[7421]= 462933398;
assign addr[7422]= 500204365;
assign addr[7423]= 537316682;
assign addr[7424]= 574258580;
assign addr[7425]= 611018340;
assign addr[7426]= 647584304;
assign addr[7427]= 683944874;
assign addr[7428]= 720088517;
assign addr[7429]= 756003771;
assign addr[7430]= 791679244;
assign addr[7431]= 827103620;
assign addr[7432]= 862265664;
assign addr[7433]= 897154224;
assign addr[7434]= 931758235;
assign addr[7435]= 966066720;
assign addr[7436]= 1000068799;
assign addr[7437]= 1033753687;
assign addr[7438]= 1067110699;
assign addr[7439]= 1100129257;
assign addr[7440]= 1132798888;
assign addr[7441]= 1165109230;
assign addr[7442]= 1197050035;
assign addr[7443]= 1228611172;
assign addr[7444]= 1259782632;
assign addr[7445]= 1290554528;
assign addr[7446]= 1320917099;
assign addr[7447]= 1350860716;
assign addr[7448]= 1380375881;
assign addr[7449]= 1409453233;
assign addr[7450]= 1438083551;
assign addr[7451]= 1466257752;
assign addr[7452]= 1493966902;
assign addr[7453]= 1521202211;
assign addr[7454]= 1547955041;
assign addr[7455]= 1574216908;
assign addr[7456]= 1599979481;
assign addr[7457]= 1625234591;
assign addr[7458]= 1649974225;
assign addr[7459]= 1674190539;
assign addr[7460]= 1697875851;
assign addr[7461]= 1721022648;
assign addr[7462]= 1743623590;
assign addr[7463]= 1765671509;
assign addr[7464]= 1787159411;
assign addr[7465]= 1808080480;
assign addr[7466]= 1828428082;
assign addr[7467]= 1848195763;
assign addr[7468]= 1867377253;
assign addr[7469]= 1885966468;
assign addr[7470]= 1903957513;
assign addr[7471]= 1921344681;
assign addr[7472]= 1938122457;
assign addr[7473]= 1954285520;
assign addr[7474]= 1969828744;
assign addr[7475]= 1984747199;
assign addr[7476]= 1999036154;
assign addr[7477]= 2012691075;
assign addr[7478]= 2025707632;
assign addr[7479]= 2038081698;
assign addr[7480]= 2049809346;
assign addr[7481]= 2060886858;
assign addr[7482]= 2071310720;
assign addr[7483]= 2081077626;
assign addr[7484]= 2090184478;
assign addr[7485]= 2098628387;
assign addr[7486]= 2106406677;
assign addr[7487]= 2113516878;
assign addr[7488]= 2119956737;
assign addr[7489]= 2125724211;
assign addr[7490]= 2130817471;
assign addr[7491]= 2135234901;
assign addr[7492]= 2138975100;
assign addr[7493]= 2142036881;
assign addr[7494]= 2144419275;
assign addr[7495]= 2146121524;
assign addr[7496]= 2147143090;
assign addr[7497]= 2147483648;
assign addr[7498]= 2147143090;
assign addr[7499]= 2146121524;
assign addr[7500]= 2144419275;
assign addr[7501]= 2142036881;
assign addr[7502]= 2138975100;
assign addr[7503]= 2135234901;
assign addr[7504]= 2130817471;
assign addr[7505]= 2125724211;
assign addr[7506]= 2119956737;
assign addr[7507]= 2113516878;
assign addr[7508]= 2106406677;
assign addr[7509]= 2098628387;
assign addr[7510]= 2090184478;
assign addr[7511]= 2081077626;
assign addr[7512]= 2071310720;
assign addr[7513]= 2060886858;
assign addr[7514]= 2049809346;
assign addr[7515]= 2038081698;
assign addr[7516]= 2025707632;
assign addr[7517]= 2012691075;
assign addr[7518]= 1999036154;
assign addr[7519]= 1984747199;
assign addr[7520]= 1969828744;
assign addr[7521]= 1954285520;
assign addr[7522]= 1938122457;
assign addr[7523]= 1921344681;
assign addr[7524]= 1903957513;
assign addr[7525]= 1885966468;
assign addr[7526]= 1867377253;
assign addr[7527]= 1848195763;
assign addr[7528]= 1828428082;
assign addr[7529]= 1808080480;
assign addr[7530]= 1787159411;
assign addr[7531]= 1765671509;
assign addr[7532]= 1743623590;
assign addr[7533]= 1721022648;
assign addr[7534]= 1697875851;
assign addr[7535]= 1674190539;
assign addr[7536]= 1649974225;
assign addr[7537]= 1625234591;
assign addr[7538]= 1599979481;
assign addr[7539]= 1574216908;
assign addr[7540]= 1547955041;
assign addr[7541]= 1521202211;
assign addr[7542]= 1493966902;
assign addr[7543]= 1466257752;
assign addr[7544]= 1438083551;
assign addr[7545]= 1409453233;
assign addr[7546]= 1380375881;
assign addr[7547]= 1350860716;
assign addr[7548]= 1320917099;
assign addr[7549]= 1290554528;
assign addr[7550]= 1259782632;
assign addr[7551]= 1228611172;
assign addr[7552]= 1197050035;
assign addr[7553]= 1165109230;
assign addr[7554]= 1132798888;
assign addr[7555]= 1100129257;
assign addr[7556]= 1067110699;
assign addr[7557]= 1033753687;
assign addr[7558]= 1000068799;
assign addr[7559]= 966066720;
assign addr[7560]= 931758235;
assign addr[7561]= 897154224;
assign addr[7562]= 862265664;
assign addr[7563]= 827103620;
assign addr[7564]= 791679244;
assign addr[7565]= 756003771;
assign addr[7566]= 720088517;
assign addr[7567]= 683944874;
assign addr[7568]= 647584304;
assign addr[7569]= 611018340;
assign addr[7570]= 574258580;
assign addr[7571]= 537316682;
assign addr[7572]= 500204365;
assign addr[7573]= 462933398;
assign addr[7574]= 425515602;
assign addr[7575]= 387962847;
assign addr[7576]= 350287041;
assign addr[7577]= 312500135;
assign addr[7578]= 274614114;
assign addr[7579]= 236640993;
assign addr[7580]= 198592817;
assign addr[7581]= 160481654;
assign addr[7582]= 122319591;
assign addr[7583]= 84118732;
assign addr[7584]= 45891193;
assign addr[7585]= 7649098;
assign addr[7586]= -30595422;
assign addr[7587]= -68830239;
assign addr[7588]= -107043224;
assign addr[7589]= -145222259;
assign addr[7590]= -183355234;
assign addr[7591]= -221430054;
assign addr[7592]= -259434643;
assign addr[7593]= -297356948;
assign addr[7594]= -335184940;
assign addr[7595]= -372906622;
assign addr[7596]= -410510029;
assign addr[7597]= -447983235;
assign addr[7598]= -485314355;
assign addr[7599]= -522491548;
assign addr[7600]= -559503022;
assign addr[7601]= -596337040;
assign addr[7602]= -632981917;
assign addr[7603]= -669426032;
assign addr[7604]= -705657826;
assign addr[7605]= -741665807;
assign addr[7606]= -777438554;
assign addr[7607]= -812964722;
assign addr[7608]= -848233042;
assign addr[7609]= -883232329;
assign addr[7610]= -917951481;
assign addr[7611]= -952379488;
assign addr[7612]= -986505429;
assign addr[7613]= -1020318481;
assign addr[7614]= -1053807919;
assign addr[7615]= -1086963121;
assign addr[7616]= -1119773573;
assign addr[7617]= -1152228866;
assign addr[7618]= -1184318708;
assign addr[7619]= -1216032921;
assign addr[7620]= -1247361445;
assign addr[7621]= -1278294345;
assign addr[7622]= -1308821808;
assign addr[7623]= -1338934154;
assign addr[7624]= -1368621831;
assign addr[7625]= -1397875423;
assign addr[7626]= -1426685652;
assign addr[7627]= -1455043381;
assign addr[7628]= -1482939614;
assign addr[7629]= -1510365504;
assign addr[7630]= -1537312353;
assign addr[7631]= -1563771613;
assign addr[7632]= -1589734894;
assign addr[7633]= -1615193959;
assign addr[7634]= -1640140734;
assign addr[7635]= -1664567307;
assign addr[7636]= -1688465931;
assign addr[7637]= -1711829025;
assign addr[7638]= -1734649179;
assign addr[7639]= -1756919156;
assign addr[7640]= -1778631892;
assign addr[7641]= -1799780501;
assign addr[7642]= -1820358275;
assign addr[7643]= -1840358687;
assign addr[7644]= -1859775393;
assign addr[7645]= -1878602237;
assign addr[7646]= -1896833245;
assign addr[7647]= -1914462636;
assign addr[7648]= -1931484818;
assign addr[7649]= -1947894393;
assign addr[7650]= -1963686155;
assign addr[7651]= -1978855097;
assign addr[7652]= -1993396407;
assign addr[7653]= -2007305472;
assign addr[7654]= -2020577882;
assign addr[7655]= -2033209426;
assign addr[7656]= -2045196100;
assign addr[7657]= -2056534099;
assign addr[7658]= -2067219829;
assign addr[7659]= -2077249901;
assign addr[7660]= -2086621133;
assign addr[7661]= -2095330553;
assign addr[7662]= -2103375398;
assign addr[7663]= -2110753117;
assign addr[7664]= -2117461370;
assign addr[7665]= -2123498030;
assign addr[7666]= -2128861181;
assign addr[7667]= -2133549123;
assign addr[7668]= -2137560369;
assign addr[7669]= -2140893646;
assign addr[7670]= -2143547897;
assign addr[7671]= -2145522281;
assign addr[7672]= -2146816171;
assign addr[7673]= -2147429158;
assign addr[7674]= -2147361045;
assign addr[7675]= -2146611856;
assign addr[7676]= -2145181827;
assign addr[7677]= -2143071413;
assign addr[7678]= -2140281282;
assign addr[7679]= -2136812319;
assign addr[7680]= -2132665626;
assign addr[7681]= -2127842516;
assign addr[7682]= -2122344521;
assign addr[7683]= -2116173382;
assign addr[7684]= -2109331059;
assign addr[7685]= -2101819720;
assign addr[7686]= -2093641749;
assign addr[7687]= -2084799740;
assign addr[7688]= -2075296495;
assign addr[7689]= -2065135031;
assign addr[7690]= -2054318569;
assign addr[7691]= -2042850540;
assign addr[7692]= -2030734582;
assign addr[7693]= -2017974537;
assign addr[7694]= -2004574453;
assign addr[7695]= -1990538579;
assign addr[7696]= -1975871368;
assign addr[7697]= -1960577471;
assign addr[7698]= -1944661739;
assign addr[7699]= -1928129220;
assign addr[7700]= -1910985158;
assign addr[7701]= -1893234990;
assign addr[7702]= -1874884346;
assign addr[7703]= -1855939047;
assign addr[7704]= -1836405100;
assign addr[7705]= -1816288703;
assign addr[7706]= -1795596234;
assign addr[7707]= -1774334257;
assign addr[7708]= -1752509516;
assign addr[7709]= -1730128933;
assign addr[7710]= -1707199606;
assign addr[7711]= -1683728808;
assign addr[7712]= -1659723983;
assign addr[7713]= -1635192744;
assign addr[7714]= -1610142873;
assign addr[7715]= -1584582314;
assign addr[7716]= -1558519173;
assign addr[7717]= -1531961719;
assign addr[7718]= -1504918373;
assign addr[7719]= -1477397714;
assign addr[7720]= -1449408469;
assign addr[7721]= -1420959516;
assign addr[7722]= -1392059879;
assign addr[7723]= -1362718723;
assign addr[7724]= -1332945355;
assign addr[7725]= -1302749217;
assign addr[7726]= -1272139887;
assign addr[7727]= -1241127074;
assign addr[7728]= -1209720613;
assign addr[7729]= -1177930466;
assign addr[7730]= -1145766716;
assign addr[7731]= -1113239564;
assign addr[7732]= -1080359326;
assign addr[7733]= -1047136432;
assign addr[7734]= -1013581418;
assign addr[7735]= -979704927;
assign addr[7736]= -945517704;
assign addr[7737]= -911030591;
assign addr[7738]= -876254528;
assign addr[7739]= -841200544;
assign addr[7740]= -805879757;
assign addr[7741]= -770303369;
assign addr[7742]= -734482665;
assign addr[7743]= -698429006;
assign addr[7744]= -662153826;
assign addr[7745]= -625668632;
assign addr[7746]= -588984994;
assign addr[7747]= -552114549;
assign addr[7748]= -515068990;
assign addr[7749]= -477860067;
assign addr[7750]= -440499581;
assign addr[7751]= -402999383;
assign addr[7752]= -365371365;
assign addr[7753]= -327627463;
assign addr[7754]= -289779648;
assign addr[7755]= -251839923;
assign addr[7756]= -213820322;
assign addr[7757]= -175732905;
assign addr[7758]= -137589750;
assign addr[7759]= -99402956;
assign addr[7760]= -61184634;
assign addr[7761]= -22946906;
assign addr[7762]= 15298099;
assign addr[7763]= 53538253;
assign addr[7764]= 91761426;
assign addr[7765]= 129955495;
assign addr[7766]= 168108346;
assign addr[7767]= 206207878;
assign addr[7768]= 244242007;
assign addr[7769]= 282198671;
assign addr[7770]= 320065829;
assign addr[7771]= 357831473;
assign addr[7772]= 395483624;
assign addr[7773]= 433010339;
assign addr[7774]= 470399716;
assign addr[7775]= 507639898;
assign addr[7776]= 544719071;
assign addr[7777]= 581625477;
assign addr[7778]= 618347408;
assign addr[7779]= 654873219;
assign addr[7780]= 691191324;
assign addr[7781]= 727290205;
assign addr[7782]= 763158411;
assign addr[7783]= 798784567;
assign addr[7784]= 834157373;
assign addr[7785]= 869265610;
assign addr[7786]= 904098143;
assign addr[7787]= 938643924;
assign addr[7788]= 972891995;
assign addr[7789]= 1006831495;
assign addr[7790]= 1040451659;
assign addr[7791]= 1073741824;
assign addr[7792]= 1106691431;
assign addr[7793]= 1139290029;
assign addr[7794]= 1171527280;
assign addr[7795]= 1203392958;
assign addr[7796]= 1234876957;
assign addr[7797]= 1265969291;
assign addr[7798]= 1296660098;
assign addr[7799]= 1326939644;
assign addr[7800]= 1356798326;
assign addr[7801]= 1386226674;
assign addr[7802]= 1415215352;
assign addr[7803]= 1443755168;
assign addr[7804]= 1471837070;
assign addr[7805]= 1499452149;
assign addr[7806]= 1526591649;
assign addr[7807]= 1553246960;
assign addr[7808]= 1579409630;
assign addr[7809]= 1605071359;
assign addr[7810]= 1630224009;
assign addr[7811]= 1654859602;
assign addr[7812]= 1678970324;
assign addr[7813]= 1702548529;
assign addr[7814]= 1725586737;
assign addr[7815]= 1748077642;
assign addr[7816]= 1770014111;
assign addr[7817]= 1791389186;
assign addr[7818]= 1812196087;
assign addr[7819]= 1832428215;
assign addr[7820]= 1852079154;
assign addr[7821]= 1871142669;
assign addr[7822]= 1889612716;
assign addr[7823]= 1907483436;
assign addr[7824]= 1924749160;
assign addr[7825]= 1941404413;
assign addr[7826]= 1957443913;
assign addr[7827]= 1972862571;
assign addr[7828]= 1987655498;
assign addr[7829]= 2001818002;
assign addr[7830]= 2015345591;
assign addr[7831]= 2028233973;
assign addr[7832]= 2040479063;
assign addr[7833]= 2052076975;
assign addr[7834]= 2063024031;
assign addr[7835]= 2073316760;
assign addr[7836]= 2082951896;
assign addr[7837]= 2091926384;
assign addr[7838]= 2100237377;
assign addr[7839]= 2107882239;
assign addr[7840]= 2114858546;
assign addr[7841]= 2121164085;
assign addr[7842]= 2126796855;
assign addr[7843]= 2131755071;
assign addr[7844]= 2136037160;
assign addr[7845]= 2139641764;
assign addr[7846]= 2142567738;
assign addr[7847]= 2144814157;
assign addr[7848]= 2146380306;
assign addr[7849]= 2147265689;
assign addr[7850]= 2147470025;
assign addr[7851]= 2146993250;
assign addr[7852]= 2145835515;
assign addr[7853]= 2143997187;
assign addr[7854]= 2141478848;
assign addr[7855]= 2138281298;
assign addr[7856]= 2134405552;
assign addr[7857]= 2129852837;
assign addr[7858]= 2124624598;
assign addr[7859]= 2118722494;
assign addr[7860]= 2112148396;
assign addr[7861]= 2104904390;
assign addr[7862]= 2096992772;
assign addr[7863]= 2088416053;
assign addr[7864]= 2079176953;
assign addr[7865]= 2069278401;
assign addr[7866]= 2058723538;
assign addr[7867]= 2047515711;
assign addr[7868]= 2035658475;
assign addr[7869]= 2023155591;
assign addr[7870]= 2010011024;
assign addr[7871]= 1996228943;
assign addr[7872]= 1981813720;
assign addr[7873]= 1966769926;
assign addr[7874]= 1951102334;
assign addr[7875]= 1934815911;
assign addr[7876]= 1917915825;
assign addr[7877]= 1900407434;
assign addr[7878]= 1882296293;
assign addr[7879]= 1863588145;
assign addr[7880]= 1844288924;
assign addr[7881]= 1824404752;
assign addr[7882]= 1803941934;
assign addr[7883]= 1782906961;
assign addr[7884]= 1761306505;
assign addr[7885]= 1739147417;
assign addr[7886]= 1716436725;
assign addr[7887]= 1693181631;
assign addr[7888]= 1669389513;
assign addr[7889]= 1645067915;
assign addr[7890]= 1620224553;
assign addr[7891]= 1594867305;
assign addr[7892]= 1569004214;
assign addr[7893]= 1542643483;
assign addr[7894]= 1515793473;
assign addr[7895]= 1488462700;
assign addr[7896]= 1460659832;
assign addr[7897]= 1432393688;
assign addr[7898]= 1403673233;
assign addr[7899]= 1374507575;
assign addr[7900]= 1344905966;
assign addr[7901]= 1314877795;
assign addr[7902]= 1284432584;
assign addr[7903]= 1253579991;
assign addr[7904]= 1222329801;
assign addr[7905]= 1190691925;
assign addr[7906]= 1158676398;
assign addr[7907]= 1126293375;
assign addr[7908]= 1093553126;
assign addr[7909]= 1060466036;
assign addr[7910]= 1027042599;
assign addr[7911]= 993293415;
assign addr[7912]= 959229189;
assign addr[7913]= 924860725;
assign addr[7914]= 890198924;
assign addr[7915]= 855254778;
assign addr[7916]= 820039373;
assign addr[7917]= 784563876;
assign addr[7918]= 748839539;
assign addr[7919]= 712877694;
assign addr[7920]= 676689746;
assign addr[7921]= 640287172;
assign addr[7922]= 603681519;
assign addr[7923]= 566884397;
assign addr[7924]= 529907477;
assign addr[7925]= 492762486;
assign addr[7926]= 455461206;
assign addr[7927]= 418015468;
assign addr[7928]= 380437148;
assign addr[7929]= 342738165;
assign addr[7930]= 304930476;
assign addr[7931]= 267026072;
assign addr[7932]= 229036977;
assign addr[7933]= 190975237;
assign addr[7934]= 152852926;
assign addr[7935]= 114682135;
assign addr[7936]= 76474970;
assign addr[7937]= 38243550;
assign addr[7938]= 0;
assign addr[7939]= -38243550;
assign addr[7940]= -76474970;
assign addr[7941]= -114682135;
assign addr[7942]= -152852926;
assign addr[7943]= -190975237;
assign addr[7944]= -229036977;
assign addr[7945]= -267026072;
assign addr[7946]= -304930476;
assign addr[7947]= -342738165;
assign addr[7948]= -380437148;
assign addr[7949]= -418015468;
assign addr[7950]= -455461206;
assign addr[7951]= -492762486;
assign addr[7952]= -529907477;
assign addr[7953]= -566884397;
assign addr[7954]= -603681519;
assign addr[7955]= -640287172;
assign addr[7956]= -676689746;
assign addr[7957]= -712877694;
assign addr[7958]= -748839539;
assign addr[7959]= -784563876;
assign addr[7960]= -820039373;
assign addr[7961]= -855254778;
assign addr[7962]= -890198924;
assign addr[7963]= -924860725;
assign addr[7964]= -959229189;
assign addr[7965]= -993293415;
assign addr[7966]= -1027042599;
assign addr[7967]= -1060466036;
assign addr[7968]= -1093553126;
assign addr[7969]= -1126293375;
assign addr[7970]= -1158676398;
assign addr[7971]= -1190691925;
assign addr[7972]= -1222329801;
assign addr[7973]= -1253579991;
assign addr[7974]= -1284432584;
assign addr[7975]= -1314877795;
assign addr[7976]= -1344905966;
assign addr[7977]= -1374507575;
assign addr[7978]= -1403673233;
assign addr[7979]= -1432393688;
assign addr[7980]= -1460659832;
assign addr[7981]= -1488462700;
assign addr[7982]= -1515793473;
assign addr[7983]= -1542643483;
assign addr[7984]= -1569004214;
assign addr[7985]= -1594867305;
assign addr[7986]= -1620224553;
assign addr[7987]= -1645067915;
assign addr[7988]= -1669389513;
assign addr[7989]= -1693181631;
assign addr[7990]= -1716436725;
assign addr[7991]= -1739147417;
assign addr[7992]= -1761306505;
assign addr[7993]= -1782906961;
assign addr[7994]= -1803941934;
assign addr[7995]= -1824404752;
assign addr[7996]= -1844288924;
assign addr[7997]= -1863588145;
assign addr[7998]= -1882296293;
assign addr[7999]= -1900407434;
assign addr[8000]= -1917915825;
assign addr[8001]= -1934815911;
assign addr[8002]= -1951102334;
assign addr[8003]= -1966769926;
assign addr[8004]= -1981813720;
assign addr[8005]= -1996228943;
assign addr[8006]= -2010011024;
assign addr[8007]= -2023155591;
assign addr[8008]= -2035658475;
assign addr[8009]= -2047515711;
assign addr[8010]= -2058723538;
assign addr[8011]= -2069278401;
assign addr[8012]= -2079176953;
assign addr[8013]= -2088416053;
assign addr[8014]= -2096992772;
assign addr[8015]= -2104904390;
assign addr[8016]= -2112148396;
assign addr[8017]= -2118722494;
assign addr[8018]= -2124624598;
assign addr[8019]= -2129852837;
assign addr[8020]= -2134405552;
assign addr[8021]= -2138281298;
assign addr[8022]= -2141478848;
assign addr[8023]= -2143997187;
assign addr[8024]= -2145835515;
assign addr[8025]= -2146993250;
assign addr[8026]= -2147470025;
assign addr[8027]= -2147265689;
assign addr[8028]= -2146380306;
assign addr[8029]= -2144814157;
assign addr[8030]= -2142567738;
assign addr[8031]= -2139641764;
assign addr[8032]= -2136037160;
assign addr[8033]= -2131755071;
assign addr[8034]= -2126796855;
assign addr[8035]= -2121164085;
assign addr[8036]= -2114858546;
assign addr[8037]= -2107882239;
assign addr[8038]= -2100237377;
assign addr[8039]= -2091926384;
assign addr[8040]= -2082951896;
assign addr[8041]= -2073316760;
assign addr[8042]= -2063024031;
assign addr[8043]= -2052076975;
assign addr[8044]= -2040479063;
assign addr[8045]= -2028233973;
assign addr[8046]= -2015345591;
assign addr[8047]= -2001818002;
assign addr[8048]= -1987655498;
assign addr[8049]= -1972862571;
assign addr[8050]= -1957443913;
assign addr[8051]= -1941404413;
assign addr[8052]= -1924749160;
assign addr[8053]= -1907483436;
assign addr[8054]= -1889612716;
assign addr[8055]= -1871142669;
assign addr[8056]= -1852079154;
assign addr[8057]= -1832428215;
assign addr[8058]= -1812196087;
assign addr[8059]= -1791389186;
assign addr[8060]= -1770014111;
assign addr[8061]= -1748077642;
assign addr[8062]= -1725586737;
assign addr[8063]= -1702548529;
assign addr[8064]= -1678970324;
assign addr[8065]= -1654859602;
assign addr[8066]= -1630224009;
assign addr[8067]= -1605071359;
assign addr[8068]= -1579409630;
assign addr[8069]= -1553246960;
assign addr[8070]= -1526591649;
assign addr[8071]= -1499452149;
assign addr[8072]= -1471837070;
assign addr[8073]= -1443755168;
assign addr[8074]= -1415215352;
assign addr[8075]= -1386226674;
assign addr[8076]= -1356798326;
assign addr[8077]= -1326939644;
assign addr[8078]= -1296660098;
assign addr[8079]= -1265969291;
assign addr[8080]= -1234876957;
assign addr[8081]= -1203392958;
assign addr[8082]= -1171527280;
assign addr[8083]= -1139290029;
assign addr[8084]= -1106691431;
assign addr[8085]= -1073741824;
assign addr[8086]= -1040451659;
assign addr[8087]= -1006831495;
assign addr[8088]= -972891995;
assign addr[8089]= -938643924;
assign addr[8090]= -904098143;
assign addr[8091]= -869265610;
assign addr[8092]= -834157373;
assign addr[8093]= -798784567;
assign addr[8094]= -763158411;
assign addr[8095]= -727290205;
assign addr[8096]= -691191324;
assign addr[8097]= -654873219;
assign addr[8098]= -618347408;
assign addr[8099]= -581625477;
assign addr[8100]= -544719071;
assign addr[8101]= -507639898;
assign addr[8102]= -470399716;
assign addr[8103]= -433010339;
assign addr[8104]= -395483624;
assign addr[8105]= -357831473;
assign addr[8106]= -320065829;
assign addr[8107]= -282198671;
assign addr[8108]= -244242007;
assign addr[8109]= -206207878;
assign addr[8110]= -168108346;
assign addr[8111]= -129955495;
assign addr[8112]= -91761426;
assign addr[8113]= -53538253;
assign addr[8114]= -15298099;
assign addr[8115]= 22946906;
assign addr[8116]= 61184634;
assign addr[8117]= 99402956;
assign addr[8118]= 137589750;
assign addr[8119]= 175732905;
assign addr[8120]= 213820322;
assign addr[8121]= 251839923;
assign addr[8122]= 289779648;
assign addr[8123]= 327627463;
assign addr[8124]= 365371365;
assign addr[8125]= 402999383;
assign addr[8126]= 440499581;
assign addr[8127]= 477860067;
assign addr[8128]= 515068990;
assign addr[8129]= 552114549;
assign addr[8130]= 588984994;
assign addr[8131]= 625668632;
assign addr[8132]= 662153826;
assign addr[8133]= 698429006;
assign addr[8134]= 734482665;
assign addr[8135]= 770303369;
assign addr[8136]= 805879757;
assign addr[8137]= 841200544;
assign addr[8138]= 876254528;
assign addr[8139]= 911030591;
assign addr[8140]= 945517704;
assign addr[8141]= 979704927;
assign addr[8142]= 1013581418;
assign addr[8143]= 1047136432;
assign addr[8144]= 1080359326;
assign addr[8145]= 1113239564;
assign addr[8146]= 1145766716;
assign addr[8147]= 1177930466;
assign addr[8148]= 1209720613;
assign addr[8149]= 1241127074;
assign addr[8150]= 1272139887;
assign addr[8151]= 1302749217;
assign addr[8152]= 1332945355;
assign addr[8153]= 1362718723;
assign addr[8154]= 1392059879;
assign addr[8155]= 1420959516;
assign addr[8156]= 1449408469;
assign addr[8157]= 1477397714;
assign addr[8158]= 1504918373;
assign addr[8159]= 1531961719;
assign addr[8160]= 1558519173;
assign addr[8161]= 1584582314;
assign addr[8162]= 1610142873;
assign addr[8163]= 1635192744;
assign addr[8164]= 1659723983;
assign addr[8165]= 1683728808;
assign addr[8166]= 1707199606;
assign addr[8167]= 1730128933;
assign addr[8168]= 1752509516;
assign addr[8169]= 1774334257;
assign addr[8170]= 1795596234;
assign addr[8171]= 1816288703;
assign addr[8172]= 1836405100;
assign addr[8173]= 1855939047;
assign addr[8174]= 1874884346;
assign addr[8175]= 1893234990;
assign addr[8176]= 1910985158;
assign addr[8177]= 1928129220;
assign addr[8178]= 1944661739;
assign addr[8179]= 1960577471;
assign addr[8180]= 1975871368;
assign addr[8181]= 1990538579;
assign addr[8182]= 2004574453;
assign addr[8183]= 2017974537;
assign addr[8184]= 2030734582;
assign addr[8185]= 2042850540;
assign addr[8186]= 2054318569;
assign addr[8187]= 2065135031;
assign addr[8188]= 2075296495;
assign addr[8189]= 2084799740;
assign addr[8190]= 2093641749;
assign addr[8191]= 2101819720;
assign addr[8192]= 2109331059;
assign addr[8193]= 2116173382;
assign addr[8194]= 2122344521;
assign addr[8195]= 2127842516;
assign addr[8196]= 2132665626;
assign addr[8197]= 2136812319;
assign addr[8198]= 2140281282;
assign addr[8199]= 2143071413;
assign addr[8200]= 2145181827;
assign addr[8201]= 2146611856;
assign addr[8202]= 2147361045;
assign addr[8203]= 2147429158;
assign addr[8204]= 2146816171;
assign addr[8205]= 2145522281;
assign addr[8206]= 2143547897;
assign addr[8207]= 2140893646;
assign addr[8208]= 2137560369;
assign addr[8209]= 2133549123;
assign addr[8210]= 2128861181;
assign addr[8211]= 2123498030;
assign addr[8212]= 2117461370;
assign addr[8213]= 2110753117;
assign addr[8214]= 2103375398;
assign addr[8215]= 2095330553;
assign addr[8216]= 2086621133;
assign addr[8217]= 2077249901;
assign addr[8218]= 2067219829;
assign addr[8219]= 2056534099;
assign addr[8220]= 2045196100;
assign addr[8221]= 2033209426;
assign addr[8222]= 2020577882;
assign addr[8223]= 2007305472;
assign addr[8224]= 1993396407;
assign addr[8225]= 1978855097;
assign addr[8226]= 1963686155;
assign addr[8227]= 1947894393;
assign addr[8228]= 1931484818;
assign addr[8229]= 1914462636;
assign addr[8230]= 1896833245;
assign addr[8231]= 1878602237;
assign addr[8232]= 1859775393;
assign addr[8233]= 1840358687;
assign addr[8234]= 1820358275;
assign addr[8235]= 1799780501;
assign addr[8236]= 1778631892;
assign addr[8237]= 1756919156;
assign addr[8238]= 1734649179;
assign addr[8239]= 1711829025;
assign addr[8240]= 1688465931;
assign addr[8241]= 1664567307;
assign addr[8242]= 1640140734;
assign addr[8243]= 1615193959;
assign addr[8244]= 1589734894;
assign addr[8245]= 1563771613;
assign addr[8246]= 1537312353;
assign addr[8247]= 1510365504;
assign addr[8248]= 1482939614;
assign addr[8249]= 1455043381;
assign addr[8250]= 1426685652;
assign addr[8251]= 1397875423;
assign addr[8252]= 1368621831;
assign addr[8253]= 1338934154;
assign addr[8254]= 1308821808;
assign addr[8255]= 1278294345;
assign addr[8256]= 1247361445;
assign addr[8257]= 1216032921;
assign addr[8258]= 1184318708;
assign addr[8259]= 1152228866;
assign addr[8260]= 1119773573;
assign addr[8261]= 1086963121;
assign addr[8262]= 1053807919;
assign addr[8263]= 1020318481;
assign addr[8264]= 986505429;
assign addr[8265]= 952379488;
assign addr[8266]= 917951481;
assign addr[8267]= 883232329;
assign addr[8268]= 848233042;
assign addr[8269]= 812964722;
assign addr[8270]= 777438554;
assign addr[8271]= 741665807;
assign addr[8272]= 705657826;
assign addr[8273]= 669426032;
assign addr[8274]= 632981917;
assign addr[8275]= 596337040;
assign addr[8276]= 559503022;
assign addr[8277]= 522491548;
assign addr[8278]= 485314355;
assign addr[8279]= 447983235;
assign addr[8280]= 410510029;
assign addr[8281]= 372906622;
assign addr[8282]= 335184940;
assign addr[8283]= 297356948;
assign addr[8284]= 259434643;
assign addr[8285]= 221430054;
assign addr[8286]= 183355234;
assign addr[8287]= 145222259;
assign addr[8288]= 107043224;
assign addr[8289]= 68830239;
assign addr[8290]= 30595422;
assign addr[8291]= -7649098;
assign addr[8292]= -45891193;
assign addr[8293]= -84118732;
assign addr[8294]= -122319591;
assign addr[8295]= -160481654;
assign addr[8296]= -198592817;
assign addr[8297]= -236640993;
assign addr[8298]= -274614114;
assign addr[8299]= -312500135;
assign addr[8300]= -350287041;
assign addr[8301]= -387962847;
assign addr[8302]= -425515602;
assign addr[8303]= -462933398;
assign addr[8304]= -500204365;
assign addr[8305]= -537316682;
assign addr[8306]= -574258580;
assign addr[8307]= -611018340;
assign addr[8308]= -647584304;
assign addr[8309]= -683944874;
assign addr[8310]= -720088517;
assign addr[8311]= -756003771;
assign addr[8312]= -791679244;
assign addr[8313]= -827103620;
assign addr[8314]= -862265664;
assign addr[8315]= -897154224;
assign addr[8316]= -931758235;
assign addr[8317]= -966066720;
assign addr[8318]= -1000068799;
assign addr[8319]= -1033753687;
assign addr[8320]= -1067110699;
assign addr[8321]= -1100129257;
assign addr[8322]= -1132798888;
assign addr[8323]= -1165109230;
assign addr[8324]= -1197050035;
assign addr[8325]= -1228611172;
assign addr[8326]= -1259782632;
assign addr[8327]= -1290554528;
assign addr[8328]= -1320917099;
assign addr[8329]= -1350860716;
assign addr[8330]= -1380375881;
assign addr[8331]= -1409453233;
assign addr[8332]= -1438083551;
assign addr[8333]= -1466257752;
assign addr[8334]= -1493966902;
assign addr[8335]= -1521202211;
assign addr[8336]= -1547955041;
assign addr[8337]= -1574216908;
assign addr[8338]= -1599979481;
assign addr[8339]= -1625234591;
assign addr[8340]= -1649974225;
assign addr[8341]= -1674190539;
assign addr[8342]= -1697875851;
assign addr[8343]= -1721022648;
assign addr[8344]= -1743623590;
assign addr[8345]= -1765671509;
assign addr[8346]= -1787159411;
assign addr[8347]= -1808080480;
assign addr[8348]= -1828428082;
assign addr[8349]= -1848195763;
assign addr[8350]= -1867377253;
assign addr[8351]= -1885966468;
assign addr[8352]= -1903957513;
assign addr[8353]= -1921344681;
assign addr[8354]= -1938122457;
assign addr[8355]= -1954285520;
assign addr[8356]= -1969828744;
assign addr[8357]= -1984747199;
assign addr[8358]= -1999036154;
assign addr[8359]= -2012691075;
assign addr[8360]= -2025707632;
assign addr[8361]= -2038081698;
assign addr[8362]= -2049809346;
assign addr[8363]= -2060886858;
assign addr[8364]= -2071310720;
assign addr[8365]= -2081077626;
assign addr[8366]= -2090184478;
assign addr[8367]= -2098628387;
assign addr[8368]= -2106406677;
assign addr[8369]= -2113516878;
assign addr[8370]= -2119956737;
assign addr[8371]= -2125724211;
assign addr[8372]= -2130817471;
assign addr[8373]= -2135234901;
assign addr[8374]= -2138975100;
assign addr[8375]= -2142036881;
assign addr[8376]= -2144419275;
assign addr[8377]= -2146121524;
assign addr[8378]= -2147143090;
assign addr[8379]= -2147483648;
assign addr[8380]= -2147143090;
assign addr[8381]= -2146121524;
assign addr[8382]= -2144419275;
assign addr[8383]= -2142036881;
assign addr[8384]= -2138975100;
assign addr[8385]= -2135234901;
assign addr[8386]= -2130817471;
assign addr[8387]= -2125724211;
assign addr[8388]= -2119956737;
assign addr[8389]= -2113516878;
assign addr[8390]= -2106406677;
assign addr[8391]= -2098628387;
assign addr[8392]= -2090184478;
assign addr[8393]= -2081077626;
assign addr[8394]= -2071310720;
assign addr[8395]= -2060886858;
assign addr[8396]= -2049809346;
assign addr[8397]= -2038081698;
assign addr[8398]= -2025707632;
assign addr[8399]= -2012691075;
assign addr[8400]= -1999036154;
assign addr[8401]= -1984747199;
assign addr[8402]= -1969828744;
assign addr[8403]= -1954285520;
assign addr[8404]= -1938122457;
assign addr[8405]= -1921344681;
assign addr[8406]= -1903957513;
assign addr[8407]= -1885966468;
assign addr[8408]= -1867377253;
assign addr[8409]= -1848195763;
assign addr[8410]= -1828428082;
assign addr[8411]= -1808080480;
assign addr[8412]= -1787159411;
assign addr[8413]= -1765671509;
assign addr[8414]= -1743623590;
assign addr[8415]= -1721022648;
assign addr[8416]= -1697875851;
assign addr[8417]= -1674190539;
assign addr[8418]= -1649974225;
assign addr[8419]= -1625234591;
assign addr[8420]= -1599979481;
assign addr[8421]= -1574216908;
assign addr[8422]= -1547955041;
assign addr[8423]= -1521202211;
assign addr[8424]= -1493966902;
assign addr[8425]= -1466257752;
assign addr[8426]= -1438083551;
assign addr[8427]= -1409453233;
assign addr[8428]= -1380375881;
assign addr[8429]= -1350860716;
assign addr[8430]= -1320917099;
assign addr[8431]= -1290554528;
assign addr[8432]= -1259782632;
assign addr[8433]= -1228611172;
assign addr[8434]= -1197050035;
assign addr[8435]= -1165109230;
assign addr[8436]= -1132798888;
assign addr[8437]= -1100129257;
assign addr[8438]= -1067110699;
assign addr[8439]= -1033753687;
assign addr[8440]= -1000068799;
assign addr[8441]= -966066720;
assign addr[8442]= -931758235;
assign addr[8443]= -897154224;
assign addr[8444]= -862265664;
assign addr[8445]= -827103620;
assign addr[8446]= -791679244;
assign addr[8447]= -756003771;
assign addr[8448]= -720088517;
assign addr[8449]= -683944874;
assign addr[8450]= -647584304;
assign addr[8451]= -611018340;
assign addr[8452]= -574258580;
assign addr[8453]= -537316682;
assign addr[8454]= -500204365;
assign addr[8455]= -462933398;
assign addr[8456]= -425515602;
assign addr[8457]= -387962847;
assign addr[8458]= -350287041;
assign addr[8459]= -312500135;
assign addr[8460]= -274614114;
assign addr[8461]= -236640993;
assign addr[8462]= -198592817;
assign addr[8463]= -160481654;
assign addr[8464]= -122319591;
assign addr[8465]= -84118732;
assign addr[8466]= -45891193;
assign addr[8467]= -7649098;
assign addr[8468]= 30595422;
assign addr[8469]= 68830239;
assign addr[8470]= 107043224;
assign addr[8471]= 145222259;
assign addr[8472]= 183355234;
assign addr[8473]= 221430054;
assign addr[8474]= 259434643;
assign addr[8475]= 297356948;
assign addr[8476]= 335184940;
assign addr[8477]= 372906622;
assign addr[8478]= 410510029;
assign addr[8479]= 447983235;
assign addr[8480]= 485314355;
assign addr[8481]= 522491548;
assign addr[8482]= 559503022;
assign addr[8483]= 596337040;
assign addr[8484]= 632981917;
assign addr[8485]= 669426032;
assign addr[8486]= 705657826;
assign addr[8487]= 741665807;
assign addr[8488]= 777438554;
assign addr[8489]= 812964722;
assign addr[8490]= 848233042;
assign addr[8491]= 883232329;
assign addr[8492]= 917951481;
assign addr[8493]= 952379488;
assign addr[8494]= 986505429;
assign addr[8495]= 1020318481;
assign addr[8496]= 1053807919;
assign addr[8497]= 1086963121;
assign addr[8498]= 1119773573;
assign addr[8499]= 1152228866;
assign addr[8500]= 1184318708;
assign addr[8501]= 1216032921;
assign addr[8502]= 1247361445;
assign addr[8503]= 1278294345;
assign addr[8504]= 1308821808;
assign addr[8505]= 1338934154;
assign addr[8506]= 1368621831;
assign addr[8507]= 1397875423;
assign addr[8508]= 1426685652;
assign addr[8509]= 1455043381;
assign addr[8510]= 1482939614;
assign addr[8511]= 1510365504;
assign addr[8512]= 1537312353;
assign addr[8513]= 1563771613;
assign addr[8514]= 1589734894;
assign addr[8515]= 1615193959;
assign addr[8516]= 1640140734;
assign addr[8517]= 1664567307;
assign addr[8518]= 1688465931;
assign addr[8519]= 1711829025;
assign addr[8520]= 1734649179;
assign addr[8521]= 1756919156;
assign addr[8522]= 1778631892;
assign addr[8523]= 1799780501;
assign addr[8524]= 1820358275;
assign addr[8525]= 1840358687;
assign addr[8526]= 1859775393;
assign addr[8527]= 1878602237;
assign addr[8528]= 1896833245;
assign addr[8529]= 1914462636;
assign addr[8530]= 1931484818;
assign addr[8531]= 1947894393;
assign addr[8532]= 1963686155;
assign addr[8533]= 1978855097;
assign addr[8534]= 1993396407;
assign addr[8535]= 2007305472;
assign addr[8536]= 2020577882;
assign addr[8537]= 2033209426;
assign addr[8538]= 2045196100;
assign addr[8539]= 2056534099;
assign addr[8540]= 2067219829;
assign addr[8541]= 2077249901;
assign addr[8542]= 2086621133;
assign addr[8543]= 2095330553;
assign addr[8544]= 2103375398;
assign addr[8545]= 2110753117;
assign addr[8546]= 2117461370;
assign addr[8547]= 2123498030;
assign addr[8548]= 2128861181;
assign addr[8549]= 2133549123;
assign addr[8550]= 2137560369;
assign addr[8551]= 2140893646;
assign addr[8552]= 2143547897;
assign addr[8553]= 2145522281;
assign addr[8554]= 2146816171;
assign addr[8555]= 2147429158;
assign addr[8556]= 2147361045;
assign addr[8557]= 2146611856;
assign addr[8558]= 2145181827;
assign addr[8559]= 2143071413;
assign addr[8560]= 2140281282;
assign addr[8561]= 2136812319;
assign addr[8562]= 2132665626;
assign addr[8563]= 2127842516;
assign addr[8564]= 2122344521;
assign addr[8565]= 2116173382;
assign addr[8566]= 2109331059;
assign addr[8567]= 2101819720;
assign addr[8568]= 2093641749;
assign addr[8569]= 2084799740;
assign addr[8570]= 2075296495;
assign addr[8571]= 2065135031;
assign addr[8572]= 2054318569;
assign addr[8573]= 2042850540;
assign addr[8574]= 2030734582;
assign addr[8575]= 2017974537;
assign addr[8576]= 2004574453;
assign addr[8577]= 1990538579;
assign addr[8578]= 1975871368;
assign addr[8579]= 1960577471;
assign addr[8580]= 1944661739;
assign addr[8581]= 1928129220;
assign addr[8582]= 1910985158;
assign addr[8583]= 1893234990;
assign addr[8584]= 1874884346;
assign addr[8585]= 1855939047;
assign addr[8586]= 1836405100;
assign addr[8587]= 1816288703;
assign addr[8588]= 1795596234;
assign addr[8589]= 1774334257;
assign addr[8590]= 1752509516;
assign addr[8591]= 1730128933;
assign addr[8592]= 1707199606;
assign addr[8593]= 1683728808;
assign addr[8594]= 1659723983;
assign addr[8595]= 1635192744;
assign addr[8596]= 1610142873;
assign addr[8597]= 1584582314;
assign addr[8598]= 1558519173;
assign addr[8599]= 1531961719;
assign addr[8600]= 1504918373;
assign addr[8601]= 1477397714;
assign addr[8602]= 1449408469;
assign addr[8603]= 1420959516;
assign addr[8604]= 1392059879;
assign addr[8605]= 1362718723;
assign addr[8606]= 1332945355;
assign addr[8607]= 1302749217;
assign addr[8608]= 1272139887;
assign addr[8609]= 1241127074;
assign addr[8610]= 1209720613;
assign addr[8611]= 1177930466;
assign addr[8612]= 1145766716;
assign addr[8613]= 1113239564;
assign addr[8614]= 1080359326;
assign addr[8615]= 1047136432;
assign addr[8616]= 1013581418;
assign addr[8617]= 979704927;
assign addr[8618]= 945517704;
assign addr[8619]= 911030591;
assign addr[8620]= 876254528;
assign addr[8621]= 841200544;
assign addr[8622]= 805879757;
assign addr[8623]= 770303369;
assign addr[8624]= 734482665;
assign addr[8625]= 698429006;
assign addr[8626]= 662153826;
assign addr[8627]= 625668632;
assign addr[8628]= 588984994;
assign addr[8629]= 552114549;
assign addr[8630]= 515068990;
assign addr[8631]= 477860067;
assign addr[8632]= 440499581;
assign addr[8633]= 402999383;
assign addr[8634]= 365371365;
assign addr[8635]= 327627463;
assign addr[8636]= 289779648;
assign addr[8637]= 251839923;
assign addr[8638]= 213820322;
assign addr[8639]= 175732905;
assign addr[8640]= 137589750;
assign addr[8641]= 99402956;
assign addr[8642]= 61184634;
assign addr[8643]= 22946906;
assign addr[8644]= -15298099;
assign addr[8645]= -53538253;
assign addr[8646]= -91761426;
assign addr[8647]= -129955495;
assign addr[8648]= -168108346;
assign addr[8649]= -206207878;
assign addr[8650]= -244242007;
assign addr[8651]= -282198671;
assign addr[8652]= -320065829;
assign addr[8653]= -357831473;
assign addr[8654]= -395483624;
assign addr[8655]= -433010339;
assign addr[8656]= -470399716;
assign addr[8657]= -507639898;
assign addr[8658]= -544719071;
assign addr[8659]= -581625477;
assign addr[8660]= -618347408;
assign addr[8661]= -654873219;
assign addr[8662]= -691191324;
assign addr[8663]= -727290205;
assign addr[8664]= -763158411;
assign addr[8665]= -798784567;
assign addr[8666]= -834157373;
assign addr[8667]= -869265610;
assign addr[8668]= -904098143;
assign addr[8669]= -938643924;
assign addr[8670]= -972891995;
assign addr[8671]= -1006831495;
assign addr[8672]= -1040451659;
assign addr[8673]= -1073741824;
assign addr[8674]= -1106691431;
assign addr[8675]= -1139290029;
assign addr[8676]= -1171527280;
assign addr[8677]= -1203392958;
assign addr[8678]= -1234876957;
assign addr[8679]= -1265969291;
assign addr[8680]= -1296660098;
assign addr[8681]= -1326939644;
assign addr[8682]= -1356798326;
assign addr[8683]= -1386226674;
assign addr[8684]= -1415215352;
assign addr[8685]= -1443755168;
assign addr[8686]= -1471837070;
assign addr[8687]= -1499452149;
assign addr[8688]= -1526591649;
assign addr[8689]= -1553246960;
assign addr[8690]= -1579409630;
assign addr[8691]= -1605071359;
assign addr[8692]= -1630224009;
assign addr[8693]= -1654859602;
assign addr[8694]= -1678970324;
assign addr[8695]= -1702548529;
assign addr[8696]= -1725586737;
assign addr[8697]= -1748077642;
assign addr[8698]= -1770014111;
assign addr[8699]= -1791389186;
assign addr[8700]= -1812196087;
assign addr[8701]= -1832428215;
assign addr[8702]= -1852079154;
assign addr[8703]= -1871142669;
assign addr[8704]= -1889612716;
assign addr[8705]= -1907483436;
assign addr[8706]= -1924749160;
assign addr[8707]= -1941404413;
assign addr[8708]= -1957443913;
assign addr[8709]= -1972862571;
assign addr[8710]= -1987655498;
assign addr[8711]= -2001818002;
assign addr[8712]= -2015345591;
assign addr[8713]= -2028233973;
assign addr[8714]= -2040479063;
assign addr[8715]= -2052076975;
assign addr[8716]= -2063024031;
assign addr[8717]= -2073316760;
assign addr[8718]= -2082951896;
assign addr[8719]= -2091926384;
assign addr[8720]= -2100237377;
assign addr[8721]= -2107882239;
assign addr[8722]= -2114858546;
assign addr[8723]= -2121164085;
assign addr[8724]= -2126796855;
assign addr[8725]= -2131755071;
assign addr[8726]= -2136037160;
assign addr[8727]= -2139641764;
assign addr[8728]= -2142567738;
assign addr[8729]= -2144814157;
assign addr[8730]= -2146380306;
assign addr[8731]= -2147265689;
assign addr[8732]= -2147470025;
assign addr[8733]= -2146993250;
assign addr[8734]= -2145835515;
assign addr[8735]= -2143997187;
assign addr[8736]= -2141478848;
assign addr[8737]= -2138281298;
assign addr[8738]= -2134405552;
assign addr[8739]= -2129852837;
assign addr[8740]= -2124624598;
assign addr[8741]= -2118722494;
assign addr[8742]= -2112148396;
assign addr[8743]= -2104904390;
assign addr[8744]= -2096992772;
assign addr[8745]= -2088416053;
assign addr[8746]= -2079176953;
assign addr[8747]= -2069278401;
assign addr[8748]= -2058723538;
assign addr[8749]= -2047515711;
assign addr[8750]= -2035658475;
assign addr[8751]= -2023155591;
assign addr[8752]= -2010011024;
assign addr[8753]= -1996228943;
assign addr[8754]= -1981813720;
assign addr[8755]= -1966769926;
assign addr[8756]= -1951102334;
assign addr[8757]= -1934815911;
assign addr[8758]= -1917915825;
assign addr[8759]= -1900407434;
assign addr[8760]= -1882296293;
assign addr[8761]= -1863588145;
assign addr[8762]= -1844288924;
assign addr[8763]= -1824404752;
assign addr[8764]= -1803941934;
assign addr[8765]= -1782906961;
assign addr[8766]= -1761306505;
assign addr[8767]= -1739147417;
assign addr[8768]= -1716436725;
assign addr[8769]= -1693181631;
assign addr[8770]= -1669389513;
assign addr[8771]= -1645067915;
assign addr[8772]= -1620224553;
assign addr[8773]= -1594867305;
assign addr[8774]= -1569004214;
assign addr[8775]= -1542643483;
assign addr[8776]= -1515793473;
assign addr[8777]= -1488462700;
assign addr[8778]= -1460659832;
assign addr[8779]= -1432393688;
assign addr[8780]= -1403673233;
assign addr[8781]= -1374507575;
assign addr[8782]= -1344905966;
assign addr[8783]= -1314877795;
assign addr[8784]= -1284432584;
assign addr[8785]= -1253579991;
assign addr[8786]= -1222329801;
assign addr[8787]= -1190691925;
assign addr[8788]= -1158676398;
assign addr[8789]= -1126293375;
assign addr[8790]= -1093553126;
assign addr[8791]= -1060466036;
assign addr[8792]= -1027042599;
assign addr[8793]= -993293415;
assign addr[8794]= -959229189;
assign addr[8795]= -924860725;
assign addr[8796]= -890198924;
assign addr[8797]= -855254778;
assign addr[8798]= -820039373;
assign addr[8799]= -784563876;
assign addr[8800]= -748839539;
assign addr[8801]= -712877694;
assign addr[8802]= -676689746;
assign addr[8803]= -640287172;
assign addr[8804]= -603681519;
assign addr[8805]= -566884397;
assign addr[8806]= -529907477;
assign addr[8807]= -492762486;
assign addr[8808]= -455461206;
assign addr[8809]= -418015468;
assign addr[8810]= -380437148;
assign addr[8811]= -342738165;
assign addr[8812]= -304930476;
assign addr[8813]= -267026072;
assign addr[8814]= -229036977;
assign addr[8815]= -190975237;
assign addr[8816]= -152852926;
assign addr[8817]= -114682135;
assign addr[8818]= -76474970;
assign addr[8819]= -38243550;
assign addr[8820]= 0;
assign addr[8821]= 38243550;
assign addr[8822]= 76474970;
assign addr[8823]= 114682135;
assign addr[8824]= 152852926;
assign addr[8825]= 190975237;
assign addr[8826]= 229036977;
assign addr[8827]= 267026072;
assign addr[8828]= 304930476;
assign addr[8829]= 342738165;
assign addr[8830]= 380437148;
assign addr[8831]= 418015468;
assign addr[8832]= 455461206;
assign addr[8833]= 492762486;
assign addr[8834]= 529907477;
assign addr[8835]= 566884397;
assign addr[8836]= 603681519;
assign addr[8837]= 640287172;
assign addr[8838]= 676689746;
assign addr[8839]= 712877694;
assign addr[8840]= 748839539;
assign addr[8841]= 784563876;
assign addr[8842]= 820039373;
assign addr[8843]= 855254778;
assign addr[8844]= 890198924;
assign addr[8845]= 924860725;
assign addr[8846]= 959229189;
assign addr[8847]= 993293415;
assign addr[8848]= 1027042599;
assign addr[8849]= 1060466036;
assign addr[8850]= 1093553126;
assign addr[8851]= 1126293375;
assign addr[8852]= 1158676398;
assign addr[8853]= 1190691925;
assign addr[8854]= 1222329801;
assign addr[8855]= 1253579991;
assign addr[8856]= 1284432584;
assign addr[8857]= 1314877795;
assign addr[8858]= 1344905966;
assign addr[8859]= 1374507575;
assign addr[8860]= 1403673233;
assign addr[8861]= 1432393688;
assign addr[8862]= 1460659832;
assign addr[8863]= 1488462700;
assign addr[8864]= 1515793473;
assign addr[8865]= 1542643483;
assign addr[8866]= 1569004214;
assign addr[8867]= 1594867305;
assign addr[8868]= 1620224553;
assign addr[8869]= 1645067915;
assign addr[8870]= 1669389513;
assign addr[8871]= 1693181631;
assign addr[8872]= 1716436725;
assign addr[8873]= 1739147417;
assign addr[8874]= 1761306505;
assign addr[8875]= 1782906961;
assign addr[8876]= 1803941934;
assign addr[8877]= 1824404752;
assign addr[8878]= 1844288924;
assign addr[8879]= 1863588145;
assign addr[8880]= 1882296293;
assign addr[8881]= 1900407434;
assign addr[8882]= 1917915825;
assign addr[8883]= 1934815911;
assign addr[8884]= 1951102334;
assign addr[8885]= 1966769926;
assign addr[8886]= 1981813720;
assign addr[8887]= 1996228943;
assign addr[8888]= 2010011024;
assign addr[8889]= 2023155591;
assign addr[8890]= 2035658475;
assign addr[8891]= 2047515711;
assign addr[8892]= 2058723538;
assign addr[8893]= 2069278401;
assign addr[8894]= 2079176953;
assign addr[8895]= 2088416053;
assign addr[8896]= 2096992772;
assign addr[8897]= 2104904390;
assign addr[8898]= 2112148396;
assign addr[8899]= 2118722494;
assign addr[8900]= 2124624598;
assign addr[8901]= 2129852837;
assign addr[8902]= 2134405552;
assign addr[8903]= 2138281298;
assign addr[8904]= 2141478848;
assign addr[8905]= 2143997187;
assign addr[8906]= 2145835515;
assign addr[8907]= 2146993250;
assign addr[8908]= 2147470025;
assign addr[8909]= 2147265689;
assign addr[8910]= 2146380306;
assign addr[8911]= 2144814157;
assign addr[8912]= 2142567738;
assign addr[8913]= 2139641764;
assign addr[8914]= 2136037160;
assign addr[8915]= 2131755071;
assign addr[8916]= 2126796855;
assign addr[8917]= 2121164085;
assign addr[8918]= 2114858546;
assign addr[8919]= 2107882239;
assign addr[8920]= 2100237377;
assign addr[8921]= 2091926384;
assign addr[8922]= 2082951896;
assign addr[8923]= 2073316760;
assign addr[8924]= 2063024031;
assign addr[8925]= 2052076975;
assign addr[8926]= 2040479063;
assign addr[8927]= 2028233973;
assign addr[8928]= 2015345591;
assign addr[8929]= 2001818002;
assign addr[8930]= 1987655498;
assign addr[8931]= 1972862571;
assign addr[8932]= 1957443913;
assign addr[8933]= 1941404413;
assign addr[8934]= 1924749160;
assign addr[8935]= 1907483436;
assign addr[8936]= 1889612716;
assign addr[8937]= 1871142669;
assign addr[8938]= 1852079154;
assign addr[8939]= 1832428215;
assign addr[8940]= 1812196087;
assign addr[8941]= 1791389186;
assign addr[8942]= 1770014111;
assign addr[8943]= 1748077642;
assign addr[8944]= 1725586737;
assign addr[8945]= 1702548529;
assign addr[8946]= 1678970324;
assign addr[8947]= 1654859602;
assign addr[8948]= 1630224009;
assign addr[8949]= 1605071359;
assign addr[8950]= 1579409630;
assign addr[8951]= 1553246960;
assign addr[8952]= 1526591649;
assign addr[8953]= 1499452149;
assign addr[8954]= 1471837070;
assign addr[8955]= 1443755168;
assign addr[8956]= 1415215352;
assign addr[8957]= 1386226674;
assign addr[8958]= 1356798326;
assign addr[8959]= 1326939644;
assign addr[8960]= 1296660098;
assign addr[8961]= 1265969291;
assign addr[8962]= 1234876957;
assign addr[8963]= 1203392958;
assign addr[8964]= 1171527280;
assign addr[8965]= 1139290029;
assign addr[8966]= 1106691431;
assign addr[8967]= 1073741824;
assign addr[8968]= 1040451659;
assign addr[8969]= 1006831495;
assign addr[8970]= 972891995;
assign addr[8971]= 938643924;
assign addr[8972]= 904098143;
assign addr[8973]= 869265610;
assign addr[8974]= 834157373;
assign addr[8975]= 798784567;
assign addr[8976]= 763158411;
assign addr[8977]= 727290205;
assign addr[8978]= 691191324;
assign addr[8979]= 654873219;
assign addr[8980]= 618347408;
assign addr[8981]= 581625477;
assign addr[8982]= 544719071;
assign addr[8983]= 507639898;
assign addr[8984]= 470399716;
assign addr[8985]= 433010339;
assign addr[8986]= 395483624;
assign addr[8987]= 357831473;
assign addr[8988]= 320065829;
assign addr[8989]= 282198671;
assign addr[8990]= 244242007;
assign addr[8991]= 206207878;
assign addr[8992]= 168108346;
assign addr[8993]= 129955495;
assign addr[8994]= 91761426;
assign addr[8995]= 53538253;
assign addr[8996]= 15298099;
assign addr[8997]= -22946906;
assign addr[8998]= -61184634;
assign addr[8999]= -99402956;
assign addr[9000]= -137589750;
assign addr[9001]= -175732905;
assign addr[9002]= -213820322;
assign addr[9003]= -251839923;
assign addr[9004]= -289779648;
assign addr[9005]= -327627463;
assign addr[9006]= -365371365;
assign addr[9007]= -402999383;
assign addr[9008]= -440499581;
assign addr[9009]= -477860067;
assign addr[9010]= -515068990;
assign addr[9011]= -552114549;
assign addr[9012]= -588984994;
assign addr[9013]= -625668632;
assign addr[9014]= -662153826;
assign addr[9015]= -698429006;
assign addr[9016]= -734482665;
assign addr[9017]= -770303369;
assign addr[9018]= -805879757;
assign addr[9019]= -841200544;
assign addr[9020]= -876254528;
assign addr[9021]= -911030591;
assign addr[9022]= -945517704;
assign addr[9023]= -979704927;
assign addr[9024]= -1013581418;
assign addr[9025]= -1047136432;
assign addr[9026]= -1080359326;
assign addr[9027]= -1113239564;
assign addr[9028]= -1145766716;
assign addr[9029]= -1177930466;
assign addr[9030]= -1209720613;
assign addr[9031]= -1241127074;
assign addr[9032]= -1272139887;
assign addr[9033]= -1302749217;
assign addr[9034]= -1332945355;
assign addr[9035]= -1362718723;
assign addr[9036]= -1392059879;
assign addr[9037]= -1420959516;
assign addr[9038]= -1449408469;
assign addr[9039]= -1477397714;
assign addr[9040]= -1504918373;
assign addr[9041]= -1531961719;
assign addr[9042]= -1558519173;
assign addr[9043]= -1584582314;
assign addr[9044]= -1610142873;
assign addr[9045]= -1635192744;
assign addr[9046]= -1659723983;
assign addr[9047]= -1683728808;
assign addr[9048]= -1707199606;
assign addr[9049]= -1730128933;
assign addr[9050]= -1752509516;
assign addr[9051]= -1774334257;
assign addr[9052]= -1795596234;
assign addr[9053]= -1816288703;
assign addr[9054]= -1836405100;
assign addr[9055]= -1855939047;
assign addr[9056]= -1874884346;
assign addr[9057]= -1893234990;
assign addr[9058]= -1910985158;
assign addr[9059]= -1928129220;
assign addr[9060]= -1944661739;
assign addr[9061]= -1960577471;
assign addr[9062]= -1975871368;
assign addr[9063]= -1990538579;
assign addr[9064]= -2004574453;
assign addr[9065]= -2017974537;
assign addr[9066]= -2030734582;
assign addr[9067]= -2042850540;
assign addr[9068]= -2054318569;
assign addr[9069]= -2065135031;
assign addr[9070]= -2075296495;
assign addr[9071]= -2084799740;
assign addr[9072]= -2093641749;
assign addr[9073]= -2101819720;
assign addr[9074]= -2109331059;
assign addr[9075]= -2116173382;
assign addr[9076]= -2122344521;
assign addr[9077]= -2127842516;
assign addr[9078]= -2132665626;
assign addr[9079]= -2136812319;
assign addr[9080]= -2140281282;
assign addr[9081]= -2143071413;
assign addr[9082]= -2145181827;
assign addr[9083]= -2146611856;
assign addr[9084]= -2147361045;
assign addr[9085]= -2147429158;
assign addr[9086]= -2146816171;
assign addr[9087]= -2145522281;
assign addr[9088]= -2143547897;
assign addr[9089]= -2140893646;
assign addr[9090]= -2137560369;
assign addr[9091]= -2133549123;
assign addr[9092]= -2128861181;
assign addr[9093]= -2123498030;
assign addr[9094]= -2117461370;
assign addr[9095]= -2110753117;
assign addr[9096]= -2103375398;
assign addr[9097]= -2095330553;
assign addr[9098]= -2086621133;
assign addr[9099]= -2077249901;
assign addr[9100]= -2067219829;
assign addr[9101]= -2056534099;
assign addr[9102]= -2045196100;
assign addr[9103]= -2033209426;
assign addr[9104]= -2020577882;
assign addr[9105]= -2007305472;
assign addr[9106]= -1993396407;
assign addr[9107]= -1978855097;
assign addr[9108]= -1963686155;
assign addr[9109]= -1947894393;
assign addr[9110]= -1931484818;
assign addr[9111]= -1914462636;
assign addr[9112]= -1896833245;
assign addr[9113]= -1878602237;
assign addr[9114]= -1859775393;
assign addr[9115]= -1840358687;
assign addr[9116]= -1820358275;
assign addr[9117]= -1799780501;
assign addr[9118]= -1778631892;
assign addr[9119]= -1756919156;
assign addr[9120]= -1734649179;
assign addr[9121]= -1711829025;
assign addr[9122]= -1688465931;
assign addr[9123]= -1664567307;
assign addr[9124]= -1640140734;
assign addr[9125]= -1615193959;
assign addr[9126]= -1589734894;
assign addr[9127]= -1563771613;
assign addr[9128]= -1537312353;
assign addr[9129]= -1510365504;
assign addr[9130]= -1482939614;
assign addr[9131]= -1455043381;
assign addr[9132]= -1426685652;
assign addr[9133]= -1397875423;
assign addr[9134]= -1368621831;
assign addr[9135]= -1338934154;
assign addr[9136]= -1308821808;
assign addr[9137]= -1278294345;
assign addr[9138]= -1247361445;
assign addr[9139]= -1216032921;
assign addr[9140]= -1184318708;
assign addr[9141]= -1152228866;
assign addr[9142]= -1119773573;
assign addr[9143]= -1086963121;
assign addr[9144]= -1053807919;
assign addr[9145]= -1020318481;
assign addr[9146]= -986505429;
assign addr[9147]= -952379488;
assign addr[9148]= -917951481;
assign addr[9149]= -883232329;
assign addr[9150]= -848233042;
assign addr[9151]= -812964722;
assign addr[9152]= -777438554;
assign addr[9153]= -741665807;
assign addr[9154]= -705657826;
assign addr[9155]= -669426032;
assign addr[9156]= -632981917;
assign addr[9157]= -596337040;
assign addr[9158]= -559503022;
assign addr[9159]= -522491548;
assign addr[9160]= -485314355;
assign addr[9161]= -447983235;
assign addr[9162]= -410510029;
assign addr[9163]= -372906622;
assign addr[9164]= -335184940;
assign addr[9165]= -297356948;
assign addr[9166]= -259434643;
assign addr[9167]= -221430054;
assign addr[9168]= -183355234;
assign addr[9169]= -145222259;
assign addr[9170]= -107043224;
assign addr[9171]= -68830239;
assign addr[9172]= -30595422;
assign addr[9173]= 7649098;
assign addr[9174]= 45891193;
assign addr[9175]= 84118732;
assign addr[9176]= 122319591;
assign addr[9177]= 160481654;
assign addr[9178]= 198592817;
assign addr[9179]= 236640993;
assign addr[9180]= 274614114;
assign addr[9181]= 312500135;
assign addr[9182]= 350287041;
assign addr[9183]= 387962847;
assign addr[9184]= 425515602;
assign addr[9185]= 462933398;
assign addr[9186]= 500204365;
assign addr[9187]= 537316682;
assign addr[9188]= 574258580;
assign addr[9189]= 611018340;
assign addr[9190]= 647584304;
assign addr[9191]= 683944874;
assign addr[9192]= 720088517;
assign addr[9193]= 756003771;
assign addr[9194]= 791679244;
assign addr[9195]= 827103620;
assign addr[9196]= 862265664;
assign addr[9197]= 897154224;
assign addr[9198]= 931758235;
assign addr[9199]= 966066720;
assign addr[9200]= 1000068799;
assign addr[9201]= 1033753687;
assign addr[9202]= 1067110699;
assign addr[9203]= 1100129257;
assign addr[9204]= 1132798888;
assign addr[9205]= 1165109230;
assign addr[9206]= 1197050035;
assign addr[9207]= 1228611172;
assign addr[9208]= 1259782632;
assign addr[9209]= 1290554528;
assign addr[9210]= 1320917099;
assign addr[9211]= 1350860716;
assign addr[9212]= 1380375881;
assign addr[9213]= 1409453233;
assign addr[9214]= 1438083551;
assign addr[9215]= 1466257752;
assign addr[9216]= 1493966902;
assign addr[9217]= 1521202211;
assign addr[9218]= 1547955041;
assign addr[9219]= 1574216908;
assign addr[9220]= 1599979481;
assign addr[9221]= 1625234591;
assign addr[9222]= 1649974225;
assign addr[9223]= 1674190539;
assign addr[9224]= 1697875851;
assign addr[9225]= 1721022648;
assign addr[9226]= 1743623590;
assign addr[9227]= 1765671509;
assign addr[9228]= 1787159411;
assign addr[9229]= 1808080480;
assign addr[9230]= 1828428082;
assign addr[9231]= 1848195763;
assign addr[9232]= 1867377253;
assign addr[9233]= 1885966468;
assign addr[9234]= 1903957513;
assign addr[9235]= 1921344681;
assign addr[9236]= 1938122457;
assign addr[9237]= 1954285520;
assign addr[9238]= 1969828744;
assign addr[9239]= 1984747199;
assign addr[9240]= 1999036154;
assign addr[9241]= 2012691075;
assign addr[9242]= 2025707632;
assign addr[9243]= 2038081698;
assign addr[9244]= 2049809346;
assign addr[9245]= 2060886858;
assign addr[9246]= 2071310720;
assign addr[9247]= 2081077626;
assign addr[9248]= 2090184478;
assign addr[9249]= 2098628387;
assign addr[9250]= 2106406677;
assign addr[9251]= 2113516878;
assign addr[9252]= 2119956737;
assign addr[9253]= 2125724211;
assign addr[9254]= 2130817471;
assign addr[9255]= 2135234901;
assign addr[9256]= 2138975100;
assign addr[9257]= 2142036881;
assign addr[9258]= 2144419275;
assign addr[9259]= 2146121524;
assign addr[9260]= 2147143090;
assign addr[9261]= 2147483648;
assign addr[9262]= 2147143090;
assign addr[9263]= 2146121524;
assign addr[9264]= 2144419275;
assign addr[9265]= 2142036881;
assign addr[9266]= 2138975100;
assign addr[9267]= 2135234901;
assign addr[9268]= 2130817471;
assign addr[9269]= 2125724211;
assign addr[9270]= 2119956737;
assign addr[9271]= 2113516878;
assign addr[9272]= 2106406677;
assign addr[9273]= 2098628387;
assign addr[9274]= 2090184478;
assign addr[9275]= 2081077626;
assign addr[9276]= 2071310720;
assign addr[9277]= 2060886858;
assign addr[9278]= 2049809346;
assign addr[9279]= 2038081698;
assign addr[9280]= 2025707632;
assign addr[9281]= 2012691075;
assign addr[9282]= 1999036154;
assign addr[9283]= 1984747199;
assign addr[9284]= 1969828744;
assign addr[9285]= 1954285520;
assign addr[9286]= 1938122457;
assign addr[9287]= 1921344681;
assign addr[9288]= 1903957513;
assign addr[9289]= 1885966468;
assign addr[9290]= 1867377253;
assign addr[9291]= 1848195763;
assign addr[9292]= 1828428082;
assign addr[9293]= 1808080480;
assign addr[9294]= 1787159411;
assign addr[9295]= 1765671509;
assign addr[9296]= 1743623590;
assign addr[9297]= 1721022648;
assign addr[9298]= 1697875851;
assign addr[9299]= 1674190539;
assign addr[9300]= 1649974225;
assign addr[9301]= 1625234591;
assign addr[9302]= 1599979481;
assign addr[9303]= 1574216908;
assign addr[9304]= 1547955041;
assign addr[9305]= 1521202211;
assign addr[9306]= 1493966902;
assign addr[9307]= 1466257752;
assign addr[9308]= 1438083551;
assign addr[9309]= 1409453233;
assign addr[9310]= 1380375881;
assign addr[9311]= 1350860716;
assign addr[9312]= 1320917099;
assign addr[9313]= 1290554528;
assign addr[9314]= 1259782632;
assign addr[9315]= 1228611172;
assign addr[9316]= 1197050035;
assign addr[9317]= 1165109230;
assign addr[9318]= 1132798888;
assign addr[9319]= 1100129257;
assign addr[9320]= 1067110699;
assign addr[9321]= 1033753687;
assign addr[9322]= 1000068799;
assign addr[9323]= 966066720;
assign addr[9324]= 931758235;
assign addr[9325]= 897154224;
assign addr[9326]= 862265664;
assign addr[9327]= 827103620;
assign addr[9328]= 791679244;
assign addr[9329]= 756003771;
assign addr[9330]= 720088517;
assign addr[9331]= 683944874;
assign addr[9332]= 647584304;
assign addr[9333]= 611018340;
assign addr[9334]= 574258580;
assign addr[9335]= 537316682;
assign addr[9336]= 500204365;
assign addr[9337]= 462933398;
assign addr[9338]= 425515602;
assign addr[9339]= 387962847;
assign addr[9340]= 350287041;
assign addr[9341]= 312500135;
assign addr[9342]= 274614114;
assign addr[9343]= 236640993;
assign addr[9344]= 198592817;
assign addr[9345]= 160481654;
assign addr[9346]= 122319591;
assign addr[9347]= 84118732;
assign addr[9348]= 45891193;
assign addr[9349]= 7649098;
assign addr[9350]= -30595422;
assign addr[9351]= -68830239;
assign addr[9352]= -107043224;
assign addr[9353]= -145222259;
assign addr[9354]= -183355234;
assign addr[9355]= -221430054;
assign addr[9356]= -259434643;
assign addr[9357]= -297356948;
assign addr[9358]= -335184940;
assign addr[9359]= -372906622;
assign addr[9360]= -410510029;
assign addr[9361]= -447983235;
assign addr[9362]= -485314355;
assign addr[9363]= -522491548;
assign addr[9364]= -559503022;
assign addr[9365]= -596337040;
assign addr[9366]= -632981917;
assign addr[9367]= -669426032;
assign addr[9368]= -705657826;
assign addr[9369]= -741665807;
assign addr[9370]= -777438554;
assign addr[9371]= -812964722;
assign addr[9372]= -848233042;
assign addr[9373]= -883232329;
assign addr[9374]= -917951481;
assign addr[9375]= -952379488;
assign addr[9376]= -986505429;
assign addr[9377]= -1020318481;
assign addr[9378]= -1053807919;
assign addr[9379]= -1086963121;
assign addr[9380]= -1119773573;
assign addr[9381]= -1152228866;
assign addr[9382]= -1184318708;
assign addr[9383]= -1216032921;
assign addr[9384]= -1247361445;
assign addr[9385]= -1278294345;
assign addr[9386]= -1308821808;
assign addr[9387]= -1338934154;
assign addr[9388]= -1368621831;
assign addr[9389]= -1397875423;
assign addr[9390]= -1426685652;
assign addr[9391]= -1455043381;
assign addr[9392]= -1482939614;
assign addr[9393]= -1510365504;
assign addr[9394]= -1537312353;
assign addr[9395]= -1563771613;
assign addr[9396]= -1589734894;
assign addr[9397]= -1615193959;
assign addr[9398]= -1640140734;
assign addr[9399]= -1664567307;
assign addr[9400]= -1688465931;
assign addr[9401]= -1711829025;
assign addr[9402]= -1734649179;
assign addr[9403]= -1756919156;
assign addr[9404]= -1778631892;
assign addr[9405]= -1799780501;
assign addr[9406]= -1820358275;
assign addr[9407]= -1840358687;
assign addr[9408]= -1859775393;
assign addr[9409]= -1878602237;
assign addr[9410]= -1896833245;
assign addr[9411]= -1914462636;
assign addr[9412]= -1931484818;
assign addr[9413]= -1947894393;
assign addr[9414]= -1963686155;
assign addr[9415]= -1978855097;
assign addr[9416]= -1993396407;
assign addr[9417]= -2007305472;
assign addr[9418]= -2020577882;
assign addr[9419]= -2033209426;
assign addr[9420]= -2045196100;
assign addr[9421]= -2056534099;
assign addr[9422]= -2067219829;
assign addr[9423]= -2077249901;
assign addr[9424]= -2086621133;
assign addr[9425]= -2095330553;
assign addr[9426]= -2103375398;
assign addr[9427]= -2110753117;
assign addr[9428]= -2117461370;
assign addr[9429]= -2123498030;
assign addr[9430]= -2128861181;
assign addr[9431]= -2133549123;
assign addr[9432]= -2137560369;
assign addr[9433]= -2140893646;
assign addr[9434]= -2143547897;
assign addr[9435]= -2145522281;
assign addr[9436]= -2146816171;
assign addr[9437]= -2147429158;
assign addr[9438]= -2147361045;
assign addr[9439]= -2146611856;
assign addr[9440]= -2145181827;
assign addr[9441]= -2143071413;
assign addr[9442]= -2140281282;
assign addr[9443]= -2136812319;
assign addr[9444]= -2132665626;
assign addr[9445]= -2127842516;
assign addr[9446]= -2122344521;
assign addr[9447]= -2116173382;
assign addr[9448]= -2109331059;
assign addr[9449]= -2101819720;
assign addr[9450]= -2093641749;
assign addr[9451]= -2084799740;
assign addr[9452]= -2075296495;
assign addr[9453]= -2065135031;
assign addr[9454]= -2054318569;
assign addr[9455]= -2042850540;
assign addr[9456]= -2030734582;
assign addr[9457]= -2017974537;
assign addr[9458]= -2004574453;
assign addr[9459]= -1990538579;
assign addr[9460]= -1975871368;
assign addr[9461]= -1960577471;
assign addr[9462]= -1944661739;
assign addr[9463]= -1928129220;
assign addr[9464]= -1910985158;
assign addr[9465]= -1893234990;
assign addr[9466]= -1874884346;
assign addr[9467]= -1855939047;
assign addr[9468]= -1836405100;
assign addr[9469]= -1816288703;
assign addr[9470]= -1795596234;
assign addr[9471]= -1774334257;
assign addr[9472]= -1752509516;
assign addr[9473]= -1730128933;
assign addr[9474]= -1707199606;
assign addr[9475]= -1683728808;
assign addr[9476]= -1659723983;
assign addr[9477]= -1635192744;
assign addr[9478]= -1610142873;
assign addr[9479]= -1584582314;
assign addr[9480]= -1558519173;
assign addr[9481]= -1531961719;
assign addr[9482]= -1504918373;
assign addr[9483]= -1477397714;
assign addr[9484]= -1449408469;
assign addr[9485]= -1420959516;
assign addr[9486]= -1392059879;
assign addr[9487]= -1362718723;
assign addr[9488]= -1332945355;
assign addr[9489]= -1302749217;
assign addr[9490]= -1272139887;
assign addr[9491]= -1241127074;
assign addr[9492]= -1209720613;
assign addr[9493]= -1177930466;
assign addr[9494]= -1145766716;
assign addr[9495]= -1113239564;
assign addr[9496]= -1080359326;
assign addr[9497]= -1047136432;
assign addr[9498]= -1013581418;
assign addr[9499]= -979704927;
assign addr[9500]= -945517704;
assign addr[9501]= -911030591;
assign addr[9502]= -876254528;
assign addr[9503]= -841200544;
assign addr[9504]= -805879757;
assign addr[9505]= -770303369;
assign addr[9506]= -734482665;
assign addr[9507]= -698429006;
assign addr[9508]= -662153826;
assign addr[9509]= -625668632;
assign addr[9510]= -588984994;
assign addr[9511]= -552114549;
assign addr[9512]= -515068990;
assign addr[9513]= -477860067;
assign addr[9514]= -440499581;
assign addr[9515]= -402999383;
assign addr[9516]= -365371365;
assign addr[9517]= -327627463;
assign addr[9518]= -289779648;
assign addr[9519]= -251839923;
assign addr[9520]= -213820322;
assign addr[9521]= -175732905;
assign addr[9522]= -137589750;
assign addr[9523]= -99402956;
assign addr[9524]= -61184634;
assign addr[9525]= -22946906;
assign addr[9526]= 15298099;
assign addr[9527]= 53538253;
assign addr[9528]= 91761426;
assign addr[9529]= 129955495;
assign addr[9530]= 168108346;
assign addr[9531]= 206207878;
assign addr[9532]= 244242007;
assign addr[9533]= 282198671;
assign addr[9534]= 320065829;
assign addr[9535]= 357831473;
assign addr[9536]= 395483624;
assign addr[9537]= 433010339;
assign addr[9538]= 470399716;
assign addr[9539]= 507639898;
assign addr[9540]= 544719071;
assign addr[9541]= 581625477;
assign addr[9542]= 618347408;
assign addr[9543]= 654873219;
assign addr[9544]= 691191324;
assign addr[9545]= 727290205;
assign addr[9546]= 763158411;
assign addr[9547]= 798784567;
assign addr[9548]= 834157373;
assign addr[9549]= 869265610;
assign addr[9550]= 904098143;
assign addr[9551]= 938643924;
assign addr[9552]= 972891995;
assign addr[9553]= 1006831495;
assign addr[9554]= 1040451659;
assign addr[9555]= 1073741824;
assign addr[9556]= 1106691431;
assign addr[9557]= 1139290029;
assign addr[9558]= 1171527280;
assign addr[9559]= 1203392958;
assign addr[9560]= 1234876957;
assign addr[9561]= 1265969291;
assign addr[9562]= 1296660098;
assign addr[9563]= 1326939644;
assign addr[9564]= 1356798326;
assign addr[9565]= 1386226674;
assign addr[9566]= 1415215352;
assign addr[9567]= 1443755168;
assign addr[9568]= 1471837070;
assign addr[9569]= 1499452149;
assign addr[9570]= 1526591649;
assign addr[9571]= 1553246960;
assign addr[9572]= 1579409630;
assign addr[9573]= 1605071359;
assign addr[9574]= 1630224009;
assign addr[9575]= 1654859602;
assign addr[9576]= 1678970324;
assign addr[9577]= 1702548529;
assign addr[9578]= 1725586737;
assign addr[9579]= 1748077642;
assign addr[9580]= 1770014111;
assign addr[9581]= 1791389186;
assign addr[9582]= 1812196087;
assign addr[9583]= 1832428215;
assign addr[9584]= 1852079154;
assign addr[9585]= 1871142669;
assign addr[9586]= 1889612716;
assign addr[9587]= 1907483436;
assign addr[9588]= 1924749160;
assign addr[9589]= 1941404413;
assign addr[9590]= 1957443913;
assign addr[9591]= 1972862571;
assign addr[9592]= 1987655498;
assign addr[9593]= 2001818002;
assign addr[9594]= 2015345591;
assign addr[9595]= 2028233973;
assign addr[9596]= 2040479063;
assign addr[9597]= 2052076975;
assign addr[9598]= 2063024031;
assign addr[9599]= 2073316760;
assign addr[9600]= 2082951896;
assign addr[9601]= 2091926384;
assign addr[9602]= 2100237377;
assign addr[9603]= 2107882239;
assign addr[9604]= 2114858546;
assign addr[9605]= 2121164085;
assign addr[9606]= 2126796855;
assign addr[9607]= 2131755071;
assign addr[9608]= 2136037160;
assign addr[9609]= 2139641764;
assign addr[9610]= 2142567738;
assign addr[9611]= 2144814157;
assign addr[9612]= 2146380306;
assign addr[9613]= 2147265689;
assign addr[9614]= 2147470025;
assign addr[9615]= 2146993250;
assign addr[9616]= 2145835515;
assign addr[9617]= 2143997187;
assign addr[9618]= 2141478848;
assign addr[9619]= 2138281298;
assign addr[9620]= 2134405552;
assign addr[9621]= 2129852837;
assign addr[9622]= 2124624598;
assign addr[9623]= 2118722494;
assign addr[9624]= 2112148396;
assign addr[9625]= 2104904390;
assign addr[9626]= 2096992772;
assign addr[9627]= 2088416053;
assign addr[9628]= 2079176953;
assign addr[9629]= 2069278401;
assign addr[9630]= 2058723538;
assign addr[9631]= 2047515711;
assign addr[9632]= 2035658475;
assign addr[9633]= 2023155591;
assign addr[9634]= 2010011024;
assign addr[9635]= 1996228943;
assign addr[9636]= 1981813720;
assign addr[9637]= 1966769926;
assign addr[9638]= 1951102334;
assign addr[9639]= 1934815911;
assign addr[9640]= 1917915825;
assign addr[9641]= 1900407434;
assign addr[9642]= 1882296293;
assign addr[9643]= 1863588145;
assign addr[9644]= 1844288924;
assign addr[9645]= 1824404752;
assign addr[9646]= 1803941934;
assign addr[9647]= 1782906961;
assign addr[9648]= 1761306505;
assign addr[9649]= 1739147417;
assign addr[9650]= 1716436725;
assign addr[9651]= 1693181631;
assign addr[9652]= 1669389513;
assign addr[9653]= 1645067915;
assign addr[9654]= 1620224553;
assign addr[9655]= 1594867305;
assign addr[9656]= 1569004214;
assign addr[9657]= 1542643483;
assign addr[9658]= 1515793473;
assign addr[9659]= 1488462700;
assign addr[9660]= 1460659832;
assign addr[9661]= 1432393688;
assign addr[9662]= 1403673233;
assign addr[9663]= 1374507575;
assign addr[9664]= 1344905966;
assign addr[9665]= 1314877795;
assign addr[9666]= 1284432584;
assign addr[9667]= 1253579991;
assign addr[9668]= 1222329801;
assign addr[9669]= 1190691925;
assign addr[9670]= 1158676398;
assign addr[9671]= 1126293375;
assign addr[9672]= 1093553126;
assign addr[9673]= 1060466036;
assign addr[9674]= 1027042599;
assign addr[9675]= 993293415;
assign addr[9676]= 959229189;
assign addr[9677]= 924860725;
assign addr[9678]= 890198924;
assign addr[9679]= 855254778;
assign addr[9680]= 820039373;
assign addr[9681]= 784563876;
assign addr[9682]= 748839539;
assign addr[9683]= 712877694;
assign addr[9684]= 676689746;
assign addr[9685]= 640287172;
assign addr[9686]= 603681519;
assign addr[9687]= 566884397;
assign addr[9688]= 529907477;
assign addr[9689]= 492762486;
assign addr[9690]= 455461206;
assign addr[9691]= 418015468;
assign addr[9692]= 380437148;
assign addr[9693]= 342738165;
assign addr[9694]= 304930476;
assign addr[9695]= 267026072;
assign addr[9696]= 229036977;
assign addr[9697]= 190975237;
assign addr[9698]= 152852926;
assign addr[9699]= 114682135;
assign addr[9700]= 76474970;
assign addr[9701]= 38243550;
assign addr[9702]= 0;
assign addr[9703]= -38243550;
assign addr[9704]= -76474970;
assign addr[9705]= -114682135;
assign addr[9706]= -152852926;
assign addr[9707]= -190975237;
assign addr[9708]= -229036977;
assign addr[9709]= -267026072;
assign addr[9710]= -304930476;
assign addr[9711]= -342738165;
assign addr[9712]= -380437148;
assign addr[9713]= -418015468;
assign addr[9714]= -455461206;
assign addr[9715]= -492762486;
assign addr[9716]= -529907477;
assign addr[9717]= -566884397;
assign addr[9718]= -603681519;
assign addr[9719]= -640287172;
assign addr[9720]= -676689746;
assign addr[9721]= -712877694;
assign addr[9722]= -748839539;
assign addr[9723]= -784563876;
assign addr[9724]= -820039373;
assign addr[9725]= -855254778;
assign addr[9726]= -890198924;
assign addr[9727]= -924860725;
assign addr[9728]= -959229189;
assign addr[9729]= -993293415;
assign addr[9730]= -1027042599;
assign addr[9731]= -1060466036;
assign addr[9732]= -1093553126;
assign addr[9733]= -1126293375;
assign addr[9734]= -1158676398;
assign addr[9735]= -1190691925;
assign addr[9736]= -1222329801;
assign addr[9737]= -1253579991;
assign addr[9738]= -1284432584;
assign addr[9739]= -1314877795;
assign addr[9740]= -1344905966;
assign addr[9741]= -1374507575;
assign addr[9742]= -1403673233;
assign addr[9743]= -1432393688;
assign addr[9744]= -1460659832;
assign addr[9745]= -1488462700;
assign addr[9746]= -1515793473;
assign addr[9747]= -1542643483;
assign addr[9748]= -1569004214;
assign addr[9749]= -1594867305;
assign addr[9750]= -1620224553;
assign addr[9751]= -1645067915;
assign addr[9752]= -1669389513;
assign addr[9753]= -1693181631;
assign addr[9754]= -1716436725;
assign addr[9755]= -1739147417;
assign addr[9756]= -1761306505;
assign addr[9757]= -1782906961;
assign addr[9758]= -1803941934;
assign addr[9759]= -1824404752;
assign addr[9760]= -1844288924;
assign addr[9761]= -1863588145;
assign addr[9762]= -1882296293;
assign addr[9763]= -1900407434;
assign addr[9764]= -1917915825;
assign addr[9765]= -1934815911;
assign addr[9766]= -1951102334;
assign addr[9767]= -1966769926;
assign addr[9768]= -1981813720;
assign addr[9769]= -1996228943;
assign addr[9770]= -2010011024;
assign addr[9771]= -2023155591;
assign addr[9772]= -2035658475;
assign addr[9773]= -2047515711;
assign addr[9774]= -2058723538;
assign addr[9775]= -2069278401;
assign addr[9776]= -2079176953;
assign addr[9777]= -2088416053;
assign addr[9778]= -2096992772;
assign addr[9779]= -2104904390;
assign addr[9780]= -2112148396;
assign addr[9781]= -2118722494;
assign addr[9782]= -2124624598;
assign addr[9783]= -2129852837;
assign addr[9784]= -2134405552;
assign addr[9785]= -2138281298;
assign addr[9786]= -2141478848;
assign addr[9787]= -2143997187;
assign addr[9788]= -2145835515;
assign addr[9789]= -2146993250;
assign addr[9790]= -2147470025;
assign addr[9791]= -2147265689;
assign addr[9792]= -2146380306;
assign addr[9793]= -2144814157;
assign addr[9794]= -2142567738;
assign addr[9795]= -2139641764;
assign addr[9796]= -2136037160;
assign addr[9797]= -2131755071;
assign addr[9798]= -2126796855;
assign addr[9799]= -2121164085;
assign addr[9800]= -2114858546;
assign addr[9801]= -2107882239;
assign addr[9802]= -2100237377;
assign addr[9803]= -2091926384;
assign addr[9804]= -2082951896;
assign addr[9805]= -2073316760;
assign addr[9806]= -2063024031;
assign addr[9807]= -2052076975;
assign addr[9808]= -2040479063;
assign addr[9809]= -2028233973;
assign addr[9810]= -2015345591;
assign addr[9811]= -2001818002;
assign addr[9812]= -1987655498;
assign addr[9813]= -1972862571;
assign addr[9814]= -1957443913;
assign addr[9815]= -1941404413;
assign addr[9816]= -1924749160;
assign addr[9817]= -1907483436;
assign addr[9818]= -1889612716;
assign addr[9819]= -1871142669;
assign addr[9820]= -1852079154;
assign addr[9821]= -1832428215;
assign addr[9822]= -1812196087;
assign addr[9823]= -1791389186;
assign addr[9824]= -1770014111;
assign addr[9825]= -1748077642;
assign addr[9826]= -1725586737;
assign addr[9827]= -1702548529;
assign addr[9828]= -1678970324;
assign addr[9829]= -1654859602;
assign addr[9830]= -1630224009;
assign addr[9831]= -1605071359;
assign addr[9832]= -1579409630;
assign addr[9833]= -1553246960;
assign addr[9834]= -1526591649;
assign addr[9835]= -1499452149;
assign addr[9836]= -1471837070;
assign addr[9837]= -1443755168;
assign addr[9838]= -1415215352;
assign addr[9839]= -1386226674;
assign addr[9840]= -1356798326;
assign addr[9841]= -1326939644;
assign addr[9842]= -1296660098;
assign addr[9843]= -1265969291;
assign addr[9844]= -1234876957;
assign addr[9845]= -1203392958;
assign addr[9846]= -1171527280;
assign addr[9847]= -1139290029;
assign addr[9848]= -1106691431;
assign addr[9849]= -1073741824;
assign addr[9850]= -1040451659;
assign addr[9851]= -1006831495;
assign addr[9852]= -972891995;
assign addr[9853]= -938643924;
assign addr[9854]= -904098143;
assign addr[9855]= -869265610;
assign addr[9856]= -834157373;
assign addr[9857]= -798784567;
assign addr[9858]= -763158411;
assign addr[9859]= -727290205;
assign addr[9860]= -691191324;
assign addr[9861]= -654873219;
assign addr[9862]= -618347408;
assign addr[9863]= -581625477;
assign addr[9864]= -544719071;
assign addr[9865]= -507639898;
assign addr[9866]= -470399716;
assign addr[9867]= -433010339;
assign addr[9868]= -395483624;
assign addr[9869]= -357831473;
assign addr[9870]= -320065829;
assign addr[9871]= -282198671;
assign addr[9872]= -244242007;
assign addr[9873]= -206207878;
assign addr[9874]= -168108346;
assign addr[9875]= -129955495;
assign addr[9876]= -91761426;
assign addr[9877]= -53538253;
assign addr[9878]= -15298099;
assign addr[9879]= 22946906;
assign addr[9880]= 61184634;
assign addr[9881]= 99402956;
assign addr[9882]= 137589750;
assign addr[9883]= 175732905;
assign addr[9884]= 213820322;
assign addr[9885]= 251839923;
assign addr[9886]= 289779648;
assign addr[9887]= 327627463;
assign addr[9888]= 365371365;
assign addr[9889]= 402999383;
assign addr[9890]= 440499581;
assign addr[9891]= 477860067;
assign addr[9892]= 515068990;
assign addr[9893]= 552114549;
assign addr[9894]= 588984994;
assign addr[9895]= 625668632;
assign addr[9896]= 662153826;
assign addr[9897]= 698429006;
assign addr[9898]= 734482665;
assign addr[9899]= 770303369;
assign addr[9900]= 805879757;
assign addr[9901]= 841200544;
assign addr[9902]= 876254528;
assign addr[9903]= 911030591;
assign addr[9904]= 945517704;
assign addr[9905]= 979704927;
assign addr[9906]= 1013581418;
assign addr[9907]= 1047136432;
assign addr[9908]= 1080359326;
assign addr[9909]= 1113239564;
assign addr[9910]= 1145766716;
assign addr[9911]= 1177930466;
assign addr[9912]= 1209720613;
assign addr[9913]= 1241127074;
assign addr[9914]= 1272139887;
assign addr[9915]= 1302749217;
assign addr[9916]= 1332945355;
assign addr[9917]= 1362718723;
assign addr[9918]= 1392059879;
assign addr[9919]= 1420959516;
assign addr[9920]= 1449408469;
assign addr[9921]= 1477397714;
assign addr[9922]= 1504918373;
assign addr[9923]= 1531961719;
assign addr[9924]= 1558519173;
assign addr[9925]= 1584582314;
assign addr[9926]= 1610142873;
assign addr[9927]= 1635192744;
assign addr[9928]= 1659723983;
assign addr[9929]= 1683728808;
assign addr[9930]= 1707199606;
assign addr[9931]= 1730128933;
assign addr[9932]= 1752509516;
assign addr[9933]= 1774334257;
assign addr[9934]= 1795596234;
assign addr[9935]= 1816288703;
assign addr[9936]= 1836405100;
assign addr[9937]= 1855939047;
assign addr[9938]= 1874884346;
assign addr[9939]= 1893234990;
assign addr[9940]= 1910985158;
assign addr[9941]= 1928129220;
assign addr[9942]= 1944661739;
assign addr[9943]= 1960577471;
assign addr[9944]= 1975871368;
assign addr[9945]= 1990538579;
assign addr[9946]= 2004574453;
assign addr[9947]= 2017974537;
assign addr[9948]= 2030734582;
assign addr[9949]= 2042850540;
assign addr[9950]= 2054318569;
assign addr[9951]= 2065135031;
assign addr[9952]= 2075296495;
assign addr[9953]= 2084799740;
assign addr[9954]= 2093641749;
assign addr[9955]= 2101819720;
assign addr[9956]= 2109331059;
assign addr[9957]= 2116173382;
assign addr[9958]= 2122344521;
assign addr[9959]= 2127842516;
assign addr[9960]= 2132665626;
assign addr[9961]= 2136812319;
assign addr[9962]= 2140281282;
assign addr[9963]= 2143071413;
assign addr[9964]= 2145181827;
assign addr[9965]= 2146611856;
assign addr[9966]= 2147361045;
assign addr[9967]= 2147429158;
assign addr[9968]= 2146816171;
assign addr[9969]= 2145522281;
assign addr[9970]= 2143547897;
assign addr[9971]= 2140893646;
assign addr[9972]= 2137560369;
assign addr[9973]= 2133549123;
assign addr[9974]= 2128861181;
assign addr[9975]= 2123498030;
assign addr[9976]= 2117461370;
assign addr[9977]= 2110753117;
assign addr[9978]= 2103375398;
assign addr[9979]= 2095330553;
assign addr[9980]= 2086621133;
assign addr[9981]= 2077249901;
assign addr[9982]= 2067219829;
assign addr[9983]= 2056534099;
assign addr[9984]= 2045196100;
assign addr[9985]= 2033209426;
assign addr[9986]= 2020577882;
assign addr[9987]= 2007305472;
assign addr[9988]= 1993396407;
assign addr[9989]= 1978855097;
assign addr[9990]= 1963686155;
assign addr[9991]= 1947894393;
assign addr[9992]= 1931484818;
assign addr[9993]= 1914462636;
assign addr[9994]= 1896833245;
assign addr[9995]= 1878602237;
assign addr[9996]= 1859775393;
assign addr[9997]= 1840358687;
assign addr[9998]= 1820358275;
assign addr[9999]= 1799780501;
assign addr[10000]= 1778631892;
assign addr[10001]= 1756919156;
assign addr[10002]= 1734649179;
assign addr[10003]= 1711829025;
assign addr[10004]= 1688465931;
assign addr[10005]= 1664567307;
assign addr[10006]= 1640140734;
assign addr[10007]= 1615193959;
assign addr[10008]= 1589734894;
assign addr[10009]= 1563771613;
assign addr[10010]= 1537312353;
assign addr[10011]= 1510365504;
assign addr[10012]= 1482939614;
assign addr[10013]= 1455043381;
assign addr[10014]= 1426685652;
assign addr[10015]= 1397875423;
assign addr[10016]= 1368621831;
assign addr[10017]= 1338934154;
assign addr[10018]= 1308821808;
assign addr[10019]= 1278294345;
assign addr[10020]= 1247361445;
assign addr[10021]= 1216032921;
assign addr[10022]= 1184318708;
assign addr[10023]= 1152228866;
assign addr[10024]= 1119773573;
assign addr[10025]= 1086963121;
assign addr[10026]= 1053807919;
assign addr[10027]= 1020318481;
assign addr[10028]= 986505429;
assign addr[10029]= 952379488;
assign addr[10030]= 917951481;
assign addr[10031]= 883232329;
assign addr[10032]= 848233042;
assign addr[10033]= 812964722;
assign addr[10034]= 777438554;
assign addr[10035]= 741665807;
assign addr[10036]= 705657826;
assign addr[10037]= 669426032;
assign addr[10038]= 632981917;
assign addr[10039]= 596337040;
assign addr[10040]= 559503022;
assign addr[10041]= 522491548;
assign addr[10042]= 485314355;
assign addr[10043]= 447983235;
assign addr[10044]= 410510029;
assign addr[10045]= 372906622;
assign addr[10046]= 335184940;
assign addr[10047]= 297356948;
assign addr[10048]= 259434643;
assign addr[10049]= 221430054;
assign addr[10050]= 183355234;
assign addr[10051]= 145222259;
assign addr[10052]= 107043224;
assign addr[10053]= 68830239;
assign addr[10054]= 30595422;
assign addr[10055]= -7649098;
assign addr[10056]= -45891193;
assign addr[10057]= -84118732;
assign addr[10058]= -122319591;
assign addr[10059]= -160481654;
assign addr[10060]= -198592817;
assign addr[10061]= -236640993;
assign addr[10062]= -274614114;
assign addr[10063]= -312500135;
assign addr[10064]= -350287041;
assign addr[10065]= -387962847;
assign addr[10066]= -425515602;
assign addr[10067]= -462933398;
assign addr[10068]= -500204365;
assign addr[10069]= -537316682;
assign addr[10070]= -574258580;
assign addr[10071]= -611018340;
assign addr[10072]= -647584304;
assign addr[10073]= -683944874;
assign addr[10074]= -720088517;
assign addr[10075]= -756003771;
assign addr[10076]= -791679244;
assign addr[10077]= -827103620;
assign addr[10078]= -862265664;
assign addr[10079]= -897154224;
assign addr[10080]= -931758235;
assign addr[10081]= -966066720;
assign addr[10082]= -1000068799;
assign addr[10083]= -1033753687;
assign addr[10084]= -1067110699;
assign addr[10085]= -1100129257;
assign addr[10086]= -1132798888;
assign addr[10087]= -1165109230;
assign addr[10088]= -1197050035;
assign addr[10089]= -1228611172;
assign addr[10090]= -1259782632;
assign addr[10091]= -1290554528;
assign addr[10092]= -1320917099;
assign addr[10093]= -1350860716;
assign addr[10094]= -1380375881;
assign addr[10095]= -1409453233;
assign addr[10096]= -1438083551;
assign addr[10097]= -1466257752;
assign addr[10098]= -1493966902;
assign addr[10099]= -1521202211;
assign addr[10100]= -1547955041;
assign addr[10101]= -1574216908;
assign addr[10102]= -1599979481;
assign addr[10103]= -1625234591;
assign addr[10104]= -1649974225;
assign addr[10105]= -1674190539;
assign addr[10106]= -1697875851;
assign addr[10107]= -1721022648;
assign addr[10108]= -1743623590;
assign addr[10109]= -1765671509;
assign addr[10110]= -1787159411;
assign addr[10111]= -1808080480;
assign addr[10112]= -1828428082;
assign addr[10113]= -1848195763;
assign addr[10114]= -1867377253;
assign addr[10115]= -1885966468;
assign addr[10116]= -1903957513;
assign addr[10117]= -1921344681;
assign addr[10118]= -1938122457;
assign addr[10119]= -1954285520;
assign addr[10120]= -1969828744;
assign addr[10121]= -1984747199;
assign addr[10122]= -1999036154;
assign addr[10123]= -2012691075;
assign addr[10124]= -2025707632;
assign addr[10125]= -2038081698;
assign addr[10126]= -2049809346;
assign addr[10127]= -2060886858;
assign addr[10128]= -2071310720;
assign addr[10129]= -2081077626;
assign addr[10130]= -2090184478;
assign addr[10131]= -2098628387;
assign addr[10132]= -2106406677;
assign addr[10133]= -2113516878;
assign addr[10134]= -2119956737;
assign addr[10135]= -2125724211;
assign addr[10136]= -2130817471;
assign addr[10137]= -2135234901;
assign addr[10138]= -2138975100;
assign addr[10139]= -2142036881;
assign addr[10140]= -2144419275;
assign addr[10141]= -2146121524;
assign addr[10142]= -2147143090;
assign addr[10143]= -2147483648;
assign addr[10144]= -2147143090;
assign addr[10145]= -2146121524;
assign addr[10146]= -2144419275;
assign addr[10147]= -2142036881;
assign addr[10148]= -2138975100;
assign addr[10149]= -2135234901;
assign addr[10150]= -2130817471;
assign addr[10151]= -2125724211;
assign addr[10152]= -2119956737;
assign addr[10153]= -2113516878;
assign addr[10154]= -2106406677;
assign addr[10155]= -2098628387;
assign addr[10156]= -2090184478;
assign addr[10157]= -2081077626;
assign addr[10158]= -2071310720;
assign addr[10159]= -2060886858;
assign addr[10160]= -2049809346;
assign addr[10161]= -2038081698;
assign addr[10162]= -2025707632;
assign addr[10163]= -2012691075;
assign addr[10164]= -1999036154;
assign addr[10165]= -1984747199;
assign addr[10166]= -1969828744;
assign addr[10167]= -1954285520;
assign addr[10168]= -1938122457;
assign addr[10169]= -1921344681;
assign addr[10170]= -1903957513;
assign addr[10171]= -1885966468;
assign addr[10172]= -1867377253;
assign addr[10173]= -1848195763;
assign addr[10174]= -1828428082;
assign addr[10175]= -1808080480;
assign addr[10176]= -1787159411;
assign addr[10177]= -1765671509;
assign addr[10178]= -1743623590;
assign addr[10179]= -1721022648;
assign addr[10180]= -1697875851;
assign addr[10181]= -1674190539;
assign addr[10182]= -1649974225;
assign addr[10183]= -1625234591;
assign addr[10184]= -1599979481;
assign addr[10185]= -1574216908;
assign addr[10186]= -1547955041;
assign addr[10187]= -1521202211;
assign addr[10188]= -1493966902;
assign addr[10189]= -1466257752;
assign addr[10190]= -1438083551;
assign addr[10191]= -1409453233;
assign addr[10192]= -1380375881;
assign addr[10193]= -1350860716;
assign addr[10194]= -1320917099;
assign addr[10195]= -1290554528;
assign addr[10196]= -1259782632;
assign addr[10197]= -1228611172;
assign addr[10198]= -1197050035;
assign addr[10199]= -1165109230;
assign addr[10200]= -1132798888;
assign addr[10201]= -1100129257;
assign addr[10202]= -1067110699;
assign addr[10203]= -1033753687;
assign addr[10204]= -1000068799;
assign addr[10205]= -966066720;
assign addr[10206]= -931758235;
assign addr[10207]= -897154224;
assign addr[10208]= -862265664;
assign addr[10209]= -827103620;
assign addr[10210]= -791679244;
assign addr[10211]= -756003771;
assign addr[10212]= -720088517;
assign addr[10213]= -683944874;
assign addr[10214]= -647584304;
assign addr[10215]= -611018340;
assign addr[10216]= -574258580;
assign addr[10217]= -537316682;
assign addr[10218]= -500204365;
assign addr[10219]= -462933398;
assign addr[10220]= -425515602;
assign addr[10221]= -387962847;
assign addr[10222]= -350287041;
assign addr[10223]= -312500135;
assign addr[10224]= -274614114;
assign addr[10225]= -236640993;
assign addr[10226]= -198592817;
assign addr[10227]= -160481654;
assign addr[10228]= -122319591;
assign addr[10229]= -84118732;
assign addr[10230]= -45891193;
assign addr[10231]= -7649098;
assign addr[10232]= 30595422;
assign addr[10233]= 68830239;
assign addr[10234]= 107043224;
assign addr[10235]= 145222259;
assign addr[10236]= 183355234;
assign addr[10237]= 221430054;
assign addr[10238]= 259434643;
assign addr[10239]= 297356948;
assign addr[10240]= 335184940;
assign addr[10241]= 372906622;
assign addr[10242]= 410510029;
assign addr[10243]= 447983235;
assign addr[10244]= 485314355;
assign addr[10245]= 522491548;
assign addr[10246]= 559503022;
assign addr[10247]= 596337040;
assign addr[10248]= 632981917;
assign addr[10249]= 669426032;
assign addr[10250]= 705657826;
assign addr[10251]= 741665807;
assign addr[10252]= 777438554;
assign addr[10253]= 812964722;
assign addr[10254]= 848233042;
assign addr[10255]= 883232329;
assign addr[10256]= 917951481;
assign addr[10257]= 952379488;
assign addr[10258]= 986505429;
assign addr[10259]= 1020318481;
assign addr[10260]= 1053807919;
assign addr[10261]= 1086963121;
assign addr[10262]= 1119773573;
assign addr[10263]= 1152228866;
assign addr[10264]= 1184318708;
assign addr[10265]= 1216032921;
assign addr[10266]= 1247361445;
assign addr[10267]= 1278294345;
assign addr[10268]= 1308821808;
assign addr[10269]= 1338934154;
assign addr[10270]= 1368621831;
assign addr[10271]= 1397875423;
assign addr[10272]= 1426685652;
assign addr[10273]= 1455043381;
assign addr[10274]= 1482939614;
assign addr[10275]= 1510365504;
assign addr[10276]= 1537312353;
assign addr[10277]= 1563771613;
assign addr[10278]= 1589734894;
assign addr[10279]= 1615193959;
assign addr[10280]= 1640140734;
assign addr[10281]= 1664567307;
assign addr[10282]= 1688465931;
assign addr[10283]= 1711829025;
assign addr[10284]= 1734649179;
assign addr[10285]= 1756919156;
assign addr[10286]= 1778631892;
assign addr[10287]= 1799780501;
assign addr[10288]= 1820358275;
assign addr[10289]= 1840358687;
assign addr[10290]= 1859775393;
assign addr[10291]= 1878602237;
assign addr[10292]= 1896833245;
assign addr[10293]= 1914462636;
assign addr[10294]= 1931484818;
assign addr[10295]= 1947894393;
assign addr[10296]= 1963686155;
assign addr[10297]= 1978855097;
assign addr[10298]= 1993396407;
assign addr[10299]= 2007305472;
assign addr[10300]= 2020577882;
assign addr[10301]= 2033209426;
assign addr[10302]= 2045196100;
assign addr[10303]= 2056534099;
assign addr[10304]= 2067219829;
assign addr[10305]= 2077249901;
assign addr[10306]= 2086621133;
assign addr[10307]= 2095330553;
assign addr[10308]= 2103375398;
assign addr[10309]= 2110753117;
assign addr[10310]= 2117461370;
assign addr[10311]= 2123498030;
assign addr[10312]= 2128861181;
assign addr[10313]= 2133549123;
assign addr[10314]= 2137560369;
assign addr[10315]= 2140893646;
assign addr[10316]= 2143547897;
assign addr[10317]= 2145522281;
assign addr[10318]= 2146816171;
assign addr[10319]= 2147429158;
assign addr[10320]= 2147361045;
assign addr[10321]= 2146611856;
assign addr[10322]= 2145181827;
assign addr[10323]= 2143071413;
assign addr[10324]= 2140281282;
assign addr[10325]= 2136812319;
assign addr[10326]= 2132665626;
assign addr[10327]= 2127842516;
assign addr[10328]= 2122344521;
assign addr[10329]= 2116173382;
assign addr[10330]= 2109331059;
assign addr[10331]= 2101819720;
assign addr[10332]= 2093641749;
assign addr[10333]= 2084799740;
assign addr[10334]= 2075296495;
assign addr[10335]= 2065135031;
assign addr[10336]= 2054318569;
assign addr[10337]= 2042850540;
assign addr[10338]= 2030734582;
assign addr[10339]= 2017974537;
assign addr[10340]= 2004574453;
assign addr[10341]= 1990538579;
assign addr[10342]= 1975871368;
assign addr[10343]= 1960577471;
assign addr[10344]= 1944661739;
assign addr[10345]= 1928129220;
assign addr[10346]= 1910985158;
assign addr[10347]= 1893234990;
assign addr[10348]= 1874884346;
assign addr[10349]= 1855939047;
assign addr[10350]= 1836405100;
assign addr[10351]= 1816288703;
assign addr[10352]= 1795596234;
assign addr[10353]= 1774334257;
assign addr[10354]= 1752509516;
assign addr[10355]= 1730128933;
assign addr[10356]= 1707199606;
assign addr[10357]= 1683728808;
assign addr[10358]= 1659723983;
assign addr[10359]= 1635192744;
assign addr[10360]= 1610142873;
assign addr[10361]= 1584582314;
assign addr[10362]= 1558519173;
assign addr[10363]= 1531961719;
assign addr[10364]= 1504918373;
assign addr[10365]= 1477397714;
assign addr[10366]= 1449408469;
assign addr[10367]= 1420959516;
assign addr[10368]= 1392059879;
assign addr[10369]= 1362718723;
assign addr[10370]= 1332945355;
assign addr[10371]= 1302749217;
assign addr[10372]= 1272139887;
assign addr[10373]= 1241127074;
assign addr[10374]= 1209720613;
assign addr[10375]= 1177930466;
assign addr[10376]= 1145766716;
assign addr[10377]= 1113239564;
assign addr[10378]= 1080359326;
assign addr[10379]= 1047136432;
assign addr[10380]= 1013581418;
assign addr[10381]= 979704927;
assign addr[10382]= 945517704;
assign addr[10383]= 911030591;
assign addr[10384]= 876254528;
assign addr[10385]= 841200544;
assign addr[10386]= 805879757;
assign addr[10387]= 770303369;
assign addr[10388]= 734482665;
assign addr[10389]= 698429006;
assign addr[10390]= 662153826;
assign addr[10391]= 625668632;
assign addr[10392]= 588984994;
assign addr[10393]= 552114549;
assign addr[10394]= 515068990;
assign addr[10395]= 477860067;
assign addr[10396]= 440499581;
assign addr[10397]= 402999383;
assign addr[10398]= 365371365;
assign addr[10399]= 327627463;
assign addr[10400]= 289779648;
assign addr[10401]= 251839923;
assign addr[10402]= 213820322;
assign addr[10403]= 175732905;
assign addr[10404]= 137589750;
assign addr[10405]= 99402956;
assign addr[10406]= 61184634;
assign addr[10407]= 22946906;
assign addr[10408]= -15298099;
assign addr[10409]= -53538253;
assign addr[10410]= -91761426;
assign addr[10411]= -129955495;
assign addr[10412]= -168108346;
assign addr[10413]= -206207878;
assign addr[10414]= -244242007;
assign addr[10415]= -282198671;
assign addr[10416]= -320065829;
assign addr[10417]= -357831473;
assign addr[10418]= -395483624;
assign addr[10419]= -433010339;
assign addr[10420]= -470399716;
assign addr[10421]= -507639898;
assign addr[10422]= -544719071;
assign addr[10423]= -581625477;
assign addr[10424]= -618347408;
assign addr[10425]= -654873219;
assign addr[10426]= -691191324;
assign addr[10427]= -727290205;
assign addr[10428]= -763158411;
assign addr[10429]= -798784567;
assign addr[10430]= -834157373;
assign addr[10431]= -869265610;
assign addr[10432]= -904098143;
assign addr[10433]= -938643924;
assign addr[10434]= -972891995;
assign addr[10435]= -1006831495;
assign addr[10436]= -1040451659;
assign addr[10437]= -1073741824;
assign addr[10438]= -1106691431;
assign addr[10439]= -1139290029;
assign addr[10440]= -1171527280;
assign addr[10441]= -1203392958;
assign addr[10442]= -1234876957;
assign addr[10443]= -1265969291;
assign addr[10444]= -1296660098;
assign addr[10445]= -1326939644;
assign addr[10446]= -1356798326;
assign addr[10447]= -1386226674;
assign addr[10448]= -1415215352;
assign addr[10449]= -1443755168;
assign addr[10450]= -1471837070;
assign addr[10451]= -1499452149;
assign addr[10452]= -1526591649;
assign addr[10453]= -1553246960;
assign addr[10454]= -1579409630;
assign addr[10455]= -1605071359;
assign addr[10456]= -1630224009;
assign addr[10457]= -1654859602;
assign addr[10458]= -1678970324;
assign addr[10459]= -1702548529;
assign addr[10460]= -1725586737;
assign addr[10461]= -1748077642;
assign addr[10462]= -1770014111;
assign addr[10463]= -1791389186;
assign addr[10464]= -1812196087;
assign addr[10465]= -1832428215;
assign addr[10466]= -1852079154;
assign addr[10467]= -1871142669;
assign addr[10468]= -1889612716;
assign addr[10469]= -1907483436;
assign addr[10470]= -1924749160;
assign addr[10471]= -1941404413;
assign addr[10472]= -1957443913;
assign addr[10473]= -1972862571;
assign addr[10474]= -1987655498;
assign addr[10475]= -2001818002;
assign addr[10476]= -2015345591;
assign addr[10477]= -2028233973;
assign addr[10478]= -2040479063;
assign addr[10479]= -2052076975;
assign addr[10480]= -2063024031;
assign addr[10481]= -2073316760;
assign addr[10482]= -2082951896;
assign addr[10483]= -2091926384;
assign addr[10484]= -2100237377;
assign addr[10485]= -2107882239;
assign addr[10486]= -2114858546;
assign addr[10487]= -2121164085;
assign addr[10488]= -2126796855;
assign addr[10489]= -2131755071;
assign addr[10490]= -2136037160;
assign addr[10491]= -2139641764;
assign addr[10492]= -2142567738;
assign addr[10493]= -2144814157;
assign addr[10494]= -2146380306;
assign addr[10495]= -2147265689;
assign addr[10496]= -2147470025;
assign addr[10497]= -2146993250;
assign addr[10498]= -2145835515;
assign addr[10499]= -2143997187;
assign addr[10500]= -2141478848;
assign addr[10501]= -2138281298;
assign addr[10502]= -2134405552;
assign addr[10503]= -2129852837;
assign addr[10504]= -2124624598;
assign addr[10505]= -2118722494;
assign addr[10506]= -2112148396;
assign addr[10507]= -2104904390;
assign addr[10508]= -2096992772;
assign addr[10509]= -2088416053;
assign addr[10510]= -2079176953;
assign addr[10511]= -2069278401;
assign addr[10512]= -2058723538;
assign addr[10513]= -2047515711;
assign addr[10514]= -2035658475;
assign addr[10515]= -2023155591;
assign addr[10516]= -2010011024;
assign addr[10517]= -1996228943;
assign addr[10518]= -1981813720;
assign addr[10519]= -1966769926;
assign addr[10520]= -1951102334;
assign addr[10521]= -1934815911;
assign addr[10522]= -1917915825;
assign addr[10523]= -1900407434;
assign addr[10524]= -1882296293;
assign addr[10525]= -1863588145;
assign addr[10526]= -1844288924;
assign addr[10527]= -1824404752;
assign addr[10528]= -1803941934;
assign addr[10529]= -1782906961;
assign addr[10530]= -1761306505;
assign addr[10531]= -1739147417;
assign addr[10532]= -1716436725;
assign addr[10533]= -1693181631;
assign addr[10534]= -1669389513;
assign addr[10535]= -1645067915;
assign addr[10536]= -1620224553;
assign addr[10537]= -1594867305;
assign addr[10538]= -1569004214;
assign addr[10539]= -1542643483;
assign addr[10540]= -1515793473;
assign addr[10541]= -1488462700;
assign addr[10542]= -1460659832;
assign addr[10543]= -1432393688;
assign addr[10544]= -1403673233;
assign addr[10545]= -1374507575;
assign addr[10546]= -1344905966;
assign addr[10547]= -1314877795;
assign addr[10548]= -1284432584;
assign addr[10549]= -1253579991;
assign addr[10550]= -1222329801;
assign addr[10551]= -1190691925;
assign addr[10552]= -1158676398;
assign addr[10553]= -1126293375;
assign addr[10554]= -1093553126;
assign addr[10555]= -1060466036;
assign addr[10556]= -1027042599;
assign addr[10557]= -993293415;
assign addr[10558]= -959229189;
assign addr[10559]= -924860725;
assign addr[10560]= -890198924;
assign addr[10561]= -855254778;
assign addr[10562]= -820039373;
assign addr[10563]= -784563876;
assign addr[10564]= -748839539;
assign addr[10565]= -712877694;
assign addr[10566]= -676689746;
assign addr[10567]= -640287172;
assign addr[10568]= -603681519;
assign addr[10569]= -566884397;
assign addr[10570]= -529907477;
assign addr[10571]= -492762486;
assign addr[10572]= -455461206;
assign addr[10573]= -418015468;
assign addr[10574]= -380437148;
assign addr[10575]= -342738165;
assign addr[10576]= -304930476;
assign addr[10577]= -267026072;
assign addr[10578]= -229036977;
assign addr[10579]= -190975237;
assign addr[10580]= -152852926;
assign addr[10581]= -114682135;
assign addr[10582]= -76474970;
assign addr[10583]= -38243550;
assign addr[10584]= 0;
assign addr[10585]= 38243550;
assign addr[10586]= 76474970;
assign addr[10587]= 114682135;
assign addr[10588]= 152852926;
assign addr[10589]= 190975237;
assign addr[10590]= 229036977;
assign addr[10591]= 267026072;
assign addr[10592]= 304930476;
assign addr[10593]= 342738165;
assign addr[10594]= 380437148;
assign addr[10595]= 418015468;
assign addr[10596]= 455461206;
assign addr[10597]= 492762486;
assign addr[10598]= 529907477;
assign addr[10599]= 566884397;
assign addr[10600]= 603681519;
assign addr[10601]= 640287172;
assign addr[10602]= 676689746;
assign addr[10603]= 712877694;
assign addr[10604]= 748839539;
assign addr[10605]= 784563876;
assign addr[10606]= 820039373;
assign addr[10607]= 855254778;
assign addr[10608]= 890198924;
assign addr[10609]= 924860725;
assign addr[10610]= 959229189;
assign addr[10611]= 993293415;
assign addr[10612]= 1027042599;
assign addr[10613]= 1060466036;
assign addr[10614]= 1093553126;
assign addr[10615]= 1126293375;
assign addr[10616]= 1158676398;
assign addr[10617]= 1190691925;
assign addr[10618]= 1222329801;
assign addr[10619]= 1253579991;
assign addr[10620]= 1284432584;
assign addr[10621]= 1314877795;
assign addr[10622]= 1344905966;
assign addr[10623]= 1374507575;
assign addr[10624]= 1403673233;
assign addr[10625]= 1432393688;
assign addr[10626]= 1460659832;
assign addr[10627]= 1488462700;
assign addr[10628]= 1515793473;
assign addr[10629]= 1542643483;
assign addr[10630]= 1569004214;
assign addr[10631]= 1594867305;
assign addr[10632]= 1620224553;
assign addr[10633]= 1645067915;
assign addr[10634]= 1669389513;
assign addr[10635]= 1693181631;
assign addr[10636]= 1716436725;
assign addr[10637]= 1739147417;
assign addr[10638]= 1761306505;
assign addr[10639]= 1782906961;
assign addr[10640]= 1803941934;
assign addr[10641]= 1824404752;
assign addr[10642]= 1844288924;
assign addr[10643]= 1863588145;
assign addr[10644]= 1882296293;
assign addr[10645]= 1900407434;
assign addr[10646]= 1917915825;
assign addr[10647]= 1934815911;
assign addr[10648]= 1951102334;
assign addr[10649]= 1966769926;
assign addr[10650]= 1981813720;
assign addr[10651]= 1996228943;
assign addr[10652]= 2010011024;
assign addr[10653]= 2023155591;
assign addr[10654]= 2035658475;
assign addr[10655]= 2047515711;
assign addr[10656]= 2058723538;
assign addr[10657]= 2069278401;
assign addr[10658]= 2079176953;
assign addr[10659]= 2088416053;
assign addr[10660]= 2096992772;
assign addr[10661]= 2104904390;
assign addr[10662]= 2112148396;
assign addr[10663]= 2118722494;
assign addr[10664]= 2124624598;
assign addr[10665]= 2129852837;
assign addr[10666]= 2134405552;
assign addr[10667]= 2138281298;
assign addr[10668]= 2141478848;
assign addr[10669]= 2143997187;
assign addr[10670]= 2145835515;
assign addr[10671]= 2146993250;
assign addr[10672]= 2147470025;
assign addr[10673]= 2147265689;
assign addr[10674]= 2146380306;
assign addr[10675]= 2144814157;
assign addr[10676]= 2142567738;
assign addr[10677]= 2139641764;
assign addr[10678]= 2136037160;
assign addr[10679]= 2131755071;
assign addr[10680]= 2126796855;
assign addr[10681]= 2121164085;
assign addr[10682]= 2114858546;
assign addr[10683]= 2107882239;
assign addr[10684]= 2100237377;
assign addr[10685]= 2091926384;
assign addr[10686]= 2082951896;
assign addr[10687]= 2073316760;
assign addr[10688]= 2063024031;
assign addr[10689]= 2052076975;
assign addr[10690]= 2040479063;
assign addr[10691]= 2028233973;
assign addr[10692]= 2015345591;
assign addr[10693]= 2001818002;
assign addr[10694]= 1987655498;
assign addr[10695]= 1972862571;
assign addr[10696]= 1957443913;
assign addr[10697]= 1941404413;
assign addr[10698]= 1924749160;
assign addr[10699]= 1907483436;
assign addr[10700]= 1889612716;
assign addr[10701]= 1871142669;
assign addr[10702]= 1852079154;
assign addr[10703]= 1832428215;
assign addr[10704]= 1812196087;
assign addr[10705]= 1791389186;
assign addr[10706]= 1770014111;
assign addr[10707]= 1748077642;
assign addr[10708]= 1725586737;
assign addr[10709]= 1702548529;
assign addr[10710]= 1678970324;
assign addr[10711]= 1654859602;
assign addr[10712]= 1630224009;
assign addr[10713]= 1605071359;
assign addr[10714]= 1579409630;
assign addr[10715]= 1553246960;
assign addr[10716]= 1526591649;
assign addr[10717]= 1499452149;
assign addr[10718]= 1471837070;
assign addr[10719]= 1443755168;
assign addr[10720]= 1415215352;
assign addr[10721]= 1386226674;
assign addr[10722]= 1356798326;
assign addr[10723]= 1326939644;
assign addr[10724]= 1296660098;
assign addr[10725]= 1265969291;
assign addr[10726]= 1234876957;
assign addr[10727]= 1203392958;
assign addr[10728]= 1171527280;
assign addr[10729]= 1139290029;
assign addr[10730]= 1106691431;
assign addr[10731]= 1073741824;
assign addr[10732]= 1040451659;
assign addr[10733]= 1006831495;
assign addr[10734]= 972891995;
assign addr[10735]= 938643924;
assign addr[10736]= 904098143;
assign addr[10737]= 869265610;
assign addr[10738]= 834157373;
assign addr[10739]= 798784567;
assign addr[10740]= 763158411;
assign addr[10741]= 727290205;
assign addr[10742]= 691191324;
assign addr[10743]= 654873219;
assign addr[10744]= 618347408;
assign addr[10745]= 581625477;
assign addr[10746]= 544719071;
assign addr[10747]= 507639898;
assign addr[10748]= 470399716;
assign addr[10749]= 433010339;
assign addr[10750]= 395483624;
assign addr[10751]= 357831473;
assign addr[10752]= 320065829;
assign addr[10753]= 282198671;
assign addr[10754]= 244242007;
assign addr[10755]= 206207878;
assign addr[10756]= 168108346;
assign addr[10757]= 129955495;
assign addr[10758]= 91761426;
assign addr[10759]= 53538253;
assign addr[10760]= 15298099;
assign addr[10761]= -22946906;
assign addr[10762]= -61184634;
assign addr[10763]= -99402956;
assign addr[10764]= -137589750;
assign addr[10765]= -175732905;
assign addr[10766]= -213820322;
assign addr[10767]= -251839923;
assign addr[10768]= -289779648;
assign addr[10769]= -327627463;
assign addr[10770]= -365371365;
assign addr[10771]= -402999383;
assign addr[10772]= -440499581;
assign addr[10773]= -477860067;
assign addr[10774]= -515068990;
assign addr[10775]= -552114549;
assign addr[10776]= -588984994;
assign addr[10777]= -625668632;
assign addr[10778]= -662153826;
assign addr[10779]= -698429006;
assign addr[10780]= -734482665;
assign addr[10781]= -770303369;
assign addr[10782]= -805879757;
assign addr[10783]= -841200544;
assign addr[10784]= -876254528;
assign addr[10785]= -911030591;
assign addr[10786]= -945517704;
assign addr[10787]= -979704927;
assign addr[10788]= -1013581418;
assign addr[10789]= -1047136432;
assign addr[10790]= -1080359326;
assign addr[10791]= -1113239564;
assign addr[10792]= -1145766716;
assign addr[10793]= -1177930466;
assign addr[10794]= -1209720613;
assign addr[10795]= -1241127074;
assign addr[10796]= -1272139887;
assign addr[10797]= -1302749217;
assign addr[10798]= -1332945355;
assign addr[10799]= -1362718723;
assign addr[10800]= -1392059879;
assign addr[10801]= -1420959516;
assign addr[10802]= -1449408469;
assign addr[10803]= -1477397714;
assign addr[10804]= -1504918373;
assign addr[10805]= -1531961719;
assign addr[10806]= -1558519173;
assign addr[10807]= -1584582314;
assign addr[10808]= -1610142873;
assign addr[10809]= -1635192744;
assign addr[10810]= -1659723983;
assign addr[10811]= -1683728808;
assign addr[10812]= -1707199606;
assign addr[10813]= -1730128933;
assign addr[10814]= -1752509516;
assign addr[10815]= -1774334257;
assign addr[10816]= -1795596234;
assign addr[10817]= -1816288703;
assign addr[10818]= -1836405100;
assign addr[10819]= -1855939047;
assign addr[10820]= -1874884346;
assign addr[10821]= -1893234990;
assign addr[10822]= -1910985158;
assign addr[10823]= -1928129220;
assign addr[10824]= -1944661739;
assign addr[10825]= -1960577471;
assign addr[10826]= -1975871368;
assign addr[10827]= -1990538579;
assign addr[10828]= -2004574453;
assign addr[10829]= -2017974537;
assign addr[10830]= -2030734582;
assign addr[10831]= -2042850540;
assign addr[10832]= -2054318569;
assign addr[10833]= -2065135031;
assign addr[10834]= -2075296495;
assign addr[10835]= -2084799740;
assign addr[10836]= -2093641749;
assign addr[10837]= -2101819720;
assign addr[10838]= -2109331059;
assign addr[10839]= -2116173382;
assign addr[10840]= -2122344521;
assign addr[10841]= -2127842516;
assign addr[10842]= -2132665626;
assign addr[10843]= -2136812319;
assign addr[10844]= -2140281282;
assign addr[10845]= -2143071413;
assign addr[10846]= -2145181827;
assign addr[10847]= -2146611856;
assign addr[10848]= -2147361045;
assign addr[10849]= -2147429158;
assign addr[10850]= -2146816171;
assign addr[10851]= -2145522281;
assign addr[10852]= -2143547897;
assign addr[10853]= -2140893646;
assign addr[10854]= -2137560369;
assign addr[10855]= -2133549123;
assign addr[10856]= -2128861181;
assign addr[10857]= -2123498030;
assign addr[10858]= -2117461370;
assign addr[10859]= -2110753117;
assign addr[10860]= -2103375398;
assign addr[10861]= -2095330553;
assign addr[10862]= -2086621133;
assign addr[10863]= -2077249901;
assign addr[10864]= -2067219829;
assign addr[10865]= -2056534099;
assign addr[10866]= -2045196100;
assign addr[10867]= -2033209426;
assign addr[10868]= -2020577882;
assign addr[10869]= -2007305472;
assign addr[10870]= -1993396407;
assign addr[10871]= -1978855097;
assign addr[10872]= -1963686155;
assign addr[10873]= -1947894393;
assign addr[10874]= -1931484818;
assign addr[10875]= -1914462636;
assign addr[10876]= -1896833245;
assign addr[10877]= -1878602237;
assign addr[10878]= -1859775393;
assign addr[10879]= -1840358687;
assign addr[10880]= -1820358275;
assign addr[10881]= -1799780501;
assign addr[10882]= -1778631892;
assign addr[10883]= -1756919156;
assign addr[10884]= -1734649179;
assign addr[10885]= -1711829025;
assign addr[10886]= -1688465931;
assign addr[10887]= -1664567307;
assign addr[10888]= -1640140734;
assign addr[10889]= -1615193959;
assign addr[10890]= -1589734894;
assign addr[10891]= -1563771613;
assign addr[10892]= -1537312353;
assign addr[10893]= -1510365504;
assign addr[10894]= -1482939614;
assign addr[10895]= -1455043381;
assign addr[10896]= -1426685652;
assign addr[10897]= -1397875423;
assign addr[10898]= -1368621831;
assign addr[10899]= -1338934154;
assign addr[10900]= -1308821808;
assign addr[10901]= -1278294345;
assign addr[10902]= -1247361445;
assign addr[10903]= -1216032921;
assign addr[10904]= -1184318708;
assign addr[10905]= -1152228866;
assign addr[10906]= -1119773573;
assign addr[10907]= -1086963121;
assign addr[10908]= -1053807919;
assign addr[10909]= -1020318481;
assign addr[10910]= -986505429;
assign addr[10911]= -952379488;
assign addr[10912]= -917951481;
assign addr[10913]= -883232329;
assign addr[10914]= -848233042;
assign addr[10915]= -812964722;
assign addr[10916]= -777438554;
assign addr[10917]= -741665807;
assign addr[10918]= -705657826;
assign addr[10919]= -669426032;
assign addr[10920]= -632981917;
assign addr[10921]= -596337040;
assign addr[10922]= -559503022;
assign addr[10923]= -522491548;
assign addr[10924]= -485314355;
assign addr[10925]= -447983235;
assign addr[10926]= -410510029;
assign addr[10927]= -372906622;
assign addr[10928]= -335184940;
assign addr[10929]= -297356948;
assign addr[10930]= -259434643;
assign addr[10931]= -221430054;
assign addr[10932]= -183355234;
assign addr[10933]= -145222259;
assign addr[10934]= -107043224;
assign addr[10935]= -68830239;
assign addr[10936]= -30595422;
assign addr[10937]= 7649098;
assign addr[10938]= 45891193;
assign addr[10939]= 84118732;
assign addr[10940]= 122319591;
assign addr[10941]= 160481654;
assign addr[10942]= 198592817;
assign addr[10943]= 236640993;
assign addr[10944]= 274614114;
assign addr[10945]= 312500135;
assign addr[10946]= 350287041;
assign addr[10947]= 387962847;
assign addr[10948]= 425515602;
assign addr[10949]= 462933398;
assign addr[10950]= 500204365;
assign addr[10951]= 537316682;
assign addr[10952]= 574258580;
assign addr[10953]= 611018340;
assign addr[10954]= 647584304;
assign addr[10955]= 683944874;
assign addr[10956]= 720088517;
assign addr[10957]= 756003771;
assign addr[10958]= 791679244;
assign addr[10959]= 827103620;
assign addr[10960]= 862265664;
assign addr[10961]= 897154224;
assign addr[10962]= 931758235;
assign addr[10963]= 966066720;
assign addr[10964]= 1000068799;
assign addr[10965]= 1033753687;
assign addr[10966]= 1067110699;
assign addr[10967]= 1100129257;
assign addr[10968]= 1132798888;
assign addr[10969]= 1165109230;
assign addr[10970]= 1197050035;
assign addr[10971]= 1228611172;
assign addr[10972]= 1259782632;
assign addr[10973]= 1290554528;
assign addr[10974]= 1320917099;
assign addr[10975]= 1350860716;
assign addr[10976]= 1380375881;
assign addr[10977]= 1409453233;
assign addr[10978]= 1438083551;
assign addr[10979]= 1466257752;
assign addr[10980]= 1493966902;
assign addr[10981]= 1521202211;
assign addr[10982]= 1547955041;
assign addr[10983]= 1574216908;
assign addr[10984]= 1599979481;
assign addr[10985]= 1625234591;
assign addr[10986]= 1649974225;
assign addr[10987]= 1674190539;
assign addr[10988]= 1697875851;
assign addr[10989]= 1721022648;
assign addr[10990]= 1743623590;
assign addr[10991]= 1765671509;
assign addr[10992]= 1787159411;
assign addr[10993]= 1808080480;
assign addr[10994]= 1828428082;
assign addr[10995]= 1848195763;
assign addr[10996]= 1867377253;
assign addr[10997]= 1885966468;
assign addr[10998]= 1903957513;
assign addr[10999]= 1921344681;
assign addr[11000]= 1938122457;
assign addr[11001]= 1954285520;
assign addr[11002]= 1969828744;
assign addr[11003]= 1984747199;
assign addr[11004]= 1999036154;
assign addr[11005]= 2012691075;
assign addr[11006]= 2025707632;
assign addr[11007]= 2038081698;
assign addr[11008]= 2049809346;
assign addr[11009]= 2060886858;
assign addr[11010]= 2071310720;
assign addr[11011]= 2081077626;
assign addr[11012]= 2090184478;
assign addr[11013]= 2098628387;
assign addr[11014]= 2106406677;
assign addr[11015]= 2113516878;
assign addr[11016]= 2119956737;
assign addr[11017]= 2125724211;
assign addr[11018]= 2130817471;
assign addr[11019]= 2135234901;
assign addr[11020]= 2138975100;
assign addr[11021]= 2142036881;
assign addr[11022]= 2144419275;
assign addr[11023]= 2146121524;
assign addr[11024]= 2147143090;
assign addr[11025]= 2147483648;
assign addr[11026]= 2147143090;
assign addr[11027]= 2146121524;
assign addr[11028]= 2144419275;
assign addr[11029]= 2142036881;
assign addr[11030]= 2138975100;
assign addr[11031]= 2135234901;
assign addr[11032]= 2130817471;
assign addr[11033]= 2125724211;
assign addr[11034]= 2119956737;
assign addr[11035]= 2113516878;
assign addr[11036]= 2106406677;
assign addr[11037]= 2098628387;
assign addr[11038]= 2090184478;
assign addr[11039]= 2081077626;
assign addr[11040]= 2071310720;
assign addr[11041]= 2060886858;
assign addr[11042]= 2049809346;
assign addr[11043]= 2038081698;
assign addr[11044]= 2025707632;
assign addr[11045]= 2012691075;
assign addr[11046]= 1999036154;
assign addr[11047]= 1984747199;
assign addr[11048]= 1969828744;
assign addr[11049]= 1954285520;
assign addr[11050]= 1938122457;
assign addr[11051]= 1921344681;
assign addr[11052]= 1903957513;
assign addr[11053]= 1885966468;
assign addr[11054]= 1867377253;
assign addr[11055]= 1848195763;
assign addr[11056]= 1828428082;
assign addr[11057]= 1808080480;
assign addr[11058]= 1787159411;
assign addr[11059]= 1765671509;
assign addr[11060]= 1743623590;
assign addr[11061]= 1721022648;
assign addr[11062]= 1697875851;
assign addr[11063]= 1674190539;
assign addr[11064]= 1649974225;
assign addr[11065]= 1625234591;
assign addr[11066]= 1599979481;
assign addr[11067]= 1574216908;
assign addr[11068]= 1547955041;
assign addr[11069]= 1521202211;
assign addr[11070]= 1493966902;
assign addr[11071]= 1466257752;
assign addr[11072]= 1438083551;
assign addr[11073]= 1409453233;
assign addr[11074]= 1380375881;
assign addr[11075]= 1350860716;
assign addr[11076]= 1320917099;
assign addr[11077]= 1290554528;
assign addr[11078]= 1259782632;
assign addr[11079]= 1228611172;
assign addr[11080]= 1197050035;
assign addr[11081]= 1165109230;
assign addr[11082]= 1132798888;
assign addr[11083]= 1100129257;
assign addr[11084]= 1067110699;
assign addr[11085]= 1033753687;
assign addr[11086]= 1000068799;
assign addr[11087]= 966066720;
assign addr[11088]= 931758235;
assign addr[11089]= 897154224;
assign addr[11090]= 862265664;
assign addr[11091]= 827103620;
assign addr[11092]= 791679244;
assign addr[11093]= 756003771;
assign addr[11094]= 720088517;
assign addr[11095]= 683944874;
assign addr[11096]= 647584304;
assign addr[11097]= 611018340;
assign addr[11098]= 574258580;
assign addr[11099]= 537316682;
assign addr[11100]= 500204365;
assign addr[11101]= 462933398;
assign addr[11102]= 425515602;
assign addr[11103]= 387962847;
assign addr[11104]= 350287041;
assign addr[11105]= 312500135;
assign addr[11106]= 274614114;
assign addr[11107]= 236640993;
assign addr[11108]= 198592817;
assign addr[11109]= 160481654;
assign addr[11110]= 122319591;
assign addr[11111]= 84118732;
assign addr[11112]= 45891193;
assign addr[11113]= 7649098;
assign addr[11114]= -30595422;
assign addr[11115]= -68830239;
assign addr[11116]= -107043224;
assign addr[11117]= -145222259;
assign addr[11118]= -183355234;
assign addr[11119]= -221430054;
assign addr[11120]= -259434643;
assign addr[11121]= -297356948;
assign addr[11122]= -335184940;
assign addr[11123]= -372906622;
assign addr[11124]= -410510029;
assign addr[11125]= -447983235;
assign addr[11126]= -485314355;
assign addr[11127]= -522491548;
assign addr[11128]= -559503022;
assign addr[11129]= -596337040;
assign addr[11130]= -632981917;
assign addr[11131]= -669426032;
assign addr[11132]= -705657826;
assign addr[11133]= -741665807;
assign addr[11134]= -777438554;
assign addr[11135]= -812964722;
assign addr[11136]= -848233042;
assign addr[11137]= -883232329;
assign addr[11138]= -917951481;
assign addr[11139]= -952379488;
assign addr[11140]= -986505429;
assign addr[11141]= -1020318481;
assign addr[11142]= -1053807919;
assign addr[11143]= -1086963121;
assign addr[11144]= -1119773573;
assign addr[11145]= -1152228866;
assign addr[11146]= -1184318708;
assign addr[11147]= -1216032921;
assign addr[11148]= -1247361445;
assign addr[11149]= -1278294345;
assign addr[11150]= -1308821808;
assign addr[11151]= -1338934154;
assign addr[11152]= -1368621831;
assign addr[11153]= -1397875423;
assign addr[11154]= -1426685652;
assign addr[11155]= -1455043381;
assign addr[11156]= -1482939614;
assign addr[11157]= -1510365504;
assign addr[11158]= -1537312353;
assign addr[11159]= -1563771613;
assign addr[11160]= -1589734894;
assign addr[11161]= -1615193959;
assign addr[11162]= -1640140734;
assign addr[11163]= -1664567307;
assign addr[11164]= -1688465931;
assign addr[11165]= -1711829025;
assign addr[11166]= -1734649179;
assign addr[11167]= -1756919156;
assign addr[11168]= -1778631892;
assign addr[11169]= -1799780501;
assign addr[11170]= -1820358275;
assign addr[11171]= -1840358687;
assign addr[11172]= -1859775393;
assign addr[11173]= -1878602237;
assign addr[11174]= -1896833245;
assign addr[11175]= -1914462636;
assign addr[11176]= -1931484818;
assign addr[11177]= -1947894393;
assign addr[11178]= -1963686155;
assign addr[11179]= -1978855097;
assign addr[11180]= -1993396407;
assign addr[11181]= -2007305472;
assign addr[11182]= -2020577882;
assign addr[11183]= -2033209426;
assign addr[11184]= -2045196100;
assign addr[11185]= -2056534099;
assign addr[11186]= -2067219829;
assign addr[11187]= -2077249901;
assign addr[11188]= -2086621133;
assign addr[11189]= -2095330553;
assign addr[11190]= -2103375398;
assign addr[11191]= -2110753117;
assign addr[11192]= -2117461370;
assign addr[11193]= -2123498030;
assign addr[11194]= -2128861181;
assign addr[11195]= -2133549123;
assign addr[11196]= -2137560369;
assign addr[11197]= -2140893646;
assign addr[11198]= -2143547897;
assign addr[11199]= -2145522281;
assign addr[11200]= -2146816171;
assign addr[11201]= -2147429158;
assign addr[11202]= -2147361045;
assign addr[11203]= -2146611856;
assign addr[11204]= -2145181827;
assign addr[11205]= -2143071413;
assign addr[11206]= -2140281282;
assign addr[11207]= -2136812319;
assign addr[11208]= -2132665626;
assign addr[11209]= -2127842516;
assign addr[11210]= -2122344521;
assign addr[11211]= -2116173382;
assign addr[11212]= -2109331059;
assign addr[11213]= -2101819720;
assign addr[11214]= -2093641749;
assign addr[11215]= -2084799740;
assign addr[11216]= -2075296495;
assign addr[11217]= -2065135031;
assign addr[11218]= -2054318569;
assign addr[11219]= -2042850540;
assign addr[11220]= -2030734582;
assign addr[11221]= -2017974537;
assign addr[11222]= -2004574453;
assign addr[11223]= -1990538579;
assign addr[11224]= -1975871368;
assign addr[11225]= -1960577471;
assign addr[11226]= -1944661739;
assign addr[11227]= -1928129220;
assign addr[11228]= -1910985158;
assign addr[11229]= -1893234990;
assign addr[11230]= -1874884346;
assign addr[11231]= -1855939047;
assign addr[11232]= -1836405100;
assign addr[11233]= -1816288703;
assign addr[11234]= -1795596234;
assign addr[11235]= -1774334257;
assign addr[11236]= -1752509516;
assign addr[11237]= -1730128933;
assign addr[11238]= -1707199606;
assign addr[11239]= -1683728808;
assign addr[11240]= -1659723983;
assign addr[11241]= -1635192744;
assign addr[11242]= -1610142873;
assign addr[11243]= -1584582314;
assign addr[11244]= -1558519173;
assign addr[11245]= -1531961719;
assign addr[11246]= -1504918373;
assign addr[11247]= -1477397714;
assign addr[11248]= -1449408469;
assign addr[11249]= -1420959516;
assign addr[11250]= -1392059879;
assign addr[11251]= -1362718723;
assign addr[11252]= -1332945355;
assign addr[11253]= -1302749217;
assign addr[11254]= -1272139887;
assign addr[11255]= -1241127074;
assign addr[11256]= -1209720613;
assign addr[11257]= -1177930466;
assign addr[11258]= -1145766716;
assign addr[11259]= -1113239564;
assign addr[11260]= -1080359326;
assign addr[11261]= -1047136432;
assign addr[11262]= -1013581418;
assign addr[11263]= -979704927;
assign addr[11264]= -945517704;
assign addr[11265]= -911030591;
assign addr[11266]= -876254528;
assign addr[11267]= -841200544;
assign addr[11268]= -805879757;
assign addr[11269]= -770303369;
assign addr[11270]= -734482665;
assign addr[11271]= -698429006;
assign addr[11272]= -662153826;
assign addr[11273]= -625668632;
assign addr[11274]= -588984994;
assign addr[11275]= -552114549;
assign addr[11276]= -515068990;
assign addr[11277]= -477860067;
assign addr[11278]= -440499581;
assign addr[11279]= -402999383;
assign addr[11280]= -365371365;
assign addr[11281]= -327627463;
assign addr[11282]= -289779648;
assign addr[11283]= -251839923;
assign addr[11284]= -213820322;
assign addr[11285]= -175732905;
assign addr[11286]= -137589750;
assign addr[11287]= -99402956;
assign addr[11288]= -61184634;
assign addr[11289]= -22946906;
assign addr[11290]= 15298099;
assign addr[11291]= 53538253;
assign addr[11292]= 91761426;
assign addr[11293]= 129955495;
assign addr[11294]= 168108346;
assign addr[11295]= 206207878;
assign addr[11296]= 244242007;
assign addr[11297]= 282198671;
assign addr[11298]= 320065829;
assign addr[11299]= 357831473;
assign addr[11300]= 395483624;
assign addr[11301]= 433010339;
assign addr[11302]= 470399716;
assign addr[11303]= 507639898;
assign addr[11304]= 544719071;
assign addr[11305]= 581625477;
assign addr[11306]= 618347408;
assign addr[11307]= 654873219;
assign addr[11308]= 691191324;
assign addr[11309]= 727290205;
assign addr[11310]= 763158411;
assign addr[11311]= 798784567;
assign addr[11312]= 834157373;
assign addr[11313]= 869265610;
assign addr[11314]= 904098143;
assign addr[11315]= 938643924;
assign addr[11316]= 972891995;
assign addr[11317]= 1006831495;
assign addr[11318]= 1040451659;
assign addr[11319]= 1073741824;
assign addr[11320]= 1106691431;
assign addr[11321]= 1139290029;
assign addr[11322]= 1171527280;
assign addr[11323]= 1203392958;
assign addr[11324]= 1234876957;
assign addr[11325]= 1265969291;
assign addr[11326]= 1296660098;
assign addr[11327]= 1326939644;
assign addr[11328]= 1356798326;
assign addr[11329]= 1386226674;
assign addr[11330]= 1415215352;
assign addr[11331]= 1443755168;
assign addr[11332]= 1471837070;
assign addr[11333]= 1499452149;
assign addr[11334]= 1526591649;
assign addr[11335]= 1553246960;
assign addr[11336]= 1579409630;
assign addr[11337]= 1605071359;
assign addr[11338]= 1630224009;
assign addr[11339]= 1654859602;
assign addr[11340]= 1678970324;
assign addr[11341]= 1702548529;
assign addr[11342]= 1725586737;
assign addr[11343]= 1748077642;
assign addr[11344]= 1770014111;
assign addr[11345]= 1791389186;
assign addr[11346]= 1812196087;
assign addr[11347]= 1832428215;
assign addr[11348]= 1852079154;
assign addr[11349]= 1871142669;
assign addr[11350]= 1889612716;
assign addr[11351]= 1907483436;
assign addr[11352]= 1924749160;
assign addr[11353]= 1941404413;
assign addr[11354]= 1957443913;
assign addr[11355]= 1972862571;
assign addr[11356]= 1987655498;
assign addr[11357]= 2001818002;
assign addr[11358]= 2015345591;
assign addr[11359]= 2028233973;
assign addr[11360]= 2040479063;
assign addr[11361]= 2052076975;
assign addr[11362]= 2063024031;
assign addr[11363]= 2073316760;
assign addr[11364]= 2082951896;
assign addr[11365]= 2091926384;
assign addr[11366]= 2100237377;
assign addr[11367]= 2107882239;
assign addr[11368]= 2114858546;
assign addr[11369]= 2121164085;
assign addr[11370]= 2126796855;
assign addr[11371]= 2131755071;
assign addr[11372]= 2136037160;
assign addr[11373]= 2139641764;
assign addr[11374]= 2142567738;
assign addr[11375]= 2144814157;
assign addr[11376]= 2146380306;
assign addr[11377]= 2147265689;
assign addr[11378]= 2147470025;
assign addr[11379]= 2146993250;
assign addr[11380]= 2145835515;
assign addr[11381]= 2143997187;
assign addr[11382]= 2141478848;
assign addr[11383]= 2138281298;
assign addr[11384]= 2134405552;
assign addr[11385]= 2129852837;
assign addr[11386]= 2124624598;
assign addr[11387]= 2118722494;
assign addr[11388]= 2112148396;
assign addr[11389]= 2104904390;
assign addr[11390]= 2096992772;
assign addr[11391]= 2088416053;
assign addr[11392]= 2079176953;
assign addr[11393]= 2069278401;
assign addr[11394]= 2058723538;
assign addr[11395]= 2047515711;
assign addr[11396]= 2035658475;
assign addr[11397]= 2023155591;
assign addr[11398]= 2010011024;
assign addr[11399]= 1996228943;
assign addr[11400]= 1981813720;
assign addr[11401]= 1966769926;
assign addr[11402]= 1951102334;
assign addr[11403]= 1934815911;
assign addr[11404]= 1917915825;
assign addr[11405]= 1900407434;
assign addr[11406]= 1882296293;
assign addr[11407]= 1863588145;
assign addr[11408]= 1844288924;
assign addr[11409]= 1824404752;
assign addr[11410]= 1803941934;
assign addr[11411]= 1782906961;
assign addr[11412]= 1761306505;
assign addr[11413]= 1739147417;
assign addr[11414]= 1716436725;
assign addr[11415]= 1693181631;
assign addr[11416]= 1669389513;
assign addr[11417]= 1645067915;
assign addr[11418]= 1620224553;
assign addr[11419]= 1594867305;
assign addr[11420]= 1569004214;
assign addr[11421]= 1542643483;
assign addr[11422]= 1515793473;
assign addr[11423]= 1488462700;
assign addr[11424]= 1460659832;
assign addr[11425]= 1432393688;
assign addr[11426]= 1403673233;
assign addr[11427]= 1374507575;
assign addr[11428]= 1344905966;
assign addr[11429]= 1314877795;
assign addr[11430]= 1284432584;
assign addr[11431]= 1253579991;
assign addr[11432]= 1222329801;
assign addr[11433]= 1190691925;
assign addr[11434]= 1158676398;
assign addr[11435]= 1126293375;
assign addr[11436]= 1093553126;
assign addr[11437]= 1060466036;
assign addr[11438]= 1027042599;
assign addr[11439]= 993293415;
assign addr[11440]= 959229189;
assign addr[11441]= 924860725;
assign addr[11442]= 890198924;
assign addr[11443]= 855254778;
assign addr[11444]= 820039373;
assign addr[11445]= 784563876;
assign addr[11446]= 748839539;
assign addr[11447]= 712877694;
assign addr[11448]= 676689746;
assign addr[11449]= 640287172;
assign addr[11450]= 603681519;
assign addr[11451]= 566884397;
assign addr[11452]= 529907477;
assign addr[11453]= 492762486;
assign addr[11454]= 455461206;
assign addr[11455]= 418015468;
assign addr[11456]= 380437148;
assign addr[11457]= 342738165;
assign addr[11458]= 304930476;
assign addr[11459]= 267026072;
assign addr[11460]= 229036977;
assign addr[11461]= 190975237;
assign addr[11462]= 152852926;
assign addr[11463]= 114682135;
assign addr[11464]= 76474970;
assign addr[11465]= 38243550;
assign addr[11466]= 0;
assign addr[11467]= -38243550;
assign addr[11468]= -76474970;
assign addr[11469]= -114682135;
assign addr[11470]= -152852926;
assign addr[11471]= -190975237;
assign addr[11472]= -229036977;
assign addr[11473]= -267026072;
assign addr[11474]= -304930476;
assign addr[11475]= -342738165;
assign addr[11476]= -380437148;
assign addr[11477]= -418015468;
assign addr[11478]= -455461206;
assign addr[11479]= -492762486;
assign addr[11480]= -529907477;
assign addr[11481]= -566884397;
assign addr[11482]= -603681519;
assign addr[11483]= -640287172;
assign addr[11484]= -676689746;
assign addr[11485]= -712877694;
assign addr[11486]= -748839539;
assign addr[11487]= -784563876;
assign addr[11488]= -820039373;
assign addr[11489]= -855254778;
assign addr[11490]= -890198924;
assign addr[11491]= -924860725;
assign addr[11492]= -959229189;
assign addr[11493]= -993293415;
assign addr[11494]= -1027042599;
assign addr[11495]= -1060466036;
assign addr[11496]= -1093553126;
assign addr[11497]= -1126293375;
assign addr[11498]= -1158676398;
assign addr[11499]= -1190691925;
assign addr[11500]= -1222329801;
assign addr[11501]= -1253579991;
assign addr[11502]= -1284432584;
assign addr[11503]= -1314877795;
assign addr[11504]= -1344905966;
assign addr[11505]= -1374507575;
assign addr[11506]= -1403673233;
assign addr[11507]= -1432393688;
assign addr[11508]= -1460659832;
assign addr[11509]= -1488462700;
assign addr[11510]= -1515793473;
assign addr[11511]= -1542643483;
assign addr[11512]= -1569004214;
assign addr[11513]= -1594867305;
assign addr[11514]= -1620224553;
assign addr[11515]= -1645067915;
assign addr[11516]= -1669389513;
assign addr[11517]= -1693181631;
assign addr[11518]= -1716436725;
assign addr[11519]= -1739147417;
assign addr[11520]= -1761306505;
assign addr[11521]= -1782906961;
assign addr[11522]= -1803941934;
assign addr[11523]= -1824404752;
assign addr[11524]= -1844288924;
assign addr[11525]= -1863588145;
assign addr[11526]= -1882296293;
assign addr[11527]= -1900407434;
assign addr[11528]= -1917915825;
assign addr[11529]= -1934815911;
assign addr[11530]= -1951102334;
assign addr[11531]= -1966769926;
assign addr[11532]= -1981813720;
assign addr[11533]= -1996228943;
assign addr[11534]= -2010011024;
assign addr[11535]= -2023155591;
assign addr[11536]= -2035658475;
assign addr[11537]= -2047515711;
assign addr[11538]= -2058723538;
assign addr[11539]= -2069278401;
assign addr[11540]= -2079176953;
assign addr[11541]= -2088416053;
assign addr[11542]= -2096992772;
assign addr[11543]= -2104904390;
assign addr[11544]= -2112148396;
assign addr[11545]= -2118722494;
assign addr[11546]= -2124624598;
assign addr[11547]= -2129852837;
assign addr[11548]= -2134405552;
assign addr[11549]= -2138281298;
assign addr[11550]= -2141478848;
assign addr[11551]= -2143997187;
assign addr[11552]= -2145835515;
assign addr[11553]= -2146993250;
assign addr[11554]= -2147470025;
assign addr[11555]= -2147265689;
assign addr[11556]= -2146380306;
assign addr[11557]= -2144814157;
assign addr[11558]= -2142567738;
assign addr[11559]= -2139641764;
assign addr[11560]= -2136037160;
assign addr[11561]= -2131755071;
assign addr[11562]= -2126796855;
assign addr[11563]= -2121164085;
assign addr[11564]= -2114858546;
assign addr[11565]= -2107882239;
assign addr[11566]= -2100237377;
assign addr[11567]= -2091926384;
assign addr[11568]= -2082951896;
assign addr[11569]= -2073316760;
assign addr[11570]= -2063024031;
assign addr[11571]= -2052076975;
assign addr[11572]= -2040479063;
assign addr[11573]= -2028233973;
assign addr[11574]= -2015345591;
assign addr[11575]= -2001818002;
assign addr[11576]= -1987655498;
assign addr[11577]= -1972862571;
assign addr[11578]= -1957443913;
assign addr[11579]= -1941404413;
assign addr[11580]= -1924749160;
assign addr[11581]= -1907483436;
assign addr[11582]= -1889612716;
assign addr[11583]= -1871142669;
assign addr[11584]= -1852079154;
assign addr[11585]= -1832428215;
assign addr[11586]= -1812196087;
assign addr[11587]= -1791389186;
assign addr[11588]= -1770014111;
assign addr[11589]= -1748077642;
assign addr[11590]= -1725586737;
assign addr[11591]= -1702548529;
assign addr[11592]= -1678970324;
assign addr[11593]= -1654859602;
assign addr[11594]= -1630224009;
assign addr[11595]= -1605071359;
assign addr[11596]= -1579409630;
assign addr[11597]= -1553246960;
assign addr[11598]= -1526591649;
assign addr[11599]= -1499452149;
assign addr[11600]= -1471837070;
assign addr[11601]= -1443755168;
assign addr[11602]= -1415215352;
assign addr[11603]= -1386226674;
assign addr[11604]= -1356798326;
assign addr[11605]= -1326939644;
assign addr[11606]= -1296660098;
assign addr[11607]= -1265969291;
assign addr[11608]= -1234876957;
assign addr[11609]= -1203392958;
assign addr[11610]= -1171527280;
assign addr[11611]= -1139290029;
assign addr[11612]= -1106691431;
assign addr[11613]= -1073741824;
assign addr[11614]= -1040451659;
assign addr[11615]= -1006831495;
assign addr[11616]= -972891995;
assign addr[11617]= -938643924;
assign addr[11618]= -904098143;
assign addr[11619]= -869265610;
assign addr[11620]= -834157373;
assign addr[11621]= -798784567;
assign addr[11622]= -763158411;
assign addr[11623]= -727290205;
assign addr[11624]= -691191324;
assign addr[11625]= -654873219;
assign addr[11626]= -618347408;
assign addr[11627]= -581625477;
assign addr[11628]= -544719071;
assign addr[11629]= -507639898;
assign addr[11630]= -470399716;
assign addr[11631]= -433010339;
assign addr[11632]= -395483624;
assign addr[11633]= -357831473;
assign addr[11634]= -320065829;
assign addr[11635]= -282198671;
assign addr[11636]= -244242007;
assign addr[11637]= -206207878;
assign addr[11638]= -168108346;
assign addr[11639]= -129955495;
assign addr[11640]= -91761426;
assign addr[11641]= -53538253;
assign addr[11642]= -15298099;
assign addr[11643]= 22946906;
assign addr[11644]= 61184634;
assign addr[11645]= 99402956;
assign addr[11646]= 137589750;
assign addr[11647]= 175732905;
assign addr[11648]= 213820322;
assign addr[11649]= 251839923;
assign addr[11650]= 289779648;
assign addr[11651]= 327627463;
assign addr[11652]= 365371365;
assign addr[11653]= 402999383;
assign addr[11654]= 440499581;
assign addr[11655]= 477860067;
assign addr[11656]= 515068990;
assign addr[11657]= 552114549;
assign addr[11658]= 588984994;
assign addr[11659]= 625668632;
assign addr[11660]= 662153826;
assign addr[11661]= 698429006;
assign addr[11662]= 734482665;
assign addr[11663]= 770303369;
assign addr[11664]= 805879757;
assign addr[11665]= 841200544;
assign addr[11666]= 876254528;
assign addr[11667]= 911030591;
assign addr[11668]= 945517704;
assign addr[11669]= 979704927;
assign addr[11670]= 1013581418;
assign addr[11671]= 1047136432;
assign addr[11672]= 1080359326;
assign addr[11673]= 1113239564;
assign addr[11674]= 1145766716;
assign addr[11675]= 1177930466;
assign addr[11676]= 1209720613;
assign addr[11677]= 1241127074;
assign addr[11678]= 1272139887;
assign addr[11679]= 1302749217;
assign addr[11680]= 1332945355;
assign addr[11681]= 1362718723;
assign addr[11682]= 1392059879;
assign addr[11683]= 1420959516;
assign addr[11684]= 1449408469;
assign addr[11685]= 1477397714;
assign addr[11686]= 1504918373;
assign addr[11687]= 1531961719;
assign addr[11688]= 1558519173;
assign addr[11689]= 1584582314;
assign addr[11690]= 1610142873;
assign addr[11691]= 1635192744;
assign addr[11692]= 1659723983;
assign addr[11693]= 1683728808;
assign addr[11694]= 1707199606;
assign addr[11695]= 1730128933;
assign addr[11696]= 1752509516;
assign addr[11697]= 1774334257;
assign addr[11698]= 1795596234;
assign addr[11699]= 1816288703;
assign addr[11700]= 1836405100;
assign addr[11701]= 1855939047;
assign addr[11702]= 1874884346;
assign addr[11703]= 1893234990;
assign addr[11704]= 1910985158;
assign addr[11705]= 1928129220;
assign addr[11706]= 1944661739;
assign addr[11707]= 1960577471;
assign addr[11708]= 1975871368;
assign addr[11709]= 1990538579;
assign addr[11710]= 2004574453;
assign addr[11711]= 2017974537;
assign addr[11712]= 2030734582;
assign addr[11713]= 2042850540;
assign addr[11714]= 2054318569;
assign addr[11715]= 2065135031;
assign addr[11716]= 2075296495;
assign addr[11717]= 2084799740;
assign addr[11718]= 2093641749;
assign addr[11719]= 2101819720;
assign addr[11720]= 2109331059;
assign addr[11721]= 2116173382;
assign addr[11722]= 2122344521;
assign addr[11723]= 2127842516;
assign addr[11724]= 2132665626;
assign addr[11725]= 2136812319;
assign addr[11726]= 2140281282;
assign addr[11727]= 2143071413;
assign addr[11728]= 2145181827;
assign addr[11729]= 2146611856;
assign addr[11730]= 2147361045;
assign addr[11731]= 2147429158;
assign addr[11732]= 2146816171;
assign addr[11733]= 2145522281;
assign addr[11734]= 2143547897;
assign addr[11735]= 2140893646;
assign addr[11736]= 2137560369;
assign addr[11737]= 2133549123;
assign addr[11738]= 2128861181;
assign addr[11739]= 2123498030;
assign addr[11740]= 2117461370;
assign addr[11741]= 2110753117;
assign addr[11742]= 2103375398;
assign addr[11743]= 2095330553;
assign addr[11744]= 2086621133;
assign addr[11745]= 2077249901;
assign addr[11746]= 2067219829;
assign addr[11747]= 2056534099;
assign addr[11748]= 2045196100;
assign addr[11749]= 2033209426;
assign addr[11750]= 2020577882;
assign addr[11751]= 2007305472;
assign addr[11752]= 1993396407;
assign addr[11753]= 1978855097;
assign addr[11754]= 1963686155;
assign addr[11755]= 1947894393;
assign addr[11756]= 1931484818;
assign addr[11757]= 1914462636;
assign addr[11758]= 1896833245;
assign addr[11759]= 1878602237;
assign addr[11760]= 1859775393;
assign addr[11761]= 1840358687;
assign addr[11762]= 1820358275;
assign addr[11763]= 1799780501;
assign addr[11764]= 1778631892;
assign addr[11765]= 1756919156;
assign addr[11766]= 1734649179;
assign addr[11767]= 1711829025;
assign addr[11768]= 1688465931;
assign addr[11769]= 1664567307;
assign addr[11770]= 1640140734;
assign addr[11771]= 1615193959;
assign addr[11772]= 1589734894;
assign addr[11773]= 1563771613;
assign addr[11774]= 1537312353;
assign addr[11775]= 1510365504;
assign addr[11776]= 1482939614;
assign addr[11777]= 1455043381;
assign addr[11778]= 1426685652;
assign addr[11779]= 1397875423;
assign addr[11780]= 1368621831;
assign addr[11781]= 1338934154;
assign addr[11782]= 1308821808;
assign addr[11783]= 1278294345;
assign addr[11784]= 1247361445;
assign addr[11785]= 1216032921;
assign addr[11786]= 1184318708;
assign addr[11787]= 1152228866;
assign addr[11788]= 1119773573;
assign addr[11789]= 1086963121;
assign addr[11790]= 1053807919;
assign addr[11791]= 1020318481;
assign addr[11792]= 986505429;
assign addr[11793]= 952379488;
assign addr[11794]= 917951481;
assign addr[11795]= 883232329;
assign addr[11796]= 848233042;
assign addr[11797]= 812964722;
assign addr[11798]= 777438554;
assign addr[11799]= 741665807;
assign addr[11800]= 705657826;
assign addr[11801]= 669426032;
assign addr[11802]= 632981917;
assign addr[11803]= 596337040;
assign addr[11804]= 559503022;
assign addr[11805]= 522491548;
assign addr[11806]= 485314355;
assign addr[11807]= 447983235;
assign addr[11808]= 410510029;
assign addr[11809]= 372906622;
assign addr[11810]= 335184940;
assign addr[11811]= 297356948;
assign addr[11812]= 259434643;
assign addr[11813]= 221430054;
assign addr[11814]= 183355234;
assign addr[11815]= 145222259;
assign addr[11816]= 107043224;
assign addr[11817]= 68830239;
assign addr[11818]= 30595422;
assign addr[11819]= -7649098;
assign addr[11820]= -45891193;
assign addr[11821]= -84118732;
assign addr[11822]= -122319591;
assign addr[11823]= -160481654;
assign addr[11824]= -198592817;
assign addr[11825]= -236640993;
assign addr[11826]= -274614114;
assign addr[11827]= -312500135;
assign addr[11828]= -350287041;
assign addr[11829]= -387962847;
assign addr[11830]= -425515602;
assign addr[11831]= -462933398;
assign addr[11832]= -500204365;
assign addr[11833]= -537316682;
assign addr[11834]= -574258580;
assign addr[11835]= -611018340;
assign addr[11836]= -647584304;
assign addr[11837]= -683944874;
assign addr[11838]= -720088517;
assign addr[11839]= -756003771;
assign addr[11840]= -791679244;
assign addr[11841]= -827103620;
assign addr[11842]= -862265664;
assign addr[11843]= -897154224;
assign addr[11844]= -931758235;
assign addr[11845]= -966066720;
assign addr[11846]= -1000068799;
assign addr[11847]= -1033753687;
assign addr[11848]= -1067110699;
assign addr[11849]= -1100129257;
assign addr[11850]= -1132798888;
assign addr[11851]= -1165109230;
assign addr[11852]= -1197050035;
assign addr[11853]= -1228611172;
assign addr[11854]= -1259782632;
assign addr[11855]= -1290554528;
assign addr[11856]= -1320917099;
assign addr[11857]= -1350860716;
assign addr[11858]= -1380375881;
assign addr[11859]= -1409453233;
assign addr[11860]= -1438083551;
assign addr[11861]= -1466257752;
assign addr[11862]= -1493966902;
assign addr[11863]= -1521202211;
assign addr[11864]= -1547955041;
assign addr[11865]= -1574216908;
assign addr[11866]= -1599979481;
assign addr[11867]= -1625234591;
assign addr[11868]= -1649974225;
assign addr[11869]= -1674190539;
assign addr[11870]= -1697875851;
assign addr[11871]= -1721022648;
assign addr[11872]= -1743623590;
assign addr[11873]= -1765671509;
assign addr[11874]= -1787159411;
assign addr[11875]= -1808080480;
assign addr[11876]= -1828428082;
assign addr[11877]= -1848195763;
assign addr[11878]= -1867377253;
assign addr[11879]= -1885966468;
assign addr[11880]= -1903957513;
assign addr[11881]= -1921344681;
assign addr[11882]= -1938122457;
assign addr[11883]= -1954285520;
assign addr[11884]= -1969828744;
assign addr[11885]= -1984747199;
assign addr[11886]= -1999036154;
assign addr[11887]= -2012691075;
assign addr[11888]= -2025707632;
assign addr[11889]= -2038081698;
assign addr[11890]= -2049809346;
assign addr[11891]= -2060886858;
assign addr[11892]= -2071310720;
assign addr[11893]= -2081077626;
assign addr[11894]= -2090184478;
assign addr[11895]= -2098628387;
assign addr[11896]= -2106406677;
assign addr[11897]= -2113516878;
assign addr[11898]= -2119956737;
assign addr[11899]= -2125724211;
assign addr[11900]= -2130817471;
assign addr[11901]= -2135234901;
assign addr[11902]= -2138975100;
assign addr[11903]= -2142036881;
assign addr[11904]= -2144419275;
assign addr[11905]= -2146121524;
assign addr[11906]= -2147143090;
assign addr[11907]= -2147483648;
assign addr[11908]= -2147143090;
assign addr[11909]= -2146121524;
assign addr[11910]= -2144419275;
assign addr[11911]= -2142036881;
assign addr[11912]= -2138975100;
assign addr[11913]= -2135234901;
assign addr[11914]= -2130817471;
assign addr[11915]= -2125724211;
assign addr[11916]= -2119956737;
assign addr[11917]= -2113516878;
assign addr[11918]= -2106406677;
assign addr[11919]= -2098628387;
assign addr[11920]= -2090184478;
assign addr[11921]= -2081077626;
assign addr[11922]= -2071310720;
assign addr[11923]= -2060886858;
assign addr[11924]= -2049809346;
assign addr[11925]= -2038081698;
assign addr[11926]= -2025707632;
assign addr[11927]= -2012691075;
assign addr[11928]= -1999036154;
assign addr[11929]= -1984747199;
assign addr[11930]= -1969828744;
assign addr[11931]= -1954285520;
assign addr[11932]= -1938122457;
assign addr[11933]= -1921344681;
assign addr[11934]= -1903957513;
assign addr[11935]= -1885966468;
assign addr[11936]= -1867377253;
assign addr[11937]= -1848195763;
assign addr[11938]= -1828428082;
assign addr[11939]= -1808080480;
assign addr[11940]= -1787159411;
assign addr[11941]= -1765671509;
assign addr[11942]= -1743623590;
assign addr[11943]= -1721022648;
assign addr[11944]= -1697875851;
assign addr[11945]= -1674190539;
assign addr[11946]= -1649974225;
assign addr[11947]= -1625234591;
assign addr[11948]= -1599979481;
assign addr[11949]= -1574216908;
assign addr[11950]= -1547955041;
assign addr[11951]= -1521202211;
assign addr[11952]= -1493966902;
assign addr[11953]= -1466257752;
assign addr[11954]= -1438083551;
assign addr[11955]= -1409453233;
assign addr[11956]= -1380375881;
assign addr[11957]= -1350860716;
assign addr[11958]= -1320917099;
assign addr[11959]= -1290554528;
assign addr[11960]= -1259782632;
assign addr[11961]= -1228611172;
assign addr[11962]= -1197050035;
assign addr[11963]= -1165109230;
assign addr[11964]= -1132798888;
assign addr[11965]= -1100129257;
assign addr[11966]= -1067110699;
assign addr[11967]= -1033753687;
assign addr[11968]= -1000068799;
assign addr[11969]= -966066720;
assign addr[11970]= -931758235;
assign addr[11971]= -897154224;
assign addr[11972]= -862265664;
assign addr[11973]= -827103620;
assign addr[11974]= -791679244;
assign addr[11975]= -756003771;
assign addr[11976]= -720088517;
assign addr[11977]= -683944874;
assign addr[11978]= -647584304;
assign addr[11979]= -611018340;
assign addr[11980]= -574258580;
assign addr[11981]= -537316682;
assign addr[11982]= -500204365;
assign addr[11983]= -462933398;
assign addr[11984]= -425515602;
assign addr[11985]= -387962847;
assign addr[11986]= -350287041;
assign addr[11987]= -312500135;
assign addr[11988]= -274614114;
assign addr[11989]= -236640993;
assign addr[11990]= -198592817;
assign addr[11991]= -160481654;
assign addr[11992]= -122319591;
assign addr[11993]= -84118732;
assign addr[11994]= -45891193;
assign addr[11995]= -7649098;
assign addr[11996]= 30595422;
assign addr[11997]= 68830239;
assign addr[11998]= 107043224;
assign addr[11999]= 145222259;
assign addr[12000]= 183355234;
assign addr[12001]= 221430054;
assign addr[12002]= 259434643;
assign addr[12003]= 297356948;
assign addr[12004]= 335184940;
assign addr[12005]= 372906622;
assign addr[12006]= 410510029;
assign addr[12007]= 447983235;
assign addr[12008]= 485314355;
assign addr[12009]= 522491548;
assign addr[12010]= 559503022;
assign addr[12011]= 596337040;
assign addr[12012]= 632981917;
assign addr[12013]= 669426032;
assign addr[12014]= 705657826;
assign addr[12015]= 741665807;
assign addr[12016]= 777438554;
assign addr[12017]= 812964722;
assign addr[12018]= 848233042;
assign addr[12019]= 883232329;
assign addr[12020]= 917951481;
assign addr[12021]= 952379488;
assign addr[12022]= 986505429;
assign addr[12023]= 1020318481;
assign addr[12024]= 1053807919;
assign addr[12025]= 1086963121;
assign addr[12026]= 1119773573;
assign addr[12027]= 1152228866;
assign addr[12028]= 1184318708;
assign addr[12029]= 1216032921;
assign addr[12030]= 1247361445;
assign addr[12031]= 1278294345;
assign addr[12032]= 1308821808;
assign addr[12033]= 1338934154;
assign addr[12034]= 1368621831;
assign addr[12035]= 1397875423;
assign addr[12036]= 1426685652;
assign addr[12037]= 1455043381;
assign addr[12038]= 1482939614;
assign addr[12039]= 1510365504;
assign addr[12040]= 1537312353;
assign addr[12041]= 1563771613;
assign addr[12042]= 1589734894;
assign addr[12043]= 1615193959;
assign addr[12044]= 1640140734;
assign addr[12045]= 1664567307;
assign addr[12046]= 1688465931;
assign addr[12047]= 1711829025;
assign addr[12048]= 1734649179;
assign addr[12049]= 1756919156;
assign addr[12050]= 1778631892;
assign addr[12051]= 1799780501;
assign addr[12052]= 1820358275;
assign addr[12053]= 1840358687;
assign addr[12054]= 1859775393;
assign addr[12055]= 1878602237;
assign addr[12056]= 1896833245;
assign addr[12057]= 1914462636;
assign addr[12058]= 1931484818;
assign addr[12059]= 1947894393;
assign addr[12060]= 1963686155;
assign addr[12061]= 1978855097;
assign addr[12062]= 1993396407;
assign addr[12063]= 2007305472;
assign addr[12064]= 2020577882;
assign addr[12065]= 2033209426;
assign addr[12066]= 2045196100;
assign addr[12067]= 2056534099;
assign addr[12068]= 2067219829;
assign addr[12069]= 2077249901;
assign addr[12070]= 2086621133;
assign addr[12071]= 2095330553;
assign addr[12072]= 2103375398;
assign addr[12073]= 2110753117;
assign addr[12074]= 2117461370;
assign addr[12075]= 2123498030;
assign addr[12076]= 2128861181;
assign addr[12077]= 2133549123;
assign addr[12078]= 2137560369;
assign addr[12079]= 2140893646;
assign addr[12080]= 2143547897;
assign addr[12081]= 2145522281;
assign addr[12082]= 2146816171;
assign addr[12083]= 2147429158;
assign addr[12084]= 2147361045;
assign addr[12085]= 2146611856;
assign addr[12086]= 2145181827;
assign addr[12087]= 2143071413;
assign addr[12088]= 2140281282;
assign addr[12089]= 2136812319;
assign addr[12090]= 2132665626;
assign addr[12091]= 2127842516;
assign addr[12092]= 2122344521;
assign addr[12093]= 2116173382;
assign addr[12094]= 2109331059;
assign addr[12095]= 2101819720;
assign addr[12096]= 2093641749;
assign addr[12097]= 2084799740;
assign addr[12098]= 2075296495;
assign addr[12099]= 2065135031;
assign addr[12100]= 2054318569;
assign addr[12101]= 2042850540;
assign addr[12102]= 2030734582;
assign addr[12103]= 2017974537;
assign addr[12104]= 2004574453;
assign addr[12105]= 1990538579;
assign addr[12106]= 1975871368;
assign addr[12107]= 1960577471;
assign addr[12108]= 1944661739;
assign addr[12109]= 1928129220;
assign addr[12110]= 1910985158;
assign addr[12111]= 1893234990;
assign addr[12112]= 1874884346;
assign addr[12113]= 1855939047;
assign addr[12114]= 1836405100;
assign addr[12115]= 1816288703;
assign addr[12116]= 1795596234;
assign addr[12117]= 1774334257;
assign addr[12118]= 1752509516;
assign addr[12119]= 1730128933;
assign addr[12120]= 1707199606;
assign addr[12121]= 1683728808;
assign addr[12122]= 1659723983;
assign addr[12123]= 1635192744;
assign addr[12124]= 1610142873;
assign addr[12125]= 1584582314;
assign addr[12126]= 1558519173;
assign addr[12127]= 1531961719;
assign addr[12128]= 1504918373;
assign addr[12129]= 1477397714;
assign addr[12130]= 1449408469;
assign addr[12131]= 1420959516;
assign addr[12132]= 1392059879;
assign addr[12133]= 1362718723;
assign addr[12134]= 1332945355;
assign addr[12135]= 1302749217;
assign addr[12136]= 1272139887;
assign addr[12137]= 1241127074;
assign addr[12138]= 1209720613;
assign addr[12139]= 1177930466;
assign addr[12140]= 1145766716;
assign addr[12141]= 1113239564;
assign addr[12142]= 1080359326;
assign addr[12143]= 1047136432;
assign addr[12144]= 1013581418;
assign addr[12145]= 979704927;
assign addr[12146]= 945517704;
assign addr[12147]= 911030591;
assign addr[12148]= 876254528;
assign addr[12149]= 841200544;
assign addr[12150]= 805879757;
assign addr[12151]= 770303369;
assign addr[12152]= 734482665;
assign addr[12153]= 698429006;
assign addr[12154]= 662153826;
assign addr[12155]= 625668632;
assign addr[12156]= 588984994;
assign addr[12157]= 552114549;
assign addr[12158]= 515068990;
assign addr[12159]= 477860067;
assign addr[12160]= 440499581;
assign addr[12161]= 402999383;
assign addr[12162]= 365371365;
assign addr[12163]= 327627463;
assign addr[12164]= 289779648;
assign addr[12165]= 251839923;
assign addr[12166]= 213820322;
assign addr[12167]= 175732905;
assign addr[12168]= 137589750;
assign addr[12169]= 99402956;
assign addr[12170]= 61184634;
assign addr[12171]= 22946906;
assign addr[12172]= -15298099;
assign addr[12173]= -53538253;
assign addr[12174]= -91761426;
assign addr[12175]= -129955495;
assign addr[12176]= -168108346;
assign addr[12177]= -206207878;
assign addr[12178]= -244242007;
assign addr[12179]= -282198671;
assign addr[12180]= -320065829;
assign addr[12181]= -357831473;
assign addr[12182]= -395483624;
assign addr[12183]= -433010339;
assign addr[12184]= -470399716;
assign addr[12185]= -507639898;
assign addr[12186]= -544719071;
assign addr[12187]= -581625477;
assign addr[12188]= -618347408;
assign addr[12189]= -654873219;
assign addr[12190]= -691191324;
assign addr[12191]= -727290205;
assign addr[12192]= -763158411;
assign addr[12193]= -798784567;
assign addr[12194]= -834157373;
assign addr[12195]= -869265610;
assign addr[12196]= -904098143;
assign addr[12197]= -938643924;
assign addr[12198]= -972891995;
assign addr[12199]= -1006831495;
assign addr[12200]= -1040451659;
assign addr[12201]= -1073741824;
assign addr[12202]= -1106691431;
assign addr[12203]= -1139290029;
assign addr[12204]= -1171527280;
assign addr[12205]= -1203392958;
assign addr[12206]= -1234876957;
assign addr[12207]= -1265969291;
assign addr[12208]= -1296660098;
assign addr[12209]= -1326939644;
assign addr[12210]= -1356798326;
assign addr[12211]= -1386226674;
assign addr[12212]= -1415215352;
assign addr[12213]= -1443755168;
assign addr[12214]= -1471837070;
assign addr[12215]= -1499452149;
assign addr[12216]= -1526591649;
assign addr[12217]= -1553246960;
assign addr[12218]= -1579409630;
assign addr[12219]= -1605071359;
assign addr[12220]= -1630224009;
assign addr[12221]= -1654859602;
assign addr[12222]= -1678970324;
assign addr[12223]= -1702548529;
assign addr[12224]= -1725586737;
assign addr[12225]= -1748077642;
assign addr[12226]= -1770014111;
assign addr[12227]= -1791389186;
assign addr[12228]= -1812196087;
assign addr[12229]= -1832428215;
assign addr[12230]= -1852079154;
assign addr[12231]= -1871142669;
assign addr[12232]= -1889612716;
assign addr[12233]= -1907483436;
assign addr[12234]= -1924749160;
assign addr[12235]= -1941404413;
assign addr[12236]= -1957443913;
assign addr[12237]= -1972862571;
assign addr[12238]= -1987655498;
assign addr[12239]= -2001818002;
assign addr[12240]= -2015345591;
assign addr[12241]= -2028233973;
assign addr[12242]= -2040479063;
assign addr[12243]= -2052076975;
assign addr[12244]= -2063024031;
assign addr[12245]= -2073316760;
assign addr[12246]= -2082951896;
assign addr[12247]= -2091926384;
assign addr[12248]= -2100237377;
assign addr[12249]= -2107882239;
assign addr[12250]= -2114858546;
assign addr[12251]= -2121164085;
assign addr[12252]= -2126796855;
assign addr[12253]= -2131755071;
assign addr[12254]= -2136037160;
assign addr[12255]= -2139641764;
assign addr[12256]= -2142567738;
assign addr[12257]= -2144814157;
assign addr[12258]= -2146380306;
assign addr[12259]= -2147265689;
assign addr[12260]= -2147470025;
assign addr[12261]= -2146993250;
assign addr[12262]= -2145835515;
assign addr[12263]= -2143997187;
assign addr[12264]= -2141478848;
assign addr[12265]= -2138281298;
assign addr[12266]= -2134405552;
assign addr[12267]= -2129852837;
assign addr[12268]= -2124624598;
assign addr[12269]= -2118722494;
assign addr[12270]= -2112148396;
assign addr[12271]= -2104904390;
assign addr[12272]= -2096992772;
assign addr[12273]= -2088416053;
assign addr[12274]= -2079176953;
assign addr[12275]= -2069278401;
assign addr[12276]= -2058723538;
assign addr[12277]= -2047515711;
assign addr[12278]= -2035658475;
assign addr[12279]= -2023155591;
assign addr[12280]= -2010011024;
assign addr[12281]= -1996228943;
assign addr[12282]= -1981813720;
assign addr[12283]= -1966769926;
assign addr[12284]= -1951102334;
assign addr[12285]= -1934815911;
assign addr[12286]= -1917915825;
assign addr[12287]= -1900407434;
assign addr[12288]= -1882296293;
assign addr[12289]= -1863588145;
assign addr[12290]= -1844288924;
assign addr[12291]= -1824404752;
assign addr[12292]= -1803941934;
assign addr[12293]= -1782906961;
assign addr[12294]= -1761306505;
assign addr[12295]= -1739147417;
assign addr[12296]= -1716436725;
assign addr[12297]= -1693181631;
assign addr[12298]= -1669389513;
assign addr[12299]= -1645067915;
assign addr[12300]= -1620224553;
assign addr[12301]= -1594867305;
assign addr[12302]= -1569004214;
assign addr[12303]= -1542643483;
assign addr[12304]= -1515793473;
assign addr[12305]= -1488462700;
assign addr[12306]= -1460659832;
assign addr[12307]= -1432393688;
assign addr[12308]= -1403673233;
assign addr[12309]= -1374507575;
assign addr[12310]= -1344905966;
assign addr[12311]= -1314877795;
assign addr[12312]= -1284432584;
assign addr[12313]= -1253579991;
assign addr[12314]= -1222329801;
assign addr[12315]= -1190691925;
assign addr[12316]= -1158676398;
assign addr[12317]= -1126293375;
assign addr[12318]= -1093553126;
assign addr[12319]= -1060466036;
assign addr[12320]= -1027042599;
assign addr[12321]= -993293415;
assign addr[12322]= -959229189;
assign addr[12323]= -924860725;
assign addr[12324]= -890198924;
assign addr[12325]= -855254778;
assign addr[12326]= -820039373;
assign addr[12327]= -784563876;
assign addr[12328]= -748839539;
assign addr[12329]= -712877694;
assign addr[12330]= -676689746;
assign addr[12331]= -640287172;
assign addr[12332]= -603681519;
assign addr[12333]= -566884397;
assign addr[12334]= -529907477;
assign addr[12335]= -492762486;
assign addr[12336]= -455461206;
assign addr[12337]= -418015468;
assign addr[12338]= -380437148;
assign addr[12339]= -342738165;
assign addr[12340]= -304930476;
assign addr[12341]= -267026072;
assign addr[12342]= -229036977;
assign addr[12343]= -190975237;
assign addr[12344]= -152852926;
assign addr[12345]= -114682135;
assign addr[12346]= -76474970;
assign addr[12347]= -38243550;
assign addr[12348]= 0;
assign addr[12349]= 38243550;
assign addr[12350]= 76474970;
assign addr[12351]= 114682135;
assign addr[12352]= 152852926;
assign addr[12353]= 190975237;
assign addr[12354]= 229036977;
assign addr[12355]= 267026072;
assign addr[12356]= 304930476;
assign addr[12357]= 342738165;
assign addr[12358]= 380437148;
assign addr[12359]= 418015468;
assign addr[12360]= 455461206;
assign addr[12361]= 492762486;
assign addr[12362]= 529907477;
assign addr[12363]= 566884397;
assign addr[12364]= 603681519;
assign addr[12365]= 640287172;
assign addr[12366]= 676689746;
assign addr[12367]= 712877694;
assign addr[12368]= 748839539;
assign addr[12369]= 784563876;
assign addr[12370]= 820039373;
assign addr[12371]= 855254778;
assign addr[12372]= 890198924;
assign addr[12373]= 924860725;
assign addr[12374]= 959229189;
assign addr[12375]= 993293415;
assign addr[12376]= 1027042599;
assign addr[12377]= 1060466036;
assign addr[12378]= 1093553126;
assign addr[12379]= 1126293375;
assign addr[12380]= 1158676398;
assign addr[12381]= 1190691925;
assign addr[12382]= 1222329801;
assign addr[12383]= 1253579991;
assign addr[12384]= 1284432584;
assign addr[12385]= 1314877795;
assign addr[12386]= 1344905966;
assign addr[12387]= 1374507575;
assign addr[12388]= 1403673233;
assign addr[12389]= 1432393688;
assign addr[12390]= 1460659832;
assign addr[12391]= 1488462700;
assign addr[12392]= 1515793473;
assign addr[12393]= 1542643483;
assign addr[12394]= 1569004214;
assign addr[12395]= 1594867305;
assign addr[12396]= 1620224553;
assign addr[12397]= 1645067915;
assign addr[12398]= 1669389513;
assign addr[12399]= 1693181631;
assign addr[12400]= 1716436725;
assign addr[12401]= 1739147417;
assign addr[12402]= 1761306505;
assign addr[12403]= 1782906961;
assign addr[12404]= 1803941934;
assign addr[12405]= 1824404752;
assign addr[12406]= 1844288924;
assign addr[12407]= 1863588145;
assign addr[12408]= 1882296293;
assign addr[12409]= 1900407434;
assign addr[12410]= 1917915825;
assign addr[12411]= 1934815911;
assign addr[12412]= 1951102334;
assign addr[12413]= 1966769926;
assign addr[12414]= 1981813720;
assign addr[12415]= 1996228943;
assign addr[12416]= 2010011024;
assign addr[12417]= 2023155591;
assign addr[12418]= 2035658475;
assign addr[12419]= 2047515711;
assign addr[12420]= 2058723538;
assign addr[12421]= 2069278401;
assign addr[12422]= 2079176953;
assign addr[12423]= 2088416053;
assign addr[12424]= 2096992772;
assign addr[12425]= 2104904390;
assign addr[12426]= 2112148396;
assign addr[12427]= 2118722494;
assign addr[12428]= 2124624598;
assign addr[12429]= 2129852837;
assign addr[12430]= 2134405552;
assign addr[12431]= 2138281298;
assign addr[12432]= 2141478848;
assign addr[12433]= 2143997187;
assign addr[12434]= 2145835515;
assign addr[12435]= 2146993250;
assign addr[12436]= 2147470025;
assign addr[12437]= 2147265689;
assign addr[12438]= 2146380306;
assign addr[12439]= 2144814157;
assign addr[12440]= 2142567738;
assign addr[12441]= 2139641764;
assign addr[12442]= 2136037160;
assign addr[12443]= 2131755071;
assign addr[12444]= 2126796855;
assign addr[12445]= 2121164085;
assign addr[12446]= 2114858546;
assign addr[12447]= 2107882239;
assign addr[12448]= 2100237377;
assign addr[12449]= 2091926384;
assign addr[12450]= 2082951896;
assign addr[12451]= 2073316760;
assign addr[12452]= 2063024031;
assign addr[12453]= 2052076975;
assign addr[12454]= 2040479063;
assign addr[12455]= 2028233973;
assign addr[12456]= 2015345591;
assign addr[12457]= 2001818002;
assign addr[12458]= 1987655498;
assign addr[12459]= 1972862571;
assign addr[12460]= 1957443913;
assign addr[12461]= 1941404413;
assign addr[12462]= 1924749160;
assign addr[12463]= 1907483436;
assign addr[12464]= 1889612716;
assign addr[12465]= 1871142669;
assign addr[12466]= 1852079154;
assign addr[12467]= 1832428215;
assign addr[12468]= 1812196087;
assign addr[12469]= 1791389186;
assign addr[12470]= 1770014111;
assign addr[12471]= 1748077642;
assign addr[12472]= 1725586737;
assign addr[12473]= 1702548529;
assign addr[12474]= 1678970324;
assign addr[12475]= 1654859602;
assign addr[12476]= 1630224009;
assign addr[12477]= 1605071359;
assign addr[12478]= 1579409630;
assign addr[12479]= 1553246960;
assign addr[12480]= 1526591649;
assign addr[12481]= 1499452149;
assign addr[12482]= 1471837070;
assign addr[12483]= 1443755168;
assign addr[12484]= 1415215352;
assign addr[12485]= 1386226674;
assign addr[12486]= 1356798326;
assign addr[12487]= 1326939644;
assign addr[12488]= 1296660098;
assign addr[12489]= 1265969291;
assign addr[12490]= 1234876957;
assign addr[12491]= 1203392958;
assign addr[12492]= 1171527280;
assign addr[12493]= 1139290029;
assign addr[12494]= 1106691431;
assign addr[12495]= 1073741824;
assign addr[12496]= 1040451659;
assign addr[12497]= 1006831495;
assign addr[12498]= 972891995;
assign addr[12499]= 938643924;
assign addr[12500]= 904098143;
assign addr[12501]= 869265610;
assign addr[12502]= 834157373;
assign addr[12503]= 798784567;
assign addr[12504]= 763158411;
assign addr[12505]= 727290205;
assign addr[12506]= 691191324;
assign addr[12507]= 654873219;
assign addr[12508]= 618347408;
assign addr[12509]= 581625477;
assign addr[12510]= 544719071;
assign addr[12511]= 507639898;
assign addr[12512]= 470399716;
assign addr[12513]= 433010339;
assign addr[12514]= 395483624;
assign addr[12515]= 357831473;
assign addr[12516]= 320065829;
assign addr[12517]= 282198671;
assign addr[12518]= 244242007;
assign addr[12519]= 206207878;
assign addr[12520]= 168108346;
assign addr[12521]= 129955495;
assign addr[12522]= 91761426;
assign addr[12523]= 53538253;
assign addr[12524]= 15298099;
assign addr[12525]= -22946906;
assign addr[12526]= -61184634;
assign addr[12527]= -99402956;
assign addr[12528]= -137589750;
assign addr[12529]= -175732905;
assign addr[12530]= -213820322;
assign addr[12531]= -251839923;
assign addr[12532]= -289779648;
assign addr[12533]= -327627463;
assign addr[12534]= -365371365;
assign addr[12535]= -402999383;
assign addr[12536]= -440499581;
assign addr[12537]= -477860067;
assign addr[12538]= -515068990;
assign addr[12539]= -552114549;
assign addr[12540]= -588984994;
assign addr[12541]= -625668632;
assign addr[12542]= -662153826;
assign addr[12543]= -698429006;
assign addr[12544]= -734482665;
assign addr[12545]= -770303369;
assign addr[12546]= -805879757;
assign addr[12547]= -841200544;
assign addr[12548]= -876254528;
assign addr[12549]= -911030591;
assign addr[12550]= -945517704;
assign addr[12551]= -979704927;
assign addr[12552]= -1013581418;
assign addr[12553]= -1047136432;
assign addr[12554]= -1080359326;
assign addr[12555]= -1113239564;
assign addr[12556]= -1145766716;
assign addr[12557]= -1177930466;
assign addr[12558]= -1209720613;
assign addr[12559]= -1241127074;
assign addr[12560]= -1272139887;
assign addr[12561]= -1302749217;
assign addr[12562]= -1332945355;
assign addr[12563]= -1362718723;
assign addr[12564]= -1392059879;
assign addr[12565]= -1420959516;
assign addr[12566]= -1449408469;
assign addr[12567]= -1477397714;
assign addr[12568]= -1504918373;
assign addr[12569]= -1531961719;
assign addr[12570]= -1558519173;
assign addr[12571]= -1584582314;
assign addr[12572]= -1610142873;
assign addr[12573]= -1635192744;
assign addr[12574]= -1659723983;
assign addr[12575]= -1683728808;
assign addr[12576]= -1707199606;
assign addr[12577]= -1730128933;
assign addr[12578]= -1752509516;
assign addr[12579]= -1774334257;
assign addr[12580]= -1795596234;
assign addr[12581]= -1816288703;
assign addr[12582]= -1836405100;
assign addr[12583]= -1855939047;
assign addr[12584]= -1874884346;
assign addr[12585]= -1893234990;
assign addr[12586]= -1910985158;
assign addr[12587]= -1928129220;
assign addr[12588]= -1944661739;
assign addr[12589]= -1960577471;
assign addr[12590]= -1975871368;
assign addr[12591]= -1990538579;
assign addr[12592]= -2004574453;
assign addr[12593]= -2017974537;
assign addr[12594]= -2030734582;
assign addr[12595]= -2042850540;
assign addr[12596]= -2054318569;
assign addr[12597]= -2065135031;
assign addr[12598]= -2075296495;
assign addr[12599]= -2084799740;
assign addr[12600]= -2093641749;
assign addr[12601]= -2101819720;
assign addr[12602]= -2109331059;
assign addr[12603]= -2116173382;
assign addr[12604]= -2122344521;
assign addr[12605]= -2127842516;
assign addr[12606]= -2132665626;
assign addr[12607]= -2136812319;
assign addr[12608]= -2140281282;
assign addr[12609]= -2143071413;
assign addr[12610]= -2145181827;
assign addr[12611]= -2146611856;
assign addr[12612]= -2147361045;
assign addr[12613]= -2147429158;
assign addr[12614]= -2146816171;
assign addr[12615]= -2145522281;
assign addr[12616]= -2143547897;
assign addr[12617]= -2140893646;
assign addr[12618]= -2137560369;
assign addr[12619]= -2133549123;
assign addr[12620]= -2128861181;
assign addr[12621]= -2123498030;
assign addr[12622]= -2117461370;
assign addr[12623]= -2110753117;
assign addr[12624]= -2103375398;
assign addr[12625]= -2095330553;
assign addr[12626]= -2086621133;
assign addr[12627]= -2077249901;
assign addr[12628]= -2067219829;
assign addr[12629]= -2056534099;
assign addr[12630]= -2045196100;
assign addr[12631]= -2033209426;
assign addr[12632]= -2020577882;
assign addr[12633]= -2007305472;
assign addr[12634]= -1993396407;
assign addr[12635]= -1978855097;
assign addr[12636]= -1963686155;
assign addr[12637]= -1947894393;
assign addr[12638]= -1931484818;
assign addr[12639]= -1914462636;
assign addr[12640]= -1896833245;
assign addr[12641]= -1878602237;
assign addr[12642]= -1859775393;
assign addr[12643]= -1840358687;
assign addr[12644]= -1820358275;
assign addr[12645]= -1799780501;
assign addr[12646]= -1778631892;
assign addr[12647]= -1756919156;
assign addr[12648]= -1734649179;
assign addr[12649]= -1711829025;
assign addr[12650]= -1688465931;
assign addr[12651]= -1664567307;
assign addr[12652]= -1640140734;
assign addr[12653]= -1615193959;
assign addr[12654]= -1589734894;
assign addr[12655]= -1563771613;
assign addr[12656]= -1537312353;
assign addr[12657]= -1510365504;
assign addr[12658]= -1482939614;
assign addr[12659]= -1455043381;
assign addr[12660]= -1426685652;
assign addr[12661]= -1397875423;
assign addr[12662]= -1368621831;
assign addr[12663]= -1338934154;
assign addr[12664]= -1308821808;
assign addr[12665]= -1278294345;
assign addr[12666]= -1247361445;
assign addr[12667]= -1216032921;
assign addr[12668]= -1184318708;
assign addr[12669]= -1152228866;
assign addr[12670]= -1119773573;
assign addr[12671]= -1086963121;
assign addr[12672]= -1053807919;
assign addr[12673]= -1020318481;
assign addr[12674]= -986505429;
assign addr[12675]= -952379488;
assign addr[12676]= -917951481;
assign addr[12677]= -883232329;
assign addr[12678]= -848233042;
assign addr[12679]= -812964722;
assign addr[12680]= -777438554;
assign addr[12681]= -741665807;
assign addr[12682]= -705657826;
assign addr[12683]= -669426032;
assign addr[12684]= -632981917;
assign addr[12685]= -596337040;
assign addr[12686]= -559503022;
assign addr[12687]= -522491548;
assign addr[12688]= -485314355;
assign addr[12689]= -447983235;
assign addr[12690]= -410510029;
assign addr[12691]= -372906622;
assign addr[12692]= -335184940;
assign addr[12693]= -297356948;
assign addr[12694]= -259434643;
assign addr[12695]= -221430054;
assign addr[12696]= -183355234;
assign addr[12697]= -145222259;
assign addr[12698]= -107043224;
assign addr[12699]= -68830239;
assign addr[12700]= -30595422;
assign addr[12701]= 7649098;
assign addr[12702]= 45891193;
assign addr[12703]= 84118732;
assign addr[12704]= 122319591;
assign addr[12705]= 160481654;
assign addr[12706]= 198592817;
assign addr[12707]= 236640993;
assign addr[12708]= 274614114;
assign addr[12709]= 312500135;
assign addr[12710]= 350287041;
assign addr[12711]= 387962847;
assign addr[12712]= 425515602;
assign addr[12713]= 462933398;
assign addr[12714]= 500204365;
assign addr[12715]= 537316682;
assign addr[12716]= 574258580;
assign addr[12717]= 611018340;
assign addr[12718]= 647584304;
assign addr[12719]= 683944874;
assign addr[12720]= 720088517;
assign addr[12721]= 756003771;
assign addr[12722]= 791679244;
assign addr[12723]= 827103620;
assign addr[12724]= 862265664;
assign addr[12725]= 897154224;
assign addr[12726]= 931758235;
assign addr[12727]= 966066720;
assign addr[12728]= 1000068799;
assign addr[12729]= 1033753687;
assign addr[12730]= 1067110699;
assign addr[12731]= 1100129257;
assign addr[12732]= 1132798888;
assign addr[12733]= 1165109230;
assign addr[12734]= 1197050035;
assign addr[12735]= 1228611172;
assign addr[12736]= 1259782632;
assign addr[12737]= 1290554528;
assign addr[12738]= 1320917099;
assign addr[12739]= 1350860716;
assign addr[12740]= 1380375881;
assign addr[12741]= 1409453233;
assign addr[12742]= 1438083551;
assign addr[12743]= 1466257752;
assign addr[12744]= 1493966902;
assign addr[12745]= 1521202211;
assign addr[12746]= 1547955041;
assign addr[12747]= 1574216908;
assign addr[12748]= 1599979481;
assign addr[12749]= 1625234591;
assign addr[12750]= 1649974225;
assign addr[12751]= 1674190539;
assign addr[12752]= 1697875851;
assign addr[12753]= 1721022648;
assign addr[12754]= 1743623590;
assign addr[12755]= 1765671509;
assign addr[12756]= 1787159411;
assign addr[12757]= 1808080480;
assign addr[12758]= 1828428082;
assign addr[12759]= 1848195763;
assign addr[12760]= 1867377253;
assign addr[12761]= 1885966468;
assign addr[12762]= 1903957513;
assign addr[12763]= 1921344681;
assign addr[12764]= 1938122457;
assign addr[12765]= 1954285520;
assign addr[12766]= 1969828744;
assign addr[12767]= 1984747199;
assign addr[12768]= 1999036154;
assign addr[12769]= 2012691075;
assign addr[12770]= 2025707632;
assign addr[12771]= 2038081698;
assign addr[12772]= 2049809346;
assign addr[12773]= 2060886858;
assign addr[12774]= 2071310720;
assign addr[12775]= 2081077626;
assign addr[12776]= 2090184478;
assign addr[12777]= 2098628387;
assign addr[12778]= 2106406677;
assign addr[12779]= 2113516878;
assign addr[12780]= 2119956737;
assign addr[12781]= 2125724211;
assign addr[12782]= 2130817471;
assign addr[12783]= 2135234901;
assign addr[12784]= 2138975100;
assign addr[12785]= 2142036881;
assign addr[12786]= 2144419275;
assign addr[12787]= 2146121524;
assign addr[12788]= 2147143090;
assign addr[12789]= 2147483648;
assign addr[12790]= 2147143090;
assign addr[12791]= 2146121524;
assign addr[12792]= 2144419275;
assign addr[12793]= 2142036881;
assign addr[12794]= 2138975100;
assign addr[12795]= 2135234901;
assign addr[12796]= 2130817471;
assign addr[12797]= 2125724211;
assign addr[12798]= 2119956737;
assign addr[12799]= 2113516878;
assign addr[12800]= 2106406677;
assign addr[12801]= 2098628387;
assign addr[12802]= 2090184478;
assign addr[12803]= 2081077626;
assign addr[12804]= 2071310720;
assign addr[12805]= 2060886858;
assign addr[12806]= 2049809346;
assign addr[12807]= 2038081698;
assign addr[12808]= 2025707632;
assign addr[12809]= 2012691075;
assign addr[12810]= 1999036154;
assign addr[12811]= 1984747199;
assign addr[12812]= 1969828744;
assign addr[12813]= 1954285520;
assign addr[12814]= 1938122457;
assign addr[12815]= 1921344681;
assign addr[12816]= 1903957513;
assign addr[12817]= 1885966468;
assign addr[12818]= 1867377253;
assign addr[12819]= 1848195763;
assign addr[12820]= 1828428082;
assign addr[12821]= 1808080480;
assign addr[12822]= 1787159411;
assign addr[12823]= 1765671509;
assign addr[12824]= 1743623590;
assign addr[12825]= 1721022648;
assign addr[12826]= 1697875851;
assign addr[12827]= 1674190539;
assign addr[12828]= 1649974225;
assign addr[12829]= 1625234591;
assign addr[12830]= 1599979481;
assign addr[12831]= 1574216908;
assign addr[12832]= 1547955041;
assign addr[12833]= 1521202211;
assign addr[12834]= 1493966902;
assign addr[12835]= 1466257752;
assign addr[12836]= 1438083551;
assign addr[12837]= 1409453233;
assign addr[12838]= 1380375881;
assign addr[12839]= 1350860716;
assign addr[12840]= 1320917099;
assign addr[12841]= 1290554528;
assign addr[12842]= 1259782632;
assign addr[12843]= 1228611172;
assign addr[12844]= 1197050035;
assign addr[12845]= 1165109230;
assign addr[12846]= 1132798888;
assign addr[12847]= 1100129257;
assign addr[12848]= 1067110699;
assign addr[12849]= 1033753687;
assign addr[12850]= 1000068799;
assign addr[12851]= 966066720;
assign addr[12852]= 931758235;
assign addr[12853]= 897154224;
assign addr[12854]= 862265664;
assign addr[12855]= 827103620;
assign addr[12856]= 791679244;
assign addr[12857]= 756003771;
assign addr[12858]= 720088517;
assign addr[12859]= 683944874;
assign addr[12860]= 647584304;
assign addr[12861]= 611018340;
assign addr[12862]= 574258580;
assign addr[12863]= 537316682;
assign addr[12864]= 500204365;
assign addr[12865]= 462933398;
assign addr[12866]= 425515602;
assign addr[12867]= 387962847;
assign addr[12868]= 350287041;
assign addr[12869]= 312500135;
assign addr[12870]= 274614114;
assign addr[12871]= 236640993;
assign addr[12872]= 198592817;
assign addr[12873]= 160481654;
assign addr[12874]= 122319591;
assign addr[12875]= 84118732;
assign addr[12876]= 45891193;
assign addr[12877]= 7649098;
assign addr[12878]= -30595422;
assign addr[12879]= -68830239;
assign addr[12880]= -107043224;
assign addr[12881]= -145222259;
assign addr[12882]= -183355234;
assign addr[12883]= -221430054;
assign addr[12884]= -259434643;
assign addr[12885]= -297356948;
assign addr[12886]= -335184940;
assign addr[12887]= -372906622;
assign addr[12888]= -410510029;
assign addr[12889]= -447983235;
assign addr[12890]= -485314355;
assign addr[12891]= -522491548;
assign addr[12892]= -559503022;
assign addr[12893]= -596337040;
assign addr[12894]= -632981917;
assign addr[12895]= -669426032;
assign addr[12896]= -705657826;
assign addr[12897]= -741665807;
assign addr[12898]= -777438554;
assign addr[12899]= -812964722;
assign addr[12900]= -848233042;
assign addr[12901]= -883232329;
assign addr[12902]= -917951481;
assign addr[12903]= -952379488;
assign addr[12904]= -986505429;
assign addr[12905]= -1020318481;
assign addr[12906]= -1053807919;
assign addr[12907]= -1086963121;
assign addr[12908]= -1119773573;
assign addr[12909]= -1152228866;
assign addr[12910]= -1184318708;
assign addr[12911]= -1216032921;
assign addr[12912]= -1247361445;
assign addr[12913]= -1278294345;
assign addr[12914]= -1308821808;
assign addr[12915]= -1338934154;
assign addr[12916]= -1368621831;
assign addr[12917]= -1397875423;
assign addr[12918]= -1426685652;
assign addr[12919]= -1455043381;
assign addr[12920]= -1482939614;
assign addr[12921]= -1510365504;
assign addr[12922]= -1537312353;
assign addr[12923]= -1563771613;
assign addr[12924]= -1589734894;
assign addr[12925]= -1615193959;
assign addr[12926]= -1640140734;
assign addr[12927]= -1664567307;
assign addr[12928]= -1688465931;
assign addr[12929]= -1711829025;
assign addr[12930]= -1734649179;
assign addr[12931]= -1756919156;
assign addr[12932]= -1778631892;
assign addr[12933]= -1799780501;
assign addr[12934]= -1820358275;
assign addr[12935]= -1840358687;
assign addr[12936]= -1859775393;
assign addr[12937]= -1878602237;
assign addr[12938]= -1896833245;
assign addr[12939]= -1914462636;
assign addr[12940]= -1931484818;
assign addr[12941]= -1947894393;
assign addr[12942]= -1963686155;
assign addr[12943]= -1978855097;
assign addr[12944]= -1993396407;
assign addr[12945]= -2007305472;
assign addr[12946]= -2020577882;
assign addr[12947]= -2033209426;
assign addr[12948]= -2045196100;
assign addr[12949]= -2056534099;
assign addr[12950]= -2067219829;
assign addr[12951]= -2077249901;
assign addr[12952]= -2086621133;
assign addr[12953]= -2095330553;
assign addr[12954]= -2103375398;
assign addr[12955]= -2110753117;
assign addr[12956]= -2117461370;
assign addr[12957]= -2123498030;
assign addr[12958]= -2128861181;
assign addr[12959]= -2133549123;
assign addr[12960]= -2137560369;
assign addr[12961]= -2140893646;
assign addr[12962]= -2143547897;
assign addr[12963]= -2145522281;
assign addr[12964]= -2146816171;
assign addr[12965]= -2147429158;
assign addr[12966]= -2147361045;
assign addr[12967]= -2146611856;
assign addr[12968]= -2145181827;
assign addr[12969]= -2143071413;
assign addr[12970]= -2140281282;
assign addr[12971]= -2136812319;
assign addr[12972]= -2132665626;
assign addr[12973]= -2127842516;
assign addr[12974]= -2122344521;
assign addr[12975]= -2116173382;
assign addr[12976]= -2109331059;
assign addr[12977]= -2101819720;
assign addr[12978]= -2093641749;
assign addr[12979]= -2084799740;
assign addr[12980]= -2075296495;
assign addr[12981]= -2065135031;
assign addr[12982]= -2054318569;
assign addr[12983]= -2042850540;
assign addr[12984]= -2030734582;
assign addr[12985]= -2017974537;
assign addr[12986]= -2004574453;
assign addr[12987]= -1990538579;
assign addr[12988]= -1975871368;
assign addr[12989]= -1960577471;
assign addr[12990]= -1944661739;
assign addr[12991]= -1928129220;
assign addr[12992]= -1910985158;
assign addr[12993]= -1893234990;
assign addr[12994]= -1874884346;
assign addr[12995]= -1855939047;
assign addr[12996]= -1836405100;
assign addr[12997]= -1816288703;
assign addr[12998]= -1795596234;
assign addr[12999]= -1774334257;
assign addr[13000]= -1752509516;
assign addr[13001]= -1730128933;
assign addr[13002]= -1707199606;
assign addr[13003]= -1683728808;
assign addr[13004]= -1659723983;
assign addr[13005]= -1635192744;
assign addr[13006]= -1610142873;
assign addr[13007]= -1584582314;
assign addr[13008]= -1558519173;
assign addr[13009]= -1531961719;
assign addr[13010]= -1504918373;
assign addr[13011]= -1477397714;
assign addr[13012]= -1449408469;
assign addr[13013]= -1420959516;
assign addr[13014]= -1392059879;
assign addr[13015]= -1362718723;
assign addr[13016]= -1332945355;
assign addr[13017]= -1302749217;
assign addr[13018]= -1272139887;
assign addr[13019]= -1241127074;
assign addr[13020]= -1209720613;
assign addr[13021]= -1177930466;
assign addr[13022]= -1145766716;
assign addr[13023]= -1113239564;
assign addr[13024]= -1080359326;
assign addr[13025]= -1047136432;
assign addr[13026]= -1013581418;
assign addr[13027]= -979704927;
assign addr[13028]= -945517704;
assign addr[13029]= -911030591;
assign addr[13030]= -876254528;
assign addr[13031]= -841200544;
assign addr[13032]= -805879757;
assign addr[13033]= -770303369;
assign addr[13034]= -734482665;
assign addr[13035]= -698429006;
assign addr[13036]= -662153826;
assign addr[13037]= -625668632;
assign addr[13038]= -588984994;
assign addr[13039]= -552114549;
assign addr[13040]= -515068990;
assign addr[13041]= -477860067;
assign addr[13042]= -440499581;
assign addr[13043]= -402999383;
assign addr[13044]= -365371365;
assign addr[13045]= -327627463;
assign addr[13046]= -289779648;
assign addr[13047]= -251839923;
assign addr[13048]= -213820322;
assign addr[13049]= -175732905;
assign addr[13050]= -137589750;
assign addr[13051]= -99402956;
assign addr[13052]= -61184634;
assign addr[13053]= -22946906;
assign addr[13054]= 15298099;
assign addr[13055]= 53538253;
assign addr[13056]= 91761426;
assign addr[13057]= 129955495;
assign addr[13058]= 168108346;
assign addr[13059]= 206207878;
assign addr[13060]= 244242007;
assign addr[13061]= 282198671;
assign addr[13062]= 320065829;
assign addr[13063]= 357831473;
assign addr[13064]= 395483624;
assign addr[13065]= 433010339;
assign addr[13066]= 470399716;
assign addr[13067]= 507639898;
assign addr[13068]= 544719071;
assign addr[13069]= 581625477;
assign addr[13070]= 618347408;
assign addr[13071]= 654873219;
assign addr[13072]= 691191324;
assign addr[13073]= 727290205;
assign addr[13074]= 763158411;
assign addr[13075]= 798784567;
assign addr[13076]= 834157373;
assign addr[13077]= 869265610;
assign addr[13078]= 904098143;
assign addr[13079]= 938643924;
assign addr[13080]= 972891995;
assign addr[13081]= 1006831495;
assign addr[13082]= 1040451659;
assign addr[13083]= 1073741824;
assign addr[13084]= 1106691431;
assign addr[13085]= 1139290029;
assign addr[13086]= 1171527280;
assign addr[13087]= 1203392958;
assign addr[13088]= 1234876957;
assign addr[13089]= 1265969291;
assign addr[13090]= 1296660098;
assign addr[13091]= 1326939644;
assign addr[13092]= 1356798326;
assign addr[13093]= 1386226674;
assign addr[13094]= 1415215352;
assign addr[13095]= 1443755168;
assign addr[13096]= 1471837070;
assign addr[13097]= 1499452149;
assign addr[13098]= 1526591649;
assign addr[13099]= 1553246960;
assign addr[13100]= 1579409630;
assign addr[13101]= 1605071359;
assign addr[13102]= 1630224009;
assign addr[13103]= 1654859602;
assign addr[13104]= 1678970324;
assign addr[13105]= 1702548529;
assign addr[13106]= 1725586737;
assign addr[13107]= 1748077642;
assign addr[13108]= 1770014111;
assign addr[13109]= 1791389186;
assign addr[13110]= 1812196087;
assign addr[13111]= 1832428215;
assign addr[13112]= 1852079154;
assign addr[13113]= 1871142669;
assign addr[13114]= 1889612716;
assign addr[13115]= 1907483436;
assign addr[13116]= 1924749160;
assign addr[13117]= 1941404413;
assign addr[13118]= 1957443913;
assign addr[13119]= 1972862571;
assign addr[13120]= 1987655498;
assign addr[13121]= 2001818002;
assign addr[13122]= 2015345591;
assign addr[13123]= 2028233973;
assign addr[13124]= 2040479063;
assign addr[13125]= 2052076975;
assign addr[13126]= 2063024031;
assign addr[13127]= 2073316760;
assign addr[13128]= 2082951896;
assign addr[13129]= 2091926384;
assign addr[13130]= 2100237377;
assign addr[13131]= 2107882239;
assign addr[13132]= 2114858546;
assign addr[13133]= 2121164085;
assign addr[13134]= 2126796855;
assign addr[13135]= 2131755071;
assign addr[13136]= 2136037160;
assign addr[13137]= 2139641764;
assign addr[13138]= 2142567738;
assign addr[13139]= 2144814157;
assign addr[13140]= 2146380306;
assign addr[13141]= 2147265689;
assign addr[13142]= 2147470025;
assign addr[13143]= 2146993250;
assign addr[13144]= 2145835515;
assign addr[13145]= 2143997187;
assign addr[13146]= 2141478848;
assign addr[13147]= 2138281298;
assign addr[13148]= 2134405552;
assign addr[13149]= 2129852837;
assign addr[13150]= 2124624598;
assign addr[13151]= 2118722494;
assign addr[13152]= 2112148396;
assign addr[13153]= 2104904390;
assign addr[13154]= 2096992772;
assign addr[13155]= 2088416053;
assign addr[13156]= 2079176953;
assign addr[13157]= 2069278401;
assign addr[13158]= 2058723538;
assign addr[13159]= 2047515711;
assign addr[13160]= 2035658475;
assign addr[13161]= 2023155591;
assign addr[13162]= 2010011024;
assign addr[13163]= 1996228943;
assign addr[13164]= 1981813720;
assign addr[13165]= 1966769926;
assign addr[13166]= 1951102334;
assign addr[13167]= 1934815911;
assign addr[13168]= 1917915825;
assign addr[13169]= 1900407434;
assign addr[13170]= 1882296293;
assign addr[13171]= 1863588145;
assign addr[13172]= 1844288924;
assign addr[13173]= 1824404752;
assign addr[13174]= 1803941934;
assign addr[13175]= 1782906961;
assign addr[13176]= 1761306505;
assign addr[13177]= 1739147417;
assign addr[13178]= 1716436725;
assign addr[13179]= 1693181631;
assign addr[13180]= 1669389513;
assign addr[13181]= 1645067915;
assign addr[13182]= 1620224553;
assign addr[13183]= 1594867305;
assign addr[13184]= 1569004214;
assign addr[13185]= 1542643483;
assign addr[13186]= 1515793473;
assign addr[13187]= 1488462700;
assign addr[13188]= 1460659832;
assign addr[13189]= 1432393688;
assign addr[13190]= 1403673233;
assign addr[13191]= 1374507575;
assign addr[13192]= 1344905966;
assign addr[13193]= 1314877795;
assign addr[13194]= 1284432584;
assign addr[13195]= 1253579991;
assign addr[13196]= 1222329801;
assign addr[13197]= 1190691925;
assign addr[13198]= 1158676398;
assign addr[13199]= 1126293375;
assign addr[13200]= 1093553126;
assign addr[13201]= 1060466036;
assign addr[13202]= 1027042599;
assign addr[13203]= 993293415;
assign addr[13204]= 959229189;
assign addr[13205]= 924860725;
assign addr[13206]= 890198924;
assign addr[13207]= 855254778;
assign addr[13208]= 820039373;
assign addr[13209]= 784563876;
assign addr[13210]= 748839539;
assign addr[13211]= 712877694;
assign addr[13212]= 676689746;
assign addr[13213]= 640287172;
assign addr[13214]= 603681519;
assign addr[13215]= 566884397;
assign addr[13216]= 529907477;
assign addr[13217]= 492762486;
assign addr[13218]= 455461206;
assign addr[13219]= 418015468;
assign addr[13220]= 380437148;
assign addr[13221]= 342738165;
assign addr[13222]= 304930476;
assign addr[13223]= 267026072;
assign addr[13224]= 229036977;
assign addr[13225]= 190975237;
assign addr[13226]= 152852926;
assign addr[13227]= 114682135;
assign addr[13228]= 76474970;
assign addr[13229]= 38243550;
assign addr[13230]= 0;
assign addr[13231]= -38243550;
assign addr[13232]= -76474970;
assign addr[13233]= -114682135;
assign addr[13234]= -152852926;
assign addr[13235]= -190975237;
assign addr[13236]= -229036977;
assign addr[13237]= -267026072;
assign addr[13238]= -304930476;
assign addr[13239]= -342738165;
assign addr[13240]= -380437148;
assign addr[13241]= -418015468;
assign addr[13242]= -455461206;
assign addr[13243]= -492762486;
assign addr[13244]= -529907477;
assign addr[13245]= -566884397;
assign addr[13246]= -603681519;
assign addr[13247]= -640287172;
assign addr[13248]= -676689746;
assign addr[13249]= -712877694;
assign addr[13250]= -748839539;
assign addr[13251]= -784563876;
assign addr[13252]= -820039373;
assign addr[13253]= -855254778;
assign addr[13254]= -890198924;
assign addr[13255]= -924860725;
assign addr[13256]= -959229189;
assign addr[13257]= -993293415;
assign addr[13258]= -1027042599;
assign addr[13259]= -1060466036;
assign addr[13260]= -1093553126;
assign addr[13261]= -1126293375;
assign addr[13262]= -1158676398;
assign addr[13263]= -1190691925;
assign addr[13264]= -1222329801;
assign addr[13265]= -1253579991;
assign addr[13266]= -1284432584;
assign addr[13267]= -1314877795;
assign addr[13268]= -1344905966;
assign addr[13269]= -1374507575;
assign addr[13270]= -1403673233;
assign addr[13271]= -1432393688;
assign addr[13272]= -1460659832;
assign addr[13273]= -1488462700;
assign addr[13274]= -1515793473;
assign addr[13275]= -1542643483;
assign addr[13276]= -1569004214;
assign addr[13277]= -1594867305;
assign addr[13278]= -1620224553;
assign addr[13279]= -1645067915;
assign addr[13280]= -1669389513;
assign addr[13281]= -1693181631;
assign addr[13282]= -1716436725;
assign addr[13283]= -1739147417;
assign addr[13284]= -1761306505;
assign addr[13285]= -1782906961;
assign addr[13286]= -1803941934;
assign addr[13287]= -1824404752;
assign addr[13288]= -1844288924;
assign addr[13289]= -1863588145;
assign addr[13290]= -1882296293;
assign addr[13291]= -1900407434;
assign addr[13292]= -1917915825;
assign addr[13293]= -1934815911;
assign addr[13294]= -1951102334;
assign addr[13295]= -1966769926;
assign addr[13296]= -1981813720;
assign addr[13297]= -1996228943;
assign addr[13298]= -2010011024;
assign addr[13299]= -2023155591;
assign addr[13300]= -2035658475;
assign addr[13301]= -2047515711;
assign addr[13302]= -2058723538;
assign addr[13303]= -2069278401;
assign addr[13304]= -2079176953;
assign addr[13305]= -2088416053;
assign addr[13306]= -2096992772;
assign addr[13307]= -2104904390;
assign addr[13308]= -2112148396;
assign addr[13309]= -2118722494;
assign addr[13310]= -2124624598;
assign addr[13311]= -2129852837;
assign addr[13312]= -2134405552;
assign addr[13313]= -2138281298;
assign addr[13314]= -2141478848;
assign addr[13315]= -2143997187;
assign addr[13316]= -2145835515;
assign addr[13317]= -2146993250;
assign addr[13318]= -2147470025;
assign addr[13319]= -2147265689;
assign addr[13320]= -2146380306;
assign addr[13321]= -2144814157;
assign addr[13322]= -2142567738;
assign addr[13323]= -2139641764;
assign addr[13324]= -2136037160;
assign addr[13325]= -2131755071;
assign addr[13326]= -2126796855;
assign addr[13327]= -2121164085;
assign addr[13328]= -2114858546;
assign addr[13329]= -2107882239;
assign addr[13330]= -2100237377;
assign addr[13331]= -2091926384;
assign addr[13332]= -2082951896;
assign addr[13333]= -2073316760;
assign addr[13334]= -2063024031;
assign addr[13335]= -2052076975;
assign addr[13336]= -2040479063;
assign addr[13337]= -2028233973;
assign addr[13338]= -2015345591;
assign addr[13339]= -2001818002;
assign addr[13340]= -1987655498;
assign addr[13341]= -1972862571;
assign addr[13342]= -1957443913;
assign addr[13343]= -1941404413;
assign addr[13344]= -1924749160;
assign addr[13345]= -1907483436;
assign addr[13346]= -1889612716;
assign addr[13347]= -1871142669;
assign addr[13348]= -1852079154;
assign addr[13349]= -1832428215;
assign addr[13350]= -1812196087;
assign addr[13351]= -1791389186;
assign addr[13352]= -1770014111;
assign addr[13353]= -1748077642;
assign addr[13354]= -1725586737;
assign addr[13355]= -1702548529;
assign addr[13356]= -1678970324;
assign addr[13357]= -1654859602;
assign addr[13358]= -1630224009;
assign addr[13359]= -1605071359;
assign addr[13360]= -1579409630;
assign addr[13361]= -1553246960;
assign addr[13362]= -1526591649;
assign addr[13363]= -1499452149;
assign addr[13364]= -1471837070;
assign addr[13365]= -1443755168;
assign addr[13366]= -1415215352;
assign addr[13367]= -1386226674;
assign addr[13368]= -1356798326;
assign addr[13369]= -1326939644;
assign addr[13370]= -1296660098;
assign addr[13371]= -1265969291;
assign addr[13372]= -1234876957;
assign addr[13373]= -1203392958;
assign addr[13374]= -1171527280;
assign addr[13375]= -1139290029;
assign addr[13376]= -1106691431;
assign addr[13377]= -1073741824;
assign addr[13378]= -1040451659;
assign addr[13379]= -1006831495;
assign addr[13380]= -972891995;
assign addr[13381]= -938643924;
assign addr[13382]= -904098143;
assign addr[13383]= -869265610;
assign addr[13384]= -834157373;
assign addr[13385]= -798784567;
assign addr[13386]= -763158411;
assign addr[13387]= -727290205;
assign addr[13388]= -691191324;
assign addr[13389]= -654873219;
assign addr[13390]= -618347408;
assign addr[13391]= -581625477;
assign addr[13392]= -544719071;
assign addr[13393]= -507639898;
assign addr[13394]= -470399716;
assign addr[13395]= -433010339;
assign addr[13396]= -395483624;
assign addr[13397]= -357831473;
assign addr[13398]= -320065829;
assign addr[13399]= -282198671;
assign addr[13400]= -244242007;
assign addr[13401]= -206207878;
assign addr[13402]= -168108346;
assign addr[13403]= -129955495;
assign addr[13404]= -91761426;
assign addr[13405]= -53538253;
assign addr[13406]= -15298099;
assign addr[13407]= 22946906;
assign addr[13408]= 61184634;
assign addr[13409]= 99402956;
assign addr[13410]= 137589750;
assign addr[13411]= 175732905;
assign addr[13412]= 213820322;
assign addr[13413]= 251839923;
assign addr[13414]= 289779648;
assign addr[13415]= 327627463;
assign addr[13416]= 365371365;
assign addr[13417]= 402999383;
assign addr[13418]= 440499581;
assign addr[13419]= 477860067;
assign addr[13420]= 515068990;
assign addr[13421]= 552114549;
assign addr[13422]= 588984994;
assign addr[13423]= 625668632;
assign addr[13424]= 662153826;
assign addr[13425]= 698429006;
assign addr[13426]= 734482665;
assign addr[13427]= 770303369;
assign addr[13428]= 805879757;
assign addr[13429]= 841200544;
assign addr[13430]= 876254528;
assign addr[13431]= 911030591;
assign addr[13432]= 945517704;
assign addr[13433]= 979704927;
assign addr[13434]= 1013581418;
assign addr[13435]= 1047136432;
assign addr[13436]= 1080359326;
assign addr[13437]= 1113239564;
assign addr[13438]= 1145766716;
assign addr[13439]= 1177930466;
assign addr[13440]= 1209720613;
assign addr[13441]= 1241127074;
assign addr[13442]= 1272139887;
assign addr[13443]= 1302749217;
assign addr[13444]= 1332945355;
assign addr[13445]= 1362718723;
assign addr[13446]= 1392059879;
assign addr[13447]= 1420959516;
assign addr[13448]= 1449408469;
assign addr[13449]= 1477397714;
assign addr[13450]= 1504918373;
assign addr[13451]= 1531961719;
assign addr[13452]= 1558519173;
assign addr[13453]= 1584582314;
assign addr[13454]= 1610142873;
assign addr[13455]= 1635192744;
assign addr[13456]= 1659723983;
assign addr[13457]= 1683728808;
assign addr[13458]= 1707199606;
assign addr[13459]= 1730128933;
assign addr[13460]= 1752509516;
assign addr[13461]= 1774334257;
assign addr[13462]= 1795596234;
assign addr[13463]= 1816288703;
assign addr[13464]= 1836405100;
assign addr[13465]= 1855939047;
assign addr[13466]= 1874884346;
assign addr[13467]= 1893234990;
assign addr[13468]= 1910985158;
assign addr[13469]= 1928129220;
assign addr[13470]= 1944661739;
assign addr[13471]= 1960577471;
assign addr[13472]= 1975871368;
assign addr[13473]= 1990538579;
assign addr[13474]= 2004574453;
assign addr[13475]= 2017974537;
assign addr[13476]= 2030734582;
assign addr[13477]= 2042850540;
assign addr[13478]= 2054318569;
assign addr[13479]= 2065135031;
assign addr[13480]= 2075296495;
assign addr[13481]= 2084799740;
assign addr[13482]= 2093641749;
assign addr[13483]= 2101819720;
assign addr[13484]= 2109331059;
assign addr[13485]= 2116173382;
assign addr[13486]= 2122344521;
assign addr[13487]= 2127842516;
assign addr[13488]= 2132665626;
assign addr[13489]= 2136812319;
assign addr[13490]= 2140281282;
assign addr[13491]= 2143071413;
assign addr[13492]= 2145181827;
assign addr[13493]= 2146611856;
assign addr[13494]= 2147361045;
assign addr[13495]= 2147429158;
assign addr[13496]= 2146816171;
assign addr[13497]= 2145522281;
assign addr[13498]= 2143547897;
assign addr[13499]= 2140893646;
assign addr[13500]= 2137560369;
assign addr[13501]= 2133549123;
assign addr[13502]= 2128861181;
assign addr[13503]= 2123498030;
assign addr[13504]= 2117461370;
assign addr[13505]= 2110753117;
assign addr[13506]= 2103375398;
assign addr[13507]= 2095330553;
assign addr[13508]= 2086621133;
assign addr[13509]= 2077249901;
assign addr[13510]= 2067219829;
assign addr[13511]= 2056534099;
assign addr[13512]= 2045196100;
assign addr[13513]= 2033209426;
assign addr[13514]= 2020577882;
assign addr[13515]= 2007305472;
assign addr[13516]= 1993396407;
assign addr[13517]= 1978855097;
assign addr[13518]= 1963686155;
assign addr[13519]= 1947894393;
assign addr[13520]= 1931484818;
assign addr[13521]= 1914462636;
assign addr[13522]= 1896833245;
assign addr[13523]= 1878602237;
assign addr[13524]= 1859775393;
assign addr[13525]= 1840358687;
assign addr[13526]= 1820358275;
assign addr[13527]= 1799780501;
assign addr[13528]= 1778631892;
assign addr[13529]= 1756919156;
assign addr[13530]= 1734649179;
assign addr[13531]= 1711829025;
assign addr[13532]= 1688465931;
assign addr[13533]= 1664567307;
assign addr[13534]= 1640140734;
assign addr[13535]= 1615193959;
assign addr[13536]= 1589734894;
assign addr[13537]= 1563771613;
assign addr[13538]= 1537312353;
assign addr[13539]= 1510365504;
assign addr[13540]= 1482939614;
assign addr[13541]= 1455043381;
assign addr[13542]= 1426685652;
assign addr[13543]= 1397875423;
assign addr[13544]= 1368621831;
assign addr[13545]= 1338934154;
assign addr[13546]= 1308821808;
assign addr[13547]= 1278294345;
assign addr[13548]= 1247361445;
assign addr[13549]= 1216032921;
assign addr[13550]= 1184318708;
assign addr[13551]= 1152228866;
assign addr[13552]= 1119773573;
assign addr[13553]= 1086963121;
assign addr[13554]= 1053807919;
assign addr[13555]= 1020318481;
assign addr[13556]= 986505429;
assign addr[13557]= 952379488;
assign addr[13558]= 917951481;
assign addr[13559]= 883232329;
assign addr[13560]= 848233042;
assign addr[13561]= 812964722;
assign addr[13562]= 777438554;
assign addr[13563]= 741665807;
assign addr[13564]= 705657826;
assign addr[13565]= 669426032;
assign addr[13566]= 632981917;
assign addr[13567]= 596337040;
assign addr[13568]= 559503022;
assign addr[13569]= 522491548;
assign addr[13570]= 485314355;
assign addr[13571]= 447983235;
assign addr[13572]= 410510029;
assign addr[13573]= 372906622;
assign addr[13574]= 335184940;
assign addr[13575]= 297356948;
assign addr[13576]= 259434643;
assign addr[13577]= 221430054;
assign addr[13578]= 183355234;
assign addr[13579]= 145222259;
assign addr[13580]= 107043224;
assign addr[13581]= 68830239;
assign addr[13582]= 30595422;
assign addr[13583]= -7649098;
assign addr[13584]= -45891193;
assign addr[13585]= -84118732;
assign addr[13586]= -122319591;
assign addr[13587]= -160481654;
assign addr[13588]= -198592817;
assign addr[13589]= -236640993;
assign addr[13590]= -274614114;
assign addr[13591]= -312500135;
assign addr[13592]= -350287041;
assign addr[13593]= -387962847;
assign addr[13594]= -425515602;
assign addr[13595]= -462933398;
assign addr[13596]= -500204365;
assign addr[13597]= -537316682;
assign addr[13598]= -574258580;
assign addr[13599]= -611018340;
assign addr[13600]= -647584304;
assign addr[13601]= -683944874;
assign addr[13602]= -720088517;
assign addr[13603]= -756003771;
assign addr[13604]= -791679244;
assign addr[13605]= -827103620;
assign addr[13606]= -862265664;
assign addr[13607]= -897154224;
assign addr[13608]= -931758235;
assign addr[13609]= -966066720;
assign addr[13610]= -1000068799;
assign addr[13611]= -1033753687;
assign addr[13612]= -1067110699;
assign addr[13613]= -1100129257;
assign addr[13614]= -1132798888;
assign addr[13615]= -1165109230;
assign addr[13616]= -1197050035;
assign addr[13617]= -1228611172;
assign addr[13618]= -1259782632;
assign addr[13619]= -1290554528;
assign addr[13620]= -1320917099;
assign addr[13621]= -1350860716;
assign addr[13622]= -1380375881;
assign addr[13623]= -1409453233;
assign addr[13624]= -1438083551;
assign addr[13625]= -1466257752;
assign addr[13626]= -1493966902;
assign addr[13627]= -1521202211;
assign addr[13628]= -1547955041;
assign addr[13629]= -1574216908;
assign addr[13630]= -1599979481;
assign addr[13631]= -1625234591;
assign addr[13632]= -1649974225;
assign addr[13633]= -1674190539;
assign addr[13634]= -1697875851;
assign addr[13635]= -1721022648;
assign addr[13636]= -1743623590;
assign addr[13637]= -1765671509;
assign addr[13638]= -1787159411;
assign addr[13639]= -1808080480;
assign addr[13640]= -1828428082;
assign addr[13641]= -1848195763;
assign addr[13642]= -1867377253;
assign addr[13643]= -1885966468;
assign addr[13644]= -1903957513;
assign addr[13645]= -1921344681;
assign addr[13646]= -1938122457;
assign addr[13647]= -1954285520;
assign addr[13648]= -1969828744;
assign addr[13649]= -1984747199;
assign addr[13650]= -1999036154;
assign addr[13651]= -2012691075;
assign addr[13652]= -2025707632;
assign addr[13653]= -2038081698;
assign addr[13654]= -2049809346;
assign addr[13655]= -2060886858;
assign addr[13656]= -2071310720;
assign addr[13657]= -2081077626;
assign addr[13658]= -2090184478;
assign addr[13659]= -2098628387;
assign addr[13660]= -2106406677;
assign addr[13661]= -2113516878;
assign addr[13662]= -2119956737;
assign addr[13663]= -2125724211;
assign addr[13664]= -2130817471;
assign addr[13665]= -2135234901;
assign addr[13666]= -2138975100;
assign addr[13667]= -2142036881;
assign addr[13668]= -2144419275;
assign addr[13669]= -2146121524;
assign addr[13670]= -2147143090;
assign addr[13671]= -2147483648;
assign addr[13672]= -2147143090;
assign addr[13673]= -2146121524;
assign addr[13674]= -2144419275;
assign addr[13675]= -2142036881;
assign addr[13676]= -2138975100;
assign addr[13677]= -2135234901;
assign addr[13678]= -2130817471;
assign addr[13679]= -2125724211;
assign addr[13680]= -2119956737;
assign addr[13681]= -2113516878;
assign addr[13682]= -2106406677;
assign addr[13683]= -2098628387;
assign addr[13684]= -2090184478;
assign addr[13685]= -2081077626;
assign addr[13686]= -2071310720;
assign addr[13687]= -2060886858;
assign addr[13688]= -2049809346;
assign addr[13689]= -2038081698;
assign addr[13690]= -2025707632;
assign addr[13691]= -2012691075;
assign addr[13692]= -1999036154;
assign addr[13693]= -1984747199;
assign addr[13694]= -1969828744;
assign addr[13695]= -1954285520;
assign addr[13696]= -1938122457;
assign addr[13697]= -1921344681;
assign addr[13698]= -1903957513;
assign addr[13699]= -1885966468;
assign addr[13700]= -1867377253;
assign addr[13701]= -1848195763;
assign addr[13702]= -1828428082;
assign addr[13703]= -1808080480;
assign addr[13704]= -1787159411;
assign addr[13705]= -1765671509;
assign addr[13706]= -1743623590;
assign addr[13707]= -1721022648;
assign addr[13708]= -1697875851;
assign addr[13709]= -1674190539;
assign addr[13710]= -1649974225;
assign addr[13711]= -1625234591;
assign addr[13712]= -1599979481;
assign addr[13713]= -1574216908;
assign addr[13714]= -1547955041;
assign addr[13715]= -1521202211;
assign addr[13716]= -1493966902;
assign addr[13717]= -1466257752;
assign addr[13718]= -1438083551;
assign addr[13719]= -1409453233;
assign addr[13720]= -1380375881;
assign addr[13721]= -1350860716;
assign addr[13722]= -1320917099;
assign addr[13723]= -1290554528;
assign addr[13724]= -1259782632;
assign addr[13725]= -1228611172;
assign addr[13726]= -1197050035;
assign addr[13727]= -1165109230;
assign addr[13728]= -1132798888;
assign addr[13729]= -1100129257;
assign addr[13730]= -1067110699;
assign addr[13731]= -1033753687;
assign addr[13732]= -1000068799;
assign addr[13733]= -966066720;
assign addr[13734]= -931758235;
assign addr[13735]= -897154224;
assign addr[13736]= -862265664;
assign addr[13737]= -827103620;
assign addr[13738]= -791679244;
assign addr[13739]= -756003771;
assign addr[13740]= -720088517;
assign addr[13741]= -683944874;
assign addr[13742]= -647584304;
assign addr[13743]= -611018340;
assign addr[13744]= -574258580;
assign addr[13745]= -537316682;
assign addr[13746]= -500204365;
assign addr[13747]= -462933398;
assign addr[13748]= -425515602;
assign addr[13749]= -387962847;
assign addr[13750]= -350287041;
assign addr[13751]= -312500135;
assign addr[13752]= -274614114;
assign addr[13753]= -236640993;
assign addr[13754]= -198592817;
assign addr[13755]= -160481654;
assign addr[13756]= -122319591;
assign addr[13757]= -84118732;
assign addr[13758]= -45891193;
assign addr[13759]= -7649098;
assign addr[13760]= 30595422;
assign addr[13761]= 68830239;
assign addr[13762]= 107043224;
assign addr[13763]= 145222259;
assign addr[13764]= 183355234;
assign addr[13765]= 221430054;
assign addr[13766]= 259434643;
assign addr[13767]= 297356948;
assign addr[13768]= 335184940;
assign addr[13769]= 372906622;
assign addr[13770]= 410510029;
assign addr[13771]= 447983235;
assign addr[13772]= 485314355;
assign addr[13773]= 522491548;
assign addr[13774]= 559503022;
assign addr[13775]= 596337040;
assign addr[13776]= 632981917;
assign addr[13777]= 669426032;
assign addr[13778]= 705657826;
assign addr[13779]= 741665807;
assign addr[13780]= 777438554;
assign addr[13781]= 812964722;
assign addr[13782]= 848233042;
assign addr[13783]= 883232329;
assign addr[13784]= 917951481;
assign addr[13785]= 952379488;
assign addr[13786]= 986505429;
assign addr[13787]= 1020318481;
assign addr[13788]= 1053807919;
assign addr[13789]= 1086963121;
assign addr[13790]= 1119773573;
assign addr[13791]= 1152228866;
assign addr[13792]= 1184318708;
assign addr[13793]= 1216032921;
assign addr[13794]= 1247361445;
assign addr[13795]= 1278294345;
assign addr[13796]= 1308821808;
assign addr[13797]= 1338934154;
assign addr[13798]= 1368621831;
assign addr[13799]= 1397875423;
assign addr[13800]= 1426685652;
assign addr[13801]= 1455043381;
assign addr[13802]= 1482939614;
assign addr[13803]= 1510365504;
assign addr[13804]= 1537312353;
assign addr[13805]= 1563771613;
assign addr[13806]= 1589734894;
assign addr[13807]= 1615193959;
assign addr[13808]= 1640140734;
assign addr[13809]= 1664567307;
assign addr[13810]= 1688465931;
assign addr[13811]= 1711829025;
assign addr[13812]= 1734649179;
assign addr[13813]= 1756919156;
assign addr[13814]= 1778631892;
assign addr[13815]= 1799780501;
assign addr[13816]= 1820358275;
assign addr[13817]= 1840358687;
assign addr[13818]= 1859775393;
assign addr[13819]= 1878602237;
assign addr[13820]= 1896833245;
assign addr[13821]= 1914462636;
assign addr[13822]= 1931484818;
assign addr[13823]= 1947894393;
assign addr[13824]= 1963686155;
assign addr[13825]= 1978855097;
assign addr[13826]= 1993396407;
assign addr[13827]= 2007305472;
assign addr[13828]= 2020577882;
assign addr[13829]= 2033209426;
assign addr[13830]= 2045196100;
assign addr[13831]= 2056534099;
assign addr[13832]= 2067219829;
assign addr[13833]= 2077249901;
assign addr[13834]= 2086621133;
assign addr[13835]= 2095330553;
assign addr[13836]= 2103375398;
assign addr[13837]= 2110753117;
assign addr[13838]= 2117461370;
assign addr[13839]= 2123498030;
assign addr[13840]= 2128861181;
assign addr[13841]= 2133549123;
assign addr[13842]= 2137560369;
assign addr[13843]= 2140893646;
assign addr[13844]= 2143547897;
assign addr[13845]= 2145522281;
assign addr[13846]= 2146816171;
assign addr[13847]= 2147429158;
assign addr[13848]= 2147361045;
assign addr[13849]= 2146611856;
assign addr[13850]= 2145181827;
assign addr[13851]= 2143071413;
assign addr[13852]= 2140281282;
assign addr[13853]= 2136812319;
assign addr[13854]= 2132665626;
assign addr[13855]= 2127842516;
assign addr[13856]= 2122344521;
assign addr[13857]= 2116173382;
assign addr[13858]= 2109331059;
assign addr[13859]= 2101819720;
assign addr[13860]= 2093641749;
assign addr[13861]= 2084799740;
assign addr[13862]= 2075296495;
assign addr[13863]= 2065135031;
assign addr[13864]= 2054318569;
assign addr[13865]= 2042850540;
assign addr[13866]= 2030734582;
assign addr[13867]= 2017974537;
assign addr[13868]= 2004574453;
assign addr[13869]= 1990538579;
assign addr[13870]= 1975871368;
assign addr[13871]= 1960577471;
assign addr[13872]= 1944661739;
assign addr[13873]= 1928129220;
assign addr[13874]= 1910985158;
assign addr[13875]= 1893234990;
assign addr[13876]= 1874884346;
assign addr[13877]= 1855939047;
assign addr[13878]= 1836405100;
assign addr[13879]= 1816288703;
assign addr[13880]= 1795596234;
assign addr[13881]= 1774334257;
assign addr[13882]= 1752509516;
assign addr[13883]= 1730128933;
assign addr[13884]= 1707199606;
assign addr[13885]= 1683728808;
assign addr[13886]= 1659723983;
assign addr[13887]= 1635192744;
assign addr[13888]= 1610142873;
assign addr[13889]= 1584582314;
assign addr[13890]= 1558519173;
assign addr[13891]= 1531961719;
assign addr[13892]= 1504918373;
assign addr[13893]= 1477397714;
assign addr[13894]= 1449408469;
assign addr[13895]= 1420959516;
assign addr[13896]= 1392059879;
assign addr[13897]= 1362718723;
assign addr[13898]= 1332945355;
assign addr[13899]= 1302749217;
assign addr[13900]= 1272139887;
assign addr[13901]= 1241127074;
assign addr[13902]= 1209720613;
assign addr[13903]= 1177930466;
assign addr[13904]= 1145766716;
assign addr[13905]= 1113239564;
assign addr[13906]= 1080359326;
assign addr[13907]= 1047136432;
assign addr[13908]= 1013581418;
assign addr[13909]= 979704927;
assign addr[13910]= 945517704;
assign addr[13911]= 911030591;
assign addr[13912]= 876254528;
assign addr[13913]= 841200544;
assign addr[13914]= 805879757;
assign addr[13915]= 770303369;
assign addr[13916]= 734482665;
assign addr[13917]= 698429006;
assign addr[13918]= 662153826;
assign addr[13919]= 625668632;
assign addr[13920]= 588984994;
assign addr[13921]= 552114549;
assign addr[13922]= 515068990;
assign addr[13923]= 477860067;
assign addr[13924]= 440499581;
assign addr[13925]= 402999383;
assign addr[13926]= 365371365;
assign addr[13927]= 327627463;
assign addr[13928]= 289779648;
assign addr[13929]= 251839923;
assign addr[13930]= 213820322;
assign addr[13931]= 175732905;
assign addr[13932]= 137589750;
assign addr[13933]= 99402956;
assign addr[13934]= 61184634;
assign addr[13935]= 22946906;
assign addr[13936]= -15298099;
assign addr[13937]= -53538253;
assign addr[13938]= -91761426;
assign addr[13939]= -129955495;
assign addr[13940]= -168108346;
assign addr[13941]= -206207878;
assign addr[13942]= -244242007;
assign addr[13943]= -282198671;
assign addr[13944]= -320065829;
assign addr[13945]= -357831473;
assign addr[13946]= -395483624;
assign addr[13947]= -433010339;
assign addr[13948]= -470399716;
assign addr[13949]= -507639898;
assign addr[13950]= -544719071;
assign addr[13951]= -581625477;
assign addr[13952]= -618347408;
assign addr[13953]= -654873219;
assign addr[13954]= -691191324;
assign addr[13955]= -727290205;
assign addr[13956]= -763158411;
assign addr[13957]= -798784567;
assign addr[13958]= -834157373;
assign addr[13959]= -869265610;
assign addr[13960]= -904098143;
assign addr[13961]= -938643924;
assign addr[13962]= -972891995;
assign addr[13963]= -1006831495;
assign addr[13964]= -1040451659;
assign addr[13965]= -1073741824;
assign addr[13966]= -1106691431;
assign addr[13967]= -1139290029;
assign addr[13968]= -1171527280;
assign addr[13969]= -1203392958;
assign addr[13970]= -1234876957;
assign addr[13971]= -1265969291;
assign addr[13972]= -1296660098;
assign addr[13973]= -1326939644;
assign addr[13974]= -1356798326;
assign addr[13975]= -1386226674;
assign addr[13976]= -1415215352;
assign addr[13977]= -1443755168;
assign addr[13978]= -1471837070;
assign addr[13979]= -1499452149;
assign addr[13980]= -1526591649;
assign addr[13981]= -1553246960;
assign addr[13982]= -1579409630;
assign addr[13983]= -1605071359;
assign addr[13984]= -1630224009;
assign addr[13985]= -1654859602;
assign addr[13986]= -1678970324;
assign addr[13987]= -1702548529;
assign addr[13988]= -1725586737;
assign addr[13989]= -1748077642;
assign addr[13990]= -1770014111;
assign addr[13991]= -1791389186;
assign addr[13992]= -1812196087;
assign addr[13993]= -1832428215;
assign addr[13994]= -1852079154;
assign addr[13995]= -1871142669;
assign addr[13996]= -1889612716;
assign addr[13997]= -1907483436;
assign addr[13998]= -1924749160;
assign addr[13999]= -1941404413;
assign addr[14000]= -1957443913;
assign addr[14001]= -1972862571;
assign addr[14002]= -1987655498;
assign addr[14003]= -2001818002;
assign addr[14004]= -2015345591;
assign addr[14005]= -2028233973;
assign addr[14006]= -2040479063;
assign addr[14007]= -2052076975;
assign addr[14008]= -2063024031;
assign addr[14009]= -2073316760;
assign addr[14010]= -2082951896;
assign addr[14011]= -2091926384;
assign addr[14012]= -2100237377;
assign addr[14013]= -2107882239;
assign addr[14014]= -2114858546;
assign addr[14015]= -2121164085;
assign addr[14016]= -2126796855;
assign addr[14017]= -2131755071;
assign addr[14018]= -2136037160;
assign addr[14019]= -2139641764;
assign addr[14020]= -2142567738;
assign addr[14021]= -2144814157;
assign addr[14022]= -2146380306;
assign addr[14023]= -2147265689;
assign addr[14024]= -2147470025;
assign addr[14025]= -2146993250;
assign addr[14026]= -2145835515;
assign addr[14027]= -2143997187;
assign addr[14028]= -2141478848;
assign addr[14029]= -2138281298;
assign addr[14030]= -2134405552;
assign addr[14031]= -2129852837;
assign addr[14032]= -2124624598;
assign addr[14033]= -2118722494;
assign addr[14034]= -2112148396;
assign addr[14035]= -2104904390;
assign addr[14036]= -2096992772;
assign addr[14037]= -2088416053;
assign addr[14038]= -2079176953;
assign addr[14039]= -2069278401;
assign addr[14040]= -2058723538;
assign addr[14041]= -2047515711;
assign addr[14042]= -2035658475;
assign addr[14043]= -2023155591;
assign addr[14044]= -2010011024;
assign addr[14045]= -1996228943;
assign addr[14046]= -1981813720;
assign addr[14047]= -1966769926;
assign addr[14048]= -1951102334;
assign addr[14049]= -1934815911;
assign addr[14050]= -1917915825;
assign addr[14051]= -1900407434;
assign addr[14052]= -1882296293;
assign addr[14053]= -1863588145;
assign addr[14054]= -1844288924;
assign addr[14055]= -1824404752;
assign addr[14056]= -1803941934;
assign addr[14057]= -1782906961;
assign addr[14058]= -1761306505;
assign addr[14059]= -1739147417;
assign addr[14060]= -1716436725;
assign addr[14061]= -1693181631;
assign addr[14062]= -1669389513;
assign addr[14063]= -1645067915;
assign addr[14064]= -1620224553;
assign addr[14065]= -1594867305;
assign addr[14066]= -1569004214;
assign addr[14067]= -1542643483;
assign addr[14068]= -1515793473;
assign addr[14069]= -1488462700;
assign addr[14070]= -1460659832;
assign addr[14071]= -1432393688;
assign addr[14072]= -1403673233;
assign addr[14073]= -1374507575;
assign addr[14074]= -1344905966;
assign addr[14075]= -1314877795;
assign addr[14076]= -1284432584;
assign addr[14077]= -1253579991;
assign addr[14078]= -1222329801;
assign addr[14079]= -1190691925;
assign addr[14080]= -1158676398;
assign addr[14081]= -1126293375;
assign addr[14082]= -1093553126;
assign addr[14083]= -1060466036;
assign addr[14084]= -1027042599;
assign addr[14085]= -993293415;
assign addr[14086]= -959229189;
assign addr[14087]= -924860725;
assign addr[14088]= -890198924;
assign addr[14089]= -855254778;
assign addr[14090]= -820039373;
assign addr[14091]= -784563876;
assign addr[14092]= -748839539;
assign addr[14093]= -712877694;
assign addr[14094]= -676689746;
assign addr[14095]= -640287172;
assign addr[14096]= -603681519;
assign addr[14097]= -566884397;
assign addr[14098]= -529907477;
assign addr[14099]= -492762486;
assign addr[14100]= -455461206;
assign addr[14101]= -418015468;
assign addr[14102]= -380437148;
assign addr[14103]= -342738165;
assign addr[14104]= -304930476;
assign addr[14105]= -267026072;
assign addr[14106]= -229036977;
assign addr[14107]= -190975237;
assign addr[14108]= -152852926;
assign addr[14109]= -114682135;
assign addr[14110]= -76474970;
assign addr[14111]= -38243550;
assign addr[14112]= 0;
assign addr[14113]= 38243550;
assign addr[14114]= 76474970;
assign addr[14115]= 114682135;
assign addr[14116]= 152852926;
assign addr[14117]= 190975237;
assign addr[14118]= 229036977;
assign addr[14119]= 267026072;
assign addr[14120]= 304930476;
assign addr[14121]= 342738165;
assign addr[14122]= 380437148;
assign addr[14123]= 418015468;
assign addr[14124]= 455461206;
assign addr[14125]= 492762486;
assign addr[14126]= 529907477;
assign addr[14127]= 566884397;
assign addr[14128]= 603681519;
assign addr[14129]= 640287172;
assign addr[14130]= 676689746;
assign addr[14131]= 712877694;
assign addr[14132]= 748839539;
assign addr[14133]= 784563876;
assign addr[14134]= 820039373;
assign addr[14135]= 855254778;
assign addr[14136]= 890198924;
assign addr[14137]= 924860725;
assign addr[14138]= 959229189;
assign addr[14139]= 993293415;
assign addr[14140]= 1027042599;
assign addr[14141]= 1060466036;
assign addr[14142]= 1093553126;
assign addr[14143]= 1126293375;
assign addr[14144]= 1158676398;
assign addr[14145]= 1190691925;
assign addr[14146]= 1222329801;
assign addr[14147]= 1253579991;
assign addr[14148]= 1284432584;
assign addr[14149]= 1314877795;
assign addr[14150]= 1344905966;
assign addr[14151]= 1374507575;
assign addr[14152]= 1403673233;
assign addr[14153]= 1432393688;
assign addr[14154]= 1460659832;
assign addr[14155]= 1488462700;
assign addr[14156]= 1515793473;
assign addr[14157]= 1542643483;
assign addr[14158]= 1569004214;
assign addr[14159]= 1594867305;
assign addr[14160]= 1620224553;
assign addr[14161]= 1645067915;
assign addr[14162]= 1669389513;
assign addr[14163]= 1693181631;
assign addr[14164]= 1716436725;
assign addr[14165]= 1739147417;
assign addr[14166]= 1761306505;
assign addr[14167]= 1782906961;
assign addr[14168]= 1803941934;
assign addr[14169]= 1824404752;
assign addr[14170]= 1844288924;
assign addr[14171]= 1863588145;
assign addr[14172]= 1882296293;
assign addr[14173]= 1900407434;
assign addr[14174]= 1917915825;
assign addr[14175]= 1934815911;
assign addr[14176]= 1951102334;
assign addr[14177]= 1966769926;
assign addr[14178]= 1981813720;
assign addr[14179]= 1996228943;
assign addr[14180]= 2010011024;
assign addr[14181]= 2023155591;
assign addr[14182]= 2035658475;
assign addr[14183]= 2047515711;
assign addr[14184]= 2058723538;
assign addr[14185]= 2069278401;
assign addr[14186]= 2079176953;
assign addr[14187]= 2088416053;
assign addr[14188]= 2096992772;
assign addr[14189]= 2104904390;
assign addr[14190]= 2112148396;
assign addr[14191]= 2118722494;
assign addr[14192]= 2124624598;
assign addr[14193]= 2129852837;
assign addr[14194]= 2134405552;
assign addr[14195]= 2138281298;
assign addr[14196]= 2141478848;
assign addr[14197]= 2143997187;
assign addr[14198]= 2145835515;
assign addr[14199]= 2146993250;
assign addr[14200]= 2147470025;
assign addr[14201]= 2147265689;
assign addr[14202]= 2146380306;
assign addr[14203]= 2144814157;
assign addr[14204]= 2142567738;
assign addr[14205]= 2139641764;
assign addr[14206]= 2136037160;
assign addr[14207]= 2131755071;
assign addr[14208]= 2126796855;
assign addr[14209]= 2121164085;
assign addr[14210]= 2114858546;
assign addr[14211]= 2107882239;
assign addr[14212]= 2100237377;
assign addr[14213]= 2091926384;
assign addr[14214]= 2082951896;
assign addr[14215]= 2073316760;
assign addr[14216]= 2063024031;
assign addr[14217]= 2052076975;
assign addr[14218]= 2040479063;
assign addr[14219]= 2028233973;
assign addr[14220]= 2015345591;
assign addr[14221]= 2001818002;
assign addr[14222]= 1987655498;
assign addr[14223]= 1972862571;
assign addr[14224]= 1957443913;
assign addr[14225]= 1941404413;
assign addr[14226]= 1924749160;
assign addr[14227]= 1907483436;
assign addr[14228]= 1889612716;
assign addr[14229]= 1871142669;
assign addr[14230]= 1852079154;
assign addr[14231]= 1832428215;
assign addr[14232]= 1812196087;
assign addr[14233]= 1791389186;
assign addr[14234]= 1770014111;
assign addr[14235]= 1748077642;
assign addr[14236]= 1725586737;
assign addr[14237]= 1702548529;
assign addr[14238]= 1678970324;
assign addr[14239]= 1654859602;
assign addr[14240]= 1630224009;
assign addr[14241]= 1605071359;
assign addr[14242]= 1579409630;
assign addr[14243]= 1553246960;
assign addr[14244]= 1526591649;
assign addr[14245]= 1499452149;
assign addr[14246]= 1471837070;
assign addr[14247]= 1443755168;
assign addr[14248]= 1415215352;
assign addr[14249]= 1386226674;
assign addr[14250]= 1356798326;
assign addr[14251]= 1326939644;
assign addr[14252]= 1296660098;
assign addr[14253]= 1265969291;
assign addr[14254]= 1234876957;
assign addr[14255]= 1203392958;
assign addr[14256]= 1171527280;
assign addr[14257]= 1139290029;
assign addr[14258]= 1106691431;
assign addr[14259]= 1073741824;
assign addr[14260]= 1040451659;
assign addr[14261]= 1006831495;
assign addr[14262]= 972891995;
assign addr[14263]= 938643924;
assign addr[14264]= 904098143;
assign addr[14265]= 869265610;
assign addr[14266]= 834157373;
assign addr[14267]= 798784567;
assign addr[14268]= 763158411;
assign addr[14269]= 727290205;
assign addr[14270]= 691191324;
assign addr[14271]= 654873219;
assign addr[14272]= 618347408;
assign addr[14273]= 581625477;
assign addr[14274]= 544719071;
assign addr[14275]= 507639898;
assign addr[14276]= 470399716;
assign addr[14277]= 433010339;
assign addr[14278]= 395483624;
assign addr[14279]= 357831473;
assign addr[14280]= 320065829;
assign addr[14281]= 282198671;
assign addr[14282]= 244242007;
assign addr[14283]= 206207878;
assign addr[14284]= 168108346;
assign addr[14285]= 129955495;
assign addr[14286]= 91761426;
assign addr[14287]= 53538253;
assign addr[14288]= 15298099;
assign addr[14289]= -22946906;
assign addr[14290]= -61184634;
assign addr[14291]= -99402956;
assign addr[14292]= -137589750;
assign addr[14293]= -175732905;
assign addr[14294]= -213820322;
assign addr[14295]= -251839923;
assign addr[14296]= -289779648;
assign addr[14297]= -327627463;
assign addr[14298]= -365371365;
assign addr[14299]= -402999383;
assign addr[14300]= -440499581;
assign addr[14301]= -477860067;
assign addr[14302]= -515068990;
assign addr[14303]= -552114549;
assign addr[14304]= -588984994;
assign addr[14305]= -625668632;
assign addr[14306]= -662153826;
assign addr[14307]= -698429006;
assign addr[14308]= -734482665;
assign addr[14309]= -770303369;
assign addr[14310]= -805879757;
assign addr[14311]= -841200544;
assign addr[14312]= -876254528;
assign addr[14313]= -911030591;
assign addr[14314]= -945517704;
assign addr[14315]= -979704927;
assign addr[14316]= -1013581418;
assign addr[14317]= -1047136432;
assign addr[14318]= -1080359326;
assign addr[14319]= -1113239564;
assign addr[14320]= -1145766716;
assign addr[14321]= -1177930466;
assign addr[14322]= -1209720613;
assign addr[14323]= -1241127074;
assign addr[14324]= -1272139887;
assign addr[14325]= -1302749217;
assign addr[14326]= -1332945355;
assign addr[14327]= -1362718723;
assign addr[14328]= -1392059879;
assign addr[14329]= -1420959516;
assign addr[14330]= -1449408469;
assign addr[14331]= -1477397714;
assign addr[14332]= -1504918373;
assign addr[14333]= -1531961719;
assign addr[14334]= -1558519173;
assign addr[14335]= -1584582314;
assign addr[14336]= -1610142873;
assign addr[14337]= -1635192744;
assign addr[14338]= -1659723983;
assign addr[14339]= -1683728808;
assign addr[14340]= -1707199606;
assign addr[14341]= -1730128933;
assign addr[14342]= -1752509516;
assign addr[14343]= -1774334257;
assign addr[14344]= -1795596234;
assign addr[14345]= -1816288703;
assign addr[14346]= -1836405100;
assign addr[14347]= -1855939047;
assign addr[14348]= -1874884346;
assign addr[14349]= -1893234990;
assign addr[14350]= -1910985158;
assign addr[14351]= -1928129220;
assign addr[14352]= -1944661739;
assign addr[14353]= -1960577471;
assign addr[14354]= -1975871368;
assign addr[14355]= -1990538579;
assign addr[14356]= -2004574453;
assign addr[14357]= -2017974537;
assign addr[14358]= -2030734582;
assign addr[14359]= -2042850540;
assign addr[14360]= -2054318569;
assign addr[14361]= -2065135031;
assign addr[14362]= -2075296495;
assign addr[14363]= -2084799740;
assign addr[14364]= -2093641749;
assign addr[14365]= -2101819720;
assign addr[14366]= -2109331059;
assign addr[14367]= -2116173382;
assign addr[14368]= -2122344521;
assign addr[14369]= -2127842516;
assign addr[14370]= -2132665626;
assign addr[14371]= -2136812319;
assign addr[14372]= -2140281282;
assign addr[14373]= -2143071413;
assign addr[14374]= -2145181827;
assign addr[14375]= -2146611856;
assign addr[14376]= -2147361045;
assign addr[14377]= -2147429158;
assign addr[14378]= -2146816171;
assign addr[14379]= -2145522281;
assign addr[14380]= -2143547897;
assign addr[14381]= -2140893646;
assign addr[14382]= -2137560369;
assign addr[14383]= -2133549123;
assign addr[14384]= -2128861181;
assign addr[14385]= -2123498030;
assign addr[14386]= -2117461370;
assign addr[14387]= -2110753117;
assign addr[14388]= -2103375398;
assign addr[14389]= -2095330553;
assign addr[14390]= -2086621133;
assign addr[14391]= -2077249901;
assign addr[14392]= -2067219829;
assign addr[14393]= -2056534099;
assign addr[14394]= -2045196100;
assign addr[14395]= -2033209426;
assign addr[14396]= -2020577882;
assign addr[14397]= -2007305472;
assign addr[14398]= -1993396407;
assign addr[14399]= -1978855097;
assign addr[14400]= -1963686155;
assign addr[14401]= -1947894393;
assign addr[14402]= -1931484818;
assign addr[14403]= -1914462636;
assign addr[14404]= -1896833245;
assign addr[14405]= -1878602237;
assign addr[14406]= -1859775393;
assign addr[14407]= -1840358687;
assign addr[14408]= -1820358275;
assign addr[14409]= -1799780501;
assign addr[14410]= -1778631892;
assign addr[14411]= -1756919156;
assign addr[14412]= -1734649179;
assign addr[14413]= -1711829025;
assign addr[14414]= -1688465931;
assign addr[14415]= -1664567307;
assign addr[14416]= -1640140734;
assign addr[14417]= -1615193959;
assign addr[14418]= -1589734894;
assign addr[14419]= -1563771613;
assign addr[14420]= -1537312353;
assign addr[14421]= -1510365504;
assign addr[14422]= -1482939614;
assign addr[14423]= -1455043381;
assign addr[14424]= -1426685652;
assign addr[14425]= -1397875423;
assign addr[14426]= -1368621831;
assign addr[14427]= -1338934154;
assign addr[14428]= -1308821808;
assign addr[14429]= -1278294345;
assign addr[14430]= -1247361445;
assign addr[14431]= -1216032921;
assign addr[14432]= -1184318708;
assign addr[14433]= -1152228866;
assign addr[14434]= -1119773573;
assign addr[14435]= -1086963121;
assign addr[14436]= -1053807919;
assign addr[14437]= -1020318481;
assign addr[14438]= -986505429;
assign addr[14439]= -952379488;
assign addr[14440]= -917951481;
assign addr[14441]= -883232329;
assign addr[14442]= -848233042;
assign addr[14443]= -812964722;
assign addr[14444]= -777438554;
assign addr[14445]= -741665807;
assign addr[14446]= -705657826;
assign addr[14447]= -669426032;
assign addr[14448]= -632981917;
assign addr[14449]= -596337040;
assign addr[14450]= -559503022;
assign addr[14451]= -522491548;
assign addr[14452]= -485314355;
assign addr[14453]= -447983235;
assign addr[14454]= -410510029;
assign addr[14455]= -372906622;
assign addr[14456]= -335184940;
assign addr[14457]= -297356948;
assign addr[14458]= -259434643;
assign addr[14459]= -221430054;
assign addr[14460]= -183355234;
assign addr[14461]= -145222259;
assign addr[14462]= -107043224;
assign addr[14463]= -68830239;
assign addr[14464]= -30595422;
assign addr[14465]= 7649098;
assign addr[14466]= 45891193;
assign addr[14467]= 84118732;
assign addr[14468]= 122319591;
assign addr[14469]= 160481654;
assign addr[14470]= 198592817;
assign addr[14471]= 236640993;
assign addr[14472]= 274614114;
assign addr[14473]= 312500135;
assign addr[14474]= 350287041;
assign addr[14475]= 387962847;
assign addr[14476]= 425515602;
assign addr[14477]= 462933398;
assign addr[14478]= 500204365;
assign addr[14479]= 537316682;
assign addr[14480]= 574258580;
assign addr[14481]= 611018340;
assign addr[14482]= 647584304;
assign addr[14483]= 683944874;
assign addr[14484]= 720088517;
assign addr[14485]= 756003771;
assign addr[14486]= 791679244;
assign addr[14487]= 827103620;
assign addr[14488]= 862265664;
assign addr[14489]= 897154224;
assign addr[14490]= 931758235;
assign addr[14491]= 966066720;
assign addr[14492]= 1000068799;
assign addr[14493]= 1033753687;
assign addr[14494]= 1067110699;
assign addr[14495]= 1100129257;
assign addr[14496]= 1132798888;
assign addr[14497]= 1165109230;
assign addr[14498]= 1197050035;
assign addr[14499]= 1228611172;
assign addr[14500]= 1259782632;
assign addr[14501]= 1290554528;
assign addr[14502]= 1320917099;
assign addr[14503]= 1350860716;
assign addr[14504]= 1380375881;
assign addr[14505]= 1409453233;
assign addr[14506]= 1438083551;
assign addr[14507]= 1466257752;
assign addr[14508]= 1493966902;
assign addr[14509]= 1521202211;
assign addr[14510]= 1547955041;
assign addr[14511]= 1574216908;
assign addr[14512]= 1599979481;
assign addr[14513]= 1625234591;
assign addr[14514]= 1649974225;
assign addr[14515]= 1674190539;
assign addr[14516]= 1697875851;
assign addr[14517]= 1721022648;
assign addr[14518]= 1743623590;
assign addr[14519]= 1765671509;
assign addr[14520]= 1787159411;
assign addr[14521]= 1808080480;
assign addr[14522]= 1828428082;
assign addr[14523]= 1848195763;
assign addr[14524]= 1867377253;
assign addr[14525]= 1885966468;
assign addr[14526]= 1903957513;
assign addr[14527]= 1921344681;
assign addr[14528]= 1938122457;
assign addr[14529]= 1954285520;
assign addr[14530]= 1969828744;
assign addr[14531]= 1984747199;
assign addr[14532]= 1999036154;
assign addr[14533]= 2012691075;
assign addr[14534]= 2025707632;
assign addr[14535]= 2038081698;
assign addr[14536]= 2049809346;
assign addr[14537]= 2060886858;
assign addr[14538]= 2071310720;
assign addr[14539]= 2081077626;
assign addr[14540]= 2090184478;
assign addr[14541]= 2098628387;
assign addr[14542]= 2106406677;
assign addr[14543]= 2113516878;
assign addr[14544]= 2119956737;
assign addr[14545]= 2125724211;
assign addr[14546]= 2130817471;
assign addr[14547]= 2135234901;
assign addr[14548]= 2138975100;
assign addr[14549]= 2142036881;
assign addr[14550]= 2144419275;
assign addr[14551]= 2146121524;
assign addr[14552]= 2147143090;
assign addr[14553]= 2147483648;
assign addr[14554]= 2147143090;
assign addr[14555]= 2146121524;
assign addr[14556]= 2144419275;
assign addr[14557]= 2142036881;
assign addr[14558]= 2138975100;
assign addr[14559]= 2135234901;
assign addr[14560]= 2130817471;
assign addr[14561]= 2125724211;
assign addr[14562]= 2119956737;
assign addr[14563]= 2113516878;
assign addr[14564]= 2106406677;
assign addr[14565]= 2098628387;
assign addr[14566]= 2090184478;
assign addr[14567]= 2081077626;
assign addr[14568]= 2071310720;
assign addr[14569]= 2060886858;
assign addr[14570]= 2049809346;
assign addr[14571]= 2038081698;
assign addr[14572]= 2025707632;
assign addr[14573]= 2012691075;
assign addr[14574]= 1999036154;
assign addr[14575]= 1984747199;
assign addr[14576]= 1969828744;
assign addr[14577]= 1954285520;
assign addr[14578]= 1938122457;
assign addr[14579]= 1921344681;
assign addr[14580]= 1903957513;
assign addr[14581]= 1885966468;
assign addr[14582]= 1867377253;
assign addr[14583]= 1848195763;
assign addr[14584]= 1828428082;
assign addr[14585]= 1808080480;
assign addr[14586]= 1787159411;
assign addr[14587]= 1765671509;
assign addr[14588]= 1743623590;
assign addr[14589]= 1721022648;
assign addr[14590]= 1697875851;
assign addr[14591]= 1674190539;
assign addr[14592]= 1649974225;
assign addr[14593]= 1625234591;
assign addr[14594]= 1599979481;
assign addr[14595]= 1574216908;
assign addr[14596]= 1547955041;
assign addr[14597]= 1521202211;
assign addr[14598]= 1493966902;
assign addr[14599]= 1466257752;
assign addr[14600]= 1438083551;
assign addr[14601]= 1409453233;
assign addr[14602]= 1380375881;
assign addr[14603]= 1350860716;
assign addr[14604]= 1320917099;
assign addr[14605]= 1290554528;
assign addr[14606]= 1259782632;
assign addr[14607]= 1228611172;
assign addr[14608]= 1197050035;
assign addr[14609]= 1165109230;
assign addr[14610]= 1132798888;
assign addr[14611]= 1100129257;
assign addr[14612]= 1067110699;
assign addr[14613]= 1033753687;
assign addr[14614]= 1000068799;
assign addr[14615]= 966066720;
assign addr[14616]= 931758235;
assign addr[14617]= 897154224;
assign addr[14618]= 862265664;
assign addr[14619]= 827103620;
assign addr[14620]= 791679244;
assign addr[14621]= 756003771;
assign addr[14622]= 720088517;
assign addr[14623]= 683944874;
assign addr[14624]= 647584304;
assign addr[14625]= 611018340;
assign addr[14626]= 574258580;
assign addr[14627]= 537316682;
assign addr[14628]= 500204365;
assign addr[14629]= 462933398;
assign addr[14630]= 425515602;
assign addr[14631]= 387962847;
assign addr[14632]= 350287041;
assign addr[14633]= 312500135;
assign addr[14634]= 274614114;
assign addr[14635]= 236640993;
assign addr[14636]= 198592817;
assign addr[14637]= 160481654;
assign addr[14638]= 122319591;
assign addr[14639]= 84118732;
assign addr[14640]= 45891193;
assign addr[14641]= 7649098;
assign addr[14642]= -30595422;
assign addr[14643]= -68830239;
assign addr[14644]= -107043224;
assign addr[14645]= -145222259;
assign addr[14646]= -183355234;
assign addr[14647]= -221430054;
assign addr[14648]= -259434643;
assign addr[14649]= -297356948;
assign addr[14650]= -335184940;
assign addr[14651]= -372906622;
assign addr[14652]= -410510029;
assign addr[14653]= -447983235;
assign addr[14654]= -485314355;
assign addr[14655]= -522491548;
assign addr[14656]= -559503022;
assign addr[14657]= -596337040;
assign addr[14658]= -632981917;
assign addr[14659]= -669426032;
assign addr[14660]= -705657826;
assign addr[14661]= -741665807;
assign addr[14662]= -777438554;
assign addr[14663]= -812964722;
assign addr[14664]= -848233042;
assign addr[14665]= -883232329;
assign addr[14666]= -917951481;
assign addr[14667]= -952379488;
assign addr[14668]= -986505429;
assign addr[14669]= -1020318481;
assign addr[14670]= -1053807919;
assign addr[14671]= -1086963121;
assign addr[14672]= -1119773573;
assign addr[14673]= -1152228866;
assign addr[14674]= -1184318708;
assign addr[14675]= -1216032921;
assign addr[14676]= -1247361445;
assign addr[14677]= -1278294345;
assign addr[14678]= -1308821808;
assign addr[14679]= -1338934154;
assign addr[14680]= -1368621831;
assign addr[14681]= -1397875423;
assign addr[14682]= -1426685652;
assign addr[14683]= -1455043381;
assign addr[14684]= -1482939614;
assign addr[14685]= -1510365504;
assign addr[14686]= -1537312353;
assign addr[14687]= -1563771613;
assign addr[14688]= -1589734894;
assign addr[14689]= -1615193959;
assign addr[14690]= -1640140734;
assign addr[14691]= -1664567307;
assign addr[14692]= -1688465931;
assign addr[14693]= -1711829025;
assign addr[14694]= -1734649179;
assign addr[14695]= -1756919156;
assign addr[14696]= -1778631892;
assign addr[14697]= -1799780501;
assign addr[14698]= -1820358275;
assign addr[14699]= -1840358687;
assign addr[14700]= -1859775393;
assign addr[14701]= -1878602237;
assign addr[14702]= -1896833245;
assign addr[14703]= -1914462636;
assign addr[14704]= -1931484818;
assign addr[14705]= -1947894393;
assign addr[14706]= -1963686155;
assign addr[14707]= -1978855097;
assign addr[14708]= -1993396407;
assign addr[14709]= -2007305472;
assign addr[14710]= -2020577882;
assign addr[14711]= -2033209426;
assign addr[14712]= -2045196100;
assign addr[14713]= -2056534099;
assign addr[14714]= -2067219829;
assign addr[14715]= -2077249901;
assign addr[14716]= -2086621133;
assign addr[14717]= -2095330553;
assign addr[14718]= -2103375398;
assign addr[14719]= -2110753117;
assign addr[14720]= -2117461370;
assign addr[14721]= -2123498030;
assign addr[14722]= -2128861181;
assign addr[14723]= -2133549123;
assign addr[14724]= -2137560369;
assign addr[14725]= -2140893646;
assign addr[14726]= -2143547897;
assign addr[14727]= -2145522281;
assign addr[14728]= -2146816171;
assign addr[14729]= -2147429158;
assign addr[14730]= -2147361045;
assign addr[14731]= -2146611856;
assign addr[14732]= -2145181827;
assign addr[14733]= -2143071413;
assign addr[14734]= -2140281282;
assign addr[14735]= -2136812319;
assign addr[14736]= -2132665626;
assign addr[14737]= -2127842516;
assign addr[14738]= -2122344521;
assign addr[14739]= -2116173382;
assign addr[14740]= -2109331059;
assign addr[14741]= -2101819720;
assign addr[14742]= -2093641749;
assign addr[14743]= -2084799740;
assign addr[14744]= -2075296495;
assign addr[14745]= -2065135031;
assign addr[14746]= -2054318569;
assign addr[14747]= -2042850540;
assign addr[14748]= -2030734582;
assign addr[14749]= -2017974537;
assign addr[14750]= -2004574453;
assign addr[14751]= -1990538579;
assign addr[14752]= -1975871368;
assign addr[14753]= -1960577471;
assign addr[14754]= -1944661739;
assign addr[14755]= -1928129220;
assign addr[14756]= -1910985158;
assign addr[14757]= -1893234990;
assign addr[14758]= -1874884346;
assign addr[14759]= -1855939047;
assign addr[14760]= -1836405100;
assign addr[14761]= -1816288703;
assign addr[14762]= -1795596234;
assign addr[14763]= -1774334257;
assign addr[14764]= -1752509516;
assign addr[14765]= -1730128933;
assign addr[14766]= -1707199606;
assign addr[14767]= -1683728808;
assign addr[14768]= -1659723983;
assign addr[14769]= -1635192744;
assign addr[14770]= -1610142873;
assign addr[14771]= -1584582314;
assign addr[14772]= -1558519173;
assign addr[14773]= -1531961719;
assign addr[14774]= -1504918373;
assign addr[14775]= -1477397714;
assign addr[14776]= -1449408469;
assign addr[14777]= -1420959516;
assign addr[14778]= -1392059879;
assign addr[14779]= -1362718723;
assign addr[14780]= -1332945355;
assign addr[14781]= -1302749217;
assign addr[14782]= -1272139887;
assign addr[14783]= -1241127074;
assign addr[14784]= -1209720613;
assign addr[14785]= -1177930466;
assign addr[14786]= -1145766716;
assign addr[14787]= -1113239564;
assign addr[14788]= -1080359326;
assign addr[14789]= -1047136432;
assign addr[14790]= -1013581418;
assign addr[14791]= -979704927;
assign addr[14792]= -945517704;
assign addr[14793]= -911030591;
assign addr[14794]= -876254528;
assign addr[14795]= -841200544;
assign addr[14796]= -805879757;
assign addr[14797]= -770303369;
assign addr[14798]= -734482665;
assign addr[14799]= -698429006;
assign addr[14800]= -662153826;
assign addr[14801]= -625668632;
assign addr[14802]= -588984994;
assign addr[14803]= -552114549;
assign addr[14804]= -515068990;
assign addr[14805]= -477860067;
assign addr[14806]= -440499581;
assign addr[14807]= -402999383;
assign addr[14808]= -365371365;
assign addr[14809]= -327627463;
assign addr[14810]= -289779648;
assign addr[14811]= -251839923;
assign addr[14812]= -213820322;
assign addr[14813]= -175732905;
assign addr[14814]= -137589750;
assign addr[14815]= -99402956;
assign addr[14816]= -61184634;
assign addr[14817]= -22946906;
assign addr[14818]= 15298099;
assign addr[14819]= 53538253;
assign addr[14820]= 91761426;
assign addr[14821]= 129955495;
assign addr[14822]= 168108346;
assign addr[14823]= 206207878;
assign addr[14824]= 244242007;
assign addr[14825]= 282198671;
assign addr[14826]= 320065829;
assign addr[14827]= 357831473;
assign addr[14828]= 395483624;
assign addr[14829]= 433010339;
assign addr[14830]= 470399716;
assign addr[14831]= 507639898;
assign addr[14832]= 544719071;
assign addr[14833]= 581625477;
assign addr[14834]= 618347408;
assign addr[14835]= 654873219;
assign addr[14836]= 691191324;
assign addr[14837]= 727290205;
assign addr[14838]= 763158411;
assign addr[14839]= 798784567;
assign addr[14840]= 834157373;
assign addr[14841]= 869265610;
assign addr[14842]= 904098143;
assign addr[14843]= 938643924;
assign addr[14844]= 972891995;
assign addr[14845]= 1006831495;
assign addr[14846]= 1040451659;
assign addr[14847]= 1073741824;
assign addr[14848]= 1106691431;
assign addr[14849]= 1139290029;
assign addr[14850]= 1171527280;
assign addr[14851]= 1203392958;
assign addr[14852]= 1234876957;
assign addr[14853]= 1265969291;
assign addr[14854]= 1296660098;
assign addr[14855]= 1326939644;
assign addr[14856]= 1356798326;
assign addr[14857]= 1386226674;
assign addr[14858]= 1415215352;
assign addr[14859]= 1443755168;
assign addr[14860]= 1471837070;
assign addr[14861]= 1499452149;
assign addr[14862]= 1526591649;
assign addr[14863]= 1553246960;
assign addr[14864]= 1579409630;
assign addr[14865]= 1605071359;
assign addr[14866]= 1630224009;
assign addr[14867]= 1654859602;
assign addr[14868]= 1678970324;
assign addr[14869]= 1702548529;
assign addr[14870]= 1725586737;
assign addr[14871]= 1748077642;
assign addr[14872]= 1770014111;
assign addr[14873]= 1791389186;
assign addr[14874]= 1812196087;
assign addr[14875]= 1832428215;
assign addr[14876]= 1852079154;
assign addr[14877]= 1871142669;
assign addr[14878]= 1889612716;
assign addr[14879]= 1907483436;
assign addr[14880]= 1924749160;
assign addr[14881]= 1941404413;
assign addr[14882]= 1957443913;
assign addr[14883]= 1972862571;
assign addr[14884]= 1987655498;
assign addr[14885]= 2001818002;
assign addr[14886]= 2015345591;
assign addr[14887]= 2028233973;
assign addr[14888]= 2040479063;
assign addr[14889]= 2052076975;
assign addr[14890]= 2063024031;
assign addr[14891]= 2073316760;
assign addr[14892]= 2082951896;
assign addr[14893]= 2091926384;
assign addr[14894]= 2100237377;
assign addr[14895]= 2107882239;
assign addr[14896]= 2114858546;
assign addr[14897]= 2121164085;
assign addr[14898]= 2126796855;
assign addr[14899]= 2131755071;
assign addr[14900]= 2136037160;
assign addr[14901]= 2139641764;
assign addr[14902]= 2142567738;
assign addr[14903]= 2144814157;
assign addr[14904]= 2146380306;
assign addr[14905]= 2147265689;
assign addr[14906]= 2147470025;
assign addr[14907]= 2146993250;
assign addr[14908]= 2145835515;
assign addr[14909]= 2143997187;
assign addr[14910]= 2141478848;
assign addr[14911]= 2138281298;
assign addr[14912]= 2134405552;
assign addr[14913]= 2129852837;
assign addr[14914]= 2124624598;
assign addr[14915]= 2118722494;
assign addr[14916]= 2112148396;
assign addr[14917]= 2104904390;
assign addr[14918]= 2096992772;
assign addr[14919]= 2088416053;
assign addr[14920]= 2079176953;
assign addr[14921]= 2069278401;
assign addr[14922]= 2058723538;
assign addr[14923]= 2047515711;
assign addr[14924]= 2035658475;
assign addr[14925]= 2023155591;
assign addr[14926]= 2010011024;
assign addr[14927]= 1996228943;
assign addr[14928]= 1981813720;
assign addr[14929]= 1966769926;
assign addr[14930]= 1951102334;
assign addr[14931]= 1934815911;
assign addr[14932]= 1917915825;
assign addr[14933]= 1900407434;
assign addr[14934]= 1882296293;
assign addr[14935]= 1863588145;
assign addr[14936]= 1844288924;
assign addr[14937]= 1824404752;
assign addr[14938]= 1803941934;
assign addr[14939]= 1782906961;
assign addr[14940]= 1761306505;
assign addr[14941]= 1739147417;
assign addr[14942]= 1716436725;
assign addr[14943]= 1693181631;
assign addr[14944]= 1669389513;
assign addr[14945]= 1645067915;
assign addr[14946]= 1620224553;
assign addr[14947]= 1594867305;
assign addr[14948]= 1569004214;
assign addr[14949]= 1542643483;
assign addr[14950]= 1515793473;
assign addr[14951]= 1488462700;
assign addr[14952]= 1460659832;
assign addr[14953]= 1432393688;
assign addr[14954]= 1403673233;
assign addr[14955]= 1374507575;
assign addr[14956]= 1344905966;
assign addr[14957]= 1314877795;
assign addr[14958]= 1284432584;
assign addr[14959]= 1253579991;
assign addr[14960]= 1222329801;
assign addr[14961]= 1190691925;
assign addr[14962]= 1158676398;
assign addr[14963]= 1126293375;
assign addr[14964]= 1093553126;
assign addr[14965]= 1060466036;
assign addr[14966]= 1027042599;
assign addr[14967]= 993293415;
assign addr[14968]= 959229189;
assign addr[14969]= 924860725;
assign addr[14970]= 890198924;
assign addr[14971]= 855254778;
assign addr[14972]= 820039373;
assign addr[14973]= 784563876;
assign addr[14974]= 748839539;
assign addr[14975]= 712877694;
assign addr[14976]= 676689746;
assign addr[14977]= 640287172;
assign addr[14978]= 603681519;
assign addr[14979]= 566884397;
assign addr[14980]= 529907477;
assign addr[14981]= 492762486;
assign addr[14982]= 455461206;
assign addr[14983]= 418015468;
assign addr[14984]= 380437148;
assign addr[14985]= 342738165;
assign addr[14986]= 304930476;
assign addr[14987]= 267026072;
assign addr[14988]= 229036977;
assign addr[14989]= 190975237;
assign addr[14990]= 152852926;
assign addr[14991]= 114682135;
assign addr[14992]= 76474970;
assign addr[14993]= 38243550;
assign addr[14994]= 0;
assign addr[14995]= -38243550;
assign addr[14996]= -76474970;
assign addr[14997]= -114682135;
assign addr[14998]= -152852926;
assign addr[14999]= -190975237;
assign addr[15000]= -229036977;
assign addr[15001]= -267026072;
assign addr[15002]= -304930476;
assign addr[15003]= -342738165;
assign addr[15004]= -380437148;
assign addr[15005]= -418015468;
assign addr[15006]= -455461206;
assign addr[15007]= -492762486;
assign addr[15008]= -529907477;
assign addr[15009]= -566884397;
assign addr[15010]= -603681519;
assign addr[15011]= -640287172;
assign addr[15012]= -676689746;
assign addr[15013]= -712877694;
assign addr[15014]= -748839539;
assign addr[15015]= -784563876;
assign addr[15016]= -820039373;
assign addr[15017]= -855254778;
assign addr[15018]= -890198924;
assign addr[15019]= -924860725;
assign addr[15020]= -959229189;
assign addr[15021]= -993293415;
assign addr[15022]= -1027042599;
assign addr[15023]= -1060466036;
assign addr[15024]= -1093553126;
assign addr[15025]= -1126293375;
assign addr[15026]= -1158676398;
assign addr[15027]= -1190691925;
assign addr[15028]= -1222329801;
assign addr[15029]= -1253579991;
assign addr[15030]= -1284432584;
assign addr[15031]= -1314877795;
assign addr[15032]= -1344905966;
assign addr[15033]= -1374507575;
assign addr[15034]= -1403673233;
assign addr[15035]= -1432393688;
assign addr[15036]= -1460659832;
assign addr[15037]= -1488462700;
assign addr[15038]= -1515793473;
assign addr[15039]= -1542643483;
assign addr[15040]= -1569004214;
assign addr[15041]= -1594867305;
assign addr[15042]= -1620224553;
assign addr[15043]= -1645067915;
assign addr[15044]= -1669389513;
assign addr[15045]= -1693181631;
assign addr[15046]= -1716436725;
assign addr[15047]= -1739147417;
assign addr[15048]= -1761306505;
assign addr[15049]= -1782906961;
assign addr[15050]= -1803941934;
assign addr[15051]= -1824404752;
assign addr[15052]= -1844288924;
assign addr[15053]= -1863588145;
assign addr[15054]= -1882296293;
assign addr[15055]= -1900407434;
assign addr[15056]= -1917915825;
assign addr[15057]= -1934815911;
assign addr[15058]= -1951102334;
assign addr[15059]= -1966769926;
assign addr[15060]= -1981813720;
assign addr[15061]= -1996228943;
assign addr[15062]= -2010011024;
assign addr[15063]= -2023155591;
assign addr[15064]= -2035658475;
assign addr[15065]= -2047515711;
assign addr[15066]= -2058723538;
assign addr[15067]= -2069278401;
assign addr[15068]= -2079176953;
assign addr[15069]= -2088416053;
assign addr[15070]= -2096992772;
assign addr[15071]= -2104904390;
assign addr[15072]= -2112148396;
assign addr[15073]= -2118722494;
assign addr[15074]= -2124624598;
assign addr[15075]= -2129852837;
assign addr[15076]= -2134405552;
assign addr[15077]= -2138281298;
assign addr[15078]= -2141478848;
assign addr[15079]= -2143997187;
assign addr[15080]= -2145835515;
assign addr[15081]= -2146993250;
assign addr[15082]= -2147470025;
assign addr[15083]= -2147265689;
assign addr[15084]= -2146380306;
assign addr[15085]= -2144814157;
assign addr[15086]= -2142567738;
assign addr[15087]= -2139641764;
assign addr[15088]= -2136037160;
assign addr[15089]= -2131755071;
assign addr[15090]= -2126796855;
assign addr[15091]= -2121164085;
assign addr[15092]= -2114858546;
assign addr[15093]= -2107882239;
assign addr[15094]= -2100237377;
assign addr[15095]= -2091926384;
assign addr[15096]= -2082951896;
assign addr[15097]= -2073316760;
assign addr[15098]= -2063024031;
assign addr[15099]= -2052076975;
assign addr[15100]= -2040479063;
assign addr[15101]= -2028233973;
assign addr[15102]= -2015345591;
assign addr[15103]= -2001818002;
assign addr[15104]= -1987655498;
assign addr[15105]= -1972862571;
assign addr[15106]= -1957443913;
assign addr[15107]= -1941404413;
assign addr[15108]= -1924749160;
assign addr[15109]= -1907483436;
assign addr[15110]= -1889612716;
assign addr[15111]= -1871142669;
assign addr[15112]= -1852079154;
assign addr[15113]= -1832428215;
assign addr[15114]= -1812196087;
assign addr[15115]= -1791389186;
assign addr[15116]= -1770014111;
assign addr[15117]= -1748077642;
assign addr[15118]= -1725586737;
assign addr[15119]= -1702548529;
assign addr[15120]= -1678970324;
assign addr[15121]= -1654859602;
assign addr[15122]= -1630224009;
assign addr[15123]= -1605071359;
assign addr[15124]= -1579409630;
assign addr[15125]= -1553246960;
assign addr[15126]= -1526591649;
assign addr[15127]= -1499452149;
assign addr[15128]= -1471837070;
assign addr[15129]= -1443755168;
assign addr[15130]= -1415215352;
assign addr[15131]= -1386226674;
assign addr[15132]= -1356798326;
assign addr[15133]= -1326939644;
assign addr[15134]= -1296660098;
assign addr[15135]= -1265969291;
assign addr[15136]= -1234876957;
assign addr[15137]= -1203392958;
assign addr[15138]= -1171527280;
assign addr[15139]= -1139290029;
assign addr[15140]= -1106691431;
assign addr[15141]= -1073741824;
assign addr[15142]= -1040451659;
assign addr[15143]= -1006831495;
assign addr[15144]= -972891995;
assign addr[15145]= -938643924;
assign addr[15146]= -904098143;
assign addr[15147]= -869265610;
assign addr[15148]= -834157373;
assign addr[15149]= -798784567;
assign addr[15150]= -763158411;
assign addr[15151]= -727290205;
assign addr[15152]= -691191324;
assign addr[15153]= -654873219;
assign addr[15154]= -618347408;
assign addr[15155]= -581625477;
assign addr[15156]= -544719071;
assign addr[15157]= -507639898;
assign addr[15158]= -470399716;
assign addr[15159]= -433010339;
assign addr[15160]= -395483624;
assign addr[15161]= -357831473;
assign addr[15162]= -320065829;
assign addr[15163]= -282198671;
assign addr[15164]= -244242007;
assign addr[15165]= -206207878;
assign addr[15166]= -168108346;
assign addr[15167]= -129955495;
assign addr[15168]= -91761426;
assign addr[15169]= -53538253;
assign addr[15170]= -15298099;
assign addr[15171]= 22946906;
assign addr[15172]= 61184634;
assign addr[15173]= 99402956;
assign addr[15174]= 137589750;
assign addr[15175]= 175732905;
assign addr[15176]= 213820322;
assign addr[15177]= 251839923;
assign addr[15178]= 289779648;
assign addr[15179]= 327627463;
assign addr[15180]= 365371365;
assign addr[15181]= 402999383;
assign addr[15182]= 440499581;
assign addr[15183]= 477860067;
assign addr[15184]= 515068990;
assign addr[15185]= 552114549;
assign addr[15186]= 588984994;
assign addr[15187]= 625668632;
assign addr[15188]= 662153826;
assign addr[15189]= 698429006;
assign addr[15190]= 734482665;
assign addr[15191]= 770303369;
assign addr[15192]= 805879757;
assign addr[15193]= 841200544;
assign addr[15194]= 876254528;
assign addr[15195]= 911030591;
assign addr[15196]= 945517704;
assign addr[15197]= 979704927;
assign addr[15198]= 1013581418;
assign addr[15199]= 1047136432;
assign addr[15200]= 1080359326;
assign addr[15201]= 1113239564;
assign addr[15202]= 1145766716;
assign addr[15203]= 1177930466;
assign addr[15204]= 1209720613;
assign addr[15205]= 1241127074;
assign addr[15206]= 1272139887;
assign addr[15207]= 1302749217;
assign addr[15208]= 1332945355;
assign addr[15209]= 1362718723;
assign addr[15210]= 1392059879;
assign addr[15211]= 1420959516;
assign addr[15212]= 1449408469;
assign addr[15213]= 1477397714;
assign addr[15214]= 1504918373;
assign addr[15215]= 1531961719;
assign addr[15216]= 1558519173;
assign addr[15217]= 1584582314;
assign addr[15218]= 1610142873;
assign addr[15219]= 1635192744;
assign addr[15220]= 1659723983;
assign addr[15221]= 1683728808;
assign addr[15222]= 1707199606;
assign addr[15223]= 1730128933;
assign addr[15224]= 1752509516;
assign addr[15225]= 1774334257;
assign addr[15226]= 1795596234;
assign addr[15227]= 1816288703;
assign addr[15228]= 1836405100;
assign addr[15229]= 1855939047;
assign addr[15230]= 1874884346;
assign addr[15231]= 1893234990;
assign addr[15232]= 1910985158;
assign addr[15233]= 1928129220;
assign addr[15234]= 1944661739;
assign addr[15235]= 1960577471;
assign addr[15236]= 1975871368;
assign addr[15237]= 1990538579;
assign addr[15238]= 2004574453;
assign addr[15239]= 2017974537;
assign addr[15240]= 2030734582;
assign addr[15241]= 2042850540;
assign addr[15242]= 2054318569;
assign addr[15243]= 2065135031;
assign addr[15244]= 2075296495;
assign addr[15245]= 2084799740;
assign addr[15246]= 2093641749;
assign addr[15247]= 2101819720;
assign addr[15248]= 2109331059;
assign addr[15249]= 2116173382;
assign addr[15250]= 2122344521;
assign addr[15251]= 2127842516;
assign addr[15252]= 2132665626;
assign addr[15253]= 2136812319;
assign addr[15254]= 2140281282;
assign addr[15255]= 2143071413;
assign addr[15256]= 2145181827;
assign addr[15257]= 2146611856;
assign addr[15258]= 2147361045;
assign addr[15259]= 2147429158;
assign addr[15260]= 2146816171;
assign addr[15261]= 2145522281;
assign addr[15262]= 2143547897;
assign addr[15263]= 2140893646;
assign addr[15264]= 2137560369;
assign addr[15265]= 2133549123;
assign addr[15266]= 2128861181;
assign addr[15267]= 2123498030;
assign addr[15268]= 2117461370;
assign addr[15269]= 2110753117;
assign addr[15270]= 2103375398;
assign addr[15271]= 2095330553;
assign addr[15272]= 2086621133;
assign addr[15273]= 2077249901;
assign addr[15274]= 2067219829;
assign addr[15275]= 2056534099;
assign addr[15276]= 2045196100;
assign addr[15277]= 2033209426;
assign addr[15278]= 2020577882;
assign addr[15279]= 2007305472;
assign addr[15280]= 1993396407;
assign addr[15281]= 1978855097;
assign addr[15282]= 1963686155;
assign addr[15283]= 1947894393;
assign addr[15284]= 1931484818;
assign addr[15285]= 1914462636;
assign addr[15286]= 1896833245;
assign addr[15287]= 1878602237;
assign addr[15288]= 1859775393;
assign addr[15289]= 1840358687;
assign addr[15290]= 1820358275;
assign addr[15291]= 1799780501;
assign addr[15292]= 1778631892;
assign addr[15293]= 1756919156;
assign addr[15294]= 1734649179;
assign addr[15295]= 1711829025;
assign addr[15296]= 1688465931;
assign addr[15297]= 1664567307;
assign addr[15298]= 1640140734;
assign addr[15299]= 1615193959;
assign addr[15300]= 1589734894;
assign addr[15301]= 1563771613;
assign addr[15302]= 1537312353;
assign addr[15303]= 1510365504;
assign addr[15304]= 1482939614;
assign addr[15305]= 1455043381;
assign addr[15306]= 1426685652;
assign addr[15307]= 1397875423;
assign addr[15308]= 1368621831;
assign addr[15309]= 1338934154;
assign addr[15310]= 1308821808;
assign addr[15311]= 1278294345;
assign addr[15312]= 1247361445;
assign addr[15313]= 1216032921;
assign addr[15314]= 1184318708;
assign addr[15315]= 1152228866;
assign addr[15316]= 1119773573;
assign addr[15317]= 1086963121;
assign addr[15318]= 1053807919;
assign addr[15319]= 1020318481;
assign addr[15320]= 986505429;
assign addr[15321]= 952379488;
assign addr[15322]= 917951481;
assign addr[15323]= 883232329;
assign addr[15324]= 848233042;
assign addr[15325]= 812964722;
assign addr[15326]= 777438554;
assign addr[15327]= 741665807;
assign addr[15328]= 705657826;
assign addr[15329]= 669426032;
assign addr[15330]= 632981917;
assign addr[15331]= 596337040;
assign addr[15332]= 559503022;
assign addr[15333]= 522491548;
assign addr[15334]= 485314355;
assign addr[15335]= 447983235;
assign addr[15336]= 410510029;
assign addr[15337]= 372906622;
assign addr[15338]= 335184940;
assign addr[15339]= 297356948;
assign addr[15340]= 259434643;
assign addr[15341]= 221430054;
assign addr[15342]= 183355234;
assign addr[15343]= 145222259;
assign addr[15344]= 107043224;
assign addr[15345]= 68830239;
assign addr[15346]= 30595422;
assign addr[15347]= -7649098;
assign addr[15348]= -45891193;
assign addr[15349]= -84118732;
assign addr[15350]= -122319591;
assign addr[15351]= -160481654;
assign addr[15352]= -198592817;
assign addr[15353]= -236640993;
assign addr[15354]= -274614114;
assign addr[15355]= -312500135;
assign addr[15356]= -350287041;
assign addr[15357]= -387962847;
assign addr[15358]= -425515602;
assign addr[15359]= -462933398;
assign addr[15360]= -500204365;
assign addr[15361]= -537316682;
assign addr[15362]= -574258580;
assign addr[15363]= -611018340;
assign addr[15364]= -647584304;
assign addr[15365]= -683944874;
assign addr[15366]= -720088517;
assign addr[15367]= -756003771;
assign addr[15368]= -791679244;
assign addr[15369]= -827103620;
assign addr[15370]= -862265664;
assign addr[15371]= -897154224;
assign addr[15372]= -931758235;
assign addr[15373]= -966066720;
assign addr[15374]= -1000068799;
assign addr[15375]= -1033753687;
assign addr[15376]= -1067110699;
assign addr[15377]= -1100129257;
assign addr[15378]= -1132798888;
assign addr[15379]= -1165109230;
assign addr[15380]= -1197050035;
assign addr[15381]= -1228611172;
assign addr[15382]= -1259782632;
assign addr[15383]= -1290554528;
assign addr[15384]= -1320917099;
assign addr[15385]= -1350860716;
assign addr[15386]= -1380375881;
assign addr[15387]= -1409453233;
assign addr[15388]= -1438083551;
assign addr[15389]= -1466257752;
assign addr[15390]= -1493966902;
assign addr[15391]= -1521202211;
assign addr[15392]= -1547955041;
assign addr[15393]= -1574216908;
assign addr[15394]= -1599979481;
assign addr[15395]= -1625234591;
assign addr[15396]= -1649974225;
assign addr[15397]= -1674190539;
assign addr[15398]= -1697875851;
assign addr[15399]= -1721022648;
assign addr[15400]= -1743623590;
assign addr[15401]= -1765671509;
assign addr[15402]= -1787159411;
assign addr[15403]= -1808080480;
assign addr[15404]= -1828428082;
assign addr[15405]= -1848195763;
assign addr[15406]= -1867377253;
assign addr[15407]= -1885966468;
assign addr[15408]= -1903957513;
assign addr[15409]= -1921344681;
assign addr[15410]= -1938122457;
assign addr[15411]= -1954285520;
assign addr[15412]= -1969828744;
assign addr[15413]= -1984747199;
assign addr[15414]= -1999036154;
assign addr[15415]= -2012691075;
assign addr[15416]= -2025707632;
assign addr[15417]= -2038081698;
assign addr[15418]= -2049809346;
assign addr[15419]= -2060886858;
assign addr[15420]= -2071310720;
assign addr[15421]= -2081077626;
assign addr[15422]= -2090184478;
assign addr[15423]= -2098628387;
assign addr[15424]= -2106406677;
assign addr[15425]= -2113516878;
assign addr[15426]= -2119956737;
assign addr[15427]= -2125724211;
assign addr[15428]= -2130817471;
assign addr[15429]= -2135234901;
assign addr[15430]= -2138975100;
assign addr[15431]= -2142036881;
assign addr[15432]= -2144419275;
assign addr[15433]= -2146121524;
assign addr[15434]= -2147143090;
assign addr[15435]= -2147483648;
assign addr[15436]= -2147143090;
assign addr[15437]= -2146121524;
assign addr[15438]= -2144419275;
assign addr[15439]= -2142036881;
assign addr[15440]= -2138975100;
assign addr[15441]= -2135234901;
assign addr[15442]= -2130817471;
assign addr[15443]= -2125724211;
assign addr[15444]= -2119956737;
assign addr[15445]= -2113516878;
assign addr[15446]= -2106406677;
assign addr[15447]= -2098628387;
assign addr[15448]= -2090184478;
assign addr[15449]= -2081077626;
assign addr[15450]= -2071310720;
assign addr[15451]= -2060886858;
assign addr[15452]= -2049809346;
assign addr[15453]= -2038081698;
assign addr[15454]= -2025707632;
assign addr[15455]= -2012691075;
assign addr[15456]= -1999036154;
assign addr[15457]= -1984747199;
assign addr[15458]= -1969828744;
assign addr[15459]= -1954285520;
assign addr[15460]= -1938122457;
assign addr[15461]= -1921344681;
assign addr[15462]= -1903957513;
assign addr[15463]= -1885966468;
assign addr[15464]= -1867377253;
assign addr[15465]= -1848195763;
assign addr[15466]= -1828428082;
assign addr[15467]= -1808080480;
assign addr[15468]= -1787159411;
assign addr[15469]= -1765671509;
assign addr[15470]= -1743623590;
assign addr[15471]= -1721022648;
assign addr[15472]= -1697875851;
assign addr[15473]= -1674190539;
assign addr[15474]= -1649974225;
assign addr[15475]= -1625234591;
assign addr[15476]= -1599979481;
assign addr[15477]= -1574216908;
assign addr[15478]= -1547955041;
assign addr[15479]= -1521202211;
assign addr[15480]= -1493966902;
assign addr[15481]= -1466257752;
assign addr[15482]= -1438083551;
assign addr[15483]= -1409453233;
assign addr[15484]= -1380375881;
assign addr[15485]= -1350860716;
assign addr[15486]= -1320917099;
assign addr[15487]= -1290554528;
assign addr[15488]= -1259782632;
assign addr[15489]= -1228611172;
assign addr[15490]= -1197050035;
assign addr[15491]= -1165109230;
assign addr[15492]= -1132798888;
assign addr[15493]= -1100129257;
assign addr[15494]= -1067110699;
assign addr[15495]= -1033753687;
assign addr[15496]= -1000068799;
assign addr[15497]= -966066720;
assign addr[15498]= -931758235;
assign addr[15499]= -897154224;
assign addr[15500]= -862265664;
assign addr[15501]= -827103620;
assign addr[15502]= -791679244;
assign addr[15503]= -756003771;
assign addr[15504]= -720088517;
assign addr[15505]= -683944874;
assign addr[15506]= -647584304;
assign addr[15507]= -611018340;
assign addr[15508]= -574258580;
assign addr[15509]= -537316682;
assign addr[15510]= -500204365;
assign addr[15511]= -462933398;
assign addr[15512]= -425515602;
assign addr[15513]= -387962847;
assign addr[15514]= -350287041;
assign addr[15515]= -312500135;
assign addr[15516]= -274614114;
assign addr[15517]= -236640993;
assign addr[15518]= -198592817;
assign addr[15519]= -160481654;
assign addr[15520]= -122319591;
assign addr[15521]= -84118732;
assign addr[15522]= -45891193;
assign addr[15523]= -7649098;
assign addr[15524]= 30595422;
assign addr[15525]= 68830239;
assign addr[15526]= 107043224;
assign addr[15527]= 145222259;
assign addr[15528]= 183355234;
assign addr[15529]= 221430054;
assign addr[15530]= 259434643;
assign addr[15531]= 297356948;
assign addr[15532]= 335184940;
assign addr[15533]= 372906622;
assign addr[15534]= 410510029;
assign addr[15535]= 447983235;
assign addr[15536]= 485314355;
assign addr[15537]= 522491548;
assign addr[15538]= 559503022;
assign addr[15539]= 596337040;
assign addr[15540]= 632981917;
assign addr[15541]= 669426032;
assign addr[15542]= 705657826;
assign addr[15543]= 741665807;
assign addr[15544]= 777438554;
assign addr[15545]= 812964722;
assign addr[15546]= 848233042;
assign addr[15547]= 883232329;
assign addr[15548]= 917951481;
assign addr[15549]= 952379488;
assign addr[15550]= 986505429;
assign addr[15551]= 1020318481;
assign addr[15552]= 1053807919;
assign addr[15553]= 1086963121;
assign addr[15554]= 1119773573;
assign addr[15555]= 1152228866;
assign addr[15556]= 1184318708;
assign addr[15557]= 1216032921;
assign addr[15558]= 1247361445;
assign addr[15559]= 1278294345;
assign addr[15560]= 1308821808;
assign addr[15561]= 1338934154;
assign addr[15562]= 1368621831;
assign addr[15563]= 1397875423;
assign addr[15564]= 1426685652;
assign addr[15565]= 1455043381;
assign addr[15566]= 1482939614;
assign addr[15567]= 1510365504;
assign addr[15568]= 1537312353;
assign addr[15569]= 1563771613;
assign addr[15570]= 1589734894;
assign addr[15571]= 1615193959;
assign addr[15572]= 1640140734;
assign addr[15573]= 1664567307;
assign addr[15574]= 1688465931;
assign addr[15575]= 1711829025;
assign addr[15576]= 1734649179;
assign addr[15577]= 1756919156;
assign addr[15578]= 1778631892;
assign addr[15579]= 1799780501;
assign addr[15580]= 1820358275;
assign addr[15581]= 1840358687;
assign addr[15582]= 1859775393;
assign addr[15583]= 1878602237;
assign addr[15584]= 1896833245;
assign addr[15585]= 1914462636;
assign addr[15586]= 1931484818;
assign addr[15587]= 1947894393;
assign addr[15588]= 1963686155;
assign addr[15589]= 1978855097;
assign addr[15590]= 1993396407;
assign addr[15591]= 2007305472;
assign addr[15592]= 2020577882;
assign addr[15593]= 2033209426;
assign addr[15594]= 2045196100;
assign addr[15595]= 2056534099;
assign addr[15596]= 2067219829;
assign addr[15597]= 2077249901;
assign addr[15598]= 2086621133;
assign addr[15599]= 2095330553;
assign addr[15600]= 2103375398;
assign addr[15601]= 2110753117;
assign addr[15602]= 2117461370;
assign addr[15603]= 2123498030;
assign addr[15604]= 2128861181;
assign addr[15605]= 2133549123;
assign addr[15606]= 2137560369;
assign addr[15607]= 2140893646;
assign addr[15608]= 2143547897;
assign addr[15609]= 2145522281;
assign addr[15610]= 2146816171;
assign addr[15611]= 2147429158;
assign addr[15612]= 2147361045;
assign addr[15613]= 2146611856;
assign addr[15614]= 2145181827;
assign addr[15615]= 2143071413;
assign addr[15616]= 2140281282;
assign addr[15617]= 2136812319;
assign addr[15618]= 2132665626;
assign addr[15619]= 2127842516;
assign addr[15620]= 2122344521;
assign addr[15621]= 2116173382;
assign addr[15622]= 2109331059;
assign addr[15623]= 2101819720;
assign addr[15624]= 2093641749;
assign addr[15625]= 2084799740;
assign addr[15626]= 2075296495;
assign addr[15627]= 2065135031;
assign addr[15628]= 2054318569;
assign addr[15629]= 2042850540;
assign addr[15630]= 2030734582;
assign addr[15631]= 2017974537;
assign addr[15632]= 2004574453;
assign addr[15633]= 1990538579;
assign addr[15634]= 1975871368;
assign addr[15635]= 1960577471;
assign addr[15636]= 1944661739;
assign addr[15637]= 1928129220;
assign addr[15638]= 1910985158;
assign addr[15639]= 1893234990;
assign addr[15640]= 1874884346;
assign addr[15641]= 1855939047;
assign addr[15642]= 1836405100;
assign addr[15643]= 1816288703;
assign addr[15644]= 1795596234;
assign addr[15645]= 1774334257;
assign addr[15646]= 1752509516;
assign addr[15647]= 1730128933;
assign addr[15648]= 1707199606;
assign addr[15649]= 1683728808;
assign addr[15650]= 1659723983;
assign addr[15651]= 1635192744;
assign addr[15652]= 1610142873;
assign addr[15653]= 1584582314;
assign addr[15654]= 1558519173;
assign addr[15655]= 1531961719;
assign addr[15656]= 1504918373;
assign addr[15657]= 1477397714;
assign addr[15658]= 1449408469;
assign addr[15659]= 1420959516;
assign addr[15660]= 1392059879;
assign addr[15661]= 1362718723;
assign addr[15662]= 1332945355;
assign addr[15663]= 1302749217;
assign addr[15664]= 1272139887;
assign addr[15665]= 1241127074;
assign addr[15666]= 1209720613;
assign addr[15667]= 1177930466;
assign addr[15668]= 1145766716;
assign addr[15669]= 1113239564;
assign addr[15670]= 1080359326;
assign addr[15671]= 1047136432;
assign addr[15672]= 1013581418;
assign addr[15673]= 979704927;
assign addr[15674]= 945517704;
assign addr[15675]= 911030591;
assign addr[15676]= 876254528;
assign addr[15677]= 841200544;
assign addr[15678]= 805879757;
assign addr[15679]= 770303369;
assign addr[15680]= 734482665;
assign addr[15681]= 698429006;
assign addr[15682]= 662153826;
assign addr[15683]= 625668632;
assign addr[15684]= 588984994;
assign addr[15685]= 552114549;
assign addr[15686]= 515068990;
assign addr[15687]= 477860067;
assign addr[15688]= 440499581;
assign addr[15689]= 402999383;
assign addr[15690]= 365371365;
assign addr[15691]= 327627463;
assign addr[15692]= 289779648;
assign addr[15693]= 251839923;
assign addr[15694]= 213820322;
assign addr[15695]= 175732905;
assign addr[15696]= 137589750;
assign addr[15697]= 99402956;
assign addr[15698]= 61184634;
assign addr[15699]= 22946906;
assign addr[15700]= -15298099;
assign addr[15701]= -53538253;
assign addr[15702]= -91761426;
assign addr[15703]= -129955495;
assign addr[15704]= -168108346;
assign addr[15705]= -206207878;
assign addr[15706]= -244242007;
assign addr[15707]= -282198671;
assign addr[15708]= -320065829;
assign addr[15709]= -357831473;
assign addr[15710]= -395483624;
assign addr[15711]= -433010339;
assign addr[15712]= -470399716;
assign addr[15713]= -507639898;
assign addr[15714]= -544719071;
assign addr[15715]= -581625477;
assign addr[15716]= -618347408;
assign addr[15717]= -654873219;
assign addr[15718]= -691191324;
assign addr[15719]= -727290205;
assign addr[15720]= -763158411;
assign addr[15721]= -798784567;
assign addr[15722]= -834157373;
assign addr[15723]= -869265610;
assign addr[15724]= -904098143;
assign addr[15725]= -938643924;
assign addr[15726]= -972891995;
assign addr[15727]= -1006831495;
assign addr[15728]= -1040451659;
assign addr[15729]= -1073741824;
assign addr[15730]= -1106691431;
assign addr[15731]= -1139290029;
assign addr[15732]= -1171527280;
assign addr[15733]= -1203392958;
assign addr[15734]= -1234876957;
assign addr[15735]= -1265969291;
assign addr[15736]= -1296660098;
assign addr[15737]= -1326939644;
assign addr[15738]= -1356798326;
assign addr[15739]= -1386226674;
assign addr[15740]= -1415215352;
assign addr[15741]= -1443755168;
assign addr[15742]= -1471837070;
assign addr[15743]= -1499452149;
assign addr[15744]= -1526591649;
assign addr[15745]= -1553246960;
assign addr[15746]= -1579409630;
assign addr[15747]= -1605071359;
assign addr[15748]= -1630224009;
assign addr[15749]= -1654859602;
assign addr[15750]= -1678970324;
assign addr[15751]= -1702548529;
assign addr[15752]= -1725586737;
assign addr[15753]= -1748077642;
assign addr[15754]= -1770014111;
assign addr[15755]= -1791389186;
assign addr[15756]= -1812196087;
assign addr[15757]= -1832428215;
assign addr[15758]= -1852079154;
assign addr[15759]= -1871142669;
assign addr[15760]= -1889612716;
assign addr[15761]= -1907483436;
assign addr[15762]= -1924749160;
assign addr[15763]= -1941404413;
assign addr[15764]= -1957443913;
assign addr[15765]= -1972862571;
assign addr[15766]= -1987655498;
assign addr[15767]= -2001818002;
assign addr[15768]= -2015345591;
assign addr[15769]= -2028233973;
assign addr[15770]= -2040479063;
assign addr[15771]= -2052076975;
assign addr[15772]= -2063024031;
assign addr[15773]= -2073316760;
assign addr[15774]= -2082951896;
assign addr[15775]= -2091926384;
assign addr[15776]= -2100237377;
assign addr[15777]= -2107882239;
assign addr[15778]= -2114858546;
assign addr[15779]= -2121164085;
assign addr[15780]= -2126796855;
assign addr[15781]= -2131755071;
assign addr[15782]= -2136037160;
assign addr[15783]= -2139641764;
assign addr[15784]= -2142567738;
assign addr[15785]= -2144814157;
assign addr[15786]= -2146380306;
assign addr[15787]= -2147265689;
assign addr[15788]= -2147470025;
assign addr[15789]= -2146993250;
assign addr[15790]= -2145835515;
assign addr[15791]= -2143997187;
assign addr[15792]= -2141478848;
assign addr[15793]= -2138281298;
assign addr[15794]= -2134405552;
assign addr[15795]= -2129852837;
assign addr[15796]= -2124624598;
assign addr[15797]= -2118722494;
assign addr[15798]= -2112148396;
assign addr[15799]= -2104904390;
assign addr[15800]= -2096992772;
assign addr[15801]= -2088416053;
assign addr[15802]= -2079176953;
assign addr[15803]= -2069278401;
assign addr[15804]= -2058723538;
assign addr[15805]= -2047515711;
assign addr[15806]= -2035658475;
assign addr[15807]= -2023155591;
assign addr[15808]= -2010011024;
assign addr[15809]= -1996228943;
assign addr[15810]= -1981813720;
assign addr[15811]= -1966769926;
assign addr[15812]= -1951102334;
assign addr[15813]= -1934815911;
assign addr[15814]= -1917915825;
assign addr[15815]= -1900407434;
assign addr[15816]= -1882296293;
assign addr[15817]= -1863588145;
assign addr[15818]= -1844288924;
assign addr[15819]= -1824404752;
assign addr[15820]= -1803941934;
assign addr[15821]= -1782906961;
assign addr[15822]= -1761306505;
assign addr[15823]= -1739147417;
assign addr[15824]= -1716436725;
assign addr[15825]= -1693181631;
assign addr[15826]= -1669389513;
assign addr[15827]= -1645067915;
assign addr[15828]= -1620224553;
assign addr[15829]= -1594867305;
assign addr[15830]= -1569004214;
assign addr[15831]= -1542643483;
assign addr[15832]= -1515793473;
assign addr[15833]= -1488462700;
assign addr[15834]= -1460659832;
assign addr[15835]= -1432393688;
assign addr[15836]= -1403673233;
assign addr[15837]= -1374507575;
assign addr[15838]= -1344905966;
assign addr[15839]= -1314877795;
assign addr[15840]= -1284432584;
assign addr[15841]= -1253579991;
assign addr[15842]= -1222329801;
assign addr[15843]= -1190691925;
assign addr[15844]= -1158676398;
assign addr[15845]= -1126293375;
assign addr[15846]= -1093553126;
assign addr[15847]= -1060466036;
assign addr[15848]= -1027042599;
assign addr[15849]= -993293415;
assign addr[15850]= -959229189;
assign addr[15851]= -924860725;
assign addr[15852]= -890198924;
assign addr[15853]= -855254778;
assign addr[15854]= -820039373;
assign addr[15855]= -784563876;
assign addr[15856]= -748839539;
assign addr[15857]= -712877694;
assign addr[15858]= -676689746;
assign addr[15859]= -640287172;
assign addr[15860]= -603681519;
assign addr[15861]= -566884397;
assign addr[15862]= -529907477;
assign addr[15863]= -492762486;
assign addr[15864]= -455461206;
assign addr[15865]= -418015468;
assign addr[15866]= -380437148;
assign addr[15867]= -342738165;
assign addr[15868]= -304930476;
assign addr[15869]= -267026072;
assign addr[15870]= -229036977;
assign addr[15871]= -190975237;
assign addr[15872]= -152852926;
assign addr[15873]= -114682135;
assign addr[15874]= -76474970;
assign addr[15875]= -38243550;
assign addr[15876]= 0;
assign addr[15877]= 38243550;
assign addr[15878]= 76474970;
assign addr[15879]= 114682135;
assign addr[15880]= 152852926;
assign addr[15881]= 190975237;
assign addr[15882]= 229036977;
assign addr[15883]= 267026072;
assign addr[15884]= 304930476;
assign addr[15885]= 342738165;
assign addr[15886]= 380437148;
assign addr[15887]= 418015468;
assign addr[15888]= 455461206;
assign addr[15889]= 492762486;
assign addr[15890]= 529907477;
assign addr[15891]= 566884397;
assign addr[15892]= 603681519;
assign addr[15893]= 640287172;
assign addr[15894]= 676689746;
assign addr[15895]= 712877694;
assign addr[15896]= 748839539;
assign addr[15897]= 784563876;
assign addr[15898]= 820039373;
assign addr[15899]= 855254778;
assign addr[15900]= 890198924;
assign addr[15901]= 924860725;
assign addr[15902]= 959229189;
assign addr[15903]= 993293415;
assign addr[15904]= 1027042599;
assign addr[15905]= 1060466036;
assign addr[15906]= 1093553126;
assign addr[15907]= 1126293375;
assign addr[15908]= 1158676398;
assign addr[15909]= 1190691925;
assign addr[15910]= 1222329801;
assign addr[15911]= 1253579991;
assign addr[15912]= 1284432584;
assign addr[15913]= 1314877795;
assign addr[15914]= 1344905966;
assign addr[15915]= 1374507575;
assign addr[15916]= 1403673233;
assign addr[15917]= 1432393688;
assign addr[15918]= 1460659832;
assign addr[15919]= 1488462700;
assign addr[15920]= 1515793473;
assign addr[15921]= 1542643483;
assign addr[15922]= 1569004214;
assign addr[15923]= 1594867305;
assign addr[15924]= 1620224553;
assign addr[15925]= 1645067915;
assign addr[15926]= 1669389513;
assign addr[15927]= 1693181631;
assign addr[15928]= 1716436725;
assign addr[15929]= 1739147417;
assign addr[15930]= 1761306505;
assign addr[15931]= 1782906961;
assign addr[15932]= 1803941934;
assign addr[15933]= 1824404752;
assign addr[15934]= 1844288924;
assign addr[15935]= 1863588145;
assign addr[15936]= 1882296293;
assign addr[15937]= 1900407434;
assign addr[15938]= 1917915825;
assign addr[15939]= 1934815911;
assign addr[15940]= 1951102334;
assign addr[15941]= 1966769926;
assign addr[15942]= 1981813720;
assign addr[15943]= 1996228943;
assign addr[15944]= 2010011024;
assign addr[15945]= 2023155591;
assign addr[15946]= 2035658475;
assign addr[15947]= 2047515711;
assign addr[15948]= 2058723538;
assign addr[15949]= 2069278401;
assign addr[15950]= 2079176953;
assign addr[15951]= 2088416053;
assign addr[15952]= 2096992772;
assign addr[15953]= 2104904390;
assign addr[15954]= 2112148396;
assign addr[15955]= 2118722494;
assign addr[15956]= 2124624598;
assign addr[15957]= 2129852837;
assign addr[15958]= 2134405552;
assign addr[15959]= 2138281298;
assign addr[15960]= 2141478848;
assign addr[15961]= 2143997187;
assign addr[15962]= 2145835515;
assign addr[15963]= 2146993250;
assign addr[15964]= 2147470025;
assign addr[15965]= 2147265689;
assign addr[15966]= 2146380306;
assign addr[15967]= 2144814157;
assign addr[15968]= 2142567738;
assign addr[15969]= 2139641764;
assign addr[15970]= 2136037160;
assign addr[15971]= 2131755071;
assign addr[15972]= 2126796855;
assign addr[15973]= 2121164085;
assign addr[15974]= 2114858546;
assign addr[15975]= 2107882239;
assign addr[15976]= 2100237377;
assign addr[15977]= 2091926384;
assign addr[15978]= 2082951896;
assign addr[15979]= 2073316760;
assign addr[15980]= 2063024031;
assign addr[15981]= 2052076975;
assign addr[15982]= 2040479063;
assign addr[15983]= 2028233973;
assign addr[15984]= 2015345591;
assign addr[15985]= 2001818002;
assign addr[15986]= 1987655498;
assign addr[15987]= 1972862571;
assign addr[15988]= 1957443913;
assign addr[15989]= 1941404413;
assign addr[15990]= 1924749160;
assign addr[15991]= 1907483436;
assign addr[15992]= 1889612716;
assign addr[15993]= 1871142669;
assign addr[15994]= 1852079154;
assign addr[15995]= 1832428215;
assign addr[15996]= 1812196087;
assign addr[15997]= 1791389186;
assign addr[15998]= 1770014111;
assign addr[15999]= 1748077642;
assign addr[16000]= 1725586737;
assign addr[16001]= 1702548529;
assign addr[16002]= 1678970324;
assign addr[16003]= 1654859602;
assign addr[16004]= 1630224009;
assign addr[16005]= 1605071359;
assign addr[16006]= 1579409630;
assign addr[16007]= 1553246960;
assign addr[16008]= 1526591649;
assign addr[16009]= 1499452149;
assign addr[16010]= 1471837070;
assign addr[16011]= 1443755168;
assign addr[16012]= 1415215352;
assign addr[16013]= 1386226674;
assign addr[16014]= 1356798326;
assign addr[16015]= 1326939644;
assign addr[16016]= 1296660098;
assign addr[16017]= 1265969291;
assign addr[16018]= 1234876957;
assign addr[16019]= 1203392958;
assign addr[16020]= 1171527280;
assign addr[16021]= 1139290029;
assign addr[16022]= 1106691431;
assign addr[16023]= 1073741824;
assign addr[16024]= 1040451659;
assign addr[16025]= 1006831495;
assign addr[16026]= 972891995;
assign addr[16027]= 938643924;
assign addr[16028]= 904098143;
assign addr[16029]= 869265610;
assign addr[16030]= 834157373;
assign addr[16031]= 798784567;
assign addr[16032]= 763158411;
assign addr[16033]= 727290205;
assign addr[16034]= 691191324;
assign addr[16035]= 654873219;
assign addr[16036]= 618347408;
assign addr[16037]= 581625477;
assign addr[16038]= 544719071;
assign addr[16039]= 507639898;
assign addr[16040]= 470399716;
assign addr[16041]= 433010339;
assign addr[16042]= 395483624;
assign addr[16043]= 357831473;
assign addr[16044]= 320065829;
assign addr[16045]= 282198671;
assign addr[16046]= 244242007;
assign addr[16047]= 206207878;
assign addr[16048]= 168108346;
assign addr[16049]= 129955495;
assign addr[16050]= 91761426;
assign addr[16051]= 53538253;
assign addr[16052]= 15298099;
assign addr[16053]= -22946906;
assign addr[16054]= -61184634;
assign addr[16055]= -99402956;
assign addr[16056]= -137589750;
assign addr[16057]= -175732905;
assign addr[16058]= -213820322;
assign addr[16059]= -251839923;
assign addr[16060]= -289779648;
assign addr[16061]= -327627463;
assign addr[16062]= -365371365;
assign addr[16063]= -402999383;
assign addr[16064]= -440499581;
assign addr[16065]= -477860067;
assign addr[16066]= -515068990;
assign addr[16067]= -552114549;
assign addr[16068]= -588984994;
assign addr[16069]= -625668632;
assign addr[16070]= -662153826;
assign addr[16071]= -698429006;
assign addr[16072]= -734482665;
assign addr[16073]= -770303369;
assign addr[16074]= -805879757;
assign addr[16075]= -841200544;
assign addr[16076]= -876254528;
assign addr[16077]= -911030591;
assign addr[16078]= -945517704;
assign addr[16079]= -979704927;
assign addr[16080]= -1013581418;
assign addr[16081]= -1047136432;
assign addr[16082]= -1080359326;
assign addr[16083]= -1113239564;
assign addr[16084]= -1145766716;
assign addr[16085]= -1177930466;
assign addr[16086]= -1209720613;
assign addr[16087]= -1241127074;
assign addr[16088]= -1272139887;
assign addr[16089]= -1302749217;
assign addr[16090]= -1332945355;
assign addr[16091]= -1362718723;
assign addr[16092]= -1392059879;
assign addr[16093]= -1420959516;
assign addr[16094]= -1449408469;
assign addr[16095]= -1477397714;
assign addr[16096]= -1504918373;
assign addr[16097]= -1531961719;
assign addr[16098]= -1558519173;
assign addr[16099]= -1584582314;
assign addr[16100]= -1610142873;
assign addr[16101]= -1635192744;
assign addr[16102]= -1659723983;
assign addr[16103]= -1683728808;
assign addr[16104]= -1707199606;
assign addr[16105]= -1730128933;
assign addr[16106]= -1752509516;
assign addr[16107]= -1774334257;
assign addr[16108]= -1795596234;
assign addr[16109]= -1816288703;
assign addr[16110]= -1836405100;
assign addr[16111]= -1855939047;
assign addr[16112]= -1874884346;
assign addr[16113]= -1893234990;
assign addr[16114]= -1910985158;
assign addr[16115]= -1928129220;
assign addr[16116]= -1944661739;
assign addr[16117]= -1960577471;
assign addr[16118]= -1975871368;
assign addr[16119]= -1990538579;
assign addr[16120]= -2004574453;
assign addr[16121]= -2017974537;
assign addr[16122]= -2030734582;
assign addr[16123]= -2042850540;
assign addr[16124]= -2054318569;
assign addr[16125]= -2065135031;
assign addr[16126]= -2075296495;
assign addr[16127]= -2084799740;
assign addr[16128]= -2093641749;
assign addr[16129]= -2101819720;
assign addr[16130]= -2109331059;
assign addr[16131]= -2116173382;
assign addr[16132]= -2122344521;
assign addr[16133]= -2127842516;
assign addr[16134]= -2132665626;
assign addr[16135]= -2136812319;
assign addr[16136]= -2140281282;
assign addr[16137]= -2143071413;
assign addr[16138]= -2145181827;
assign addr[16139]= -2146611856;
assign addr[16140]= -2147361045;
assign addr[16141]= -2147429158;
assign addr[16142]= -2146816171;
assign addr[16143]= -2145522281;
assign addr[16144]= -2143547897;
assign addr[16145]= -2140893646;
assign addr[16146]= -2137560369;
assign addr[16147]= -2133549123;
assign addr[16148]= -2128861181;
assign addr[16149]= -2123498030;
assign addr[16150]= -2117461370;
assign addr[16151]= -2110753117;
assign addr[16152]= -2103375398;
assign addr[16153]= -2095330553;
assign addr[16154]= -2086621133;
assign addr[16155]= -2077249901;
assign addr[16156]= -2067219829;
assign addr[16157]= -2056534099;
assign addr[16158]= -2045196100;
assign addr[16159]= -2033209426;
assign addr[16160]= -2020577882;
assign addr[16161]= -2007305472;
assign addr[16162]= -1993396407;
assign addr[16163]= -1978855097;
assign addr[16164]= -1963686155;
assign addr[16165]= -1947894393;
assign addr[16166]= -1931484818;
assign addr[16167]= -1914462636;
assign addr[16168]= -1896833245;
assign addr[16169]= -1878602237;
assign addr[16170]= -1859775393;
assign addr[16171]= -1840358687;
assign addr[16172]= -1820358275;
assign addr[16173]= -1799780501;
assign addr[16174]= -1778631892;
assign addr[16175]= -1756919156;
assign addr[16176]= -1734649179;
assign addr[16177]= -1711829025;
assign addr[16178]= -1688465931;
assign addr[16179]= -1664567307;
assign addr[16180]= -1640140734;
assign addr[16181]= -1615193959;
assign addr[16182]= -1589734894;
assign addr[16183]= -1563771613;
assign addr[16184]= -1537312353;
assign addr[16185]= -1510365504;
assign addr[16186]= -1482939614;
assign addr[16187]= -1455043381;
assign addr[16188]= -1426685652;
assign addr[16189]= -1397875423;
assign addr[16190]= -1368621831;
assign addr[16191]= -1338934154;
assign addr[16192]= -1308821808;
assign addr[16193]= -1278294345;
assign addr[16194]= -1247361445;
assign addr[16195]= -1216032921;
assign addr[16196]= -1184318708;
assign addr[16197]= -1152228866;
assign addr[16198]= -1119773573;
assign addr[16199]= -1086963121;
assign addr[16200]= -1053807919;
assign addr[16201]= -1020318481;
assign addr[16202]= -986505429;
assign addr[16203]= -952379488;
assign addr[16204]= -917951481;
assign addr[16205]= -883232329;
assign addr[16206]= -848233042;
assign addr[16207]= -812964722;
assign addr[16208]= -777438554;
assign addr[16209]= -741665807;
assign addr[16210]= -705657826;
assign addr[16211]= -669426032;
assign addr[16212]= -632981917;
assign addr[16213]= -596337040;
assign addr[16214]= -559503022;
assign addr[16215]= -522491548;
assign addr[16216]= -485314355;
assign addr[16217]= -447983235;
assign addr[16218]= -410510029;
assign addr[16219]= -372906622;
assign addr[16220]= -335184940;
assign addr[16221]= -297356948;
assign addr[16222]= -259434643;
assign addr[16223]= -221430054;
assign addr[16224]= -183355234;
assign addr[16225]= -145222259;
assign addr[16226]= -107043224;
assign addr[16227]= -68830239;
assign addr[16228]= -30595422;
assign addr[16229]= 7649098;
assign addr[16230]= 45891193;
assign addr[16231]= 84118732;
assign addr[16232]= 122319591;
assign addr[16233]= 160481654;
assign addr[16234]= 198592817;
assign addr[16235]= 236640993;
assign addr[16236]= 274614114;
assign addr[16237]= 312500135;
assign addr[16238]= 350287041;
assign addr[16239]= 387962847;
assign addr[16240]= 425515602;
assign addr[16241]= 462933398;
assign addr[16242]= 500204365;
assign addr[16243]= 537316682;
assign addr[16244]= 574258580;
assign addr[16245]= 611018340;
assign addr[16246]= 647584304;
assign addr[16247]= 683944874;
assign addr[16248]= 720088517;
assign addr[16249]= 756003771;
assign addr[16250]= 791679244;
assign addr[16251]= 827103620;
assign addr[16252]= 862265664;
assign addr[16253]= 897154224;
assign addr[16254]= 931758235;
assign addr[16255]= 966066720;
assign addr[16256]= 1000068799;
assign addr[16257]= 1033753687;
assign addr[16258]= 1067110699;
assign addr[16259]= 1100129257;
assign addr[16260]= 1132798888;
assign addr[16261]= 1165109230;
assign addr[16262]= 1197050035;
assign addr[16263]= 1228611172;
assign addr[16264]= 1259782632;
assign addr[16265]= 1290554528;
assign addr[16266]= 1320917099;
assign addr[16267]= 1350860716;
assign addr[16268]= 1380375881;
assign addr[16269]= 1409453233;
assign addr[16270]= 1438083551;
assign addr[16271]= 1466257752;
assign addr[16272]= 1493966902;
assign addr[16273]= 1521202211;
assign addr[16274]= 1547955041;
assign addr[16275]= 1574216908;
assign addr[16276]= 1599979481;
assign addr[16277]= 1625234591;
assign addr[16278]= 1649974225;
assign addr[16279]= 1674190539;
assign addr[16280]= 1697875851;
assign addr[16281]= 1721022648;
assign addr[16282]= 1743623590;
assign addr[16283]= 1765671509;
assign addr[16284]= 1787159411;
assign addr[16285]= 1808080480;
assign addr[16286]= 1828428082;
assign addr[16287]= 1848195763;
assign addr[16288]= 1867377253;
assign addr[16289]= 1885966468;
assign addr[16290]= 1903957513;
assign addr[16291]= 1921344681;
assign addr[16292]= 1938122457;
assign addr[16293]= 1954285520;
assign addr[16294]= 1969828744;
assign addr[16295]= 1984747199;
assign addr[16296]= 1999036154;
assign addr[16297]= 2012691075;
assign addr[16298]= 2025707632;
assign addr[16299]= 2038081698;
assign addr[16300]= 2049809346;
assign addr[16301]= 2060886858;
assign addr[16302]= 2071310720;
assign addr[16303]= 2081077626;
assign addr[16304]= 2090184478;
assign addr[16305]= 2098628387;
assign addr[16306]= 2106406677;
assign addr[16307]= 2113516878;
assign addr[16308]= 2119956737;
assign addr[16309]= 2125724211;
assign addr[16310]= 2130817471;
assign addr[16311]= 2135234901;
assign addr[16312]= 2138975100;
assign addr[16313]= 2142036881;
assign addr[16314]= 2144419275;
assign addr[16315]= 2146121524;
assign addr[16316]= 2147143090;
assign addr[16317]= 2147483648;
assign addr[16318]= 2147143090;
assign addr[16319]= 2146121524;
assign addr[16320]= 2144419275;
assign addr[16321]= 2142036881;
assign addr[16322]= 2138975100;
assign addr[16323]= 2135234901;
assign addr[16324]= 2130817471;
assign addr[16325]= 2125724211;
assign addr[16326]= 2119956737;
assign addr[16327]= 2113516878;
assign addr[16328]= 2106406677;
assign addr[16329]= 2098628387;
assign addr[16330]= 2090184478;
assign addr[16331]= 2081077626;
assign addr[16332]= 2071310720;
assign addr[16333]= 2060886858;
assign addr[16334]= 2049809346;
assign addr[16335]= 2038081698;
assign addr[16336]= 2025707632;
assign addr[16337]= 2012691075;
assign addr[16338]= 1999036154;
assign addr[16339]= 1984747199;
assign addr[16340]= 1969828744;
assign addr[16341]= 1954285520;
assign addr[16342]= 1938122457;
assign addr[16343]= 1921344681;
assign addr[16344]= 1903957513;
assign addr[16345]= 1885966468;
assign addr[16346]= 1867377253;
assign addr[16347]= 1848195763;
assign addr[16348]= 1828428082;
assign addr[16349]= 1808080480;
assign addr[16350]= 1787159411;
assign addr[16351]= 1765671509;
assign addr[16352]= 1743623590;
assign addr[16353]= 1721022648;
assign addr[16354]= 1697875851;
assign addr[16355]= 1674190539;
assign addr[16356]= 1649974225;
assign addr[16357]= 1625234591;
assign addr[16358]= 1599979481;
assign addr[16359]= 1574216908;
assign addr[16360]= 1547955041;
assign addr[16361]= 1521202211;
assign addr[16362]= 1493966902;
assign addr[16363]= 1466257752;
assign addr[16364]= 1438083551;
assign addr[16365]= 1409453233;
assign addr[16366]= 1380375881;
assign addr[16367]= 1350860716;
assign addr[16368]= 1320917099;
assign addr[16369]= 1290554528;
assign addr[16370]= 1259782632;
assign addr[16371]= 1228611172;
assign addr[16372]= 1197050035;
assign addr[16373]= 1165109230;
assign addr[16374]= 1132798888;
assign addr[16375]= 1100129257;
assign addr[16376]= 1067110699;
assign addr[16377]= 1033753687;
assign addr[16378]= 1000068799;
assign addr[16379]= 966066720;
assign addr[16380]= 931758235;
assign addr[16381]= 897154224;
assign addr[16382]= 862265664;
assign addr[16383]= 827103620;
assign addr[16384]= 791679244;
assign addr[16385]= 756003771;
assign addr[16386]= 720088517;
assign addr[16387]= 683944874;
assign addr[16388]= 647584304;
assign addr[16389]= 611018340;
assign addr[16390]= 574258580;
assign addr[16391]= 537316682;
assign addr[16392]= 500204365;
assign addr[16393]= 462933398;
assign addr[16394]= 425515602;
assign addr[16395]= 387962847;
assign addr[16396]= 350287041;
assign addr[16397]= 312500135;
assign addr[16398]= 274614114;
assign addr[16399]= 236640993;
assign addr[16400]= 198592817;
assign addr[16401]= 160481654;
assign addr[16402]= 122319591;
assign addr[16403]= 84118732;
assign addr[16404]= 45891193;
assign addr[16405]= 7649098;
assign addr[16406]= -30595422;
assign addr[16407]= -68830239;
assign addr[16408]= -107043224;
assign addr[16409]= -145222259;
assign addr[16410]= -183355234;
assign addr[16411]= -221430054;
assign addr[16412]= -259434643;
assign addr[16413]= -297356948;
assign addr[16414]= -335184940;
assign addr[16415]= -372906622;
assign addr[16416]= -410510029;
assign addr[16417]= -447983235;
assign addr[16418]= -485314355;
assign addr[16419]= -522491548;
assign addr[16420]= -559503022;
assign addr[16421]= -596337040;
assign addr[16422]= -632981917;
assign addr[16423]= -669426032;
assign addr[16424]= -705657826;
assign addr[16425]= -741665807;
assign addr[16426]= -777438554;
assign addr[16427]= -812964722;
assign addr[16428]= -848233042;
assign addr[16429]= -883232329;
assign addr[16430]= -917951481;
assign addr[16431]= -952379488;
assign addr[16432]= -986505429;
assign addr[16433]= -1020318481;
assign addr[16434]= -1053807919;
assign addr[16435]= -1086963121;
assign addr[16436]= -1119773573;
assign addr[16437]= -1152228866;
assign addr[16438]= -1184318708;
assign addr[16439]= -1216032921;
assign addr[16440]= -1247361445;
assign addr[16441]= -1278294345;
assign addr[16442]= -1308821808;
assign addr[16443]= -1338934154;
assign addr[16444]= -1368621831;
assign addr[16445]= -1397875423;
assign addr[16446]= -1426685652;
assign addr[16447]= -1455043381;
assign addr[16448]= -1482939614;
assign addr[16449]= -1510365504;
assign addr[16450]= -1537312353;
assign addr[16451]= -1563771613;
assign addr[16452]= -1589734894;
assign addr[16453]= -1615193959;
assign addr[16454]= -1640140734;
assign addr[16455]= -1664567307;
assign addr[16456]= -1688465931;
assign addr[16457]= -1711829025;
assign addr[16458]= -1734649179;
assign addr[16459]= -1756919156;
assign addr[16460]= -1778631892;
assign addr[16461]= -1799780501;
assign addr[16462]= -1820358275;
assign addr[16463]= -1840358687;
assign addr[16464]= -1859775393;
assign addr[16465]= -1878602237;
assign addr[16466]= -1896833245;
assign addr[16467]= -1914462636;
assign addr[16468]= -1931484818;
assign addr[16469]= -1947894393;
assign addr[16470]= -1963686155;
assign addr[16471]= -1978855097;
assign addr[16472]= -1993396407;
assign addr[16473]= -2007305472;
assign addr[16474]= -2020577882;
assign addr[16475]= -2033209426;
assign addr[16476]= -2045196100;
assign addr[16477]= -2056534099;
assign addr[16478]= -2067219829;
assign addr[16479]= -2077249901;
assign addr[16480]= -2086621133;
assign addr[16481]= -2095330553;
assign addr[16482]= -2103375398;
assign addr[16483]= -2110753117;
assign addr[16484]= -2117461370;
assign addr[16485]= -2123498030;
assign addr[16486]= -2128861181;
assign addr[16487]= -2133549123;
assign addr[16488]= -2137560369;
assign addr[16489]= -2140893646;
assign addr[16490]= -2143547897;
assign addr[16491]= -2145522281;
assign addr[16492]= -2146816171;
assign addr[16493]= -2147429158;
assign addr[16494]= -2147361045;
assign addr[16495]= -2146611856;
assign addr[16496]= -2145181827;
assign addr[16497]= -2143071413;
assign addr[16498]= -2140281282;
assign addr[16499]= -2136812319;
assign addr[16500]= -2132665626;
assign addr[16501]= -2127842516;
assign addr[16502]= -2122344521;
assign addr[16503]= -2116173382;
assign addr[16504]= -2109331059;
assign addr[16505]= -2101819720;
assign addr[16506]= -2093641749;
assign addr[16507]= -2084799740;
assign addr[16508]= -2075296495;
assign addr[16509]= -2065135031;
assign addr[16510]= -2054318569;
assign addr[16511]= -2042850540;
assign addr[16512]= -2030734582;
assign addr[16513]= -2017974537;
assign addr[16514]= -2004574453;
assign addr[16515]= -1990538579;
assign addr[16516]= -1975871368;
assign addr[16517]= -1960577471;
assign addr[16518]= -1944661739;
assign addr[16519]= -1928129220;
assign addr[16520]= -1910985158;
assign addr[16521]= -1893234990;
assign addr[16522]= -1874884346;
assign addr[16523]= -1855939047;
assign addr[16524]= -1836405100;
assign addr[16525]= -1816288703;
assign addr[16526]= -1795596234;
assign addr[16527]= -1774334257;
assign addr[16528]= -1752509516;
assign addr[16529]= -1730128933;
assign addr[16530]= -1707199606;
assign addr[16531]= -1683728808;
assign addr[16532]= -1659723983;
assign addr[16533]= -1635192744;
assign addr[16534]= -1610142873;
assign addr[16535]= -1584582314;
assign addr[16536]= -1558519173;
assign addr[16537]= -1531961719;
assign addr[16538]= -1504918373;
assign addr[16539]= -1477397714;
assign addr[16540]= -1449408469;
assign addr[16541]= -1420959516;
assign addr[16542]= -1392059879;
assign addr[16543]= -1362718723;
assign addr[16544]= -1332945355;
assign addr[16545]= -1302749217;
assign addr[16546]= -1272139887;
assign addr[16547]= -1241127074;
assign addr[16548]= -1209720613;
assign addr[16549]= -1177930466;
assign addr[16550]= -1145766716;
assign addr[16551]= -1113239564;
assign addr[16552]= -1080359326;
assign addr[16553]= -1047136432;
assign addr[16554]= -1013581418;
assign addr[16555]= -979704927;
assign addr[16556]= -945517704;
assign addr[16557]= -911030591;
assign addr[16558]= -876254528;
assign addr[16559]= -841200544;
assign addr[16560]= -805879757;
assign addr[16561]= -770303369;
assign addr[16562]= -734482665;
assign addr[16563]= -698429006;
assign addr[16564]= -662153826;
assign addr[16565]= -625668632;
assign addr[16566]= -588984994;
assign addr[16567]= -552114549;
assign addr[16568]= -515068990;
assign addr[16569]= -477860067;
assign addr[16570]= -440499581;
assign addr[16571]= -402999383;
assign addr[16572]= -365371365;
assign addr[16573]= -327627463;
assign addr[16574]= -289779648;
assign addr[16575]= -251839923;
assign addr[16576]= -213820322;
assign addr[16577]= -175732905;
assign addr[16578]= -137589750;
assign addr[16579]= -99402956;
assign addr[16580]= -61184634;
assign addr[16581]= -22946906;
assign addr[16582]= 15298099;
assign addr[16583]= 53538253;
assign addr[16584]= 91761426;
assign addr[16585]= 129955495;
assign addr[16586]= 168108346;
assign addr[16587]= 206207878;
assign addr[16588]= 244242007;
assign addr[16589]= 282198671;
assign addr[16590]= 320065829;
assign addr[16591]= 357831473;
assign addr[16592]= 395483624;
assign addr[16593]= 433010339;
assign addr[16594]= 470399716;
assign addr[16595]= 507639898;
assign addr[16596]= 544719071;
assign addr[16597]= 581625477;
assign addr[16598]= 618347408;
assign addr[16599]= 654873219;
assign addr[16600]= 691191324;
assign addr[16601]= 727290205;
assign addr[16602]= 763158411;
assign addr[16603]= 798784567;
assign addr[16604]= 834157373;
assign addr[16605]= 869265610;
assign addr[16606]= 904098143;
assign addr[16607]= 938643924;
assign addr[16608]= 972891995;
assign addr[16609]= 1006831495;
assign addr[16610]= 1040451659;
assign addr[16611]= 1073741824;
assign addr[16612]= 1106691431;
assign addr[16613]= 1139290029;
assign addr[16614]= 1171527280;
assign addr[16615]= 1203392958;
assign addr[16616]= 1234876957;
assign addr[16617]= 1265969291;
assign addr[16618]= 1296660098;
assign addr[16619]= 1326939644;
assign addr[16620]= 1356798326;
assign addr[16621]= 1386226674;
assign addr[16622]= 1415215352;
assign addr[16623]= 1443755168;
assign addr[16624]= 1471837070;
assign addr[16625]= 1499452149;
assign addr[16626]= 1526591649;
assign addr[16627]= 1553246960;
assign addr[16628]= 1579409630;
assign addr[16629]= 1605071359;
assign addr[16630]= 1630224009;
assign addr[16631]= 1654859602;
assign addr[16632]= 1678970324;
assign addr[16633]= 1702548529;
assign addr[16634]= 1725586737;
assign addr[16635]= 1748077642;
assign addr[16636]= 1770014111;
assign addr[16637]= 1791389186;
assign addr[16638]= 1812196087;
assign addr[16639]= 1832428215;
assign addr[16640]= 1852079154;
assign addr[16641]= 1871142669;
assign addr[16642]= 1889612716;
assign addr[16643]= 1907483436;
assign addr[16644]= 1924749160;
assign addr[16645]= 1941404413;
assign addr[16646]= 1957443913;
assign addr[16647]= 1972862571;
assign addr[16648]= 1987655498;
assign addr[16649]= 2001818002;
assign addr[16650]= 2015345591;
assign addr[16651]= 2028233973;
assign addr[16652]= 2040479063;
assign addr[16653]= 2052076975;
assign addr[16654]= 2063024031;
assign addr[16655]= 2073316760;
assign addr[16656]= 2082951896;
assign addr[16657]= 2091926384;
assign addr[16658]= 2100237377;
assign addr[16659]= 2107882239;
assign addr[16660]= 2114858546;
assign addr[16661]= 2121164085;
assign addr[16662]= 2126796855;
assign addr[16663]= 2131755071;
assign addr[16664]= 2136037160;
assign addr[16665]= 2139641764;
assign addr[16666]= 2142567738;
assign addr[16667]= 2144814157;
assign addr[16668]= 2146380306;
assign addr[16669]= 2147265689;
assign addr[16670]= 2147470025;
assign addr[16671]= 2146993250;
assign addr[16672]= 2145835515;
assign addr[16673]= 2143997187;
assign addr[16674]= 2141478848;
assign addr[16675]= 2138281298;
assign addr[16676]= 2134405552;
assign addr[16677]= 2129852837;
assign addr[16678]= 2124624598;
assign addr[16679]= 2118722494;
assign addr[16680]= 2112148396;
assign addr[16681]= 2104904390;
assign addr[16682]= 2096992772;
assign addr[16683]= 2088416053;
assign addr[16684]= 2079176953;
assign addr[16685]= 2069278401;
assign addr[16686]= 2058723538;
assign addr[16687]= 2047515711;
assign addr[16688]= 2035658475;
assign addr[16689]= 2023155591;
assign addr[16690]= 2010011024;
assign addr[16691]= 1996228943;
assign addr[16692]= 1981813720;
assign addr[16693]= 1966769926;
assign addr[16694]= 1951102334;
assign addr[16695]= 1934815911;
assign addr[16696]= 1917915825;
assign addr[16697]= 1900407434;
assign addr[16698]= 1882296293;
assign addr[16699]= 1863588145;
assign addr[16700]= 1844288924;
assign addr[16701]= 1824404752;
assign addr[16702]= 1803941934;
assign addr[16703]= 1782906961;
assign addr[16704]= 1761306505;
assign addr[16705]= 1739147417;
assign addr[16706]= 1716436725;
assign addr[16707]= 1693181631;
assign addr[16708]= 1669389513;
assign addr[16709]= 1645067915;
assign addr[16710]= 1620224553;
assign addr[16711]= 1594867305;
assign addr[16712]= 1569004214;
assign addr[16713]= 1542643483;
assign addr[16714]= 1515793473;
assign addr[16715]= 1488462700;
assign addr[16716]= 1460659832;
assign addr[16717]= 1432393688;
assign addr[16718]= 1403673233;
assign addr[16719]= 1374507575;
assign addr[16720]= 1344905966;
assign addr[16721]= 1314877795;
assign addr[16722]= 1284432584;
assign addr[16723]= 1253579991;
assign addr[16724]= 1222329801;
assign addr[16725]= 1190691925;
assign addr[16726]= 1158676398;
assign addr[16727]= 1126293375;
assign addr[16728]= 1093553126;
assign addr[16729]= 1060466036;
assign addr[16730]= 1027042599;
assign addr[16731]= 993293415;
assign addr[16732]= 959229189;
assign addr[16733]= 924860725;
assign addr[16734]= 890198924;
assign addr[16735]= 855254778;
assign addr[16736]= 820039373;
assign addr[16737]= 784563876;
assign addr[16738]= 748839539;
assign addr[16739]= 712877694;
assign addr[16740]= 676689746;
assign addr[16741]= 640287172;
assign addr[16742]= 603681519;
assign addr[16743]= 566884397;
assign addr[16744]= 529907477;
assign addr[16745]= 492762486;
assign addr[16746]= 455461206;
assign addr[16747]= 418015468;
assign addr[16748]= 380437148;
assign addr[16749]= 342738165;
assign addr[16750]= 304930476;
assign addr[16751]= 267026072;
assign addr[16752]= 229036977;
assign addr[16753]= 190975237;
assign addr[16754]= 152852926;
assign addr[16755]= 114682135;
assign addr[16756]= 76474970;
assign addr[16757]= 38243550;
assign addr[16758]= 0;
assign addr[16759]= -38243550;
assign addr[16760]= -76474970;
assign addr[16761]= -114682135;
assign addr[16762]= -152852926;
assign addr[16763]= -190975237;
assign addr[16764]= -229036977;
assign addr[16765]= -267026072;
assign addr[16766]= -304930476;
assign addr[16767]= -342738165;
assign addr[16768]= -380437148;
assign addr[16769]= -418015468;
assign addr[16770]= -455461206;
assign addr[16771]= -492762486;
assign addr[16772]= -529907477;
assign addr[16773]= -566884397;
assign addr[16774]= -603681519;
assign addr[16775]= -640287172;
assign addr[16776]= -676689746;
assign addr[16777]= -712877694;
assign addr[16778]= -748839539;
assign addr[16779]= -784563876;
assign addr[16780]= -820039373;
assign addr[16781]= -855254778;
assign addr[16782]= -890198924;
assign addr[16783]= -924860725;
assign addr[16784]= -959229189;
assign addr[16785]= -993293415;
assign addr[16786]= -1027042599;
assign addr[16787]= -1060466036;
assign addr[16788]= -1093553126;
assign addr[16789]= -1126293375;
assign addr[16790]= -1158676398;
assign addr[16791]= -1190691925;
assign addr[16792]= -1222329801;
assign addr[16793]= -1253579991;
assign addr[16794]= -1284432584;
assign addr[16795]= -1314877795;
assign addr[16796]= -1344905966;
assign addr[16797]= -1374507575;
assign addr[16798]= -1403673233;
assign addr[16799]= -1432393688;
assign addr[16800]= -1460659832;
assign addr[16801]= -1488462700;
assign addr[16802]= -1515793473;
assign addr[16803]= -1542643483;
assign addr[16804]= -1569004214;
assign addr[16805]= -1594867305;
assign addr[16806]= -1620224553;
assign addr[16807]= -1645067915;
assign addr[16808]= -1669389513;
assign addr[16809]= -1693181631;
assign addr[16810]= -1716436725;
assign addr[16811]= -1739147417;
assign addr[16812]= -1761306505;
assign addr[16813]= -1782906961;
assign addr[16814]= -1803941934;
assign addr[16815]= -1824404752;
assign addr[16816]= -1844288924;
assign addr[16817]= -1863588145;
assign addr[16818]= -1882296293;
assign addr[16819]= -1900407434;
assign addr[16820]= -1917915825;
assign addr[16821]= -1934815911;
assign addr[16822]= -1951102334;
assign addr[16823]= -1966769926;
assign addr[16824]= -1981813720;
assign addr[16825]= -1996228943;
assign addr[16826]= -2010011024;
assign addr[16827]= -2023155591;
assign addr[16828]= -2035658475;
assign addr[16829]= -2047515711;
assign addr[16830]= -2058723538;
assign addr[16831]= -2069278401;
assign addr[16832]= -2079176953;
assign addr[16833]= -2088416053;
assign addr[16834]= -2096992772;
assign addr[16835]= -2104904390;
assign addr[16836]= -2112148396;
assign addr[16837]= -2118722494;
assign addr[16838]= -2124624598;
assign addr[16839]= -2129852837;
assign addr[16840]= -2134405552;
assign addr[16841]= -2138281298;
assign addr[16842]= -2141478848;
assign addr[16843]= -2143997187;
assign addr[16844]= -2145835515;
assign addr[16845]= -2146993250;
assign addr[16846]= -2147470025;
assign addr[16847]= -2147265689;
assign addr[16848]= -2146380306;
assign addr[16849]= -2144814157;
assign addr[16850]= -2142567738;
assign addr[16851]= -2139641764;
assign addr[16852]= -2136037160;
assign addr[16853]= -2131755071;
assign addr[16854]= -2126796855;
assign addr[16855]= -2121164085;
assign addr[16856]= -2114858546;
assign addr[16857]= -2107882239;
assign addr[16858]= -2100237377;
assign addr[16859]= -2091926384;
assign addr[16860]= -2082951896;
assign addr[16861]= -2073316760;
assign addr[16862]= -2063024031;
assign addr[16863]= -2052076975;
assign addr[16864]= -2040479063;
assign addr[16865]= -2028233973;
assign addr[16866]= -2015345591;
assign addr[16867]= -2001818002;
assign addr[16868]= -1987655498;
assign addr[16869]= -1972862571;
assign addr[16870]= -1957443913;
assign addr[16871]= -1941404413;
assign addr[16872]= -1924749160;
assign addr[16873]= -1907483436;
assign addr[16874]= -1889612716;
assign addr[16875]= -1871142669;
assign addr[16876]= -1852079154;
assign addr[16877]= -1832428215;
assign addr[16878]= -1812196087;
assign addr[16879]= -1791389186;
assign addr[16880]= -1770014111;
assign addr[16881]= -1748077642;
assign addr[16882]= -1725586737;
assign addr[16883]= -1702548529;
assign addr[16884]= -1678970324;
assign addr[16885]= -1654859602;
assign addr[16886]= -1630224009;
assign addr[16887]= -1605071359;
assign addr[16888]= -1579409630;
assign addr[16889]= -1553246960;
assign addr[16890]= -1526591649;
assign addr[16891]= -1499452149;
assign addr[16892]= -1471837070;
assign addr[16893]= -1443755168;
assign addr[16894]= -1415215352;
assign addr[16895]= -1386226674;
assign addr[16896]= -1356798326;
assign addr[16897]= -1326939644;
assign addr[16898]= -1296660098;
assign addr[16899]= -1265969291;
assign addr[16900]= -1234876957;
assign addr[16901]= -1203392958;
assign addr[16902]= -1171527280;
assign addr[16903]= -1139290029;
assign addr[16904]= -1106691431;
assign addr[16905]= -1073741824;
assign addr[16906]= -1040451659;
assign addr[16907]= -1006831495;
assign addr[16908]= -972891995;
assign addr[16909]= -938643924;
assign addr[16910]= -904098143;
assign addr[16911]= -869265610;
assign addr[16912]= -834157373;
assign addr[16913]= -798784567;
assign addr[16914]= -763158411;
assign addr[16915]= -727290205;
assign addr[16916]= -691191324;
assign addr[16917]= -654873219;
assign addr[16918]= -618347408;
assign addr[16919]= -581625477;
assign addr[16920]= -544719071;
assign addr[16921]= -507639898;
assign addr[16922]= -470399716;
assign addr[16923]= -433010339;
assign addr[16924]= -395483624;
assign addr[16925]= -357831473;
assign addr[16926]= -320065829;
assign addr[16927]= -282198671;
assign addr[16928]= -244242007;
assign addr[16929]= -206207878;
assign addr[16930]= -168108346;
assign addr[16931]= -129955495;
assign addr[16932]= -91761426;
assign addr[16933]= -53538253;
assign addr[16934]= -15298099;
assign addr[16935]= 22946906;
assign addr[16936]= 61184634;
assign addr[16937]= 99402956;
assign addr[16938]= 137589750;
assign addr[16939]= 175732905;
assign addr[16940]= 213820322;
assign addr[16941]= 251839923;
assign addr[16942]= 289779648;
assign addr[16943]= 327627463;
assign addr[16944]= 365371365;
assign addr[16945]= 402999383;
assign addr[16946]= 440499581;
assign addr[16947]= 477860067;
assign addr[16948]= 515068990;
assign addr[16949]= 552114549;
assign addr[16950]= 588984994;
assign addr[16951]= 625668632;
assign addr[16952]= 662153826;
assign addr[16953]= 698429006;
assign addr[16954]= 734482665;
assign addr[16955]= 770303369;
assign addr[16956]= 805879757;
assign addr[16957]= 841200544;
assign addr[16958]= 876254528;
assign addr[16959]= 911030591;
assign addr[16960]= 945517704;
assign addr[16961]= 979704927;
assign addr[16962]= 1013581418;
assign addr[16963]= 1047136432;
assign addr[16964]= 1080359326;
assign addr[16965]= 1113239564;
assign addr[16966]= 1145766716;
assign addr[16967]= 1177930466;
assign addr[16968]= 1209720613;
assign addr[16969]= 1241127074;
assign addr[16970]= 1272139887;
assign addr[16971]= 1302749217;
assign addr[16972]= 1332945355;
assign addr[16973]= 1362718723;
assign addr[16974]= 1392059879;
assign addr[16975]= 1420959516;
assign addr[16976]= 1449408469;
assign addr[16977]= 1477397714;
assign addr[16978]= 1504918373;
assign addr[16979]= 1531961719;
assign addr[16980]= 1558519173;
assign addr[16981]= 1584582314;
assign addr[16982]= 1610142873;
assign addr[16983]= 1635192744;
assign addr[16984]= 1659723983;
assign addr[16985]= 1683728808;
assign addr[16986]= 1707199606;
assign addr[16987]= 1730128933;
assign addr[16988]= 1752509516;
assign addr[16989]= 1774334257;
assign addr[16990]= 1795596234;
assign addr[16991]= 1816288703;
assign addr[16992]= 1836405100;
assign addr[16993]= 1855939047;
assign addr[16994]= 1874884346;
assign addr[16995]= 1893234990;
assign addr[16996]= 1910985158;
assign addr[16997]= 1928129220;
assign addr[16998]= 1944661739;
assign addr[16999]= 1960577471;
assign addr[17000]= 1975871368;
assign addr[17001]= 1990538579;
assign addr[17002]= 2004574453;
assign addr[17003]= 2017974537;
assign addr[17004]= 2030734582;
assign addr[17005]= 2042850540;
assign addr[17006]= 2054318569;
assign addr[17007]= 2065135031;
assign addr[17008]= 2075296495;
assign addr[17009]= 2084799740;
assign addr[17010]= 2093641749;
assign addr[17011]= 2101819720;
assign addr[17012]= 2109331059;
assign addr[17013]= 2116173382;
assign addr[17014]= 2122344521;
assign addr[17015]= 2127842516;
assign addr[17016]= 2132665626;
assign addr[17017]= 2136812319;
assign addr[17018]= 2140281282;
assign addr[17019]= 2143071413;
assign addr[17020]= 2145181827;
assign addr[17021]= 2146611856;
assign addr[17022]= 2147361045;
assign addr[17023]= 2147429158;
assign addr[17024]= 2146816171;
assign addr[17025]= 2145522281;
assign addr[17026]= 2143547897;
assign addr[17027]= 2140893646;
assign addr[17028]= 2137560369;
assign addr[17029]= 2133549123;
assign addr[17030]= 2128861181;
assign addr[17031]= 2123498030;
assign addr[17032]= 2117461370;
assign addr[17033]= 2110753117;
assign addr[17034]= 2103375398;
assign addr[17035]= 2095330553;
assign addr[17036]= 2086621133;
assign addr[17037]= 2077249901;
assign addr[17038]= 2067219829;
assign addr[17039]= 2056534099;
assign addr[17040]= 2045196100;
assign addr[17041]= 2033209426;
assign addr[17042]= 2020577882;
assign addr[17043]= 2007305472;
assign addr[17044]= 1993396407;
assign addr[17045]= 1978855097;
assign addr[17046]= 1963686155;
assign addr[17047]= 1947894393;
assign addr[17048]= 1931484818;
assign addr[17049]= 1914462636;
assign addr[17050]= 1896833245;
assign addr[17051]= 1878602237;
assign addr[17052]= 1859775393;
assign addr[17053]= 1840358687;
assign addr[17054]= 1820358275;
assign addr[17055]= 1799780501;
assign addr[17056]= 1778631892;
assign addr[17057]= 1756919156;
assign addr[17058]= 1734649179;
assign addr[17059]= 1711829025;
assign addr[17060]= 1688465931;
assign addr[17061]= 1664567307;
assign addr[17062]= 1640140734;
assign addr[17063]= 1615193959;
assign addr[17064]= 1589734894;
assign addr[17065]= 1563771613;
assign addr[17066]= 1537312353;
assign addr[17067]= 1510365504;
assign addr[17068]= 1482939614;
assign addr[17069]= 1455043381;
assign addr[17070]= 1426685652;
assign addr[17071]= 1397875423;
assign addr[17072]= 1368621831;
assign addr[17073]= 1338934154;
assign addr[17074]= 1308821808;
assign addr[17075]= 1278294345;
assign addr[17076]= 1247361445;
assign addr[17077]= 1216032921;
assign addr[17078]= 1184318708;
assign addr[17079]= 1152228866;
assign addr[17080]= 1119773573;
assign addr[17081]= 1086963121;
assign addr[17082]= 1053807919;
assign addr[17083]= 1020318481;
assign addr[17084]= 986505429;
assign addr[17085]= 952379488;
assign addr[17086]= 917951481;
assign addr[17087]= 883232329;
assign addr[17088]= 848233042;
assign addr[17089]= 812964722;
assign addr[17090]= 777438554;
assign addr[17091]= 741665807;
assign addr[17092]= 705657826;
assign addr[17093]= 669426032;
assign addr[17094]= 632981917;
assign addr[17095]= 596337040;
assign addr[17096]= 559503022;
assign addr[17097]= 522491548;
assign addr[17098]= 485314355;
assign addr[17099]= 447983235;
assign addr[17100]= 410510029;
assign addr[17101]= 372906622;
assign addr[17102]= 335184940;
assign addr[17103]= 297356948;
assign addr[17104]= 259434643;
assign addr[17105]= 221430054;
assign addr[17106]= 183355234;
assign addr[17107]= 145222259;
assign addr[17108]= 107043224;
assign addr[17109]= 68830239;
assign addr[17110]= 30595422;
assign addr[17111]= -7649098;
assign addr[17112]= -45891193;
assign addr[17113]= -84118732;
assign addr[17114]= -122319591;
assign addr[17115]= -160481654;
assign addr[17116]= -198592817;
assign addr[17117]= -236640993;
assign addr[17118]= -274614114;
assign addr[17119]= -312500135;
assign addr[17120]= -350287041;
assign addr[17121]= -387962847;
assign addr[17122]= -425515602;
assign addr[17123]= -462933398;
assign addr[17124]= -500204365;
assign addr[17125]= -537316682;
assign addr[17126]= -574258580;
assign addr[17127]= -611018340;
assign addr[17128]= -647584304;
assign addr[17129]= -683944874;
assign addr[17130]= -720088517;
assign addr[17131]= -756003771;
assign addr[17132]= -791679244;
assign addr[17133]= -827103620;
assign addr[17134]= -862265664;
assign addr[17135]= -897154224;
assign addr[17136]= -931758235;
assign addr[17137]= -966066720;
assign addr[17138]= -1000068799;
assign addr[17139]= -1033753687;
assign addr[17140]= -1067110699;
assign addr[17141]= -1100129257;
assign addr[17142]= -1132798888;
assign addr[17143]= -1165109230;
assign addr[17144]= -1197050035;
assign addr[17145]= -1228611172;
assign addr[17146]= -1259782632;
assign addr[17147]= -1290554528;
assign addr[17148]= -1320917099;
assign addr[17149]= -1350860716;
assign addr[17150]= -1380375881;
assign addr[17151]= -1409453233;
assign addr[17152]= -1438083551;
assign addr[17153]= -1466257752;
assign addr[17154]= -1493966902;
assign addr[17155]= -1521202211;
assign addr[17156]= -1547955041;
assign addr[17157]= -1574216908;
assign addr[17158]= -1599979481;
assign addr[17159]= -1625234591;
assign addr[17160]= -1649974225;
assign addr[17161]= -1674190539;
assign addr[17162]= -1697875851;
assign addr[17163]= -1721022648;
assign addr[17164]= -1743623590;
assign addr[17165]= -1765671509;
assign addr[17166]= -1787159411;
assign addr[17167]= -1808080480;
assign addr[17168]= -1828428082;
assign addr[17169]= -1848195763;
assign addr[17170]= -1867377253;
assign addr[17171]= -1885966468;
assign addr[17172]= -1903957513;
assign addr[17173]= -1921344681;
assign addr[17174]= -1938122457;
assign addr[17175]= -1954285520;
assign addr[17176]= -1969828744;
assign addr[17177]= -1984747199;
assign addr[17178]= -1999036154;
assign addr[17179]= -2012691075;
assign addr[17180]= -2025707632;
assign addr[17181]= -2038081698;
assign addr[17182]= -2049809346;
assign addr[17183]= -2060886858;
assign addr[17184]= -2071310720;
assign addr[17185]= -2081077626;
assign addr[17186]= -2090184478;
assign addr[17187]= -2098628387;
assign addr[17188]= -2106406677;
assign addr[17189]= -2113516878;
assign addr[17190]= -2119956737;
assign addr[17191]= -2125724211;
assign addr[17192]= -2130817471;
assign addr[17193]= -2135234901;
assign addr[17194]= -2138975100;
assign addr[17195]= -2142036881;
assign addr[17196]= -2144419275;
assign addr[17197]= -2146121524;
assign addr[17198]= -2147143090;
assign addr[17199]= -2147483648;
assign addr[17200]= -2147143090;
assign addr[17201]= -2146121524;
assign addr[17202]= -2144419275;
assign addr[17203]= -2142036881;
assign addr[17204]= -2138975100;
assign addr[17205]= -2135234901;
assign addr[17206]= -2130817471;
assign addr[17207]= -2125724211;
assign addr[17208]= -2119956737;
assign addr[17209]= -2113516878;
assign addr[17210]= -2106406677;
assign addr[17211]= -2098628387;
assign addr[17212]= -2090184478;
assign addr[17213]= -2081077626;
assign addr[17214]= -2071310720;
assign addr[17215]= -2060886858;
assign addr[17216]= -2049809346;
assign addr[17217]= -2038081698;
assign addr[17218]= -2025707632;
assign addr[17219]= -2012691075;
assign addr[17220]= -1999036154;
assign addr[17221]= -1984747199;
assign addr[17222]= -1969828744;
assign addr[17223]= -1954285520;
assign addr[17224]= -1938122457;
assign addr[17225]= -1921344681;
assign addr[17226]= -1903957513;
assign addr[17227]= -1885966468;
assign addr[17228]= -1867377253;
assign addr[17229]= -1848195763;
assign addr[17230]= -1828428082;
assign addr[17231]= -1808080480;
assign addr[17232]= -1787159411;
assign addr[17233]= -1765671509;
assign addr[17234]= -1743623590;
assign addr[17235]= -1721022648;
assign addr[17236]= -1697875851;
assign addr[17237]= -1674190539;
assign addr[17238]= -1649974225;
assign addr[17239]= -1625234591;
assign addr[17240]= -1599979481;
assign addr[17241]= -1574216908;
assign addr[17242]= -1547955041;
assign addr[17243]= -1521202211;
assign addr[17244]= -1493966902;
assign addr[17245]= -1466257752;
assign addr[17246]= -1438083551;
assign addr[17247]= -1409453233;
assign addr[17248]= -1380375881;
assign addr[17249]= -1350860716;
assign addr[17250]= -1320917099;
assign addr[17251]= -1290554528;
assign addr[17252]= -1259782632;
assign addr[17253]= -1228611172;
assign addr[17254]= -1197050035;
assign addr[17255]= -1165109230;
assign addr[17256]= -1132798888;
assign addr[17257]= -1100129257;
assign addr[17258]= -1067110699;
assign addr[17259]= -1033753687;
assign addr[17260]= -1000068799;
assign addr[17261]= -966066720;
assign addr[17262]= -931758235;
assign addr[17263]= -897154224;
assign addr[17264]= -862265664;
assign addr[17265]= -827103620;
assign addr[17266]= -791679244;
assign addr[17267]= -756003771;
assign addr[17268]= -720088517;
assign addr[17269]= -683944874;
assign addr[17270]= -647584304;
assign addr[17271]= -611018340;
assign addr[17272]= -574258580;
assign addr[17273]= -537316682;
assign addr[17274]= -500204365;
assign addr[17275]= -462933398;
assign addr[17276]= -425515602;
assign addr[17277]= -387962847;
assign addr[17278]= -350287041;
assign addr[17279]= -312500135;
assign addr[17280]= -274614114;
assign addr[17281]= -236640993;
assign addr[17282]= -198592817;
assign addr[17283]= -160481654;
assign addr[17284]= -122319591;
assign addr[17285]= -84118732;
assign addr[17286]= -45891193;
assign addr[17287]= -7649098;
assign addr[17288]= 30595422;
assign addr[17289]= 68830239;
assign addr[17290]= 107043224;
assign addr[17291]= 145222259;
assign addr[17292]= 183355234;
assign addr[17293]= 221430054;
assign addr[17294]= 259434643;
assign addr[17295]= 297356948;
assign addr[17296]= 335184940;
assign addr[17297]= 372906622;
assign addr[17298]= 410510029;
assign addr[17299]= 447983235;
assign addr[17300]= 485314355;
assign addr[17301]= 522491548;
assign addr[17302]= 559503022;
assign addr[17303]= 596337040;
assign addr[17304]= 632981917;
assign addr[17305]= 669426032;
assign addr[17306]= 705657826;
assign addr[17307]= 741665807;
assign addr[17308]= 777438554;
assign addr[17309]= 812964722;
assign addr[17310]= 848233042;
assign addr[17311]= 883232329;
assign addr[17312]= 917951481;
assign addr[17313]= 952379488;
assign addr[17314]= 986505429;
assign addr[17315]= 1020318481;
assign addr[17316]= 1053807919;
assign addr[17317]= 1086963121;
assign addr[17318]= 1119773573;
assign addr[17319]= 1152228866;
assign addr[17320]= 1184318708;
assign addr[17321]= 1216032921;
assign addr[17322]= 1247361445;
assign addr[17323]= 1278294345;
assign addr[17324]= 1308821808;
assign addr[17325]= 1338934154;
assign addr[17326]= 1368621831;
assign addr[17327]= 1397875423;
assign addr[17328]= 1426685652;
assign addr[17329]= 1455043381;
assign addr[17330]= 1482939614;
assign addr[17331]= 1510365504;
assign addr[17332]= 1537312353;
assign addr[17333]= 1563771613;
assign addr[17334]= 1589734894;
assign addr[17335]= 1615193959;
assign addr[17336]= 1640140734;
assign addr[17337]= 1664567307;
assign addr[17338]= 1688465931;
assign addr[17339]= 1711829025;
assign addr[17340]= 1734649179;
assign addr[17341]= 1756919156;
assign addr[17342]= 1778631892;
assign addr[17343]= 1799780501;
assign addr[17344]= 1820358275;
assign addr[17345]= 1840358687;
assign addr[17346]= 1859775393;
assign addr[17347]= 1878602237;
assign addr[17348]= 1896833245;
assign addr[17349]= 1914462636;
assign addr[17350]= 1931484818;
assign addr[17351]= 1947894393;
assign addr[17352]= 1963686155;
assign addr[17353]= 1978855097;
assign addr[17354]= 1993396407;
assign addr[17355]= 2007305472;
assign addr[17356]= 2020577882;
assign addr[17357]= 2033209426;
assign addr[17358]= 2045196100;
assign addr[17359]= 2056534099;
assign addr[17360]= 2067219829;
assign addr[17361]= 2077249901;
assign addr[17362]= 2086621133;
assign addr[17363]= 2095330553;
assign addr[17364]= 2103375398;
assign addr[17365]= 2110753117;
assign addr[17366]= 2117461370;
assign addr[17367]= 2123498030;
assign addr[17368]= 2128861181;
assign addr[17369]= 2133549123;
assign addr[17370]= 2137560369;
assign addr[17371]= 2140893646;
assign addr[17372]= 2143547897;
assign addr[17373]= 2145522281;
assign addr[17374]= 2146816171;
assign addr[17375]= 2147429158;
assign addr[17376]= 2147361045;
assign addr[17377]= 2146611856;
assign addr[17378]= 2145181827;
assign addr[17379]= 2143071413;
assign addr[17380]= 2140281282;
assign addr[17381]= 2136812319;
assign addr[17382]= 2132665626;
assign addr[17383]= 2127842516;
assign addr[17384]= 2122344521;
assign addr[17385]= 2116173382;
assign addr[17386]= 2109331059;
assign addr[17387]= 2101819720;
assign addr[17388]= 2093641749;
assign addr[17389]= 2084799740;
assign addr[17390]= 2075296495;
assign addr[17391]= 2065135031;
assign addr[17392]= 2054318569;
assign addr[17393]= 2042850540;
assign addr[17394]= 2030734582;
assign addr[17395]= 2017974537;
assign addr[17396]= 2004574453;
assign addr[17397]= 1990538579;
assign addr[17398]= 1975871368;
assign addr[17399]= 1960577471;
assign addr[17400]= 1944661739;
assign addr[17401]= 1928129220;
assign addr[17402]= 1910985158;
assign addr[17403]= 1893234990;
assign addr[17404]= 1874884346;
assign addr[17405]= 1855939047;
assign addr[17406]= 1836405100;
assign addr[17407]= 1816288703;
assign addr[17408]= 1795596234;
assign addr[17409]= 1774334257;
assign addr[17410]= 1752509516;
assign addr[17411]= 1730128933;
assign addr[17412]= 1707199606;
assign addr[17413]= 1683728808;
assign addr[17414]= 1659723983;
assign addr[17415]= 1635192744;
assign addr[17416]= 1610142873;
assign addr[17417]= 1584582314;
assign addr[17418]= 1558519173;
assign addr[17419]= 1531961719;
assign addr[17420]= 1504918373;
assign addr[17421]= 1477397714;
assign addr[17422]= 1449408469;
assign addr[17423]= 1420959516;
assign addr[17424]= 1392059879;
assign addr[17425]= 1362718723;
assign addr[17426]= 1332945355;
assign addr[17427]= 1302749217;
assign addr[17428]= 1272139887;
assign addr[17429]= 1241127074;
assign addr[17430]= 1209720613;
assign addr[17431]= 1177930466;
assign addr[17432]= 1145766716;
assign addr[17433]= 1113239564;
assign addr[17434]= 1080359326;
assign addr[17435]= 1047136432;
assign addr[17436]= 1013581418;
assign addr[17437]= 979704927;
assign addr[17438]= 945517704;
assign addr[17439]= 911030591;
assign addr[17440]= 876254528;
assign addr[17441]= 841200544;
assign addr[17442]= 805879757;
assign addr[17443]= 770303369;
assign addr[17444]= 734482665;
assign addr[17445]= 698429006;
assign addr[17446]= 662153826;
assign addr[17447]= 625668632;
assign addr[17448]= 588984994;
assign addr[17449]= 552114549;
assign addr[17450]= 515068990;
assign addr[17451]= 477860067;
assign addr[17452]= 440499581;
assign addr[17453]= 402999383;
assign addr[17454]= 365371365;
assign addr[17455]= 327627463;
assign addr[17456]= 289779648;
assign addr[17457]= 251839923;
assign addr[17458]= 213820322;
assign addr[17459]= 175732905;
assign addr[17460]= 137589750;
assign addr[17461]= 99402956;
assign addr[17462]= 61184634;
assign addr[17463]= 22946906;
assign addr[17464]= -15298099;
assign addr[17465]= -53538253;
assign addr[17466]= -91761426;
assign addr[17467]= -129955495;
assign addr[17468]= -168108346;
assign addr[17469]= -206207878;
assign addr[17470]= -244242007;
assign addr[17471]= -282198671;
assign addr[17472]= -320065829;
assign addr[17473]= -357831473;
assign addr[17474]= -395483624;
assign addr[17475]= -433010339;
assign addr[17476]= -470399716;
assign addr[17477]= -507639898;
assign addr[17478]= -544719071;
assign addr[17479]= -581625477;
assign addr[17480]= -618347408;
assign addr[17481]= -654873219;
assign addr[17482]= -691191324;
assign addr[17483]= -727290205;
assign addr[17484]= -763158411;
assign addr[17485]= -798784567;
assign addr[17486]= -834157373;
assign addr[17487]= -869265610;
assign addr[17488]= -904098143;
assign addr[17489]= -938643924;
assign addr[17490]= -972891995;
assign addr[17491]= -1006831495;
assign addr[17492]= -1040451659;
assign addr[17493]= -1073741824;
assign addr[17494]= -1106691431;
assign addr[17495]= -1139290029;
assign addr[17496]= -1171527280;
assign addr[17497]= -1203392958;
assign addr[17498]= -1234876957;
assign addr[17499]= -1265969291;
assign addr[17500]= -1296660098;
assign addr[17501]= -1326939644;
assign addr[17502]= -1356798326;
assign addr[17503]= -1386226674;
assign addr[17504]= -1415215352;
assign addr[17505]= -1443755168;
assign addr[17506]= -1471837070;
assign addr[17507]= -1499452149;
assign addr[17508]= -1526591649;
assign addr[17509]= -1553246960;
assign addr[17510]= -1579409630;
assign addr[17511]= -1605071359;
assign addr[17512]= -1630224009;
assign addr[17513]= -1654859602;
assign addr[17514]= -1678970324;
assign addr[17515]= -1702548529;
assign addr[17516]= -1725586737;
assign addr[17517]= -1748077642;
assign addr[17518]= -1770014111;
assign addr[17519]= -1791389186;
assign addr[17520]= -1812196087;
assign addr[17521]= -1832428215;
assign addr[17522]= -1852079154;
assign addr[17523]= -1871142669;
assign addr[17524]= -1889612716;
assign addr[17525]= -1907483436;
assign addr[17526]= -1924749160;
assign addr[17527]= -1941404413;
assign addr[17528]= -1957443913;
assign addr[17529]= -1972862571;
assign addr[17530]= -1987655498;
assign addr[17531]= -2001818002;
assign addr[17532]= -2015345591;
assign addr[17533]= -2028233973;
assign addr[17534]= -2040479063;
assign addr[17535]= -2052076975;
assign addr[17536]= -2063024031;
assign addr[17537]= -2073316760;
assign addr[17538]= -2082951896;
assign addr[17539]= -2091926384;
assign addr[17540]= -2100237377;
assign addr[17541]= -2107882239;
assign addr[17542]= -2114858546;
assign addr[17543]= -2121164085;
assign addr[17544]= -2126796855;
assign addr[17545]= -2131755071;
assign addr[17546]= -2136037160;
assign addr[17547]= -2139641764;
assign addr[17548]= -2142567738;
assign addr[17549]= -2144814157;
assign addr[17550]= -2146380306;
assign addr[17551]= -2147265689;
assign addr[17552]= -2147470025;
assign addr[17553]= -2146993250;
assign addr[17554]= -2145835515;
assign addr[17555]= -2143997187;
assign addr[17556]= -2141478848;
assign addr[17557]= -2138281298;
assign addr[17558]= -2134405552;
assign addr[17559]= -2129852837;
assign addr[17560]= -2124624598;
assign addr[17561]= -2118722494;
assign addr[17562]= -2112148396;
assign addr[17563]= -2104904390;
assign addr[17564]= -2096992772;
assign addr[17565]= -2088416053;
assign addr[17566]= -2079176953;
assign addr[17567]= -2069278401;
assign addr[17568]= -2058723538;
assign addr[17569]= -2047515711;
assign addr[17570]= -2035658475;
assign addr[17571]= -2023155591;
assign addr[17572]= -2010011024;
assign addr[17573]= -1996228943;
assign addr[17574]= -1981813720;
assign addr[17575]= -1966769926;
assign addr[17576]= -1951102334;
assign addr[17577]= -1934815911;
assign addr[17578]= -1917915825;
assign addr[17579]= -1900407434;
assign addr[17580]= -1882296293;
assign addr[17581]= -1863588145;
assign addr[17582]= -1844288924;
assign addr[17583]= -1824404752;
assign addr[17584]= -1803941934;
assign addr[17585]= -1782906961;
assign addr[17586]= -1761306505;
assign addr[17587]= -1739147417;
assign addr[17588]= -1716436725;
assign addr[17589]= -1693181631;
assign addr[17590]= -1669389513;
assign addr[17591]= -1645067915;
assign addr[17592]= -1620224553;
assign addr[17593]= -1594867305;
assign addr[17594]= -1569004214;
assign addr[17595]= -1542643483;
assign addr[17596]= -1515793473;
assign addr[17597]= -1488462700;
assign addr[17598]= -1460659832;
assign addr[17599]= -1432393688;
assign addr[17600]= -1403673233;
assign addr[17601]= -1374507575;
assign addr[17602]= -1344905966;
assign addr[17603]= -1314877795;
assign addr[17604]= -1284432584;
assign addr[17605]= -1253579991;
assign addr[17606]= -1222329801;
assign addr[17607]= -1190691925;
assign addr[17608]= -1158676398;
assign addr[17609]= -1126293375;
assign addr[17610]= -1093553126;
assign addr[17611]= -1060466036;
assign addr[17612]= -1027042599;
assign addr[17613]= -993293415;
assign addr[17614]= -959229189;
assign addr[17615]= -924860725;
assign addr[17616]= -890198924;
assign addr[17617]= -855254778;
assign addr[17618]= -820039373;
assign addr[17619]= -784563876;
assign addr[17620]= -748839539;
assign addr[17621]= -712877694;
assign addr[17622]= -676689746;
assign addr[17623]= -640287172;
assign addr[17624]= -603681519;
assign addr[17625]= -566884397;
assign addr[17626]= -529907477;
assign addr[17627]= -492762486;
assign addr[17628]= -455461206;
assign addr[17629]= -418015468;
assign addr[17630]= -380437148;
assign addr[17631]= -342738165;
assign addr[17632]= -304930476;
assign addr[17633]= -267026072;
assign addr[17634]= -229036977;
assign addr[17635]= -190975237;
assign addr[17636]= -152852926;
assign addr[17637]= -114682135;
assign addr[17638]= -76474970;
assign addr[17639]= -38243550;
assign addr[17640]= 0;
assign addr[17641]= 38243550;
assign addr[17642]= 76474970;
assign addr[17643]= 114682135;
assign addr[17644]= 152852926;
assign addr[17645]= 190975237;
assign addr[17646]= 229036977;
assign addr[17647]= 267026072;
assign addr[17648]= 304930476;
assign addr[17649]= 342738165;
assign addr[17650]= 380437148;
assign addr[17651]= 418015468;
assign addr[17652]= 455461206;
assign addr[17653]= 492762486;
assign addr[17654]= 529907477;
assign addr[17655]= 566884397;
assign addr[17656]= 603681519;
assign addr[17657]= 640287172;
assign addr[17658]= 676689746;
assign addr[17659]= 712877694;
assign addr[17660]= 748839539;
assign addr[17661]= 784563876;
assign addr[17662]= 820039373;
assign addr[17663]= 855254778;
assign addr[17664]= 890198924;
assign addr[17665]= 924860725;
assign addr[17666]= 959229189;
assign addr[17667]= 993293415;
assign addr[17668]= 1027042599;
assign addr[17669]= 1060466036;
assign addr[17670]= 1093553126;
assign addr[17671]= 1126293375;
assign addr[17672]= 1158676398;
assign addr[17673]= 1190691925;
assign addr[17674]= 1222329801;
assign addr[17675]= 1253579991;
assign addr[17676]= 1284432584;
assign addr[17677]= 1314877795;
assign addr[17678]= 1344905966;
assign addr[17679]= 1374507575;
assign addr[17680]= 1403673233;
assign addr[17681]= 1432393688;
assign addr[17682]= 1460659832;
assign addr[17683]= 1488462700;
assign addr[17684]= 1515793473;
assign addr[17685]= 1542643483;
assign addr[17686]= 1569004214;
assign addr[17687]= 1594867305;
assign addr[17688]= 1620224553;
assign addr[17689]= 1645067915;
assign addr[17690]= 1669389513;
assign addr[17691]= 1693181631;
assign addr[17692]= 1716436725;
assign addr[17693]= 1739147417;
assign addr[17694]= 1761306505;
assign addr[17695]= 1782906961;
assign addr[17696]= 1803941934;
assign addr[17697]= 1824404752;
assign addr[17698]= 1844288924;
assign addr[17699]= 1863588145;
assign addr[17700]= 1882296293;
assign addr[17701]= 1900407434;
assign addr[17702]= 1917915825;
assign addr[17703]= 1934815911;
assign addr[17704]= 1951102334;
assign addr[17705]= 1966769926;
assign addr[17706]= 1981813720;
assign addr[17707]= 1996228943;
assign addr[17708]= 2010011024;
assign addr[17709]= 2023155591;
assign addr[17710]= 2035658475;
assign addr[17711]= 2047515711;
assign addr[17712]= 2058723538;
assign addr[17713]= 2069278401;
assign addr[17714]= 2079176953;
assign addr[17715]= 2088416053;
assign addr[17716]= 2096992772;
assign addr[17717]= 2104904390;
assign addr[17718]= 2112148396;
assign addr[17719]= 2118722494;
assign addr[17720]= 2124624598;
assign addr[17721]= 2129852837;
assign addr[17722]= 2134405552;
assign addr[17723]= 2138281298;
assign addr[17724]= 2141478848;
assign addr[17725]= 2143997187;
assign addr[17726]= 2145835515;
assign addr[17727]= 2146993250;
assign addr[17728]= 2147470025;
assign addr[17729]= 2147265689;
assign addr[17730]= 2146380306;
assign addr[17731]= 2144814157;
assign addr[17732]= 2142567738;
assign addr[17733]= 2139641764;
assign addr[17734]= 2136037160;
assign addr[17735]= 2131755071;
assign addr[17736]= 2126796855;
assign addr[17737]= 2121164085;
assign addr[17738]= 2114858546;
assign addr[17739]= 2107882239;
assign addr[17740]= 2100237377;
assign addr[17741]= 2091926384;
assign addr[17742]= 2082951896;
assign addr[17743]= 2073316760;
assign addr[17744]= 2063024031;
assign addr[17745]= 2052076975;
assign addr[17746]= 2040479063;
assign addr[17747]= 2028233973;
assign addr[17748]= 2015345591;
assign addr[17749]= 2001818002;
assign addr[17750]= 1987655498;
assign addr[17751]= 1972862571;
assign addr[17752]= 1957443913;
assign addr[17753]= 1941404413;
assign addr[17754]= 1924749160;
assign addr[17755]= 1907483436;
assign addr[17756]= 1889612716;
assign addr[17757]= 1871142669;
assign addr[17758]= 1852079154;
assign addr[17759]= 1832428215;
assign addr[17760]= 1812196087;
assign addr[17761]= 1791389186;
assign addr[17762]= 1770014111;
assign addr[17763]= 1748077642;
assign addr[17764]= 1725586737;
assign addr[17765]= 1702548529;
assign addr[17766]= 1678970324;
assign addr[17767]= 1654859602;
assign addr[17768]= 1630224009;
assign addr[17769]= 1605071359;
assign addr[17770]= 1579409630;
assign addr[17771]= 1553246960;
assign addr[17772]= 1526591649;
assign addr[17773]= 1499452149;
assign addr[17774]= 1471837070;
assign addr[17775]= 1443755168;
assign addr[17776]= 1415215352;
assign addr[17777]= 1386226674;
assign addr[17778]= 1356798326;
assign addr[17779]= 1326939644;
assign addr[17780]= 1296660098;
assign addr[17781]= 1265969291;
assign addr[17782]= 1234876957;
assign addr[17783]= 1203392958;
assign addr[17784]= 1171527280;
assign addr[17785]= 1139290029;
assign addr[17786]= 1106691431;
assign addr[17787]= 1073741824;
assign addr[17788]= 1040451659;
assign addr[17789]= 1006831495;
assign addr[17790]= 972891995;
assign addr[17791]= 938643924;
assign addr[17792]= 904098143;
assign addr[17793]= 869265610;
assign addr[17794]= 834157373;
assign addr[17795]= 798784567;
assign addr[17796]= 763158411;
assign addr[17797]= 727290205;
assign addr[17798]= 691191324;
assign addr[17799]= 654873219;
assign addr[17800]= 618347408;
assign addr[17801]= 581625477;
assign addr[17802]= 544719071;
assign addr[17803]= 507639898;
assign addr[17804]= 470399716;
assign addr[17805]= 433010339;
assign addr[17806]= 395483624;
assign addr[17807]= 357831473;
assign addr[17808]= 320065829;
assign addr[17809]= 282198671;
assign addr[17810]= 244242007;
assign addr[17811]= 206207878;
assign addr[17812]= 168108346;
assign addr[17813]= 129955495;
assign addr[17814]= 91761426;
assign addr[17815]= 53538253;
assign addr[17816]= 15298099;
assign addr[17817]= -22946906;
assign addr[17818]= -61184634;
assign addr[17819]= -99402956;
assign addr[17820]= -137589750;
assign addr[17821]= -175732905;
assign addr[17822]= -213820322;
assign addr[17823]= -251839923;
assign addr[17824]= -289779648;
assign addr[17825]= -327627463;
assign addr[17826]= -365371365;
assign addr[17827]= -402999383;
assign addr[17828]= -440499581;
assign addr[17829]= -477860067;
assign addr[17830]= -515068990;
assign addr[17831]= -552114549;
assign addr[17832]= -588984994;
assign addr[17833]= -625668632;
assign addr[17834]= -662153826;
assign addr[17835]= -698429006;
assign addr[17836]= -734482665;
assign addr[17837]= -770303369;
assign addr[17838]= -805879757;
assign addr[17839]= -841200544;
assign addr[17840]= -876254528;
assign addr[17841]= -911030591;
assign addr[17842]= -945517704;
assign addr[17843]= -979704927;
assign addr[17844]= -1013581418;
assign addr[17845]= -1047136432;
assign addr[17846]= -1080359326;
assign addr[17847]= -1113239564;
assign addr[17848]= -1145766716;
assign addr[17849]= -1177930466;
assign addr[17850]= -1209720613;
assign addr[17851]= -1241127074;
assign addr[17852]= -1272139887;
assign addr[17853]= -1302749217;
assign addr[17854]= -1332945355;
assign addr[17855]= -1362718723;
assign addr[17856]= -1392059879;
assign addr[17857]= -1420959516;
assign addr[17858]= -1449408469;
assign addr[17859]= -1477397714;
assign addr[17860]= -1504918373;
assign addr[17861]= -1531961719;
assign addr[17862]= -1558519173;
assign addr[17863]= -1584582314;
assign addr[17864]= -1610142873;
assign addr[17865]= -1635192744;
assign addr[17866]= -1659723983;
assign addr[17867]= -1683728808;
assign addr[17868]= -1707199606;
assign addr[17869]= -1730128933;
assign addr[17870]= -1752509516;
assign addr[17871]= -1774334257;
assign addr[17872]= -1795596234;
assign addr[17873]= -1816288703;
assign addr[17874]= -1836405100;
assign addr[17875]= -1855939047;
assign addr[17876]= -1874884346;
assign addr[17877]= -1893234990;
assign addr[17878]= -1910985158;
assign addr[17879]= -1928129220;
assign addr[17880]= -1944661739;
assign addr[17881]= -1960577471;
assign addr[17882]= -1975871368;
assign addr[17883]= -1990538579;
assign addr[17884]= -2004574453;
assign addr[17885]= -2017974537;
assign addr[17886]= -2030734582;
assign addr[17887]= -2042850540;
assign addr[17888]= -2054318569;
assign addr[17889]= -2065135031;
assign addr[17890]= -2075296495;
assign addr[17891]= -2084799740;
assign addr[17892]= -2093641749;
assign addr[17893]= -2101819720;
assign addr[17894]= -2109331059;
assign addr[17895]= -2116173382;
assign addr[17896]= -2122344521;
assign addr[17897]= -2127842516;
assign addr[17898]= -2132665626;
assign addr[17899]= -2136812319;
assign addr[17900]= -2140281282;
assign addr[17901]= -2143071413;
assign addr[17902]= -2145181827;
assign addr[17903]= -2146611856;
assign addr[17904]= -2147361045;
assign addr[17905]= -2147429158;
assign addr[17906]= -2146816171;
assign addr[17907]= -2145522281;
assign addr[17908]= -2143547897;
assign addr[17909]= -2140893646;
assign addr[17910]= -2137560369;
assign addr[17911]= -2133549123;
assign addr[17912]= -2128861181;
assign addr[17913]= -2123498030;
assign addr[17914]= -2117461370;
assign addr[17915]= -2110753117;
assign addr[17916]= -2103375398;
assign addr[17917]= -2095330553;
assign addr[17918]= -2086621133;
assign addr[17919]= -2077249901;
assign addr[17920]= -2067219829;
assign addr[17921]= -2056534099;
assign addr[17922]= -2045196100;
assign addr[17923]= -2033209426;
assign addr[17924]= -2020577882;
assign addr[17925]= -2007305472;
assign addr[17926]= -1993396407;
assign addr[17927]= -1978855097;
assign addr[17928]= -1963686155;
assign addr[17929]= -1947894393;
assign addr[17930]= -1931484818;
assign addr[17931]= -1914462636;
assign addr[17932]= -1896833245;
assign addr[17933]= -1878602237;
assign addr[17934]= -1859775393;
assign addr[17935]= -1840358687;
assign addr[17936]= -1820358275;
assign addr[17937]= -1799780501;
assign addr[17938]= -1778631892;
assign addr[17939]= -1756919156;
assign addr[17940]= -1734649179;
assign addr[17941]= -1711829025;
assign addr[17942]= -1688465931;
assign addr[17943]= -1664567307;
assign addr[17944]= -1640140734;
assign addr[17945]= -1615193959;
assign addr[17946]= -1589734894;
assign addr[17947]= -1563771613;
assign addr[17948]= -1537312353;
assign addr[17949]= -1510365504;
assign addr[17950]= -1482939614;
assign addr[17951]= -1455043381;
assign addr[17952]= -1426685652;
assign addr[17953]= -1397875423;
assign addr[17954]= -1368621831;
assign addr[17955]= -1338934154;
assign addr[17956]= -1308821808;
assign addr[17957]= -1278294345;
assign addr[17958]= -1247361445;
assign addr[17959]= -1216032921;
assign addr[17960]= -1184318708;
assign addr[17961]= -1152228866;
assign addr[17962]= -1119773573;
assign addr[17963]= -1086963121;
assign addr[17964]= -1053807919;
assign addr[17965]= -1020318481;
assign addr[17966]= -986505429;
assign addr[17967]= -952379488;
assign addr[17968]= -917951481;
assign addr[17969]= -883232329;
assign addr[17970]= -848233042;
assign addr[17971]= -812964722;
assign addr[17972]= -777438554;
assign addr[17973]= -741665807;
assign addr[17974]= -705657826;
assign addr[17975]= -669426032;
assign addr[17976]= -632981917;
assign addr[17977]= -596337040;
assign addr[17978]= -559503022;
assign addr[17979]= -522491548;
assign addr[17980]= -485314355;
assign addr[17981]= -447983235;
assign addr[17982]= -410510029;
assign addr[17983]= -372906622;
assign addr[17984]= -335184940;
assign addr[17985]= -297356948;
assign addr[17986]= -259434643;
assign addr[17987]= -221430054;
assign addr[17988]= -183355234;
assign addr[17989]= -145222259;
assign addr[17990]= -107043224;
assign addr[17991]= -68830239;
assign addr[17992]= -30595422;
assign addr[17993]= 7649098;
assign addr[17994]= 45891193;
assign addr[17995]= 84118732;
assign addr[17996]= 122319591;
assign addr[17997]= 160481654;
assign addr[17998]= 198592817;
assign addr[17999]= 236640993;
assign addr[18000]= 274614114;
assign addr[18001]= 312500135;
assign addr[18002]= 350287041;
assign addr[18003]= 387962847;
assign addr[18004]= 425515602;
assign addr[18005]= 462933398;
assign addr[18006]= 500204365;
assign addr[18007]= 537316682;
assign addr[18008]= 574258580;
assign addr[18009]= 611018340;
assign addr[18010]= 647584304;
assign addr[18011]= 683944874;
assign addr[18012]= 720088517;
assign addr[18013]= 756003771;
assign addr[18014]= 791679244;
assign addr[18015]= 827103620;
assign addr[18016]= 862265664;
assign addr[18017]= 897154224;
assign addr[18018]= 931758235;
assign addr[18019]= 966066720;
assign addr[18020]= 1000068799;
assign addr[18021]= 1033753687;
assign addr[18022]= 1067110699;
assign addr[18023]= 1100129257;
assign addr[18024]= 1132798888;
assign addr[18025]= 1165109230;
assign addr[18026]= 1197050035;
assign addr[18027]= 1228611172;
assign addr[18028]= 1259782632;
assign addr[18029]= 1290554528;
assign addr[18030]= 1320917099;
assign addr[18031]= 1350860716;
assign addr[18032]= 1380375881;
assign addr[18033]= 1409453233;
assign addr[18034]= 1438083551;
assign addr[18035]= 1466257752;
assign addr[18036]= 1493966902;
assign addr[18037]= 1521202211;
assign addr[18038]= 1547955041;
assign addr[18039]= 1574216908;
assign addr[18040]= 1599979481;
assign addr[18041]= 1625234591;
assign addr[18042]= 1649974225;
assign addr[18043]= 1674190539;
assign addr[18044]= 1697875851;
assign addr[18045]= 1721022648;
assign addr[18046]= 1743623590;
assign addr[18047]= 1765671509;
assign addr[18048]= 1787159411;
assign addr[18049]= 1808080480;
assign addr[18050]= 1828428082;
assign addr[18051]= 1848195763;
assign addr[18052]= 1867377253;
assign addr[18053]= 1885966468;
assign addr[18054]= 1903957513;
assign addr[18055]= 1921344681;
assign addr[18056]= 1938122457;
assign addr[18057]= 1954285520;
assign addr[18058]= 1969828744;
assign addr[18059]= 1984747199;
assign addr[18060]= 1999036154;
assign addr[18061]= 2012691075;
assign addr[18062]= 2025707632;
assign addr[18063]= 2038081698;
assign addr[18064]= 2049809346;
assign addr[18065]= 2060886858;
assign addr[18066]= 2071310720;
assign addr[18067]= 2081077626;
assign addr[18068]= 2090184478;
assign addr[18069]= 2098628387;
assign addr[18070]= 2106406677;
assign addr[18071]= 2113516878;
assign addr[18072]= 2119956737;
assign addr[18073]= 2125724211;
assign addr[18074]= 2130817471;
assign addr[18075]= 2135234901;
assign addr[18076]= 2138975100;
assign addr[18077]= 2142036881;
assign addr[18078]= 2144419275;
assign addr[18079]= 2146121524;
assign addr[18080]= 2147143090;
assign addr[18081]= 2147483648;
assign addr[18082]= 2147143090;
assign addr[18083]= 2146121524;
assign addr[18084]= 2144419275;
assign addr[18085]= 2142036881;
assign addr[18086]= 2138975100;
assign addr[18087]= 2135234901;
assign addr[18088]= 2130817471;
assign addr[18089]= 2125724211;
assign addr[18090]= 2119956737;
assign addr[18091]= 2113516878;
assign addr[18092]= 2106406677;
assign addr[18093]= 2098628387;
assign addr[18094]= 2090184478;
assign addr[18095]= 2081077626;
assign addr[18096]= 2071310720;
assign addr[18097]= 2060886858;
assign addr[18098]= 2049809346;
assign addr[18099]= 2038081698;
assign addr[18100]= 2025707632;
assign addr[18101]= 2012691075;
assign addr[18102]= 1999036154;
assign addr[18103]= 1984747199;
assign addr[18104]= 1969828744;
assign addr[18105]= 1954285520;
assign addr[18106]= 1938122457;
assign addr[18107]= 1921344681;
assign addr[18108]= 1903957513;
assign addr[18109]= 1885966468;
assign addr[18110]= 1867377253;
assign addr[18111]= 1848195763;
assign addr[18112]= 1828428082;
assign addr[18113]= 1808080480;
assign addr[18114]= 1787159411;
assign addr[18115]= 1765671509;
assign addr[18116]= 1743623590;
assign addr[18117]= 1721022648;
assign addr[18118]= 1697875851;
assign addr[18119]= 1674190539;
assign addr[18120]= 1649974225;
assign addr[18121]= 1625234591;
assign addr[18122]= 1599979481;
assign addr[18123]= 1574216908;
assign addr[18124]= 1547955041;
assign addr[18125]= 1521202211;
assign addr[18126]= 1493966902;
assign addr[18127]= 1466257752;
assign addr[18128]= 1438083551;
assign addr[18129]= 1409453233;
assign addr[18130]= 1380375881;
assign addr[18131]= 1350860716;
assign addr[18132]= 1320917099;
assign addr[18133]= 1290554528;
assign addr[18134]= 1259782632;
assign addr[18135]= 1228611172;
assign addr[18136]= 1197050035;
assign addr[18137]= 1165109230;
assign addr[18138]= 1132798888;
assign addr[18139]= 1100129257;
assign addr[18140]= 1067110699;
assign addr[18141]= 1033753687;
assign addr[18142]= 1000068799;
assign addr[18143]= 966066720;
assign addr[18144]= 931758235;
assign addr[18145]= 897154224;
assign addr[18146]= 862265664;
assign addr[18147]= 827103620;
assign addr[18148]= 791679244;
assign addr[18149]= 756003771;
assign addr[18150]= 720088517;
assign addr[18151]= 683944874;
assign addr[18152]= 647584304;
assign addr[18153]= 611018340;
assign addr[18154]= 574258580;
assign addr[18155]= 537316682;
assign addr[18156]= 500204365;
assign addr[18157]= 462933398;
assign addr[18158]= 425515602;
assign addr[18159]= 387962847;
assign addr[18160]= 350287041;
assign addr[18161]= 312500135;
assign addr[18162]= 274614114;
assign addr[18163]= 236640993;
assign addr[18164]= 198592817;
assign addr[18165]= 160481654;
assign addr[18166]= 122319591;
assign addr[18167]= 84118732;
assign addr[18168]= 45891193;
assign addr[18169]= 7649098;
assign addr[18170]= -30595422;
assign addr[18171]= -68830239;
assign addr[18172]= -107043224;
assign addr[18173]= -145222259;
assign addr[18174]= -183355234;
assign addr[18175]= -221430054;
assign addr[18176]= -259434643;
assign addr[18177]= -297356948;
assign addr[18178]= -335184940;
assign addr[18179]= -372906622;
assign addr[18180]= -410510029;
assign addr[18181]= -447983235;
assign addr[18182]= -485314355;
assign addr[18183]= -522491548;
assign addr[18184]= -559503022;
assign addr[18185]= -596337040;
assign addr[18186]= -632981917;
assign addr[18187]= -669426032;
assign addr[18188]= -705657826;
assign addr[18189]= -741665807;
assign addr[18190]= -777438554;
assign addr[18191]= -812964722;
assign addr[18192]= -848233042;
assign addr[18193]= -883232329;
assign addr[18194]= -917951481;
assign addr[18195]= -952379488;
assign addr[18196]= -986505429;
assign addr[18197]= -1020318481;
assign addr[18198]= -1053807919;
assign addr[18199]= -1086963121;
assign addr[18200]= -1119773573;
assign addr[18201]= -1152228866;
assign addr[18202]= -1184318708;
assign addr[18203]= -1216032921;
assign addr[18204]= -1247361445;
assign addr[18205]= -1278294345;
assign addr[18206]= -1308821808;
assign addr[18207]= -1338934154;
assign addr[18208]= -1368621831;
assign addr[18209]= -1397875423;
assign addr[18210]= -1426685652;
assign addr[18211]= -1455043381;
assign addr[18212]= -1482939614;
assign addr[18213]= -1510365504;
assign addr[18214]= -1537312353;
assign addr[18215]= -1563771613;
assign addr[18216]= -1589734894;
assign addr[18217]= -1615193959;
assign addr[18218]= -1640140734;
assign addr[18219]= -1664567307;
assign addr[18220]= -1688465931;
assign addr[18221]= -1711829025;
assign addr[18222]= -1734649179;
assign addr[18223]= -1756919156;
assign addr[18224]= -1778631892;
assign addr[18225]= -1799780501;
assign addr[18226]= -1820358275;
assign addr[18227]= -1840358687;
assign addr[18228]= -1859775393;
assign addr[18229]= -1878602237;
assign addr[18230]= -1896833245;
assign addr[18231]= -1914462636;
assign addr[18232]= -1931484818;
assign addr[18233]= -1947894393;
assign addr[18234]= -1963686155;
assign addr[18235]= -1978855097;
assign addr[18236]= -1993396407;
assign addr[18237]= -2007305472;
assign addr[18238]= -2020577882;
assign addr[18239]= -2033209426;
assign addr[18240]= -2045196100;
assign addr[18241]= -2056534099;
assign addr[18242]= -2067219829;
assign addr[18243]= -2077249901;
assign addr[18244]= -2086621133;
assign addr[18245]= -2095330553;
assign addr[18246]= -2103375398;
assign addr[18247]= -2110753117;
assign addr[18248]= -2117461370;
assign addr[18249]= -2123498030;
assign addr[18250]= -2128861181;
assign addr[18251]= -2133549123;
assign addr[18252]= -2137560369;
assign addr[18253]= -2140893646;
assign addr[18254]= -2143547897;
assign addr[18255]= -2145522281;
assign addr[18256]= -2146816171;
assign addr[18257]= -2147429158;
assign addr[18258]= -2147361045;
assign addr[18259]= -2146611856;
assign addr[18260]= -2145181827;
assign addr[18261]= -2143071413;
assign addr[18262]= -2140281282;
assign addr[18263]= -2136812319;
assign addr[18264]= -2132665626;
assign addr[18265]= -2127842516;
assign addr[18266]= -2122344521;
assign addr[18267]= -2116173382;
assign addr[18268]= -2109331059;
assign addr[18269]= -2101819720;
assign addr[18270]= -2093641749;
assign addr[18271]= -2084799740;
assign addr[18272]= -2075296495;
assign addr[18273]= -2065135031;
assign addr[18274]= -2054318569;
assign addr[18275]= -2042850540;
assign addr[18276]= -2030734582;
assign addr[18277]= -2017974537;
assign addr[18278]= -2004574453;
assign addr[18279]= -1990538579;
assign addr[18280]= -1975871368;
assign addr[18281]= -1960577471;
assign addr[18282]= -1944661739;
assign addr[18283]= -1928129220;
assign addr[18284]= -1910985158;
assign addr[18285]= -1893234990;
assign addr[18286]= -1874884346;
assign addr[18287]= -1855939047;
assign addr[18288]= -1836405100;
assign addr[18289]= -1816288703;
assign addr[18290]= -1795596234;
assign addr[18291]= -1774334257;
assign addr[18292]= -1752509516;
assign addr[18293]= -1730128933;
assign addr[18294]= -1707199606;
assign addr[18295]= -1683728808;
assign addr[18296]= -1659723983;
assign addr[18297]= -1635192744;
assign addr[18298]= -1610142873;
assign addr[18299]= -1584582314;
assign addr[18300]= -1558519173;
assign addr[18301]= -1531961719;
assign addr[18302]= -1504918373;
assign addr[18303]= -1477397714;
assign addr[18304]= -1449408469;
assign addr[18305]= -1420959516;
assign addr[18306]= -1392059879;
assign addr[18307]= -1362718723;
assign addr[18308]= -1332945355;
assign addr[18309]= -1302749217;
assign addr[18310]= -1272139887;
assign addr[18311]= -1241127074;
assign addr[18312]= -1209720613;
assign addr[18313]= -1177930466;
assign addr[18314]= -1145766716;
assign addr[18315]= -1113239564;
assign addr[18316]= -1080359326;
assign addr[18317]= -1047136432;
assign addr[18318]= -1013581418;
assign addr[18319]= -979704927;
assign addr[18320]= -945517704;
assign addr[18321]= -911030591;
assign addr[18322]= -876254528;
assign addr[18323]= -841200544;
assign addr[18324]= -805879757;
assign addr[18325]= -770303369;
assign addr[18326]= -734482665;
assign addr[18327]= -698429006;
assign addr[18328]= -662153826;
assign addr[18329]= -625668632;
assign addr[18330]= -588984994;
assign addr[18331]= -552114549;
assign addr[18332]= -515068990;
assign addr[18333]= -477860067;
assign addr[18334]= -440499581;
assign addr[18335]= -402999383;
assign addr[18336]= -365371365;
assign addr[18337]= -327627463;
assign addr[18338]= -289779648;
assign addr[18339]= -251839923;
assign addr[18340]= -213820322;
assign addr[18341]= -175732905;
assign addr[18342]= -137589750;
assign addr[18343]= -99402956;
assign addr[18344]= -61184634;
assign addr[18345]= -22946906;
assign addr[18346]= 15298099;
assign addr[18347]= 53538253;
assign addr[18348]= 91761426;
assign addr[18349]= 129955495;
assign addr[18350]= 168108346;
assign addr[18351]= 206207878;
assign addr[18352]= 244242007;
assign addr[18353]= 282198671;
assign addr[18354]= 320065829;
assign addr[18355]= 357831473;
assign addr[18356]= 395483624;
assign addr[18357]= 433010339;
assign addr[18358]= 470399716;
assign addr[18359]= 507639898;
assign addr[18360]= 544719071;
assign addr[18361]= 581625477;
assign addr[18362]= 618347408;
assign addr[18363]= 654873219;
assign addr[18364]= 691191324;
assign addr[18365]= 727290205;
assign addr[18366]= 763158411;
assign addr[18367]= 798784567;
assign addr[18368]= 834157373;
assign addr[18369]= 869265610;
assign addr[18370]= 904098143;
assign addr[18371]= 938643924;
assign addr[18372]= 972891995;
assign addr[18373]= 1006831495;
assign addr[18374]= 1040451659;
assign addr[18375]= 1073741824;
assign addr[18376]= 1106691431;
assign addr[18377]= 1139290029;
assign addr[18378]= 1171527280;
assign addr[18379]= 1203392958;
assign addr[18380]= 1234876957;
assign addr[18381]= 1265969291;
assign addr[18382]= 1296660098;
assign addr[18383]= 1326939644;
assign addr[18384]= 1356798326;
assign addr[18385]= 1386226674;
assign addr[18386]= 1415215352;
assign addr[18387]= 1443755168;
assign addr[18388]= 1471837070;
assign addr[18389]= 1499452149;
assign addr[18390]= 1526591649;
assign addr[18391]= 1553246960;
assign addr[18392]= 1579409630;
assign addr[18393]= 1605071359;
assign addr[18394]= 1630224009;
assign addr[18395]= 1654859602;
assign addr[18396]= 1678970324;
assign addr[18397]= 1702548529;
assign addr[18398]= 1725586737;
assign addr[18399]= 1748077642;
assign addr[18400]= 1770014111;
assign addr[18401]= 1791389186;
assign addr[18402]= 1812196087;
assign addr[18403]= 1832428215;
assign addr[18404]= 1852079154;
assign addr[18405]= 1871142669;
assign addr[18406]= 1889612716;
assign addr[18407]= 1907483436;
assign addr[18408]= 1924749160;
assign addr[18409]= 1941404413;
assign addr[18410]= 1957443913;
assign addr[18411]= 1972862571;
assign addr[18412]= 1987655498;
assign addr[18413]= 2001818002;
assign addr[18414]= 2015345591;
assign addr[18415]= 2028233973;
assign addr[18416]= 2040479063;
assign addr[18417]= 2052076975;
assign addr[18418]= 2063024031;
assign addr[18419]= 2073316760;
assign addr[18420]= 2082951896;
assign addr[18421]= 2091926384;
assign addr[18422]= 2100237377;
assign addr[18423]= 2107882239;
assign addr[18424]= 2114858546;
assign addr[18425]= 2121164085;
assign addr[18426]= 2126796855;
assign addr[18427]= 2131755071;
assign addr[18428]= 2136037160;
assign addr[18429]= 2139641764;
assign addr[18430]= 2142567738;
assign addr[18431]= 2144814157;
assign addr[18432]= 2146380306;
assign addr[18433]= 2147265689;
assign addr[18434]= 2147470025;
assign addr[18435]= 2146993250;
assign addr[18436]= 2145835515;
assign addr[18437]= 2143997187;
assign addr[18438]= 2141478848;
assign addr[18439]= 2138281298;
assign addr[18440]= 2134405552;
assign addr[18441]= 2129852837;
assign addr[18442]= 2124624598;
assign addr[18443]= 2118722494;
assign addr[18444]= 2112148396;
assign addr[18445]= 2104904390;
assign addr[18446]= 2096992772;
assign addr[18447]= 2088416053;
assign addr[18448]= 2079176953;
assign addr[18449]= 2069278401;
assign addr[18450]= 2058723538;
assign addr[18451]= 2047515711;
assign addr[18452]= 2035658475;
assign addr[18453]= 2023155591;
assign addr[18454]= 2010011024;
assign addr[18455]= 1996228943;
assign addr[18456]= 1981813720;
assign addr[18457]= 1966769926;
assign addr[18458]= 1951102334;
assign addr[18459]= 1934815911;
assign addr[18460]= 1917915825;
assign addr[18461]= 1900407434;
assign addr[18462]= 1882296293;
assign addr[18463]= 1863588145;
assign addr[18464]= 1844288924;
assign addr[18465]= 1824404752;
assign addr[18466]= 1803941934;
assign addr[18467]= 1782906961;
assign addr[18468]= 1761306505;
assign addr[18469]= 1739147417;
assign addr[18470]= 1716436725;
assign addr[18471]= 1693181631;
assign addr[18472]= 1669389513;
assign addr[18473]= 1645067915;
assign addr[18474]= 1620224553;
assign addr[18475]= 1594867305;
assign addr[18476]= 1569004214;
assign addr[18477]= 1542643483;
assign addr[18478]= 1515793473;
assign addr[18479]= 1488462700;
assign addr[18480]= 1460659832;
assign addr[18481]= 1432393688;
assign addr[18482]= 1403673233;
assign addr[18483]= 1374507575;
assign addr[18484]= 1344905966;
assign addr[18485]= 1314877795;
assign addr[18486]= 1284432584;
assign addr[18487]= 1253579991;
assign addr[18488]= 1222329801;
assign addr[18489]= 1190691925;
assign addr[18490]= 1158676398;
assign addr[18491]= 1126293375;
assign addr[18492]= 1093553126;
assign addr[18493]= 1060466036;
assign addr[18494]= 1027042599;
assign addr[18495]= 993293415;
assign addr[18496]= 959229189;
assign addr[18497]= 924860725;
assign addr[18498]= 890198924;
assign addr[18499]= 855254778;
assign addr[18500]= 820039373;
assign addr[18501]= 784563876;
assign addr[18502]= 748839539;
assign addr[18503]= 712877694;
assign addr[18504]= 676689746;
assign addr[18505]= 640287172;
assign addr[18506]= 603681519;
assign addr[18507]= 566884397;
assign addr[18508]= 529907477;
assign addr[18509]= 492762486;
assign addr[18510]= 455461206;
assign addr[18511]= 418015468;
assign addr[18512]= 380437148;
assign addr[18513]= 342738165;
assign addr[18514]= 304930476;
assign addr[18515]= 267026072;
assign addr[18516]= 229036977;
assign addr[18517]= 190975237;
assign addr[18518]= 152852926;
assign addr[18519]= 114682135;
assign addr[18520]= 76474970;
assign addr[18521]= 38243550;
assign addr[18522]= 0;
assign addr[18523]= -38243550;
assign addr[18524]= -76474970;
assign addr[18525]= -114682135;
assign addr[18526]= -152852926;
assign addr[18527]= -190975237;
assign addr[18528]= -229036977;
assign addr[18529]= -267026072;
assign addr[18530]= -304930476;
assign addr[18531]= -342738165;
assign addr[18532]= -380437148;
assign addr[18533]= -418015468;
assign addr[18534]= -455461206;
assign addr[18535]= -492762486;
assign addr[18536]= -529907477;
assign addr[18537]= -566884397;
assign addr[18538]= -603681519;
assign addr[18539]= -640287172;
assign addr[18540]= -676689746;
assign addr[18541]= -712877694;
assign addr[18542]= -748839539;
assign addr[18543]= -784563876;
assign addr[18544]= -820039373;
assign addr[18545]= -855254778;
assign addr[18546]= -890198924;
assign addr[18547]= -924860725;
assign addr[18548]= -959229189;
assign addr[18549]= -993293415;
assign addr[18550]= -1027042599;
assign addr[18551]= -1060466036;
assign addr[18552]= -1093553126;
assign addr[18553]= -1126293375;
assign addr[18554]= -1158676398;
assign addr[18555]= -1190691925;
assign addr[18556]= -1222329801;
assign addr[18557]= -1253579991;
assign addr[18558]= -1284432584;
assign addr[18559]= -1314877795;
assign addr[18560]= -1344905966;
assign addr[18561]= -1374507575;
assign addr[18562]= -1403673233;
assign addr[18563]= -1432393688;
assign addr[18564]= -1460659832;
assign addr[18565]= -1488462700;
assign addr[18566]= -1515793473;
assign addr[18567]= -1542643483;
assign addr[18568]= -1569004214;
assign addr[18569]= -1594867305;
assign addr[18570]= -1620224553;
assign addr[18571]= -1645067915;
assign addr[18572]= -1669389513;
assign addr[18573]= -1693181631;
assign addr[18574]= -1716436725;
assign addr[18575]= -1739147417;
assign addr[18576]= -1761306505;
assign addr[18577]= -1782906961;
assign addr[18578]= -1803941934;
assign addr[18579]= -1824404752;
assign addr[18580]= -1844288924;
assign addr[18581]= -1863588145;
assign addr[18582]= -1882296293;
assign addr[18583]= -1900407434;
assign addr[18584]= -1917915825;
assign addr[18585]= -1934815911;
assign addr[18586]= -1951102334;
assign addr[18587]= -1966769926;
assign addr[18588]= -1981813720;
assign addr[18589]= -1996228943;
assign addr[18590]= -2010011024;
assign addr[18591]= -2023155591;
assign addr[18592]= -2035658475;
assign addr[18593]= -2047515711;
assign addr[18594]= -2058723538;
assign addr[18595]= -2069278401;
assign addr[18596]= -2079176953;
assign addr[18597]= -2088416053;
assign addr[18598]= -2096992772;
assign addr[18599]= -2104904390;
assign addr[18600]= -2112148396;
assign addr[18601]= -2118722494;
assign addr[18602]= -2124624598;
assign addr[18603]= -2129852837;
assign addr[18604]= -2134405552;
assign addr[18605]= -2138281298;
assign addr[18606]= -2141478848;
assign addr[18607]= -2143997187;
assign addr[18608]= -2145835515;
assign addr[18609]= -2146993250;
assign addr[18610]= -2147470025;
assign addr[18611]= -2147265689;
assign addr[18612]= -2146380306;
assign addr[18613]= -2144814157;
assign addr[18614]= -2142567738;
assign addr[18615]= -2139641764;
assign addr[18616]= -2136037160;
assign addr[18617]= -2131755071;
assign addr[18618]= -2126796855;
assign addr[18619]= -2121164085;
assign addr[18620]= -2114858546;
assign addr[18621]= -2107882239;
assign addr[18622]= -2100237377;
assign addr[18623]= -2091926384;
assign addr[18624]= -2082951896;
assign addr[18625]= -2073316760;
assign addr[18626]= -2063024031;
assign addr[18627]= -2052076975;
assign addr[18628]= -2040479063;
assign addr[18629]= -2028233973;
assign addr[18630]= -2015345591;
assign addr[18631]= -2001818002;
assign addr[18632]= -1987655498;
assign addr[18633]= -1972862571;
assign addr[18634]= -1957443913;
assign addr[18635]= -1941404413;
assign addr[18636]= -1924749160;
assign addr[18637]= -1907483436;
assign addr[18638]= -1889612716;
assign addr[18639]= -1871142669;
assign addr[18640]= -1852079154;
assign addr[18641]= -1832428215;
assign addr[18642]= -1812196087;
assign addr[18643]= -1791389186;
assign addr[18644]= -1770014111;
assign addr[18645]= -1748077642;
assign addr[18646]= -1725586737;
assign addr[18647]= -1702548529;
assign addr[18648]= -1678970324;
assign addr[18649]= -1654859602;
assign addr[18650]= -1630224009;
assign addr[18651]= -1605071359;
assign addr[18652]= -1579409630;
assign addr[18653]= -1553246960;
assign addr[18654]= -1526591649;
assign addr[18655]= -1499452149;
assign addr[18656]= -1471837070;
assign addr[18657]= -1443755168;
assign addr[18658]= -1415215352;
assign addr[18659]= -1386226674;
assign addr[18660]= -1356798326;
assign addr[18661]= -1326939644;
assign addr[18662]= -1296660098;
assign addr[18663]= -1265969291;
assign addr[18664]= -1234876957;
assign addr[18665]= -1203392958;
assign addr[18666]= -1171527280;
assign addr[18667]= -1139290029;
assign addr[18668]= -1106691431;
assign addr[18669]= -1073741824;
assign addr[18670]= -1040451659;
assign addr[18671]= -1006831495;
assign addr[18672]= -972891995;
assign addr[18673]= -938643924;
assign addr[18674]= -904098143;
assign addr[18675]= -869265610;
assign addr[18676]= -834157373;
assign addr[18677]= -798784567;
assign addr[18678]= -763158411;
assign addr[18679]= -727290205;
assign addr[18680]= -691191324;
assign addr[18681]= -654873219;
assign addr[18682]= -618347408;
assign addr[18683]= -581625477;
assign addr[18684]= -544719071;
assign addr[18685]= -507639898;
assign addr[18686]= -470399716;
assign addr[18687]= -433010339;
assign addr[18688]= -395483624;
assign addr[18689]= -357831473;
assign addr[18690]= -320065829;
assign addr[18691]= -282198671;
assign addr[18692]= -244242007;
assign addr[18693]= -206207878;
assign addr[18694]= -168108346;
assign addr[18695]= -129955495;
assign addr[18696]= -91761426;
assign addr[18697]= -53538253;
assign addr[18698]= -15298099;
assign addr[18699]= 22946906;
assign addr[18700]= 61184634;
assign addr[18701]= 99402956;
assign addr[18702]= 137589750;
assign addr[18703]= 175732905;
assign addr[18704]= 213820322;
assign addr[18705]= 251839923;
assign addr[18706]= 289779648;
assign addr[18707]= 327627463;
assign addr[18708]= 365371365;
assign addr[18709]= 402999383;
assign addr[18710]= 440499581;
assign addr[18711]= 477860067;
assign addr[18712]= 515068990;
assign addr[18713]= 552114549;
assign addr[18714]= 588984994;
assign addr[18715]= 625668632;
assign addr[18716]= 662153826;
assign addr[18717]= 698429006;
assign addr[18718]= 734482665;
assign addr[18719]= 770303369;
assign addr[18720]= 805879757;
assign addr[18721]= 841200544;
assign addr[18722]= 876254528;
assign addr[18723]= 911030591;
assign addr[18724]= 945517704;
assign addr[18725]= 979704927;
assign addr[18726]= 1013581418;
assign addr[18727]= 1047136432;
assign addr[18728]= 1080359326;
assign addr[18729]= 1113239564;
assign addr[18730]= 1145766716;
assign addr[18731]= 1177930466;
assign addr[18732]= 1209720613;
assign addr[18733]= 1241127074;
assign addr[18734]= 1272139887;
assign addr[18735]= 1302749217;
assign addr[18736]= 1332945355;
assign addr[18737]= 1362718723;
assign addr[18738]= 1392059879;
assign addr[18739]= 1420959516;
assign addr[18740]= 1449408469;
assign addr[18741]= 1477397714;
assign addr[18742]= 1504918373;
assign addr[18743]= 1531961719;
assign addr[18744]= 1558519173;
assign addr[18745]= 1584582314;
assign addr[18746]= 1610142873;
assign addr[18747]= 1635192744;
assign addr[18748]= 1659723983;
assign addr[18749]= 1683728808;
assign addr[18750]= 1707199606;
assign addr[18751]= 1730128933;
assign addr[18752]= 1752509516;
assign addr[18753]= 1774334257;
assign addr[18754]= 1795596234;
assign addr[18755]= 1816288703;
assign addr[18756]= 1836405100;
assign addr[18757]= 1855939047;
assign addr[18758]= 1874884346;
assign addr[18759]= 1893234990;
assign addr[18760]= 1910985158;
assign addr[18761]= 1928129220;
assign addr[18762]= 1944661739;
assign addr[18763]= 1960577471;
assign addr[18764]= 1975871368;
assign addr[18765]= 1990538579;
assign addr[18766]= 2004574453;
assign addr[18767]= 2017974537;
assign addr[18768]= 2030734582;
assign addr[18769]= 2042850540;
assign addr[18770]= 2054318569;
assign addr[18771]= 2065135031;
assign addr[18772]= 2075296495;
assign addr[18773]= 2084799740;
assign addr[18774]= 2093641749;
assign addr[18775]= 2101819720;
assign addr[18776]= 2109331059;
assign addr[18777]= 2116173382;
assign addr[18778]= 2122344521;
assign addr[18779]= 2127842516;
assign addr[18780]= 2132665626;
assign addr[18781]= 2136812319;
assign addr[18782]= 2140281282;
assign addr[18783]= 2143071413;
assign addr[18784]= 2145181827;
assign addr[18785]= 2146611856;
assign addr[18786]= 2147361045;
assign addr[18787]= 2147429158;
assign addr[18788]= 2146816171;
assign addr[18789]= 2145522281;
assign addr[18790]= 2143547897;
assign addr[18791]= 2140893646;
assign addr[18792]= 2137560369;
assign addr[18793]= 2133549123;
assign addr[18794]= 2128861181;
assign addr[18795]= 2123498030;
assign addr[18796]= 2117461370;
assign addr[18797]= 2110753117;
assign addr[18798]= 2103375398;
assign addr[18799]= 2095330553;
assign addr[18800]= 2086621133;
assign addr[18801]= 2077249901;
assign addr[18802]= 2067219829;
assign addr[18803]= 2056534099;
assign addr[18804]= 2045196100;
assign addr[18805]= 2033209426;
assign addr[18806]= 2020577882;
assign addr[18807]= 2007305472;
assign addr[18808]= 1993396407;
assign addr[18809]= 1978855097;
assign addr[18810]= 1963686155;
assign addr[18811]= 1947894393;
assign addr[18812]= 1931484818;
assign addr[18813]= 1914462636;
assign addr[18814]= 1896833245;
assign addr[18815]= 1878602237;
assign addr[18816]= 1859775393;
assign addr[18817]= 1840358687;
assign addr[18818]= 1820358275;
assign addr[18819]= 1799780501;
assign addr[18820]= 1778631892;
assign addr[18821]= 1756919156;
assign addr[18822]= 1734649179;
assign addr[18823]= 1711829025;
assign addr[18824]= 1688465931;
assign addr[18825]= 1664567307;
assign addr[18826]= 1640140734;
assign addr[18827]= 1615193959;
assign addr[18828]= 1589734894;
assign addr[18829]= 1563771613;
assign addr[18830]= 1537312353;
assign addr[18831]= 1510365504;
assign addr[18832]= 1482939614;
assign addr[18833]= 1455043381;
assign addr[18834]= 1426685652;
assign addr[18835]= 1397875423;
assign addr[18836]= 1368621831;
assign addr[18837]= 1338934154;
assign addr[18838]= 1308821808;
assign addr[18839]= 1278294345;
assign addr[18840]= 1247361445;
assign addr[18841]= 1216032921;
assign addr[18842]= 1184318708;
assign addr[18843]= 1152228866;
assign addr[18844]= 1119773573;
assign addr[18845]= 1086963121;
assign addr[18846]= 1053807919;
assign addr[18847]= 1020318481;
assign addr[18848]= 986505429;
assign addr[18849]= 952379488;
assign addr[18850]= 917951481;
assign addr[18851]= 883232329;
assign addr[18852]= 848233042;
assign addr[18853]= 812964722;
assign addr[18854]= 777438554;
assign addr[18855]= 741665807;
assign addr[18856]= 705657826;
assign addr[18857]= 669426032;
assign addr[18858]= 632981917;
assign addr[18859]= 596337040;
assign addr[18860]= 559503022;
assign addr[18861]= 522491548;
assign addr[18862]= 485314355;
assign addr[18863]= 447983235;
assign addr[18864]= 410510029;
assign addr[18865]= 372906622;
assign addr[18866]= 335184940;
assign addr[18867]= 297356948;
assign addr[18868]= 259434643;
assign addr[18869]= 221430054;
assign addr[18870]= 183355234;
assign addr[18871]= 145222259;
assign addr[18872]= 107043224;
assign addr[18873]= 68830239;
assign addr[18874]= 30595422;
assign addr[18875]= -7649098;
assign addr[18876]= -45891193;
assign addr[18877]= -84118732;
assign addr[18878]= -122319591;
assign addr[18879]= -160481654;
assign addr[18880]= -198592817;
assign addr[18881]= -236640993;
assign addr[18882]= -274614114;
assign addr[18883]= -312500135;
assign addr[18884]= -350287041;
assign addr[18885]= -387962847;
assign addr[18886]= -425515602;
assign addr[18887]= -462933398;
assign addr[18888]= -500204365;
assign addr[18889]= -537316682;
assign addr[18890]= -574258580;
assign addr[18891]= -611018340;
assign addr[18892]= -647584304;
assign addr[18893]= -683944874;
assign addr[18894]= -720088517;
assign addr[18895]= -756003771;
assign addr[18896]= -791679244;
assign addr[18897]= -827103620;
assign addr[18898]= -862265664;
assign addr[18899]= -897154224;
assign addr[18900]= -931758235;
assign addr[18901]= -966066720;
assign addr[18902]= -1000068799;
assign addr[18903]= -1033753687;
assign addr[18904]= -1067110699;
assign addr[18905]= -1100129257;
assign addr[18906]= -1132798888;
assign addr[18907]= -1165109230;
assign addr[18908]= -1197050035;
assign addr[18909]= -1228611172;
assign addr[18910]= -1259782632;
assign addr[18911]= -1290554528;
assign addr[18912]= -1320917099;
assign addr[18913]= -1350860716;
assign addr[18914]= -1380375881;
assign addr[18915]= -1409453233;
assign addr[18916]= -1438083551;
assign addr[18917]= -1466257752;
assign addr[18918]= -1493966902;
assign addr[18919]= -1521202211;
assign addr[18920]= -1547955041;
assign addr[18921]= -1574216908;
assign addr[18922]= -1599979481;
assign addr[18923]= -1625234591;
assign addr[18924]= -1649974225;
assign addr[18925]= -1674190539;
assign addr[18926]= -1697875851;
assign addr[18927]= -1721022648;
assign addr[18928]= -1743623590;
assign addr[18929]= -1765671509;
assign addr[18930]= -1787159411;
assign addr[18931]= -1808080480;
assign addr[18932]= -1828428082;
assign addr[18933]= -1848195763;
assign addr[18934]= -1867377253;
assign addr[18935]= -1885966468;
assign addr[18936]= -1903957513;
assign addr[18937]= -1921344681;
assign addr[18938]= -1938122457;
assign addr[18939]= -1954285520;
assign addr[18940]= -1969828744;
assign addr[18941]= -1984747199;
assign addr[18942]= -1999036154;
assign addr[18943]= -2012691075;
assign addr[18944]= -2025707632;
assign addr[18945]= -2038081698;
assign addr[18946]= -2049809346;
assign addr[18947]= -2060886858;
assign addr[18948]= -2071310720;
assign addr[18949]= -2081077626;
assign addr[18950]= -2090184478;
assign addr[18951]= -2098628387;
assign addr[18952]= -2106406677;
assign addr[18953]= -2113516878;
assign addr[18954]= -2119956737;
assign addr[18955]= -2125724211;
assign addr[18956]= -2130817471;
assign addr[18957]= -2135234901;
assign addr[18958]= -2138975100;
assign addr[18959]= -2142036881;
assign addr[18960]= -2144419275;
assign addr[18961]= -2146121524;
assign addr[18962]= -2147143090;
assign addr[18963]= -2147483648;
assign addr[18964]= -2147143090;
assign addr[18965]= -2146121524;
assign addr[18966]= -2144419275;
assign addr[18967]= -2142036881;
assign addr[18968]= -2138975100;
assign addr[18969]= -2135234901;
assign addr[18970]= -2130817471;
assign addr[18971]= -2125724211;
assign addr[18972]= -2119956737;
assign addr[18973]= -2113516878;
assign addr[18974]= -2106406677;
assign addr[18975]= -2098628387;
assign addr[18976]= -2090184478;
assign addr[18977]= -2081077626;
assign addr[18978]= -2071310720;
assign addr[18979]= -2060886858;
assign addr[18980]= -2049809346;
assign addr[18981]= -2038081698;
assign addr[18982]= -2025707632;
assign addr[18983]= -2012691075;
assign addr[18984]= -1999036154;
assign addr[18985]= -1984747199;
assign addr[18986]= -1969828744;
assign addr[18987]= -1954285520;
assign addr[18988]= -1938122457;
assign addr[18989]= -1921344681;
assign addr[18990]= -1903957513;
assign addr[18991]= -1885966468;
assign addr[18992]= -1867377253;
assign addr[18993]= -1848195763;
assign addr[18994]= -1828428082;
assign addr[18995]= -1808080480;
assign addr[18996]= -1787159411;
assign addr[18997]= -1765671509;
assign addr[18998]= -1743623590;
assign addr[18999]= -1721022648;
assign addr[19000]= -1697875851;
assign addr[19001]= -1674190539;
assign addr[19002]= -1649974225;
assign addr[19003]= -1625234591;
assign addr[19004]= -1599979481;
assign addr[19005]= -1574216908;
assign addr[19006]= -1547955041;
assign addr[19007]= -1521202211;
assign addr[19008]= -1493966902;
assign addr[19009]= -1466257752;
assign addr[19010]= -1438083551;
assign addr[19011]= -1409453233;
assign addr[19012]= -1380375881;
assign addr[19013]= -1350860716;
assign addr[19014]= -1320917099;
assign addr[19015]= -1290554528;
assign addr[19016]= -1259782632;
assign addr[19017]= -1228611172;
assign addr[19018]= -1197050035;
assign addr[19019]= -1165109230;
assign addr[19020]= -1132798888;
assign addr[19021]= -1100129257;
assign addr[19022]= -1067110699;
assign addr[19023]= -1033753687;
assign addr[19024]= -1000068799;
assign addr[19025]= -966066720;
assign addr[19026]= -931758235;
assign addr[19027]= -897154224;
assign addr[19028]= -862265664;
assign addr[19029]= -827103620;
assign addr[19030]= -791679244;
assign addr[19031]= -756003771;
assign addr[19032]= -720088517;
assign addr[19033]= -683944874;
assign addr[19034]= -647584304;
assign addr[19035]= -611018340;
assign addr[19036]= -574258580;
assign addr[19037]= -537316682;
assign addr[19038]= -500204365;
assign addr[19039]= -462933398;
assign addr[19040]= -425515602;
assign addr[19041]= -387962847;
assign addr[19042]= -350287041;
assign addr[19043]= -312500135;
assign addr[19044]= -274614114;
assign addr[19045]= -236640993;
assign addr[19046]= -198592817;
assign addr[19047]= -160481654;
assign addr[19048]= -122319591;
assign addr[19049]= -84118732;
assign addr[19050]= -45891193;
assign addr[19051]= -7649098;
assign addr[19052]= 30595422;
assign addr[19053]= 68830239;
assign addr[19054]= 107043224;
assign addr[19055]= 145222259;
assign addr[19056]= 183355234;
assign addr[19057]= 221430054;
assign addr[19058]= 259434643;
assign addr[19059]= 297356948;
assign addr[19060]= 335184940;
assign addr[19061]= 372906622;
assign addr[19062]= 410510029;
assign addr[19063]= 447983235;
assign addr[19064]= 485314355;
assign addr[19065]= 522491548;
assign addr[19066]= 559503022;
assign addr[19067]= 596337040;
assign addr[19068]= 632981917;
assign addr[19069]= 669426032;
assign addr[19070]= 705657826;
assign addr[19071]= 741665807;
assign addr[19072]= 777438554;
assign addr[19073]= 812964722;
assign addr[19074]= 848233042;
assign addr[19075]= 883232329;
assign addr[19076]= 917951481;
assign addr[19077]= 952379488;
assign addr[19078]= 986505429;
assign addr[19079]= 1020318481;
assign addr[19080]= 1053807919;
assign addr[19081]= 1086963121;
assign addr[19082]= 1119773573;
assign addr[19083]= 1152228866;
assign addr[19084]= 1184318708;
assign addr[19085]= 1216032921;
assign addr[19086]= 1247361445;
assign addr[19087]= 1278294345;
assign addr[19088]= 1308821808;
assign addr[19089]= 1338934154;
assign addr[19090]= 1368621831;
assign addr[19091]= 1397875423;
assign addr[19092]= 1426685652;
assign addr[19093]= 1455043381;
assign addr[19094]= 1482939614;
assign addr[19095]= 1510365504;
assign addr[19096]= 1537312353;
assign addr[19097]= 1563771613;
assign addr[19098]= 1589734894;
assign addr[19099]= 1615193959;
assign addr[19100]= 1640140734;
assign addr[19101]= 1664567307;
assign addr[19102]= 1688465931;
assign addr[19103]= 1711829025;
assign addr[19104]= 1734649179;
assign addr[19105]= 1756919156;
assign addr[19106]= 1778631892;
assign addr[19107]= 1799780501;
assign addr[19108]= 1820358275;
assign addr[19109]= 1840358687;
assign addr[19110]= 1859775393;
assign addr[19111]= 1878602237;
assign addr[19112]= 1896833245;
assign addr[19113]= 1914462636;
assign addr[19114]= 1931484818;
assign addr[19115]= 1947894393;
assign addr[19116]= 1963686155;
assign addr[19117]= 1978855097;
assign addr[19118]= 1993396407;
assign addr[19119]= 2007305472;
assign addr[19120]= 2020577882;
assign addr[19121]= 2033209426;
assign addr[19122]= 2045196100;
assign addr[19123]= 2056534099;
assign addr[19124]= 2067219829;
assign addr[19125]= 2077249901;
assign addr[19126]= 2086621133;
assign addr[19127]= 2095330553;
assign addr[19128]= 2103375398;
assign addr[19129]= 2110753117;
assign addr[19130]= 2117461370;
assign addr[19131]= 2123498030;
assign addr[19132]= 2128861181;
assign addr[19133]= 2133549123;
assign addr[19134]= 2137560369;
assign addr[19135]= 2140893646;
assign addr[19136]= 2143547897;
assign addr[19137]= 2145522281;
assign addr[19138]= 2146816171;
assign addr[19139]= 2147429158;
assign addr[19140]= 2147361045;
assign addr[19141]= 2146611856;
assign addr[19142]= 2145181827;
assign addr[19143]= 2143071413;
assign addr[19144]= 2140281282;
assign addr[19145]= 2136812319;
assign addr[19146]= 2132665626;
assign addr[19147]= 2127842516;
assign addr[19148]= 2122344521;
assign addr[19149]= 2116173382;
assign addr[19150]= 2109331059;
assign addr[19151]= 2101819720;
assign addr[19152]= 2093641749;
assign addr[19153]= 2084799740;
assign addr[19154]= 2075296495;
assign addr[19155]= 2065135031;
assign addr[19156]= 2054318569;
assign addr[19157]= 2042850540;
assign addr[19158]= 2030734582;
assign addr[19159]= 2017974537;
assign addr[19160]= 2004574453;
assign addr[19161]= 1990538579;
assign addr[19162]= 1975871368;
assign addr[19163]= 1960577471;
assign addr[19164]= 1944661739;
assign addr[19165]= 1928129220;
assign addr[19166]= 1910985158;
assign addr[19167]= 1893234990;
assign addr[19168]= 1874884346;
assign addr[19169]= 1855939047;
assign addr[19170]= 1836405100;
assign addr[19171]= 1816288703;
assign addr[19172]= 1795596234;
assign addr[19173]= 1774334257;
assign addr[19174]= 1752509516;
assign addr[19175]= 1730128933;
assign addr[19176]= 1707199606;
assign addr[19177]= 1683728808;
assign addr[19178]= 1659723983;
assign addr[19179]= 1635192744;
assign addr[19180]= 1610142873;
assign addr[19181]= 1584582314;
assign addr[19182]= 1558519173;
assign addr[19183]= 1531961719;
assign addr[19184]= 1504918373;
assign addr[19185]= 1477397714;
assign addr[19186]= 1449408469;
assign addr[19187]= 1420959516;
assign addr[19188]= 1392059879;
assign addr[19189]= 1362718723;
assign addr[19190]= 1332945355;
assign addr[19191]= 1302749217;
assign addr[19192]= 1272139887;
assign addr[19193]= 1241127074;
assign addr[19194]= 1209720613;
assign addr[19195]= 1177930466;
assign addr[19196]= 1145766716;
assign addr[19197]= 1113239564;
assign addr[19198]= 1080359326;
assign addr[19199]= 1047136432;
assign addr[19200]= 1013581418;
assign addr[19201]= 979704927;
assign addr[19202]= 945517704;
assign addr[19203]= 911030591;
assign addr[19204]= 876254528;
assign addr[19205]= 841200544;
assign addr[19206]= 805879757;
assign addr[19207]= 770303369;
assign addr[19208]= 734482665;
assign addr[19209]= 698429006;
assign addr[19210]= 662153826;
assign addr[19211]= 625668632;
assign addr[19212]= 588984994;
assign addr[19213]= 552114549;
assign addr[19214]= 515068990;
assign addr[19215]= 477860067;
assign addr[19216]= 440499581;
assign addr[19217]= 402999383;
assign addr[19218]= 365371365;
assign addr[19219]= 327627463;
assign addr[19220]= 289779648;
assign addr[19221]= 251839923;
assign addr[19222]= 213820322;
assign addr[19223]= 175732905;
assign addr[19224]= 137589750;
assign addr[19225]= 99402956;
assign addr[19226]= 61184634;
assign addr[19227]= 22946906;
assign addr[19228]= -15298099;
assign addr[19229]= -53538253;
assign addr[19230]= -91761426;
assign addr[19231]= -129955495;
assign addr[19232]= -168108346;
assign addr[19233]= -206207878;
assign addr[19234]= -244242007;
assign addr[19235]= -282198671;
assign addr[19236]= -320065829;
assign addr[19237]= -357831473;
assign addr[19238]= -395483624;
assign addr[19239]= -433010339;
assign addr[19240]= -470399716;
assign addr[19241]= -507639898;
assign addr[19242]= -544719071;
assign addr[19243]= -581625477;
assign addr[19244]= -618347408;
assign addr[19245]= -654873219;
assign addr[19246]= -691191324;
assign addr[19247]= -727290205;
assign addr[19248]= -763158411;
assign addr[19249]= -798784567;
assign addr[19250]= -834157373;
assign addr[19251]= -869265610;
assign addr[19252]= -904098143;
assign addr[19253]= -938643924;
assign addr[19254]= -972891995;
assign addr[19255]= -1006831495;
assign addr[19256]= -1040451659;
assign addr[19257]= -1073741824;
assign addr[19258]= -1106691431;
assign addr[19259]= -1139290029;
assign addr[19260]= -1171527280;
assign addr[19261]= -1203392958;
assign addr[19262]= -1234876957;
assign addr[19263]= -1265969291;
assign addr[19264]= -1296660098;
assign addr[19265]= -1326939644;
assign addr[19266]= -1356798326;
assign addr[19267]= -1386226674;
assign addr[19268]= -1415215352;
assign addr[19269]= -1443755168;
assign addr[19270]= -1471837070;
assign addr[19271]= -1499452149;
assign addr[19272]= -1526591649;
assign addr[19273]= -1553246960;
assign addr[19274]= -1579409630;
assign addr[19275]= -1605071359;
assign addr[19276]= -1630224009;
assign addr[19277]= -1654859602;
assign addr[19278]= -1678970324;
assign addr[19279]= -1702548529;
assign addr[19280]= -1725586737;
assign addr[19281]= -1748077642;
assign addr[19282]= -1770014111;
assign addr[19283]= -1791389186;
assign addr[19284]= -1812196087;
assign addr[19285]= -1832428215;
assign addr[19286]= -1852079154;
assign addr[19287]= -1871142669;
assign addr[19288]= -1889612716;
assign addr[19289]= -1907483436;
assign addr[19290]= -1924749160;
assign addr[19291]= -1941404413;
assign addr[19292]= -1957443913;
assign addr[19293]= -1972862571;
assign addr[19294]= -1987655498;
assign addr[19295]= -2001818002;
assign addr[19296]= -2015345591;
assign addr[19297]= -2028233973;
assign addr[19298]= -2040479063;
assign addr[19299]= -2052076975;
assign addr[19300]= -2063024031;
assign addr[19301]= -2073316760;
assign addr[19302]= -2082951896;
assign addr[19303]= -2091926384;
assign addr[19304]= -2100237377;
assign addr[19305]= -2107882239;
assign addr[19306]= -2114858546;
assign addr[19307]= -2121164085;
assign addr[19308]= -2126796855;
assign addr[19309]= -2131755071;
assign addr[19310]= -2136037160;
assign addr[19311]= -2139641764;
assign addr[19312]= -2142567738;
assign addr[19313]= -2144814157;
assign addr[19314]= -2146380306;
assign addr[19315]= -2147265689;
assign addr[19316]= -2147470025;
assign addr[19317]= -2146993250;
assign addr[19318]= -2145835515;
assign addr[19319]= -2143997187;
assign addr[19320]= -2141478848;
assign addr[19321]= -2138281298;
assign addr[19322]= -2134405552;
assign addr[19323]= -2129852837;
assign addr[19324]= -2124624598;
assign addr[19325]= -2118722494;
assign addr[19326]= -2112148396;
assign addr[19327]= -2104904390;
assign addr[19328]= -2096992772;
assign addr[19329]= -2088416053;
assign addr[19330]= -2079176953;
assign addr[19331]= -2069278401;
assign addr[19332]= -2058723538;
assign addr[19333]= -2047515711;
assign addr[19334]= -2035658475;
assign addr[19335]= -2023155591;
assign addr[19336]= -2010011024;
assign addr[19337]= -1996228943;
assign addr[19338]= -1981813720;
assign addr[19339]= -1966769926;
assign addr[19340]= -1951102334;
assign addr[19341]= -1934815911;
assign addr[19342]= -1917915825;
assign addr[19343]= -1900407434;
assign addr[19344]= -1882296293;
assign addr[19345]= -1863588145;
assign addr[19346]= -1844288924;
assign addr[19347]= -1824404752;
assign addr[19348]= -1803941934;
assign addr[19349]= -1782906961;
assign addr[19350]= -1761306505;
assign addr[19351]= -1739147417;
assign addr[19352]= -1716436725;
assign addr[19353]= -1693181631;
assign addr[19354]= -1669389513;
assign addr[19355]= -1645067915;
assign addr[19356]= -1620224553;
assign addr[19357]= -1594867305;
assign addr[19358]= -1569004214;
assign addr[19359]= -1542643483;
assign addr[19360]= -1515793473;
assign addr[19361]= -1488462700;
assign addr[19362]= -1460659832;
assign addr[19363]= -1432393688;
assign addr[19364]= -1403673233;
assign addr[19365]= -1374507575;
assign addr[19366]= -1344905966;
assign addr[19367]= -1314877795;
assign addr[19368]= -1284432584;
assign addr[19369]= -1253579991;
assign addr[19370]= -1222329801;
assign addr[19371]= -1190691925;
assign addr[19372]= -1158676398;
assign addr[19373]= -1126293375;
assign addr[19374]= -1093553126;
assign addr[19375]= -1060466036;
assign addr[19376]= -1027042599;
assign addr[19377]= -993293415;
assign addr[19378]= -959229189;
assign addr[19379]= -924860725;
assign addr[19380]= -890198924;
assign addr[19381]= -855254778;
assign addr[19382]= -820039373;
assign addr[19383]= -784563876;
assign addr[19384]= -748839539;
assign addr[19385]= -712877694;
assign addr[19386]= -676689746;
assign addr[19387]= -640287172;
assign addr[19388]= -603681519;
assign addr[19389]= -566884397;
assign addr[19390]= -529907477;
assign addr[19391]= -492762486;
assign addr[19392]= -455461206;
assign addr[19393]= -418015468;
assign addr[19394]= -380437148;
assign addr[19395]= -342738165;
assign addr[19396]= -304930476;
assign addr[19397]= -267026072;
assign addr[19398]= -229036977;
assign addr[19399]= -190975237;
assign addr[19400]= -152852926;
assign addr[19401]= -114682135;
assign addr[19402]= -76474970;
assign addr[19403]= -38243550;
assign addr[19404]= 0;
assign addr[19405]= 38243550;
assign addr[19406]= 76474970;
assign addr[19407]= 114682135;
assign addr[19408]= 152852926;
assign addr[19409]= 190975237;
assign addr[19410]= 229036977;
assign addr[19411]= 267026072;
assign addr[19412]= 304930476;
assign addr[19413]= 342738165;
assign addr[19414]= 380437148;
assign addr[19415]= 418015468;
assign addr[19416]= 455461206;
assign addr[19417]= 492762486;
assign addr[19418]= 529907477;
assign addr[19419]= 566884397;
assign addr[19420]= 603681519;
assign addr[19421]= 640287172;
assign addr[19422]= 676689746;
assign addr[19423]= 712877694;
assign addr[19424]= 748839539;
assign addr[19425]= 784563876;
assign addr[19426]= 820039373;
assign addr[19427]= 855254778;
assign addr[19428]= 890198924;
assign addr[19429]= 924860725;
assign addr[19430]= 959229189;
assign addr[19431]= 993293415;
assign addr[19432]= 1027042599;
assign addr[19433]= 1060466036;
assign addr[19434]= 1093553126;
assign addr[19435]= 1126293375;
assign addr[19436]= 1158676398;
assign addr[19437]= 1190691925;
assign addr[19438]= 1222329801;
assign addr[19439]= 1253579991;
assign addr[19440]= 1284432584;
assign addr[19441]= 1314877795;
assign addr[19442]= 1344905966;
assign addr[19443]= 1374507575;
assign addr[19444]= 1403673233;
assign addr[19445]= 1432393688;
assign addr[19446]= 1460659832;
assign addr[19447]= 1488462700;
assign addr[19448]= 1515793473;
assign addr[19449]= 1542643483;
assign addr[19450]= 1569004214;
assign addr[19451]= 1594867305;
assign addr[19452]= 1620224553;
assign addr[19453]= 1645067915;
assign addr[19454]= 1669389513;
assign addr[19455]= 1693181631;
assign addr[19456]= 1716436725;
assign addr[19457]= 1739147417;
assign addr[19458]= 1761306505;
assign addr[19459]= 1782906961;
assign addr[19460]= 1803941934;
assign addr[19461]= 1824404752;
assign addr[19462]= 1844288924;
assign addr[19463]= 1863588145;
assign addr[19464]= 1882296293;
assign addr[19465]= 1900407434;
assign addr[19466]= 1917915825;
assign addr[19467]= 1934815911;
assign addr[19468]= 1951102334;
assign addr[19469]= 1966769926;
assign addr[19470]= 1981813720;
assign addr[19471]= 1996228943;
assign addr[19472]= 2010011024;
assign addr[19473]= 2023155591;
assign addr[19474]= 2035658475;
assign addr[19475]= 2047515711;
assign addr[19476]= 2058723538;
assign addr[19477]= 2069278401;
assign addr[19478]= 2079176953;
assign addr[19479]= 2088416053;
assign addr[19480]= 2096992772;
assign addr[19481]= 2104904390;
assign addr[19482]= 2112148396;
assign addr[19483]= 2118722494;
assign addr[19484]= 2124624598;
assign addr[19485]= 2129852837;
assign addr[19486]= 2134405552;
assign addr[19487]= 2138281298;
assign addr[19488]= 2141478848;
assign addr[19489]= 2143997187;
assign addr[19490]= 2145835515;
assign addr[19491]= 2146993250;
assign addr[19492]= 2147470025;
assign addr[19493]= 2147265689;
assign addr[19494]= 2146380306;
assign addr[19495]= 2144814157;
assign addr[19496]= 2142567738;
assign addr[19497]= 2139641764;
assign addr[19498]= 2136037160;
assign addr[19499]= 2131755071;
assign addr[19500]= 2126796855;
assign addr[19501]= 2121164085;
assign addr[19502]= 2114858546;
assign addr[19503]= 2107882239;
assign addr[19504]= 2100237377;
assign addr[19505]= 2091926384;
assign addr[19506]= 2082951896;
assign addr[19507]= 2073316760;
assign addr[19508]= 2063024031;
assign addr[19509]= 2052076975;
assign addr[19510]= 2040479063;
assign addr[19511]= 2028233973;
assign addr[19512]= 2015345591;
assign addr[19513]= 2001818002;
assign addr[19514]= 1987655498;
assign addr[19515]= 1972862571;
assign addr[19516]= 1957443913;
assign addr[19517]= 1941404413;
assign addr[19518]= 1924749160;
assign addr[19519]= 1907483436;
assign addr[19520]= 1889612716;
assign addr[19521]= 1871142669;
assign addr[19522]= 1852079154;
assign addr[19523]= 1832428215;
assign addr[19524]= 1812196087;
assign addr[19525]= 1791389186;
assign addr[19526]= 1770014111;
assign addr[19527]= 1748077642;
assign addr[19528]= 1725586737;
assign addr[19529]= 1702548529;
assign addr[19530]= 1678970324;
assign addr[19531]= 1654859602;
assign addr[19532]= 1630224009;
assign addr[19533]= 1605071359;
assign addr[19534]= 1579409630;
assign addr[19535]= 1553246960;
assign addr[19536]= 1526591649;
assign addr[19537]= 1499452149;
assign addr[19538]= 1471837070;
assign addr[19539]= 1443755168;
assign addr[19540]= 1415215352;
assign addr[19541]= 1386226674;
assign addr[19542]= 1356798326;
assign addr[19543]= 1326939644;
assign addr[19544]= 1296660098;
assign addr[19545]= 1265969291;
assign addr[19546]= 1234876957;
assign addr[19547]= 1203392958;
assign addr[19548]= 1171527280;
assign addr[19549]= 1139290029;
assign addr[19550]= 1106691431;
assign addr[19551]= 1073741824;
assign addr[19552]= 1040451659;
assign addr[19553]= 1006831495;
assign addr[19554]= 972891995;
assign addr[19555]= 938643924;
assign addr[19556]= 904098143;
assign addr[19557]= 869265610;
assign addr[19558]= 834157373;
assign addr[19559]= 798784567;
assign addr[19560]= 763158411;
assign addr[19561]= 727290205;
assign addr[19562]= 691191324;
assign addr[19563]= 654873219;
assign addr[19564]= 618347408;
assign addr[19565]= 581625477;
assign addr[19566]= 544719071;
assign addr[19567]= 507639898;
assign addr[19568]= 470399716;
assign addr[19569]= 433010339;
assign addr[19570]= 395483624;
assign addr[19571]= 357831473;
assign addr[19572]= 320065829;
assign addr[19573]= 282198671;
assign addr[19574]= 244242007;
assign addr[19575]= 206207878;
assign addr[19576]= 168108346;
assign addr[19577]= 129955495;
assign addr[19578]= 91761426;
assign addr[19579]= 53538253;
assign addr[19580]= 15298099;
assign addr[19581]= -22946906;
assign addr[19582]= -61184634;
assign addr[19583]= -99402956;
assign addr[19584]= -137589750;
assign addr[19585]= -175732905;
assign addr[19586]= -213820322;
assign addr[19587]= -251839923;
assign addr[19588]= -289779648;
assign addr[19589]= -327627463;
assign addr[19590]= -365371365;
assign addr[19591]= -402999383;
assign addr[19592]= -440499581;
assign addr[19593]= -477860067;
assign addr[19594]= -515068990;
assign addr[19595]= -552114549;
assign addr[19596]= -588984994;
assign addr[19597]= -625668632;
assign addr[19598]= -662153826;
assign addr[19599]= -698429006;
assign addr[19600]= -734482665;
assign addr[19601]= -770303369;
assign addr[19602]= -805879757;
assign addr[19603]= -841200544;
assign addr[19604]= -876254528;
assign addr[19605]= -911030591;
assign addr[19606]= -945517704;
assign addr[19607]= -979704927;
assign addr[19608]= -1013581418;
assign addr[19609]= -1047136432;
assign addr[19610]= -1080359326;
assign addr[19611]= -1113239564;
assign addr[19612]= -1145766716;
assign addr[19613]= -1177930466;
assign addr[19614]= -1209720613;
assign addr[19615]= -1241127074;
assign addr[19616]= -1272139887;
assign addr[19617]= -1302749217;
assign addr[19618]= -1332945355;
assign addr[19619]= -1362718723;
assign addr[19620]= -1392059879;
assign addr[19621]= -1420959516;
assign addr[19622]= -1449408469;
assign addr[19623]= -1477397714;
assign addr[19624]= -1504918373;
assign addr[19625]= -1531961719;
assign addr[19626]= -1558519173;
assign addr[19627]= -1584582314;
assign addr[19628]= -1610142873;
assign addr[19629]= -1635192744;
assign addr[19630]= -1659723983;
assign addr[19631]= -1683728808;
assign addr[19632]= -1707199606;
assign addr[19633]= -1730128933;
assign addr[19634]= -1752509516;
assign addr[19635]= -1774334257;
assign addr[19636]= -1795596234;
assign addr[19637]= -1816288703;
assign addr[19638]= -1836405100;
assign addr[19639]= -1855939047;
assign addr[19640]= -1874884346;
assign addr[19641]= -1893234990;
assign addr[19642]= -1910985158;
assign addr[19643]= -1928129220;
assign addr[19644]= -1944661739;
assign addr[19645]= -1960577471;
assign addr[19646]= -1975871368;
assign addr[19647]= -1990538579;
assign addr[19648]= -2004574453;
assign addr[19649]= -2017974537;
assign addr[19650]= -2030734582;
assign addr[19651]= -2042850540;
assign addr[19652]= -2054318569;
assign addr[19653]= -2065135031;
assign addr[19654]= -2075296495;
assign addr[19655]= -2084799740;
assign addr[19656]= -2093641749;
assign addr[19657]= -2101819720;
assign addr[19658]= -2109331059;
assign addr[19659]= -2116173382;
assign addr[19660]= -2122344521;
assign addr[19661]= -2127842516;
assign addr[19662]= -2132665626;
assign addr[19663]= -2136812319;
assign addr[19664]= -2140281282;
assign addr[19665]= -2143071413;
assign addr[19666]= -2145181827;
assign addr[19667]= -2146611856;
assign addr[19668]= -2147361045;
assign addr[19669]= -2147429158;
assign addr[19670]= -2146816171;
assign addr[19671]= -2145522281;
assign addr[19672]= -2143547897;
assign addr[19673]= -2140893646;
assign addr[19674]= -2137560369;
assign addr[19675]= -2133549123;
assign addr[19676]= -2128861181;
assign addr[19677]= -2123498030;
assign addr[19678]= -2117461370;
assign addr[19679]= -2110753117;
assign addr[19680]= -2103375398;
assign addr[19681]= -2095330553;
assign addr[19682]= -2086621133;
assign addr[19683]= -2077249901;
assign addr[19684]= -2067219829;
assign addr[19685]= -2056534099;
assign addr[19686]= -2045196100;
assign addr[19687]= -2033209426;
assign addr[19688]= -2020577882;
assign addr[19689]= -2007305472;
assign addr[19690]= -1993396407;
assign addr[19691]= -1978855097;
assign addr[19692]= -1963686155;
assign addr[19693]= -1947894393;
assign addr[19694]= -1931484818;
assign addr[19695]= -1914462636;
assign addr[19696]= -1896833245;
assign addr[19697]= -1878602237;
assign addr[19698]= -1859775393;
assign addr[19699]= -1840358687;
assign addr[19700]= -1820358275;
assign addr[19701]= -1799780501;
assign addr[19702]= -1778631892;
assign addr[19703]= -1756919156;
assign addr[19704]= -1734649179;
assign addr[19705]= -1711829025;
assign addr[19706]= -1688465931;
assign addr[19707]= -1664567307;
assign addr[19708]= -1640140734;
assign addr[19709]= -1615193959;
assign addr[19710]= -1589734894;
assign addr[19711]= -1563771613;
assign addr[19712]= -1537312353;
assign addr[19713]= -1510365504;
assign addr[19714]= -1482939614;
assign addr[19715]= -1455043381;
assign addr[19716]= -1426685652;
assign addr[19717]= -1397875423;
assign addr[19718]= -1368621831;
assign addr[19719]= -1338934154;
assign addr[19720]= -1308821808;
assign addr[19721]= -1278294345;
assign addr[19722]= -1247361445;
assign addr[19723]= -1216032921;
assign addr[19724]= -1184318708;
assign addr[19725]= -1152228866;
assign addr[19726]= -1119773573;
assign addr[19727]= -1086963121;
assign addr[19728]= -1053807919;
assign addr[19729]= -1020318481;
assign addr[19730]= -986505429;
assign addr[19731]= -952379488;
assign addr[19732]= -917951481;
assign addr[19733]= -883232329;
assign addr[19734]= -848233042;
assign addr[19735]= -812964722;
assign addr[19736]= -777438554;
assign addr[19737]= -741665807;
assign addr[19738]= -705657826;
assign addr[19739]= -669426032;
assign addr[19740]= -632981917;
assign addr[19741]= -596337040;
assign addr[19742]= -559503022;
assign addr[19743]= -522491548;
assign addr[19744]= -485314355;
assign addr[19745]= -447983235;
assign addr[19746]= -410510029;
assign addr[19747]= -372906622;
assign addr[19748]= -335184940;
assign addr[19749]= -297356948;
assign addr[19750]= -259434643;
assign addr[19751]= -221430054;
assign addr[19752]= -183355234;
assign addr[19753]= -145222259;
assign addr[19754]= -107043224;
assign addr[19755]= -68830239;
assign addr[19756]= -30595422;
assign addr[19757]= 7649098;
assign addr[19758]= 45891193;
assign addr[19759]= 84118732;
assign addr[19760]= 122319591;
assign addr[19761]= 160481654;
assign addr[19762]= 198592817;
assign addr[19763]= 236640993;
assign addr[19764]= 274614114;
assign addr[19765]= 312500135;
assign addr[19766]= 350287041;
assign addr[19767]= 387962847;
assign addr[19768]= 425515602;
assign addr[19769]= 462933398;
assign addr[19770]= 500204365;
assign addr[19771]= 537316682;
assign addr[19772]= 574258580;
assign addr[19773]= 611018340;
assign addr[19774]= 647584304;
assign addr[19775]= 683944874;
assign addr[19776]= 720088517;
assign addr[19777]= 756003771;
assign addr[19778]= 791679244;
assign addr[19779]= 827103620;
assign addr[19780]= 862265664;
assign addr[19781]= 897154224;
assign addr[19782]= 931758235;
assign addr[19783]= 966066720;
assign addr[19784]= 1000068799;
assign addr[19785]= 1033753687;
assign addr[19786]= 1067110699;
assign addr[19787]= 1100129257;
assign addr[19788]= 1132798888;
assign addr[19789]= 1165109230;
assign addr[19790]= 1197050035;
assign addr[19791]= 1228611172;
assign addr[19792]= 1259782632;
assign addr[19793]= 1290554528;
assign addr[19794]= 1320917099;
assign addr[19795]= 1350860716;
assign addr[19796]= 1380375881;
assign addr[19797]= 1409453233;
assign addr[19798]= 1438083551;
assign addr[19799]= 1466257752;
assign addr[19800]= 1493966902;
assign addr[19801]= 1521202211;
assign addr[19802]= 1547955041;
assign addr[19803]= 1574216908;
assign addr[19804]= 1599979481;
assign addr[19805]= 1625234591;
assign addr[19806]= 1649974225;
assign addr[19807]= 1674190539;
assign addr[19808]= 1697875851;
assign addr[19809]= 1721022648;
assign addr[19810]= 1743623590;
assign addr[19811]= 1765671509;
assign addr[19812]= 1787159411;
assign addr[19813]= 1808080480;
assign addr[19814]= 1828428082;
assign addr[19815]= 1848195763;
assign addr[19816]= 1867377253;
assign addr[19817]= 1885966468;
assign addr[19818]= 1903957513;
assign addr[19819]= 1921344681;
assign addr[19820]= 1938122457;
assign addr[19821]= 1954285520;
assign addr[19822]= 1969828744;
assign addr[19823]= 1984747199;
assign addr[19824]= 1999036154;
assign addr[19825]= 2012691075;
assign addr[19826]= 2025707632;
assign addr[19827]= 2038081698;
assign addr[19828]= 2049809346;
assign addr[19829]= 2060886858;
assign addr[19830]= 2071310720;
assign addr[19831]= 2081077626;
assign addr[19832]= 2090184478;
assign addr[19833]= 2098628387;
assign addr[19834]= 2106406677;
assign addr[19835]= 2113516878;
assign addr[19836]= 2119956737;
assign addr[19837]= 2125724211;
assign addr[19838]= 2130817471;
assign addr[19839]= 2135234901;
assign addr[19840]= 2138975100;
assign addr[19841]= 2142036881;
assign addr[19842]= 2144419275;
assign addr[19843]= 2146121524;
assign addr[19844]= 2147143090;
assign addr[19845]= 2147483648;
assign addr[19846]= 2147143090;
assign addr[19847]= 2146121524;
assign addr[19848]= 2144419275;
assign addr[19849]= 2142036881;
assign addr[19850]= 2138975100;
assign addr[19851]= 2135234901;
assign addr[19852]= 2130817471;
assign addr[19853]= 2125724211;
assign addr[19854]= 2119956737;
assign addr[19855]= 2113516878;
assign addr[19856]= 2106406677;
assign addr[19857]= 2098628387;
assign addr[19858]= 2090184478;
assign addr[19859]= 2081077626;
assign addr[19860]= 2071310720;
assign addr[19861]= 2060886858;
assign addr[19862]= 2049809346;
assign addr[19863]= 2038081698;
assign addr[19864]= 2025707632;
assign addr[19865]= 2012691075;
assign addr[19866]= 1999036154;
assign addr[19867]= 1984747199;
assign addr[19868]= 1969828744;
assign addr[19869]= 1954285520;
assign addr[19870]= 1938122457;
assign addr[19871]= 1921344681;
assign addr[19872]= 1903957513;
assign addr[19873]= 1885966468;
assign addr[19874]= 1867377253;
assign addr[19875]= 1848195763;
assign addr[19876]= 1828428082;
assign addr[19877]= 1808080480;
assign addr[19878]= 1787159411;
assign addr[19879]= 1765671509;
assign addr[19880]= 1743623590;
assign addr[19881]= 1721022648;
assign addr[19882]= 1697875851;
assign addr[19883]= 1674190539;
assign addr[19884]= 1649974225;
assign addr[19885]= 1625234591;
assign addr[19886]= 1599979481;
assign addr[19887]= 1574216908;
assign addr[19888]= 1547955041;
assign addr[19889]= 1521202211;
assign addr[19890]= 1493966902;
assign addr[19891]= 1466257752;
assign addr[19892]= 1438083551;
assign addr[19893]= 1409453233;
assign addr[19894]= 1380375881;
assign addr[19895]= 1350860716;
assign addr[19896]= 1320917099;
assign addr[19897]= 1290554528;
assign addr[19898]= 1259782632;
assign addr[19899]= 1228611172;
assign addr[19900]= 1197050035;
assign addr[19901]= 1165109230;
assign addr[19902]= 1132798888;
assign addr[19903]= 1100129257;
assign addr[19904]= 1067110699;
assign addr[19905]= 1033753687;
assign addr[19906]= 1000068799;
assign addr[19907]= 966066720;
assign addr[19908]= 931758235;
assign addr[19909]= 897154224;
assign addr[19910]= 862265664;
assign addr[19911]= 827103620;
assign addr[19912]= 791679244;
assign addr[19913]= 756003771;
assign addr[19914]= 720088517;
assign addr[19915]= 683944874;
assign addr[19916]= 647584304;
assign addr[19917]= 611018340;
assign addr[19918]= 574258580;
assign addr[19919]= 537316682;
assign addr[19920]= 500204365;
assign addr[19921]= 462933398;
assign addr[19922]= 425515602;
assign addr[19923]= 387962847;
assign addr[19924]= 350287041;
assign addr[19925]= 312500135;
assign addr[19926]= 274614114;
assign addr[19927]= 236640993;
assign addr[19928]= 198592817;
assign addr[19929]= 160481654;
assign addr[19930]= 122319591;
assign addr[19931]= 84118732;
assign addr[19932]= 45891193;
assign addr[19933]= 7649098;
assign addr[19934]= -30595422;
assign addr[19935]= -68830239;
assign addr[19936]= -107043224;
assign addr[19937]= -145222259;
assign addr[19938]= -183355234;
assign addr[19939]= -221430054;
assign addr[19940]= -259434643;
assign addr[19941]= -297356948;
assign addr[19942]= -335184940;
assign addr[19943]= -372906622;
assign addr[19944]= -410510029;
assign addr[19945]= -447983235;
assign addr[19946]= -485314355;
assign addr[19947]= -522491548;
assign addr[19948]= -559503022;
assign addr[19949]= -596337040;
assign addr[19950]= -632981917;
assign addr[19951]= -669426032;
assign addr[19952]= -705657826;
assign addr[19953]= -741665807;
assign addr[19954]= -777438554;
assign addr[19955]= -812964722;
assign addr[19956]= -848233042;
assign addr[19957]= -883232329;
assign addr[19958]= -917951481;
assign addr[19959]= -952379488;
assign addr[19960]= -986505429;
assign addr[19961]= -1020318481;
assign addr[19962]= -1053807919;
assign addr[19963]= -1086963121;
assign addr[19964]= -1119773573;
assign addr[19965]= -1152228866;
assign addr[19966]= -1184318708;
assign addr[19967]= -1216032921;
assign addr[19968]= -1247361445;
assign addr[19969]= -1278294345;
assign addr[19970]= -1308821808;
assign addr[19971]= -1338934154;
assign addr[19972]= -1368621831;
assign addr[19973]= -1397875423;
assign addr[19974]= -1426685652;
assign addr[19975]= -1455043381;
assign addr[19976]= -1482939614;
assign addr[19977]= -1510365504;
assign addr[19978]= -1537312353;
assign addr[19979]= -1563771613;
assign addr[19980]= -1589734894;
assign addr[19981]= -1615193959;
assign addr[19982]= -1640140734;
assign addr[19983]= -1664567307;
assign addr[19984]= -1688465931;
assign addr[19985]= -1711829025;
assign addr[19986]= -1734649179;
assign addr[19987]= -1756919156;
assign addr[19988]= -1778631892;
assign addr[19989]= -1799780501;
assign addr[19990]= -1820358275;
assign addr[19991]= -1840358687;
assign addr[19992]= -1859775393;
assign addr[19993]= -1878602237;
assign addr[19994]= -1896833245;
assign addr[19995]= -1914462636;
assign addr[19996]= -1931484818;
assign addr[19997]= -1947894393;
assign addr[19998]= -1963686155;
assign addr[19999]= -1978855097;
assign addr[20000]= -1993396407;
assign addr[20001]= -2007305472;
assign addr[20002]= -2020577882;
assign addr[20003]= -2033209426;
assign addr[20004]= -2045196100;
assign addr[20005]= -2056534099;
assign addr[20006]= -2067219829;
assign addr[20007]= -2077249901;
assign addr[20008]= -2086621133;
assign addr[20009]= -2095330553;
assign addr[20010]= -2103375398;
assign addr[20011]= -2110753117;
assign addr[20012]= -2117461370;
assign addr[20013]= -2123498030;
assign addr[20014]= -2128861181;
assign addr[20015]= -2133549123;
assign addr[20016]= -2137560369;
assign addr[20017]= -2140893646;
assign addr[20018]= -2143547897;
assign addr[20019]= -2145522281;
assign addr[20020]= -2146816171;
assign addr[20021]= -2147429158;
assign addr[20022]= -2147361045;
assign addr[20023]= -2146611856;
assign addr[20024]= -2145181827;
assign addr[20025]= -2143071413;
assign addr[20026]= -2140281282;
assign addr[20027]= -2136812319;
assign addr[20028]= -2132665626;
assign addr[20029]= -2127842516;
assign addr[20030]= -2122344521;
assign addr[20031]= -2116173382;
assign addr[20032]= -2109331059;
assign addr[20033]= -2101819720;
assign addr[20034]= -2093641749;
assign addr[20035]= -2084799740;
assign addr[20036]= -2075296495;
assign addr[20037]= -2065135031;
assign addr[20038]= -2054318569;
assign addr[20039]= -2042850540;
assign addr[20040]= -2030734582;
assign addr[20041]= -2017974537;
assign addr[20042]= -2004574453;
assign addr[20043]= -1990538579;
assign addr[20044]= -1975871368;
assign addr[20045]= -1960577471;
assign addr[20046]= -1944661739;
assign addr[20047]= -1928129220;
assign addr[20048]= -1910985158;
assign addr[20049]= -1893234990;
assign addr[20050]= -1874884346;
assign addr[20051]= -1855939047;
assign addr[20052]= -1836405100;
assign addr[20053]= -1816288703;
assign addr[20054]= -1795596234;
assign addr[20055]= -1774334257;
assign addr[20056]= -1752509516;
assign addr[20057]= -1730128933;
assign addr[20058]= -1707199606;
assign addr[20059]= -1683728808;
assign addr[20060]= -1659723983;
assign addr[20061]= -1635192744;
assign addr[20062]= -1610142873;
assign addr[20063]= -1584582314;
assign addr[20064]= -1558519173;
assign addr[20065]= -1531961719;
assign addr[20066]= -1504918373;
assign addr[20067]= -1477397714;
assign addr[20068]= -1449408469;
assign addr[20069]= -1420959516;
assign addr[20070]= -1392059879;
assign addr[20071]= -1362718723;
assign addr[20072]= -1332945355;
assign addr[20073]= -1302749217;
assign addr[20074]= -1272139887;
assign addr[20075]= -1241127074;
assign addr[20076]= -1209720613;
assign addr[20077]= -1177930466;
assign addr[20078]= -1145766716;
assign addr[20079]= -1113239564;
assign addr[20080]= -1080359326;
assign addr[20081]= -1047136432;
assign addr[20082]= -1013581418;
assign addr[20083]= -979704927;
assign addr[20084]= -945517704;
assign addr[20085]= -911030591;
assign addr[20086]= -876254528;
assign addr[20087]= -841200544;
assign addr[20088]= -805879757;
assign addr[20089]= -770303369;
assign addr[20090]= -734482665;
assign addr[20091]= -698429006;
assign addr[20092]= -662153826;
assign addr[20093]= -625668632;
assign addr[20094]= -588984994;
assign addr[20095]= -552114549;
assign addr[20096]= -515068990;
assign addr[20097]= -477860067;
assign addr[20098]= -440499581;
assign addr[20099]= -402999383;
assign addr[20100]= -365371365;
assign addr[20101]= -327627463;
assign addr[20102]= -289779648;
assign addr[20103]= -251839923;
assign addr[20104]= -213820322;
assign addr[20105]= -175732905;
assign addr[20106]= -137589750;
assign addr[20107]= -99402956;
assign addr[20108]= -61184634;
assign addr[20109]= -22946906;
assign addr[20110]= 15298099;
assign addr[20111]= 53538253;
assign addr[20112]= 91761426;
assign addr[20113]= 129955495;
assign addr[20114]= 168108346;
assign addr[20115]= 206207878;
assign addr[20116]= 244242007;
assign addr[20117]= 282198671;
assign addr[20118]= 320065829;
assign addr[20119]= 357831473;
assign addr[20120]= 395483624;
assign addr[20121]= 433010339;
assign addr[20122]= 470399716;
assign addr[20123]= 507639898;
assign addr[20124]= 544719071;
assign addr[20125]= 581625477;
assign addr[20126]= 618347408;
assign addr[20127]= 654873219;
assign addr[20128]= 691191324;
assign addr[20129]= 727290205;
assign addr[20130]= 763158411;
assign addr[20131]= 798784567;
assign addr[20132]= 834157373;
assign addr[20133]= 869265610;
assign addr[20134]= 904098143;
assign addr[20135]= 938643924;
assign addr[20136]= 972891995;
assign addr[20137]= 1006831495;
assign addr[20138]= 1040451659;
assign addr[20139]= 1073741824;
assign addr[20140]= 1106691431;
assign addr[20141]= 1139290029;
assign addr[20142]= 1171527280;
assign addr[20143]= 1203392958;
assign addr[20144]= 1234876957;
assign addr[20145]= 1265969291;
assign addr[20146]= 1296660098;
assign addr[20147]= 1326939644;
assign addr[20148]= 1356798326;
assign addr[20149]= 1386226674;
assign addr[20150]= 1415215352;
assign addr[20151]= 1443755168;
assign addr[20152]= 1471837070;
assign addr[20153]= 1499452149;
assign addr[20154]= 1526591649;
assign addr[20155]= 1553246960;
assign addr[20156]= 1579409630;
assign addr[20157]= 1605071359;
assign addr[20158]= 1630224009;
assign addr[20159]= 1654859602;
assign addr[20160]= 1678970324;
assign addr[20161]= 1702548529;
assign addr[20162]= 1725586737;
assign addr[20163]= 1748077642;
assign addr[20164]= 1770014111;
assign addr[20165]= 1791389186;
assign addr[20166]= 1812196087;
assign addr[20167]= 1832428215;
assign addr[20168]= 1852079154;
assign addr[20169]= 1871142669;
assign addr[20170]= 1889612716;
assign addr[20171]= 1907483436;
assign addr[20172]= 1924749160;
assign addr[20173]= 1941404413;
assign addr[20174]= 1957443913;
assign addr[20175]= 1972862571;
assign addr[20176]= 1987655498;
assign addr[20177]= 2001818002;
assign addr[20178]= 2015345591;
assign addr[20179]= 2028233973;
assign addr[20180]= 2040479063;
assign addr[20181]= 2052076975;
assign addr[20182]= 2063024031;
assign addr[20183]= 2073316760;
assign addr[20184]= 2082951896;
assign addr[20185]= 2091926384;
assign addr[20186]= 2100237377;
assign addr[20187]= 2107882239;
assign addr[20188]= 2114858546;
assign addr[20189]= 2121164085;
assign addr[20190]= 2126796855;
assign addr[20191]= 2131755071;
assign addr[20192]= 2136037160;
assign addr[20193]= 2139641764;
assign addr[20194]= 2142567738;
assign addr[20195]= 2144814157;
assign addr[20196]= 2146380306;
assign addr[20197]= 2147265689;
assign addr[20198]= 2147470025;
assign addr[20199]= 2146993250;
assign addr[20200]= 2145835515;
assign addr[20201]= 2143997187;
assign addr[20202]= 2141478848;
assign addr[20203]= 2138281298;
assign addr[20204]= 2134405552;
assign addr[20205]= 2129852837;
assign addr[20206]= 2124624598;
assign addr[20207]= 2118722494;
assign addr[20208]= 2112148396;
assign addr[20209]= 2104904390;
assign addr[20210]= 2096992772;
assign addr[20211]= 2088416053;
assign addr[20212]= 2079176953;
assign addr[20213]= 2069278401;
assign addr[20214]= 2058723538;
assign addr[20215]= 2047515711;
assign addr[20216]= 2035658475;
assign addr[20217]= 2023155591;
assign addr[20218]= 2010011024;
assign addr[20219]= 1996228943;
assign addr[20220]= 1981813720;
assign addr[20221]= 1966769926;
assign addr[20222]= 1951102334;
assign addr[20223]= 1934815911;
assign addr[20224]= 1917915825;
assign addr[20225]= 1900407434;
assign addr[20226]= 1882296293;
assign addr[20227]= 1863588145;
assign addr[20228]= 1844288924;
assign addr[20229]= 1824404752;
assign addr[20230]= 1803941934;
assign addr[20231]= 1782906961;
assign addr[20232]= 1761306505;
assign addr[20233]= 1739147417;
assign addr[20234]= 1716436725;
assign addr[20235]= 1693181631;
assign addr[20236]= 1669389513;
assign addr[20237]= 1645067915;
assign addr[20238]= 1620224553;
assign addr[20239]= 1594867305;
assign addr[20240]= 1569004214;
assign addr[20241]= 1542643483;
assign addr[20242]= 1515793473;
assign addr[20243]= 1488462700;
assign addr[20244]= 1460659832;
assign addr[20245]= 1432393688;
assign addr[20246]= 1403673233;
assign addr[20247]= 1374507575;
assign addr[20248]= 1344905966;
assign addr[20249]= 1314877795;
assign addr[20250]= 1284432584;
assign addr[20251]= 1253579991;
assign addr[20252]= 1222329801;
assign addr[20253]= 1190691925;
assign addr[20254]= 1158676398;
assign addr[20255]= 1126293375;
assign addr[20256]= 1093553126;
assign addr[20257]= 1060466036;
assign addr[20258]= 1027042599;
assign addr[20259]= 993293415;
assign addr[20260]= 959229189;
assign addr[20261]= 924860725;
assign addr[20262]= 890198924;
assign addr[20263]= 855254778;
assign addr[20264]= 820039373;
assign addr[20265]= 784563876;
assign addr[20266]= 748839539;
assign addr[20267]= 712877694;
assign addr[20268]= 676689746;
assign addr[20269]= 640287172;
assign addr[20270]= 603681519;
assign addr[20271]= 566884397;
assign addr[20272]= 529907477;
assign addr[20273]= 492762486;
assign addr[20274]= 455461206;
assign addr[20275]= 418015468;
assign addr[20276]= 380437148;
assign addr[20277]= 342738165;
assign addr[20278]= 304930476;
assign addr[20279]= 267026072;
assign addr[20280]= 229036977;
assign addr[20281]= 190975237;
assign addr[20282]= 152852926;
assign addr[20283]= 114682135;
assign addr[20284]= 76474970;
assign addr[20285]= 38243550;
assign addr[20286]= 0;
assign addr[20287]= -38243550;
assign addr[20288]= -76474970;
assign addr[20289]= -114682135;
assign addr[20290]= -152852926;
assign addr[20291]= -190975237;
assign addr[20292]= -229036977;
assign addr[20293]= -267026072;
assign addr[20294]= -304930476;
assign addr[20295]= -342738165;
assign addr[20296]= -380437148;
assign addr[20297]= -418015468;
assign addr[20298]= -455461206;
assign addr[20299]= -492762486;
assign addr[20300]= -529907477;
assign addr[20301]= -566884397;
assign addr[20302]= -603681519;
assign addr[20303]= -640287172;
assign addr[20304]= -676689746;
assign addr[20305]= -712877694;
assign addr[20306]= -748839539;
assign addr[20307]= -784563876;
assign addr[20308]= -820039373;
assign addr[20309]= -855254778;
assign addr[20310]= -890198924;
assign addr[20311]= -924860725;
assign addr[20312]= -959229189;
assign addr[20313]= -993293415;
assign addr[20314]= -1027042599;
assign addr[20315]= -1060466036;
assign addr[20316]= -1093553126;
assign addr[20317]= -1126293375;
assign addr[20318]= -1158676398;
assign addr[20319]= -1190691925;
assign addr[20320]= -1222329801;
assign addr[20321]= -1253579991;
assign addr[20322]= -1284432584;
assign addr[20323]= -1314877795;
assign addr[20324]= -1344905966;
assign addr[20325]= -1374507575;
assign addr[20326]= -1403673233;
assign addr[20327]= -1432393688;
assign addr[20328]= -1460659832;
assign addr[20329]= -1488462700;
assign addr[20330]= -1515793473;
assign addr[20331]= -1542643483;
assign addr[20332]= -1569004214;
assign addr[20333]= -1594867305;
assign addr[20334]= -1620224553;
assign addr[20335]= -1645067915;
assign addr[20336]= -1669389513;
assign addr[20337]= -1693181631;
assign addr[20338]= -1716436725;
assign addr[20339]= -1739147417;
assign addr[20340]= -1761306505;
assign addr[20341]= -1782906961;
assign addr[20342]= -1803941934;
assign addr[20343]= -1824404752;
assign addr[20344]= -1844288924;
assign addr[20345]= -1863588145;
assign addr[20346]= -1882296293;
assign addr[20347]= -1900407434;
assign addr[20348]= -1917915825;
assign addr[20349]= -1934815911;
assign addr[20350]= -1951102334;
assign addr[20351]= -1966769926;
assign addr[20352]= -1981813720;
assign addr[20353]= -1996228943;
assign addr[20354]= -2010011024;
assign addr[20355]= -2023155591;
assign addr[20356]= -2035658475;
assign addr[20357]= -2047515711;
assign addr[20358]= -2058723538;
assign addr[20359]= -2069278401;
assign addr[20360]= -2079176953;
assign addr[20361]= -2088416053;
assign addr[20362]= -2096992772;
assign addr[20363]= -2104904390;
assign addr[20364]= -2112148396;
assign addr[20365]= -2118722494;
assign addr[20366]= -2124624598;
assign addr[20367]= -2129852837;
assign addr[20368]= -2134405552;
assign addr[20369]= -2138281298;
assign addr[20370]= -2141478848;
assign addr[20371]= -2143997187;
assign addr[20372]= -2145835515;
assign addr[20373]= -2146993250;
assign addr[20374]= -2147470025;
assign addr[20375]= -2147265689;
assign addr[20376]= -2146380306;
assign addr[20377]= -2144814157;
assign addr[20378]= -2142567738;
assign addr[20379]= -2139641764;
assign addr[20380]= -2136037160;
assign addr[20381]= -2131755071;
assign addr[20382]= -2126796855;
assign addr[20383]= -2121164085;
assign addr[20384]= -2114858546;
assign addr[20385]= -2107882239;
assign addr[20386]= -2100237377;
assign addr[20387]= -2091926384;
assign addr[20388]= -2082951896;
assign addr[20389]= -2073316760;
assign addr[20390]= -2063024031;
assign addr[20391]= -2052076975;
assign addr[20392]= -2040479063;
assign addr[20393]= -2028233973;
assign addr[20394]= -2015345591;
assign addr[20395]= -2001818002;
assign addr[20396]= -1987655498;
assign addr[20397]= -1972862571;
assign addr[20398]= -1957443913;
assign addr[20399]= -1941404413;
assign addr[20400]= -1924749160;
assign addr[20401]= -1907483436;
assign addr[20402]= -1889612716;
assign addr[20403]= -1871142669;
assign addr[20404]= -1852079154;
assign addr[20405]= -1832428215;
assign addr[20406]= -1812196087;
assign addr[20407]= -1791389186;
assign addr[20408]= -1770014111;
assign addr[20409]= -1748077642;
assign addr[20410]= -1725586737;
assign addr[20411]= -1702548529;
assign addr[20412]= -1678970324;
assign addr[20413]= -1654859602;
assign addr[20414]= -1630224009;
assign addr[20415]= -1605071359;
assign addr[20416]= -1579409630;
assign addr[20417]= -1553246960;
assign addr[20418]= -1526591649;
assign addr[20419]= -1499452149;
assign addr[20420]= -1471837070;
assign addr[20421]= -1443755168;
assign addr[20422]= -1415215352;
assign addr[20423]= -1386226674;
assign addr[20424]= -1356798326;
assign addr[20425]= -1326939644;
assign addr[20426]= -1296660098;
assign addr[20427]= -1265969291;
assign addr[20428]= -1234876957;
assign addr[20429]= -1203392958;
assign addr[20430]= -1171527280;
assign addr[20431]= -1139290029;
assign addr[20432]= -1106691431;
assign addr[20433]= -1073741824;
assign addr[20434]= -1040451659;
assign addr[20435]= -1006831495;
assign addr[20436]= -972891995;
assign addr[20437]= -938643924;
assign addr[20438]= -904098143;
assign addr[20439]= -869265610;
assign addr[20440]= -834157373;
assign addr[20441]= -798784567;
assign addr[20442]= -763158411;
assign addr[20443]= -727290205;
assign addr[20444]= -691191324;
assign addr[20445]= -654873219;
assign addr[20446]= -618347408;
assign addr[20447]= -581625477;
assign addr[20448]= -544719071;
assign addr[20449]= -507639898;
assign addr[20450]= -470399716;
assign addr[20451]= -433010339;
assign addr[20452]= -395483624;
assign addr[20453]= -357831473;
assign addr[20454]= -320065829;
assign addr[20455]= -282198671;
assign addr[20456]= -244242007;
assign addr[20457]= -206207878;
assign addr[20458]= -168108346;
assign addr[20459]= -129955495;
assign addr[20460]= -91761426;
assign addr[20461]= -53538253;
assign addr[20462]= -15298099;
assign addr[20463]= 22946906;
assign addr[20464]= 61184634;
assign addr[20465]= 99402956;
assign addr[20466]= 137589750;
assign addr[20467]= 175732905;
assign addr[20468]= 213820322;
assign addr[20469]= 251839923;
assign addr[20470]= 289779648;
assign addr[20471]= 327627463;
assign addr[20472]= 365371365;
assign addr[20473]= 402999383;
assign addr[20474]= 440499581;
assign addr[20475]= 477860067;
assign addr[20476]= 515068990;
assign addr[20477]= 552114549;
assign addr[20478]= 588984994;
assign addr[20479]= 625668632;
assign addr[20480]= 662153826;
assign addr[20481]= 698429006;
assign addr[20482]= 734482665;
assign addr[20483]= 770303369;
assign addr[20484]= 805879757;
assign addr[20485]= 841200544;
assign addr[20486]= 876254528;
assign addr[20487]= 911030591;
assign addr[20488]= 945517704;
assign addr[20489]= 979704927;
assign addr[20490]= 1013581418;
assign addr[20491]= 1047136432;
assign addr[20492]= 1080359326;
assign addr[20493]= 1113239564;
assign addr[20494]= 1145766716;
assign addr[20495]= 1177930466;
assign addr[20496]= 1209720613;
assign addr[20497]= 1241127074;
assign addr[20498]= 1272139887;
assign addr[20499]= 1302749217;
assign addr[20500]= 1332945355;
assign addr[20501]= 1362718723;
assign addr[20502]= 1392059879;
assign addr[20503]= 1420959516;
assign addr[20504]= 1449408469;
assign addr[20505]= 1477397714;
assign addr[20506]= 1504918373;
assign addr[20507]= 1531961719;
assign addr[20508]= 1558519173;
assign addr[20509]= 1584582314;
assign addr[20510]= 1610142873;
assign addr[20511]= 1635192744;
assign addr[20512]= 1659723983;
assign addr[20513]= 1683728808;
assign addr[20514]= 1707199606;
assign addr[20515]= 1730128933;
assign addr[20516]= 1752509516;
assign addr[20517]= 1774334257;
assign addr[20518]= 1795596234;
assign addr[20519]= 1816288703;
assign addr[20520]= 1836405100;
assign addr[20521]= 1855939047;
assign addr[20522]= 1874884346;
assign addr[20523]= 1893234990;
assign addr[20524]= 1910985158;
assign addr[20525]= 1928129220;
assign addr[20526]= 1944661739;
assign addr[20527]= 1960577471;
assign addr[20528]= 1975871368;
assign addr[20529]= 1990538579;
assign addr[20530]= 2004574453;
assign addr[20531]= 2017974537;
assign addr[20532]= 2030734582;
assign addr[20533]= 2042850540;
assign addr[20534]= 2054318569;
assign addr[20535]= 2065135031;
assign addr[20536]= 2075296495;
assign addr[20537]= 2084799740;
assign addr[20538]= 2093641749;
assign addr[20539]= 2101819720;
assign addr[20540]= 2109331059;
assign addr[20541]= 2116173382;
assign addr[20542]= 2122344521;
assign addr[20543]= 2127842516;
assign addr[20544]= 2132665626;
assign addr[20545]= 2136812319;
assign addr[20546]= 2140281282;
assign addr[20547]= 2143071413;
assign addr[20548]= 2145181827;
assign addr[20549]= 2146611856;
assign addr[20550]= 2147361045;
assign addr[20551]= 2147429158;
assign addr[20552]= 2146816171;
assign addr[20553]= 2145522281;
assign addr[20554]= 2143547897;
assign addr[20555]= 2140893646;
assign addr[20556]= 2137560369;
assign addr[20557]= 2133549123;
assign addr[20558]= 2128861181;
assign addr[20559]= 2123498030;
assign addr[20560]= 2117461370;
assign addr[20561]= 2110753117;
assign addr[20562]= 2103375398;
assign addr[20563]= 2095330553;
assign addr[20564]= 2086621133;
assign addr[20565]= 2077249901;
assign addr[20566]= 2067219829;
assign addr[20567]= 2056534099;
assign addr[20568]= 2045196100;
assign addr[20569]= 2033209426;
assign addr[20570]= 2020577882;
assign addr[20571]= 2007305472;
assign addr[20572]= 1993396407;
assign addr[20573]= 1978855097;
assign addr[20574]= 1963686155;
assign addr[20575]= 1947894393;
assign addr[20576]= 1931484818;
assign addr[20577]= 1914462636;
assign addr[20578]= 1896833245;
assign addr[20579]= 1878602237;
assign addr[20580]= 1859775393;
assign addr[20581]= 1840358687;
assign addr[20582]= 1820358275;
assign addr[20583]= 1799780501;
assign addr[20584]= 1778631892;
assign addr[20585]= 1756919156;
assign addr[20586]= 1734649179;
assign addr[20587]= 1711829025;
assign addr[20588]= 1688465931;
assign addr[20589]= 1664567307;
assign addr[20590]= 1640140734;
assign addr[20591]= 1615193959;
assign addr[20592]= 1589734894;
assign addr[20593]= 1563771613;
assign addr[20594]= 1537312353;
assign addr[20595]= 1510365504;
assign addr[20596]= 1482939614;
assign addr[20597]= 1455043381;
assign addr[20598]= 1426685652;
assign addr[20599]= 1397875423;
assign addr[20600]= 1368621831;
assign addr[20601]= 1338934154;
assign addr[20602]= 1308821808;
assign addr[20603]= 1278294345;
assign addr[20604]= 1247361445;
assign addr[20605]= 1216032921;
assign addr[20606]= 1184318708;
assign addr[20607]= 1152228866;
assign addr[20608]= 1119773573;
assign addr[20609]= 1086963121;
assign addr[20610]= 1053807919;
assign addr[20611]= 1020318481;
assign addr[20612]= 986505429;
assign addr[20613]= 952379488;
assign addr[20614]= 917951481;
assign addr[20615]= 883232329;
assign addr[20616]= 848233042;
assign addr[20617]= 812964722;
assign addr[20618]= 777438554;
assign addr[20619]= 741665807;
assign addr[20620]= 705657826;
assign addr[20621]= 669426032;
assign addr[20622]= 632981917;
assign addr[20623]= 596337040;
assign addr[20624]= 559503022;
assign addr[20625]= 522491548;
assign addr[20626]= 485314355;
assign addr[20627]= 447983235;
assign addr[20628]= 410510029;
assign addr[20629]= 372906622;
assign addr[20630]= 335184940;
assign addr[20631]= 297356948;
assign addr[20632]= 259434643;
assign addr[20633]= 221430054;
assign addr[20634]= 183355234;
assign addr[20635]= 145222259;
assign addr[20636]= 107043224;
assign addr[20637]= 68830239;
assign addr[20638]= 30595422;
assign addr[20639]= -7649098;
assign addr[20640]= -45891193;
assign addr[20641]= -84118732;
assign addr[20642]= -122319591;
assign addr[20643]= -160481654;
assign addr[20644]= -198592817;
assign addr[20645]= -236640993;
assign addr[20646]= -274614114;
assign addr[20647]= -312500135;
assign addr[20648]= -350287041;
assign addr[20649]= -387962847;
assign addr[20650]= -425515602;
assign addr[20651]= -462933398;
assign addr[20652]= -500204365;
assign addr[20653]= -537316682;
assign addr[20654]= -574258580;
assign addr[20655]= -611018340;
assign addr[20656]= -647584304;
assign addr[20657]= -683944874;
assign addr[20658]= -720088517;
assign addr[20659]= -756003771;
assign addr[20660]= -791679244;
assign addr[20661]= -827103620;
assign addr[20662]= -862265664;
assign addr[20663]= -897154224;
assign addr[20664]= -931758235;
assign addr[20665]= -966066720;
assign addr[20666]= -1000068799;
assign addr[20667]= -1033753687;
assign addr[20668]= -1067110699;
assign addr[20669]= -1100129257;
assign addr[20670]= -1132798888;
assign addr[20671]= -1165109230;
assign addr[20672]= -1197050035;
assign addr[20673]= -1228611172;
assign addr[20674]= -1259782632;
assign addr[20675]= -1290554528;
assign addr[20676]= -1320917099;
assign addr[20677]= -1350860716;
assign addr[20678]= -1380375881;
assign addr[20679]= -1409453233;
assign addr[20680]= -1438083551;
assign addr[20681]= -1466257752;
assign addr[20682]= -1493966902;
assign addr[20683]= -1521202211;
assign addr[20684]= -1547955041;
assign addr[20685]= -1574216908;
assign addr[20686]= -1599979481;
assign addr[20687]= -1625234591;
assign addr[20688]= -1649974225;
assign addr[20689]= -1674190539;
assign addr[20690]= -1697875851;
assign addr[20691]= -1721022648;
assign addr[20692]= -1743623590;
assign addr[20693]= -1765671509;
assign addr[20694]= -1787159411;
assign addr[20695]= -1808080480;
assign addr[20696]= -1828428082;
assign addr[20697]= -1848195763;
assign addr[20698]= -1867377253;
assign addr[20699]= -1885966468;
assign addr[20700]= -1903957513;
assign addr[20701]= -1921344681;
assign addr[20702]= -1938122457;
assign addr[20703]= -1954285520;
assign addr[20704]= -1969828744;
assign addr[20705]= -1984747199;
assign addr[20706]= -1999036154;
assign addr[20707]= -2012691075;
assign addr[20708]= -2025707632;
assign addr[20709]= -2038081698;
assign addr[20710]= -2049809346;
assign addr[20711]= -2060886858;
assign addr[20712]= -2071310720;
assign addr[20713]= -2081077626;
assign addr[20714]= -2090184478;
assign addr[20715]= -2098628387;
assign addr[20716]= -2106406677;
assign addr[20717]= -2113516878;
assign addr[20718]= -2119956737;
assign addr[20719]= -2125724211;
assign addr[20720]= -2130817471;
assign addr[20721]= -2135234901;
assign addr[20722]= -2138975100;
assign addr[20723]= -2142036881;
assign addr[20724]= -2144419275;
assign addr[20725]= -2146121524;
assign addr[20726]= -2147143090;
assign addr[20727]= -2147483648;
assign addr[20728]= -2147143090;
assign addr[20729]= -2146121524;
assign addr[20730]= -2144419275;
assign addr[20731]= -2142036881;
assign addr[20732]= -2138975100;
assign addr[20733]= -2135234901;
assign addr[20734]= -2130817471;
assign addr[20735]= -2125724211;
assign addr[20736]= -2119956737;
assign addr[20737]= -2113516878;
assign addr[20738]= -2106406677;
assign addr[20739]= -2098628387;
assign addr[20740]= -2090184478;
assign addr[20741]= -2081077626;
assign addr[20742]= -2071310720;
assign addr[20743]= -2060886858;
assign addr[20744]= -2049809346;
assign addr[20745]= -2038081698;
assign addr[20746]= -2025707632;
assign addr[20747]= -2012691075;
assign addr[20748]= -1999036154;
assign addr[20749]= -1984747199;
assign addr[20750]= -1969828744;
assign addr[20751]= -1954285520;
assign addr[20752]= -1938122457;
assign addr[20753]= -1921344681;
assign addr[20754]= -1903957513;
assign addr[20755]= -1885966468;
assign addr[20756]= -1867377253;
assign addr[20757]= -1848195763;
assign addr[20758]= -1828428082;
assign addr[20759]= -1808080480;
assign addr[20760]= -1787159411;
assign addr[20761]= -1765671509;
assign addr[20762]= -1743623590;
assign addr[20763]= -1721022648;
assign addr[20764]= -1697875851;
assign addr[20765]= -1674190539;
assign addr[20766]= -1649974225;
assign addr[20767]= -1625234591;
assign addr[20768]= -1599979481;
assign addr[20769]= -1574216908;
assign addr[20770]= -1547955041;
assign addr[20771]= -1521202211;
assign addr[20772]= -1493966902;
assign addr[20773]= -1466257752;
assign addr[20774]= -1438083551;
assign addr[20775]= -1409453233;
assign addr[20776]= -1380375881;
assign addr[20777]= -1350860716;
assign addr[20778]= -1320917099;
assign addr[20779]= -1290554528;
assign addr[20780]= -1259782632;
assign addr[20781]= -1228611172;
assign addr[20782]= -1197050035;
assign addr[20783]= -1165109230;
assign addr[20784]= -1132798888;
assign addr[20785]= -1100129257;
assign addr[20786]= -1067110699;
assign addr[20787]= -1033753687;
assign addr[20788]= -1000068799;
assign addr[20789]= -966066720;
assign addr[20790]= -931758235;
assign addr[20791]= -897154224;
assign addr[20792]= -862265664;
assign addr[20793]= -827103620;
assign addr[20794]= -791679244;
assign addr[20795]= -756003771;
assign addr[20796]= -720088517;
assign addr[20797]= -683944874;
assign addr[20798]= -647584304;
assign addr[20799]= -611018340;
assign addr[20800]= -574258580;
assign addr[20801]= -537316682;
assign addr[20802]= -500204365;
assign addr[20803]= -462933398;
assign addr[20804]= -425515602;
assign addr[20805]= -387962847;
assign addr[20806]= -350287041;
assign addr[20807]= -312500135;
assign addr[20808]= -274614114;
assign addr[20809]= -236640993;
assign addr[20810]= -198592817;
assign addr[20811]= -160481654;
assign addr[20812]= -122319591;
assign addr[20813]= -84118732;
assign addr[20814]= -45891193;
assign addr[20815]= -7649098;
assign addr[20816]= 30595422;
assign addr[20817]= 68830239;
assign addr[20818]= 107043224;
assign addr[20819]= 145222259;
assign addr[20820]= 183355234;
assign addr[20821]= 221430054;
assign addr[20822]= 259434643;
assign addr[20823]= 297356948;
assign addr[20824]= 335184940;
assign addr[20825]= 372906622;
assign addr[20826]= 410510029;
assign addr[20827]= 447983235;
assign addr[20828]= 485314355;
assign addr[20829]= 522491548;
assign addr[20830]= 559503022;
assign addr[20831]= 596337040;
assign addr[20832]= 632981917;
assign addr[20833]= 669426032;
assign addr[20834]= 705657826;
assign addr[20835]= 741665807;
assign addr[20836]= 777438554;
assign addr[20837]= 812964722;
assign addr[20838]= 848233042;
assign addr[20839]= 883232329;
assign addr[20840]= 917951481;
assign addr[20841]= 952379488;
assign addr[20842]= 986505429;
assign addr[20843]= 1020318481;
assign addr[20844]= 1053807919;
assign addr[20845]= 1086963121;
assign addr[20846]= 1119773573;
assign addr[20847]= 1152228866;
assign addr[20848]= 1184318708;
assign addr[20849]= 1216032921;
assign addr[20850]= 1247361445;
assign addr[20851]= 1278294345;
assign addr[20852]= 1308821808;
assign addr[20853]= 1338934154;
assign addr[20854]= 1368621831;
assign addr[20855]= 1397875423;
assign addr[20856]= 1426685652;
assign addr[20857]= 1455043381;
assign addr[20858]= 1482939614;
assign addr[20859]= 1510365504;
assign addr[20860]= 1537312353;
assign addr[20861]= 1563771613;
assign addr[20862]= 1589734894;
assign addr[20863]= 1615193959;
assign addr[20864]= 1640140734;
assign addr[20865]= 1664567307;
assign addr[20866]= 1688465931;
assign addr[20867]= 1711829025;
assign addr[20868]= 1734649179;
assign addr[20869]= 1756919156;
assign addr[20870]= 1778631892;
assign addr[20871]= 1799780501;
assign addr[20872]= 1820358275;
assign addr[20873]= 1840358687;
assign addr[20874]= 1859775393;
assign addr[20875]= 1878602237;
assign addr[20876]= 1896833245;
assign addr[20877]= 1914462636;
assign addr[20878]= 1931484818;
assign addr[20879]= 1947894393;
assign addr[20880]= 1963686155;
assign addr[20881]= 1978855097;
assign addr[20882]= 1993396407;
assign addr[20883]= 2007305472;
assign addr[20884]= 2020577882;
assign addr[20885]= 2033209426;
assign addr[20886]= 2045196100;
assign addr[20887]= 2056534099;
assign addr[20888]= 2067219829;
assign addr[20889]= 2077249901;
assign addr[20890]= 2086621133;
assign addr[20891]= 2095330553;
assign addr[20892]= 2103375398;
assign addr[20893]= 2110753117;
assign addr[20894]= 2117461370;
assign addr[20895]= 2123498030;
assign addr[20896]= 2128861181;
assign addr[20897]= 2133549123;
assign addr[20898]= 2137560369;
assign addr[20899]= 2140893646;
assign addr[20900]= 2143547897;
assign addr[20901]= 2145522281;
assign addr[20902]= 2146816171;
assign addr[20903]= 2147429158;
assign addr[20904]= 2147361045;
assign addr[20905]= 2146611856;
assign addr[20906]= 2145181827;
assign addr[20907]= 2143071413;
assign addr[20908]= 2140281282;
assign addr[20909]= 2136812319;
assign addr[20910]= 2132665626;
assign addr[20911]= 2127842516;
assign addr[20912]= 2122344521;
assign addr[20913]= 2116173382;
assign addr[20914]= 2109331059;
assign addr[20915]= 2101819720;
assign addr[20916]= 2093641749;
assign addr[20917]= 2084799740;
assign addr[20918]= 2075296495;
assign addr[20919]= 2065135031;
assign addr[20920]= 2054318569;
assign addr[20921]= 2042850540;
assign addr[20922]= 2030734582;
assign addr[20923]= 2017974537;
assign addr[20924]= 2004574453;
assign addr[20925]= 1990538579;
assign addr[20926]= 1975871368;
assign addr[20927]= 1960577471;
assign addr[20928]= 1944661739;
assign addr[20929]= 1928129220;
assign addr[20930]= 1910985158;
assign addr[20931]= 1893234990;
assign addr[20932]= 1874884346;
assign addr[20933]= 1855939047;
assign addr[20934]= 1836405100;
assign addr[20935]= 1816288703;
assign addr[20936]= 1795596234;
assign addr[20937]= 1774334257;
assign addr[20938]= 1752509516;
assign addr[20939]= 1730128933;
assign addr[20940]= 1707199606;
assign addr[20941]= 1683728808;
assign addr[20942]= 1659723983;
assign addr[20943]= 1635192744;
assign addr[20944]= 1610142873;
assign addr[20945]= 1584582314;
assign addr[20946]= 1558519173;
assign addr[20947]= 1531961719;
assign addr[20948]= 1504918373;
assign addr[20949]= 1477397714;
assign addr[20950]= 1449408469;
assign addr[20951]= 1420959516;
assign addr[20952]= 1392059879;
assign addr[20953]= 1362718723;
assign addr[20954]= 1332945355;
assign addr[20955]= 1302749217;
assign addr[20956]= 1272139887;
assign addr[20957]= 1241127074;
assign addr[20958]= 1209720613;
assign addr[20959]= 1177930466;
assign addr[20960]= 1145766716;
assign addr[20961]= 1113239564;
assign addr[20962]= 1080359326;
assign addr[20963]= 1047136432;
assign addr[20964]= 1013581418;
assign addr[20965]= 979704927;
assign addr[20966]= 945517704;
assign addr[20967]= 911030591;
assign addr[20968]= 876254528;
assign addr[20969]= 841200544;
assign addr[20970]= 805879757;
assign addr[20971]= 770303369;
assign addr[20972]= 734482665;
assign addr[20973]= 698429006;
assign addr[20974]= 662153826;
assign addr[20975]= 625668632;
assign addr[20976]= 588984994;
assign addr[20977]= 552114549;
assign addr[20978]= 515068990;
assign addr[20979]= 477860067;
assign addr[20980]= 440499581;
assign addr[20981]= 402999383;
assign addr[20982]= 365371365;
assign addr[20983]= 327627463;
assign addr[20984]= 289779648;
assign addr[20985]= 251839923;
assign addr[20986]= 213820322;
assign addr[20987]= 175732905;
assign addr[20988]= 137589750;
assign addr[20989]= 99402956;
assign addr[20990]= 61184634;
assign addr[20991]= 22946906;
assign addr[20992]= -15298099;
assign addr[20993]= -53538253;
assign addr[20994]= -91761426;
assign addr[20995]= -129955495;
assign addr[20996]= -168108346;
assign addr[20997]= -206207878;
assign addr[20998]= -244242007;
assign addr[20999]= -282198671;
assign addr[21000]= -320065829;
assign addr[21001]= -357831473;
assign addr[21002]= -395483624;
assign addr[21003]= -433010339;
assign addr[21004]= -470399716;
assign addr[21005]= -507639898;
assign addr[21006]= -544719071;
assign addr[21007]= -581625477;
assign addr[21008]= -618347408;
assign addr[21009]= -654873219;
assign addr[21010]= -691191324;
assign addr[21011]= -727290205;
assign addr[21012]= -763158411;
assign addr[21013]= -798784567;
assign addr[21014]= -834157373;
assign addr[21015]= -869265610;
assign addr[21016]= -904098143;
assign addr[21017]= -938643924;
assign addr[21018]= -972891995;
assign addr[21019]= -1006831495;
assign addr[21020]= -1040451659;
assign addr[21021]= -1073741824;
assign addr[21022]= -1106691431;
assign addr[21023]= -1139290029;
assign addr[21024]= -1171527280;
assign addr[21025]= -1203392958;
assign addr[21026]= -1234876957;
assign addr[21027]= -1265969291;
assign addr[21028]= -1296660098;
assign addr[21029]= -1326939644;
assign addr[21030]= -1356798326;
assign addr[21031]= -1386226674;
assign addr[21032]= -1415215352;
assign addr[21033]= -1443755168;
assign addr[21034]= -1471837070;
assign addr[21035]= -1499452149;
assign addr[21036]= -1526591649;
assign addr[21037]= -1553246960;
assign addr[21038]= -1579409630;
assign addr[21039]= -1605071359;
assign addr[21040]= -1630224009;
assign addr[21041]= -1654859602;
assign addr[21042]= -1678970324;
assign addr[21043]= -1702548529;
assign addr[21044]= -1725586737;
assign addr[21045]= -1748077642;
assign addr[21046]= -1770014111;
assign addr[21047]= -1791389186;
assign addr[21048]= -1812196087;
assign addr[21049]= -1832428215;
assign addr[21050]= -1852079154;
assign addr[21051]= -1871142669;
assign addr[21052]= -1889612716;
assign addr[21053]= -1907483436;
assign addr[21054]= -1924749160;
assign addr[21055]= -1941404413;
assign addr[21056]= -1957443913;
assign addr[21057]= -1972862571;
assign addr[21058]= -1987655498;
assign addr[21059]= -2001818002;
assign addr[21060]= -2015345591;
assign addr[21061]= -2028233973;
assign addr[21062]= -2040479063;
assign addr[21063]= -2052076975;
assign addr[21064]= -2063024031;
assign addr[21065]= -2073316760;
assign addr[21066]= -2082951896;
assign addr[21067]= -2091926384;
assign addr[21068]= -2100237377;
assign addr[21069]= -2107882239;
assign addr[21070]= -2114858546;
assign addr[21071]= -2121164085;
assign addr[21072]= -2126796855;
assign addr[21073]= -2131755071;
assign addr[21074]= -2136037160;
assign addr[21075]= -2139641764;
assign addr[21076]= -2142567738;
assign addr[21077]= -2144814157;
assign addr[21078]= -2146380306;
assign addr[21079]= -2147265689;
assign addr[21080]= -2147470025;
assign addr[21081]= -2146993250;
assign addr[21082]= -2145835515;
assign addr[21083]= -2143997187;
assign addr[21084]= -2141478848;
assign addr[21085]= -2138281298;
assign addr[21086]= -2134405552;
assign addr[21087]= -2129852837;
assign addr[21088]= -2124624598;
assign addr[21089]= -2118722494;
assign addr[21090]= -2112148396;
assign addr[21091]= -2104904390;
assign addr[21092]= -2096992772;
assign addr[21093]= -2088416053;
assign addr[21094]= -2079176953;
assign addr[21095]= -2069278401;
assign addr[21096]= -2058723538;
assign addr[21097]= -2047515711;
assign addr[21098]= -2035658475;
assign addr[21099]= -2023155591;
assign addr[21100]= -2010011024;
assign addr[21101]= -1996228943;
assign addr[21102]= -1981813720;
assign addr[21103]= -1966769926;
assign addr[21104]= -1951102334;
assign addr[21105]= -1934815911;
assign addr[21106]= -1917915825;
assign addr[21107]= -1900407434;
assign addr[21108]= -1882296293;
assign addr[21109]= -1863588145;
assign addr[21110]= -1844288924;
assign addr[21111]= -1824404752;
assign addr[21112]= -1803941934;
assign addr[21113]= -1782906961;
assign addr[21114]= -1761306505;
assign addr[21115]= -1739147417;
assign addr[21116]= -1716436725;
assign addr[21117]= -1693181631;
assign addr[21118]= -1669389513;
assign addr[21119]= -1645067915;
assign addr[21120]= -1620224553;
assign addr[21121]= -1594867305;
assign addr[21122]= -1569004214;
assign addr[21123]= -1542643483;
assign addr[21124]= -1515793473;
assign addr[21125]= -1488462700;
assign addr[21126]= -1460659832;
assign addr[21127]= -1432393688;
assign addr[21128]= -1403673233;
assign addr[21129]= -1374507575;
assign addr[21130]= -1344905966;
assign addr[21131]= -1314877795;
assign addr[21132]= -1284432584;
assign addr[21133]= -1253579991;
assign addr[21134]= -1222329801;
assign addr[21135]= -1190691925;
assign addr[21136]= -1158676398;
assign addr[21137]= -1126293375;
assign addr[21138]= -1093553126;
assign addr[21139]= -1060466036;
assign addr[21140]= -1027042599;
assign addr[21141]= -993293415;
assign addr[21142]= -959229189;
assign addr[21143]= -924860725;
assign addr[21144]= -890198924;
assign addr[21145]= -855254778;
assign addr[21146]= -820039373;
assign addr[21147]= -784563876;
assign addr[21148]= -748839539;
assign addr[21149]= -712877694;
assign addr[21150]= -676689746;
assign addr[21151]= -640287172;
assign addr[21152]= -603681519;
assign addr[21153]= -566884397;
assign addr[21154]= -529907477;
assign addr[21155]= -492762486;
assign addr[21156]= -455461206;
assign addr[21157]= -418015468;
assign addr[21158]= -380437148;
assign addr[21159]= -342738165;
assign addr[21160]= -304930476;
assign addr[21161]= -267026072;
assign addr[21162]= -229036977;
assign addr[21163]= -190975237;
assign addr[21164]= -152852926;
assign addr[21165]= -114682135;
assign addr[21166]= -76474970;
assign addr[21167]= -38243550;
assign addr[21168]= 0;
assign addr[21169]= 38243550;
assign addr[21170]= 76474970;
assign addr[21171]= 114682135;
assign addr[21172]= 152852926;
assign addr[21173]= 190975237;
assign addr[21174]= 229036977;
assign addr[21175]= 267026072;
assign addr[21176]= 304930476;
assign addr[21177]= 342738165;
assign addr[21178]= 380437148;
assign addr[21179]= 418015468;
assign addr[21180]= 455461206;
assign addr[21181]= 492762486;
assign addr[21182]= 529907477;
assign addr[21183]= 566884397;
assign addr[21184]= 603681519;
assign addr[21185]= 640287172;
assign addr[21186]= 676689746;
assign addr[21187]= 712877694;
assign addr[21188]= 748839539;
assign addr[21189]= 784563876;
assign addr[21190]= 820039373;
assign addr[21191]= 855254778;
assign addr[21192]= 890198924;
assign addr[21193]= 924860725;
assign addr[21194]= 959229189;
assign addr[21195]= 993293415;
assign addr[21196]= 1027042599;
assign addr[21197]= 1060466036;
assign addr[21198]= 1093553126;
assign addr[21199]= 1126293375;
assign addr[21200]= 1158676398;
assign addr[21201]= 1190691925;
assign addr[21202]= 1222329801;
assign addr[21203]= 1253579991;
assign addr[21204]= 1284432584;
assign addr[21205]= 1314877795;
assign addr[21206]= 1344905966;
assign addr[21207]= 1374507575;
assign addr[21208]= 1403673233;
assign addr[21209]= 1432393688;
assign addr[21210]= 1460659832;
assign addr[21211]= 1488462700;
assign addr[21212]= 1515793473;
assign addr[21213]= 1542643483;
assign addr[21214]= 1569004214;
assign addr[21215]= 1594867305;
assign addr[21216]= 1620224553;
assign addr[21217]= 1645067915;
assign addr[21218]= 1669389513;
assign addr[21219]= 1693181631;
assign addr[21220]= 1716436725;
assign addr[21221]= 1739147417;
assign addr[21222]= 1761306505;
assign addr[21223]= 1782906961;
assign addr[21224]= 1803941934;
assign addr[21225]= 1824404752;
assign addr[21226]= 1844288924;
assign addr[21227]= 1863588145;
assign addr[21228]= 1882296293;
assign addr[21229]= 1900407434;
assign addr[21230]= 1917915825;
assign addr[21231]= 1934815911;
assign addr[21232]= 1951102334;
assign addr[21233]= 1966769926;
assign addr[21234]= 1981813720;
assign addr[21235]= 1996228943;
assign addr[21236]= 2010011024;
assign addr[21237]= 2023155591;
assign addr[21238]= 2035658475;
assign addr[21239]= 2047515711;
assign addr[21240]= 2058723538;
assign addr[21241]= 2069278401;
assign addr[21242]= 2079176953;
assign addr[21243]= 2088416053;
assign addr[21244]= 2096992772;
assign addr[21245]= 2104904390;
assign addr[21246]= 2112148396;
assign addr[21247]= 2118722494;
assign addr[21248]= 2124624598;
assign addr[21249]= 2129852837;
assign addr[21250]= 2134405552;
assign addr[21251]= 2138281298;
assign addr[21252]= 2141478848;
assign addr[21253]= 2143997187;
assign addr[21254]= 2145835515;
assign addr[21255]= 2146993250;
assign addr[21256]= 2147470025;
assign addr[21257]= 2147265689;
assign addr[21258]= 2146380306;
assign addr[21259]= 2144814157;
assign addr[21260]= 2142567738;
assign addr[21261]= 2139641764;
assign addr[21262]= 2136037160;
assign addr[21263]= 2131755071;
assign addr[21264]= 2126796855;
assign addr[21265]= 2121164085;
assign addr[21266]= 2114858546;
assign addr[21267]= 2107882239;
assign addr[21268]= 2100237377;
assign addr[21269]= 2091926384;
assign addr[21270]= 2082951896;
assign addr[21271]= 2073316760;
assign addr[21272]= 2063024031;
assign addr[21273]= 2052076975;
assign addr[21274]= 2040479063;
assign addr[21275]= 2028233973;
assign addr[21276]= 2015345591;
assign addr[21277]= 2001818002;
assign addr[21278]= 1987655498;
assign addr[21279]= 1972862571;
assign addr[21280]= 1957443913;
assign addr[21281]= 1941404413;
assign addr[21282]= 1924749160;
assign addr[21283]= 1907483436;
assign addr[21284]= 1889612716;
assign addr[21285]= 1871142669;
assign addr[21286]= 1852079154;
assign addr[21287]= 1832428215;
assign addr[21288]= 1812196087;
assign addr[21289]= 1791389186;
assign addr[21290]= 1770014111;
assign addr[21291]= 1748077642;
assign addr[21292]= 1725586737;
assign addr[21293]= 1702548529;
assign addr[21294]= 1678970324;
assign addr[21295]= 1654859602;
assign addr[21296]= 1630224009;
assign addr[21297]= 1605071359;
assign addr[21298]= 1579409630;
assign addr[21299]= 1553246960;
assign addr[21300]= 1526591649;
assign addr[21301]= 1499452149;
assign addr[21302]= 1471837070;
assign addr[21303]= 1443755168;
assign addr[21304]= 1415215352;
assign addr[21305]= 1386226674;
assign addr[21306]= 1356798326;
assign addr[21307]= 1326939644;
assign addr[21308]= 1296660098;
assign addr[21309]= 1265969291;
assign addr[21310]= 1234876957;
assign addr[21311]= 1203392958;
assign addr[21312]= 1171527280;
assign addr[21313]= 1139290029;
assign addr[21314]= 1106691431;
assign addr[21315]= 1073741824;
assign addr[21316]= 1040451659;
assign addr[21317]= 1006831495;
assign addr[21318]= 972891995;
assign addr[21319]= 938643924;
assign addr[21320]= 904098143;
assign addr[21321]= 869265610;
assign addr[21322]= 834157373;
assign addr[21323]= 798784567;
assign addr[21324]= 763158411;
assign addr[21325]= 727290205;
assign addr[21326]= 691191324;
assign addr[21327]= 654873219;
assign addr[21328]= 618347408;
assign addr[21329]= 581625477;
assign addr[21330]= 544719071;
assign addr[21331]= 507639898;
assign addr[21332]= 470399716;
assign addr[21333]= 433010339;
assign addr[21334]= 395483624;
assign addr[21335]= 357831473;
assign addr[21336]= 320065829;
assign addr[21337]= 282198671;
assign addr[21338]= 244242007;
assign addr[21339]= 206207878;
assign addr[21340]= 168108346;
assign addr[21341]= 129955495;
assign addr[21342]= 91761426;
assign addr[21343]= 53538253;
assign addr[21344]= 15298099;
assign addr[21345]= -22946906;
assign addr[21346]= -61184634;
assign addr[21347]= -99402956;
assign addr[21348]= -137589750;
assign addr[21349]= -175732905;
assign addr[21350]= -213820322;
assign addr[21351]= -251839923;
assign addr[21352]= -289779648;
assign addr[21353]= -327627463;
assign addr[21354]= -365371365;
assign addr[21355]= -402999383;
assign addr[21356]= -440499581;
assign addr[21357]= -477860067;
assign addr[21358]= -515068990;
assign addr[21359]= -552114549;
assign addr[21360]= -588984994;
assign addr[21361]= -625668632;
assign addr[21362]= -662153826;
assign addr[21363]= -698429006;
assign addr[21364]= -734482665;
assign addr[21365]= -770303369;
assign addr[21366]= -805879757;
assign addr[21367]= -841200544;
assign addr[21368]= -876254528;
assign addr[21369]= -911030591;
assign addr[21370]= -945517704;
assign addr[21371]= -979704927;
assign addr[21372]= -1013581418;
assign addr[21373]= -1047136432;
assign addr[21374]= -1080359326;
assign addr[21375]= -1113239564;
assign addr[21376]= -1145766716;
assign addr[21377]= -1177930466;
assign addr[21378]= -1209720613;
assign addr[21379]= -1241127074;
assign addr[21380]= -1272139887;
assign addr[21381]= -1302749217;
assign addr[21382]= -1332945355;
assign addr[21383]= -1362718723;
assign addr[21384]= -1392059879;
assign addr[21385]= -1420959516;
assign addr[21386]= -1449408469;
assign addr[21387]= -1477397714;
assign addr[21388]= -1504918373;
assign addr[21389]= -1531961719;
assign addr[21390]= -1558519173;
assign addr[21391]= -1584582314;
assign addr[21392]= -1610142873;
assign addr[21393]= -1635192744;
assign addr[21394]= -1659723983;
assign addr[21395]= -1683728808;
assign addr[21396]= -1707199606;
assign addr[21397]= -1730128933;
assign addr[21398]= -1752509516;
assign addr[21399]= -1774334257;
assign addr[21400]= -1795596234;
assign addr[21401]= -1816288703;
assign addr[21402]= -1836405100;
assign addr[21403]= -1855939047;
assign addr[21404]= -1874884346;
assign addr[21405]= -1893234990;
assign addr[21406]= -1910985158;
assign addr[21407]= -1928129220;
assign addr[21408]= -1944661739;
assign addr[21409]= -1960577471;
assign addr[21410]= -1975871368;
assign addr[21411]= -1990538579;
assign addr[21412]= -2004574453;
assign addr[21413]= -2017974537;
assign addr[21414]= -2030734582;
assign addr[21415]= -2042850540;
assign addr[21416]= -2054318569;
assign addr[21417]= -2065135031;
assign addr[21418]= -2075296495;
assign addr[21419]= -2084799740;
assign addr[21420]= -2093641749;
assign addr[21421]= -2101819720;
assign addr[21422]= -2109331059;
assign addr[21423]= -2116173382;
assign addr[21424]= -2122344521;
assign addr[21425]= -2127842516;
assign addr[21426]= -2132665626;
assign addr[21427]= -2136812319;
assign addr[21428]= -2140281282;
assign addr[21429]= -2143071413;
assign addr[21430]= -2145181827;
assign addr[21431]= -2146611856;
assign addr[21432]= -2147361045;
assign addr[21433]= -2147429158;
assign addr[21434]= -2146816171;
assign addr[21435]= -2145522281;
assign addr[21436]= -2143547897;
assign addr[21437]= -2140893646;
assign addr[21438]= -2137560369;
assign addr[21439]= -2133549123;
assign addr[21440]= -2128861181;
assign addr[21441]= -2123498030;
assign addr[21442]= -2117461370;
assign addr[21443]= -2110753117;
assign addr[21444]= -2103375398;
assign addr[21445]= -2095330553;
assign addr[21446]= -2086621133;
assign addr[21447]= -2077249901;
assign addr[21448]= -2067219829;
assign addr[21449]= -2056534099;
assign addr[21450]= -2045196100;
assign addr[21451]= -2033209426;
assign addr[21452]= -2020577882;
assign addr[21453]= -2007305472;
assign addr[21454]= -1993396407;
assign addr[21455]= -1978855097;
assign addr[21456]= -1963686155;
assign addr[21457]= -1947894393;
assign addr[21458]= -1931484818;
assign addr[21459]= -1914462636;
assign addr[21460]= -1896833245;
assign addr[21461]= -1878602237;
assign addr[21462]= -1859775393;
assign addr[21463]= -1840358687;
assign addr[21464]= -1820358275;
assign addr[21465]= -1799780501;
assign addr[21466]= -1778631892;
assign addr[21467]= -1756919156;
assign addr[21468]= -1734649179;
assign addr[21469]= -1711829025;
assign addr[21470]= -1688465931;
assign addr[21471]= -1664567307;
assign addr[21472]= -1640140734;
assign addr[21473]= -1615193959;
assign addr[21474]= -1589734894;
assign addr[21475]= -1563771613;
assign addr[21476]= -1537312353;
assign addr[21477]= -1510365504;
assign addr[21478]= -1482939614;
assign addr[21479]= -1455043381;
assign addr[21480]= -1426685652;
assign addr[21481]= -1397875423;
assign addr[21482]= -1368621831;
assign addr[21483]= -1338934154;
assign addr[21484]= -1308821808;
assign addr[21485]= -1278294345;
assign addr[21486]= -1247361445;
assign addr[21487]= -1216032921;
assign addr[21488]= -1184318708;
assign addr[21489]= -1152228866;
assign addr[21490]= -1119773573;
assign addr[21491]= -1086963121;
assign addr[21492]= -1053807919;
assign addr[21493]= -1020318481;
assign addr[21494]= -986505429;
assign addr[21495]= -952379488;
assign addr[21496]= -917951481;
assign addr[21497]= -883232329;
assign addr[21498]= -848233042;
assign addr[21499]= -812964722;
assign addr[21500]= -777438554;
assign addr[21501]= -741665807;
assign addr[21502]= -705657826;
assign addr[21503]= -669426032;
assign addr[21504]= -632981917;
assign addr[21505]= -596337040;
assign addr[21506]= -559503022;
assign addr[21507]= -522491548;
assign addr[21508]= -485314355;
assign addr[21509]= -447983235;
assign addr[21510]= -410510029;
assign addr[21511]= -372906622;
assign addr[21512]= -335184940;
assign addr[21513]= -297356948;
assign addr[21514]= -259434643;
assign addr[21515]= -221430054;
assign addr[21516]= -183355234;
assign addr[21517]= -145222259;
assign addr[21518]= -107043224;
assign addr[21519]= -68830239;
assign addr[21520]= -30595422;
assign addr[21521]= 7649098;
assign addr[21522]= 45891193;
assign addr[21523]= 84118732;
assign addr[21524]= 122319591;
assign addr[21525]= 160481654;
assign addr[21526]= 198592817;
assign addr[21527]= 236640993;
assign addr[21528]= 274614114;
assign addr[21529]= 312500135;
assign addr[21530]= 350287041;
assign addr[21531]= 387962847;
assign addr[21532]= 425515602;
assign addr[21533]= 462933398;
assign addr[21534]= 500204365;
assign addr[21535]= 537316682;
assign addr[21536]= 574258580;
assign addr[21537]= 611018340;
assign addr[21538]= 647584304;
assign addr[21539]= 683944874;
assign addr[21540]= 720088517;
assign addr[21541]= 756003771;
assign addr[21542]= 791679244;
assign addr[21543]= 827103620;
assign addr[21544]= 862265664;
assign addr[21545]= 897154224;
assign addr[21546]= 931758235;
assign addr[21547]= 966066720;
assign addr[21548]= 1000068799;
assign addr[21549]= 1033753687;
assign addr[21550]= 1067110699;
assign addr[21551]= 1100129257;
assign addr[21552]= 1132798888;
assign addr[21553]= 1165109230;
assign addr[21554]= 1197050035;
assign addr[21555]= 1228611172;
assign addr[21556]= 1259782632;
assign addr[21557]= 1290554528;
assign addr[21558]= 1320917099;
assign addr[21559]= 1350860716;
assign addr[21560]= 1380375881;
assign addr[21561]= 1409453233;
assign addr[21562]= 1438083551;
assign addr[21563]= 1466257752;
assign addr[21564]= 1493966902;
assign addr[21565]= 1521202211;
assign addr[21566]= 1547955041;
assign addr[21567]= 1574216908;
assign addr[21568]= 1599979481;
assign addr[21569]= 1625234591;
assign addr[21570]= 1649974225;
assign addr[21571]= 1674190539;
assign addr[21572]= 1697875851;
assign addr[21573]= 1721022648;
assign addr[21574]= 1743623590;
assign addr[21575]= 1765671509;
assign addr[21576]= 1787159411;
assign addr[21577]= 1808080480;
assign addr[21578]= 1828428082;
assign addr[21579]= 1848195763;
assign addr[21580]= 1867377253;
assign addr[21581]= 1885966468;
assign addr[21582]= 1903957513;
assign addr[21583]= 1921344681;
assign addr[21584]= 1938122457;
assign addr[21585]= 1954285520;
assign addr[21586]= 1969828744;
assign addr[21587]= 1984747199;
assign addr[21588]= 1999036154;
assign addr[21589]= 2012691075;
assign addr[21590]= 2025707632;
assign addr[21591]= 2038081698;
assign addr[21592]= 2049809346;
assign addr[21593]= 2060886858;
assign addr[21594]= 2071310720;
assign addr[21595]= 2081077626;
assign addr[21596]= 2090184478;
assign addr[21597]= 2098628387;
assign addr[21598]= 2106406677;
assign addr[21599]= 2113516878;
assign addr[21600]= 2119956737;
assign addr[21601]= 2125724211;
assign addr[21602]= 2130817471;
assign addr[21603]= 2135234901;
assign addr[21604]= 2138975100;
assign addr[21605]= 2142036881;
assign addr[21606]= 2144419275;
assign addr[21607]= 2146121524;
assign addr[21608]= 2147143090;
assign addr[21609]= 2147483648;
assign addr[21610]= 2147143090;
assign addr[21611]= 2146121524;
assign addr[21612]= 2144419275;
assign addr[21613]= 2142036881;
assign addr[21614]= 2138975100;
assign addr[21615]= 2135234901;
assign addr[21616]= 2130817471;
assign addr[21617]= 2125724211;
assign addr[21618]= 2119956737;
assign addr[21619]= 2113516878;
assign addr[21620]= 2106406677;
assign addr[21621]= 2098628387;
assign addr[21622]= 2090184478;
assign addr[21623]= 2081077626;
assign addr[21624]= 2071310720;
assign addr[21625]= 2060886858;
assign addr[21626]= 2049809346;
assign addr[21627]= 2038081698;
assign addr[21628]= 2025707632;
assign addr[21629]= 2012691075;
assign addr[21630]= 1999036154;
assign addr[21631]= 1984747199;
assign addr[21632]= 1969828744;
assign addr[21633]= 1954285520;
assign addr[21634]= 1938122457;
assign addr[21635]= 1921344681;
assign addr[21636]= 1903957513;
assign addr[21637]= 1885966468;
assign addr[21638]= 1867377253;
assign addr[21639]= 1848195763;
assign addr[21640]= 1828428082;
assign addr[21641]= 1808080480;
assign addr[21642]= 1787159411;
assign addr[21643]= 1765671509;
assign addr[21644]= 1743623590;
assign addr[21645]= 1721022648;
assign addr[21646]= 1697875851;
assign addr[21647]= 1674190539;
assign addr[21648]= 1649974225;
assign addr[21649]= 1625234591;
assign addr[21650]= 1599979481;
assign addr[21651]= 1574216908;
assign addr[21652]= 1547955041;
assign addr[21653]= 1521202211;
assign addr[21654]= 1493966902;
assign addr[21655]= 1466257752;
assign addr[21656]= 1438083551;
assign addr[21657]= 1409453233;
assign addr[21658]= 1380375881;
assign addr[21659]= 1350860716;
assign addr[21660]= 1320917099;
assign addr[21661]= 1290554528;
assign addr[21662]= 1259782632;
assign addr[21663]= 1228611172;
assign addr[21664]= 1197050035;
assign addr[21665]= 1165109230;
assign addr[21666]= 1132798888;
assign addr[21667]= 1100129257;
assign addr[21668]= 1067110699;
assign addr[21669]= 1033753687;
assign addr[21670]= 1000068799;
assign addr[21671]= 966066720;
assign addr[21672]= 931758235;
assign addr[21673]= 897154224;
assign addr[21674]= 862265664;
assign addr[21675]= 827103620;
assign addr[21676]= 791679244;
assign addr[21677]= 756003771;
assign addr[21678]= 720088517;
assign addr[21679]= 683944874;
assign addr[21680]= 647584304;
assign addr[21681]= 611018340;
assign addr[21682]= 574258580;
assign addr[21683]= 537316682;
assign addr[21684]= 500204365;
assign addr[21685]= 462933398;
assign addr[21686]= 425515602;
assign addr[21687]= 387962847;
assign addr[21688]= 350287041;
assign addr[21689]= 312500135;
assign addr[21690]= 274614114;
assign addr[21691]= 236640993;
assign addr[21692]= 198592817;
assign addr[21693]= 160481654;
assign addr[21694]= 122319591;
assign addr[21695]= 84118732;
assign addr[21696]= 45891193;
assign addr[21697]= 7649098;
assign addr[21698]= -30595422;
assign addr[21699]= -68830239;
assign addr[21700]= -107043224;
assign addr[21701]= -145222259;
assign addr[21702]= -183355234;
assign addr[21703]= -221430054;
assign addr[21704]= -259434643;
assign addr[21705]= -297356948;
assign addr[21706]= -335184940;
assign addr[21707]= -372906622;
assign addr[21708]= -410510029;
assign addr[21709]= -447983235;
assign addr[21710]= -485314355;
assign addr[21711]= -522491548;
assign addr[21712]= -559503022;
assign addr[21713]= -596337040;
assign addr[21714]= -632981917;
assign addr[21715]= -669426032;
assign addr[21716]= -705657826;
assign addr[21717]= -741665807;
assign addr[21718]= -777438554;
assign addr[21719]= -812964722;
assign addr[21720]= -848233042;
assign addr[21721]= -883232329;
assign addr[21722]= -917951481;
assign addr[21723]= -952379488;
assign addr[21724]= -986505429;
assign addr[21725]= -1020318481;
assign addr[21726]= -1053807919;
assign addr[21727]= -1086963121;
assign addr[21728]= -1119773573;
assign addr[21729]= -1152228866;
assign addr[21730]= -1184318708;
assign addr[21731]= -1216032921;
assign addr[21732]= -1247361445;
assign addr[21733]= -1278294345;
assign addr[21734]= -1308821808;
assign addr[21735]= -1338934154;
assign addr[21736]= -1368621831;
assign addr[21737]= -1397875423;
assign addr[21738]= -1426685652;
assign addr[21739]= -1455043381;
assign addr[21740]= -1482939614;
assign addr[21741]= -1510365504;
assign addr[21742]= -1537312353;
assign addr[21743]= -1563771613;
assign addr[21744]= -1589734894;
assign addr[21745]= -1615193959;
assign addr[21746]= -1640140734;
assign addr[21747]= -1664567307;
assign addr[21748]= -1688465931;
assign addr[21749]= -1711829025;
assign addr[21750]= -1734649179;
assign addr[21751]= -1756919156;
assign addr[21752]= -1778631892;
assign addr[21753]= -1799780501;
assign addr[21754]= -1820358275;
assign addr[21755]= -1840358687;
assign addr[21756]= -1859775393;
assign addr[21757]= -1878602237;
assign addr[21758]= -1896833245;
assign addr[21759]= -1914462636;
assign addr[21760]= -1931484818;
assign addr[21761]= -1947894393;
assign addr[21762]= -1963686155;
assign addr[21763]= -1978855097;
assign addr[21764]= -1993396407;
assign addr[21765]= -2007305472;
assign addr[21766]= -2020577882;
assign addr[21767]= -2033209426;
assign addr[21768]= -2045196100;
assign addr[21769]= -2056534099;
assign addr[21770]= -2067219829;
assign addr[21771]= -2077249901;
assign addr[21772]= -2086621133;
assign addr[21773]= -2095330553;
assign addr[21774]= -2103375398;
assign addr[21775]= -2110753117;
assign addr[21776]= -2117461370;
assign addr[21777]= -2123498030;
assign addr[21778]= -2128861181;
assign addr[21779]= -2133549123;
assign addr[21780]= -2137560369;
assign addr[21781]= -2140893646;
assign addr[21782]= -2143547897;
assign addr[21783]= -2145522281;
assign addr[21784]= -2146816171;
assign addr[21785]= -2147429158;
assign addr[21786]= -2147361045;
assign addr[21787]= -2146611856;
assign addr[21788]= -2145181827;
assign addr[21789]= -2143071413;
assign addr[21790]= -2140281282;
assign addr[21791]= -2136812319;
assign addr[21792]= -2132665626;
assign addr[21793]= -2127842516;
assign addr[21794]= -2122344521;
assign addr[21795]= -2116173382;
assign addr[21796]= -2109331059;
assign addr[21797]= -2101819720;
assign addr[21798]= -2093641749;
assign addr[21799]= -2084799740;
assign addr[21800]= -2075296495;
assign addr[21801]= -2065135031;
assign addr[21802]= -2054318569;
assign addr[21803]= -2042850540;
assign addr[21804]= -2030734582;
assign addr[21805]= -2017974537;
assign addr[21806]= -2004574453;
assign addr[21807]= -1990538579;
assign addr[21808]= -1975871368;
assign addr[21809]= -1960577471;
assign addr[21810]= -1944661739;
assign addr[21811]= -1928129220;
assign addr[21812]= -1910985158;
assign addr[21813]= -1893234990;
assign addr[21814]= -1874884346;
assign addr[21815]= -1855939047;
assign addr[21816]= -1836405100;
assign addr[21817]= -1816288703;
assign addr[21818]= -1795596234;
assign addr[21819]= -1774334257;
assign addr[21820]= -1752509516;
assign addr[21821]= -1730128933;
assign addr[21822]= -1707199606;
assign addr[21823]= -1683728808;
assign addr[21824]= -1659723983;
assign addr[21825]= -1635192744;
assign addr[21826]= -1610142873;
assign addr[21827]= -1584582314;
assign addr[21828]= -1558519173;
assign addr[21829]= -1531961719;
assign addr[21830]= -1504918373;
assign addr[21831]= -1477397714;
assign addr[21832]= -1449408469;
assign addr[21833]= -1420959516;
assign addr[21834]= -1392059879;
assign addr[21835]= -1362718723;
assign addr[21836]= -1332945355;
assign addr[21837]= -1302749217;
assign addr[21838]= -1272139887;
assign addr[21839]= -1241127074;
assign addr[21840]= -1209720613;
assign addr[21841]= -1177930466;
assign addr[21842]= -1145766716;
assign addr[21843]= -1113239564;
assign addr[21844]= -1080359326;
assign addr[21845]= -1047136432;
assign addr[21846]= -1013581418;
assign addr[21847]= -979704927;
assign addr[21848]= -945517704;
assign addr[21849]= -911030591;
assign addr[21850]= -876254528;
assign addr[21851]= -841200544;
assign addr[21852]= -805879757;
assign addr[21853]= -770303369;
assign addr[21854]= -734482665;
assign addr[21855]= -698429006;
assign addr[21856]= -662153826;
assign addr[21857]= -625668632;
assign addr[21858]= -588984994;
assign addr[21859]= -552114549;
assign addr[21860]= -515068990;
assign addr[21861]= -477860067;
assign addr[21862]= -440499581;
assign addr[21863]= -402999383;
assign addr[21864]= -365371365;
assign addr[21865]= -327627463;
assign addr[21866]= -289779648;
assign addr[21867]= -251839923;
assign addr[21868]= -213820322;
assign addr[21869]= -175732905;
assign addr[21870]= -137589750;
assign addr[21871]= -99402956;
assign addr[21872]= -61184634;
assign addr[21873]= -22946906;
assign addr[21874]= 15298099;
assign addr[21875]= 53538253;
assign addr[21876]= 91761426;
assign addr[21877]= 129955495;
assign addr[21878]= 168108346;
assign addr[21879]= 206207878;
assign addr[21880]= 244242007;
assign addr[21881]= 282198671;
assign addr[21882]= 320065829;
assign addr[21883]= 357831473;
assign addr[21884]= 395483624;
assign addr[21885]= 433010339;
assign addr[21886]= 470399716;
assign addr[21887]= 507639898;
assign addr[21888]= 544719071;
assign addr[21889]= 581625477;
assign addr[21890]= 618347408;
assign addr[21891]= 654873219;
assign addr[21892]= 691191324;
assign addr[21893]= 727290205;
assign addr[21894]= 763158411;
assign addr[21895]= 798784567;
assign addr[21896]= 834157373;
assign addr[21897]= 869265610;
assign addr[21898]= 904098143;
assign addr[21899]= 938643924;
assign addr[21900]= 972891995;
assign addr[21901]= 1006831495;
assign addr[21902]= 1040451659;
assign addr[21903]= 1073741824;
assign addr[21904]= 1106691431;
assign addr[21905]= 1139290029;
assign addr[21906]= 1171527280;
assign addr[21907]= 1203392958;
assign addr[21908]= 1234876957;
assign addr[21909]= 1265969291;
assign addr[21910]= 1296660098;
assign addr[21911]= 1326939644;
assign addr[21912]= 1356798326;
assign addr[21913]= 1386226674;
assign addr[21914]= 1415215352;
assign addr[21915]= 1443755168;
assign addr[21916]= 1471837070;
assign addr[21917]= 1499452149;
assign addr[21918]= 1526591649;
assign addr[21919]= 1553246960;
assign addr[21920]= 1579409630;
assign addr[21921]= 1605071359;
assign addr[21922]= 1630224009;
assign addr[21923]= 1654859602;
assign addr[21924]= 1678970324;
assign addr[21925]= 1702548529;
assign addr[21926]= 1725586737;
assign addr[21927]= 1748077642;
assign addr[21928]= 1770014111;
assign addr[21929]= 1791389186;
assign addr[21930]= 1812196087;
assign addr[21931]= 1832428215;
assign addr[21932]= 1852079154;
assign addr[21933]= 1871142669;
assign addr[21934]= 1889612716;
assign addr[21935]= 1907483436;
assign addr[21936]= 1924749160;
assign addr[21937]= 1941404413;
assign addr[21938]= 1957443913;
assign addr[21939]= 1972862571;
assign addr[21940]= 1987655498;
assign addr[21941]= 2001818002;
assign addr[21942]= 2015345591;
assign addr[21943]= 2028233973;
assign addr[21944]= 2040479063;
assign addr[21945]= 2052076975;
assign addr[21946]= 2063024031;
assign addr[21947]= 2073316760;
assign addr[21948]= 2082951896;
assign addr[21949]= 2091926384;
assign addr[21950]= 2100237377;
assign addr[21951]= 2107882239;
assign addr[21952]= 2114858546;
assign addr[21953]= 2121164085;
assign addr[21954]= 2126796855;
assign addr[21955]= 2131755071;
assign addr[21956]= 2136037160;
assign addr[21957]= 2139641764;
assign addr[21958]= 2142567738;
assign addr[21959]= 2144814157;
assign addr[21960]= 2146380306;
assign addr[21961]= 2147265689;
assign addr[21962]= 2147470025;
assign addr[21963]= 2146993250;
assign addr[21964]= 2145835515;
assign addr[21965]= 2143997187;
assign addr[21966]= 2141478848;
assign addr[21967]= 2138281298;
assign addr[21968]= 2134405552;
assign addr[21969]= 2129852837;
assign addr[21970]= 2124624598;
assign addr[21971]= 2118722494;
assign addr[21972]= 2112148396;
assign addr[21973]= 2104904390;
assign addr[21974]= 2096992772;
assign addr[21975]= 2088416053;
assign addr[21976]= 2079176953;
assign addr[21977]= 2069278401;
assign addr[21978]= 2058723538;
assign addr[21979]= 2047515711;
assign addr[21980]= 2035658475;
assign addr[21981]= 2023155591;
assign addr[21982]= 2010011024;
assign addr[21983]= 1996228943;
assign addr[21984]= 1981813720;
assign addr[21985]= 1966769926;
assign addr[21986]= 1951102334;
assign addr[21987]= 1934815911;
assign addr[21988]= 1917915825;
assign addr[21989]= 1900407434;
assign addr[21990]= 1882296293;
assign addr[21991]= 1863588145;
assign addr[21992]= 1844288924;
assign addr[21993]= 1824404752;
assign addr[21994]= 1803941934;
assign addr[21995]= 1782906961;
assign addr[21996]= 1761306505;
assign addr[21997]= 1739147417;
assign addr[21998]= 1716436725;
assign addr[21999]= 1693181631;
assign addr[22000]= 1669389513;
assign addr[22001]= 1645067915;
assign addr[22002]= 1620224553;
assign addr[22003]= 1594867305;
assign addr[22004]= 1569004214;
assign addr[22005]= 1542643483;
assign addr[22006]= 1515793473;
assign addr[22007]= 1488462700;
assign addr[22008]= 1460659832;
assign addr[22009]= 1432393688;
assign addr[22010]= 1403673233;
assign addr[22011]= 1374507575;
assign addr[22012]= 1344905966;
assign addr[22013]= 1314877795;
assign addr[22014]= 1284432584;
assign addr[22015]= 1253579991;
assign addr[22016]= 1222329801;
assign addr[22017]= 1190691925;
assign addr[22018]= 1158676398;
assign addr[22019]= 1126293375;
assign addr[22020]= 1093553126;
assign addr[22021]= 1060466036;
assign addr[22022]= 1027042599;
assign addr[22023]= 993293415;
assign addr[22024]= 959229189;
assign addr[22025]= 924860725;
assign addr[22026]= 890198924;
assign addr[22027]= 855254778;
assign addr[22028]= 820039373;
assign addr[22029]= 784563876;
assign addr[22030]= 748839539;
assign addr[22031]= 712877694;
assign addr[22032]= 676689746;
assign addr[22033]= 640287172;
assign addr[22034]= 603681519;
assign addr[22035]= 566884397;
assign addr[22036]= 529907477;
assign addr[22037]= 492762486;
assign addr[22038]= 455461206;
assign addr[22039]= 418015468;
assign addr[22040]= 380437148;
assign addr[22041]= 342738165;
assign addr[22042]= 304930476;
assign addr[22043]= 267026072;
assign addr[22044]= 229036977;
assign addr[22045]= 190975237;
assign addr[22046]= 152852926;
assign addr[22047]= 114682135;
assign addr[22048]= 76474970;
assign addr[22049]= 38243550;
assign addr[22050]= 0;
assign addr[22051]= -38243550;
assign addr[22052]= -76474970;
assign addr[22053]= -114682135;
assign addr[22054]= -152852926;
assign addr[22055]= -190975237;
assign addr[22056]= -229036977;
assign addr[22057]= -267026072;
assign addr[22058]= -304930476;
assign addr[22059]= -342738165;
assign addr[22060]= -380437148;
assign addr[22061]= -418015468;
assign addr[22062]= -455461206;
assign addr[22063]= -492762486;
assign addr[22064]= -529907477;
assign addr[22065]= -566884397;
assign addr[22066]= -603681519;
assign addr[22067]= -640287172;
assign addr[22068]= -676689746;
assign addr[22069]= -712877694;
assign addr[22070]= -748839539;
assign addr[22071]= -784563876;
assign addr[22072]= -820039373;
assign addr[22073]= -855254778;
assign addr[22074]= -890198924;
assign addr[22075]= -924860725;
assign addr[22076]= -959229189;
assign addr[22077]= -993293415;
assign addr[22078]= -1027042599;
assign addr[22079]= -1060466036;
assign addr[22080]= -1093553126;
assign addr[22081]= -1126293375;
assign addr[22082]= -1158676398;
assign addr[22083]= -1190691925;
assign addr[22084]= -1222329801;
assign addr[22085]= -1253579991;
assign addr[22086]= -1284432584;
assign addr[22087]= -1314877795;
assign addr[22088]= -1344905966;
assign addr[22089]= -1374507575;
assign addr[22090]= -1403673233;
assign addr[22091]= -1432393688;
assign addr[22092]= -1460659832;
assign addr[22093]= -1488462700;
assign addr[22094]= -1515793473;
assign addr[22095]= -1542643483;
assign addr[22096]= -1569004214;
assign addr[22097]= -1594867305;
assign addr[22098]= -1620224553;
assign addr[22099]= -1645067915;
assign addr[22100]= -1669389513;
assign addr[22101]= -1693181631;
assign addr[22102]= -1716436725;
assign addr[22103]= -1739147417;
assign addr[22104]= -1761306505;
assign addr[22105]= -1782906961;
assign addr[22106]= -1803941934;
assign addr[22107]= -1824404752;
assign addr[22108]= -1844288924;
assign addr[22109]= -1863588145;
assign addr[22110]= -1882296293;
assign addr[22111]= -1900407434;
assign addr[22112]= -1917915825;
assign addr[22113]= -1934815911;
assign addr[22114]= -1951102334;
assign addr[22115]= -1966769926;
assign addr[22116]= -1981813720;
assign addr[22117]= -1996228943;
assign addr[22118]= -2010011024;
assign addr[22119]= -2023155591;
assign addr[22120]= -2035658475;
assign addr[22121]= -2047515711;
assign addr[22122]= -2058723538;
assign addr[22123]= -2069278401;
assign addr[22124]= -2079176953;
assign addr[22125]= -2088416053;
assign addr[22126]= -2096992772;
assign addr[22127]= -2104904390;
assign addr[22128]= -2112148396;
assign addr[22129]= -2118722494;
assign addr[22130]= -2124624598;
assign addr[22131]= -2129852837;
assign addr[22132]= -2134405552;
assign addr[22133]= -2138281298;
assign addr[22134]= -2141478848;
assign addr[22135]= -2143997187;
assign addr[22136]= -2145835515;
assign addr[22137]= -2146993250;
assign addr[22138]= -2147470025;
assign addr[22139]= -2147265689;
assign addr[22140]= -2146380306;
assign addr[22141]= -2144814157;
assign addr[22142]= -2142567738;
assign addr[22143]= -2139641764;
assign addr[22144]= -2136037160;
assign addr[22145]= -2131755071;
assign addr[22146]= -2126796855;
assign addr[22147]= -2121164085;
assign addr[22148]= -2114858546;
assign addr[22149]= -2107882239;
assign addr[22150]= -2100237377;
assign addr[22151]= -2091926384;
assign addr[22152]= -2082951896;
assign addr[22153]= -2073316760;
assign addr[22154]= -2063024031;
assign addr[22155]= -2052076975;
assign addr[22156]= -2040479063;
assign addr[22157]= -2028233973;
assign addr[22158]= -2015345591;
assign addr[22159]= -2001818002;
assign addr[22160]= -1987655498;
assign addr[22161]= -1972862571;
assign addr[22162]= -1957443913;
assign addr[22163]= -1941404413;
assign addr[22164]= -1924749160;
assign addr[22165]= -1907483436;
assign addr[22166]= -1889612716;
assign addr[22167]= -1871142669;
assign addr[22168]= -1852079154;
assign addr[22169]= -1832428215;
assign addr[22170]= -1812196087;
assign addr[22171]= -1791389186;
assign addr[22172]= -1770014111;
assign addr[22173]= -1748077642;
assign addr[22174]= -1725586737;
assign addr[22175]= -1702548529;
assign addr[22176]= -1678970324;
assign addr[22177]= -1654859602;
assign addr[22178]= -1630224009;
assign addr[22179]= -1605071359;
assign addr[22180]= -1579409630;
assign addr[22181]= -1553246960;
assign addr[22182]= -1526591649;
assign addr[22183]= -1499452149;
assign addr[22184]= -1471837070;
assign addr[22185]= -1443755168;
assign addr[22186]= -1415215352;
assign addr[22187]= -1386226674;
assign addr[22188]= -1356798326;
assign addr[22189]= -1326939644;
assign addr[22190]= -1296660098;
assign addr[22191]= -1265969291;
assign addr[22192]= -1234876957;
assign addr[22193]= -1203392958;
assign addr[22194]= -1171527280;
assign addr[22195]= -1139290029;
assign addr[22196]= -1106691431;
assign addr[22197]= -1073741824;
assign addr[22198]= -1040451659;
assign addr[22199]= -1006831495;
assign addr[22200]= -972891995;
assign addr[22201]= -938643924;
assign addr[22202]= -904098143;
assign addr[22203]= -869265610;
assign addr[22204]= -834157373;
assign addr[22205]= -798784567;
assign addr[22206]= -763158411;
assign addr[22207]= -727290205;
assign addr[22208]= -691191324;
assign addr[22209]= -654873219;
assign addr[22210]= -618347408;
assign addr[22211]= -581625477;
assign addr[22212]= -544719071;
assign addr[22213]= -507639898;
assign addr[22214]= -470399716;
assign addr[22215]= -433010339;
assign addr[22216]= -395483624;
assign addr[22217]= -357831473;
assign addr[22218]= -320065829;
assign addr[22219]= -282198671;
assign addr[22220]= -244242007;
assign addr[22221]= -206207878;
assign addr[22222]= -168108346;
assign addr[22223]= -129955495;
assign addr[22224]= -91761426;
assign addr[22225]= -53538253;
assign addr[22226]= -15298099;
assign addr[22227]= 22946906;
assign addr[22228]= 61184634;
assign addr[22229]= 99402956;
assign addr[22230]= 137589750;
assign addr[22231]= 175732905;
assign addr[22232]= 213820322;
assign addr[22233]= 251839923;
assign addr[22234]= 289779648;
assign addr[22235]= 327627463;
assign addr[22236]= 365371365;
assign addr[22237]= 402999383;
assign addr[22238]= 440499581;
assign addr[22239]= 477860067;
assign addr[22240]= 515068990;
assign addr[22241]= 552114549;
assign addr[22242]= 588984994;
assign addr[22243]= 625668632;
assign addr[22244]= 662153826;
assign addr[22245]= 698429006;
assign addr[22246]= 734482665;
assign addr[22247]= 770303369;
assign addr[22248]= 805879757;
assign addr[22249]= 841200544;
assign addr[22250]= 876254528;
assign addr[22251]= 911030591;
assign addr[22252]= 945517704;
assign addr[22253]= 979704927;
assign addr[22254]= 1013581418;
assign addr[22255]= 1047136432;
assign addr[22256]= 1080359326;
assign addr[22257]= 1113239564;
assign addr[22258]= 1145766716;
assign addr[22259]= 1177930466;
assign addr[22260]= 1209720613;
assign addr[22261]= 1241127074;
assign addr[22262]= 1272139887;
assign addr[22263]= 1302749217;
assign addr[22264]= 1332945355;
assign addr[22265]= 1362718723;
assign addr[22266]= 1392059879;
assign addr[22267]= 1420959516;
assign addr[22268]= 1449408469;
assign addr[22269]= 1477397714;
assign addr[22270]= 1504918373;
assign addr[22271]= 1531961719;
assign addr[22272]= 1558519173;
assign addr[22273]= 1584582314;
assign addr[22274]= 1610142873;
assign addr[22275]= 1635192744;
assign addr[22276]= 1659723983;
assign addr[22277]= 1683728808;
assign addr[22278]= 1707199606;
assign addr[22279]= 1730128933;
assign addr[22280]= 1752509516;
assign addr[22281]= 1774334257;
assign addr[22282]= 1795596234;
assign addr[22283]= 1816288703;
assign addr[22284]= 1836405100;
assign addr[22285]= 1855939047;
assign addr[22286]= 1874884346;
assign addr[22287]= 1893234990;
assign addr[22288]= 1910985158;
assign addr[22289]= 1928129220;
assign addr[22290]= 1944661739;
assign addr[22291]= 1960577471;
assign addr[22292]= 1975871368;
assign addr[22293]= 1990538579;
assign addr[22294]= 2004574453;
assign addr[22295]= 2017974537;
assign addr[22296]= 2030734582;
assign addr[22297]= 2042850540;
assign addr[22298]= 2054318569;
assign addr[22299]= 2065135031;
assign addr[22300]= 2075296495;
assign addr[22301]= 2084799740;
assign addr[22302]= 2093641749;
assign addr[22303]= 2101819720;
assign addr[22304]= 2109331059;
assign addr[22305]= 2116173382;
assign addr[22306]= 2122344521;
assign addr[22307]= 2127842516;
assign addr[22308]= 2132665626;
assign addr[22309]= 2136812319;
assign addr[22310]= 2140281282;
assign addr[22311]= 2143071413;
assign addr[22312]= 2145181827;
assign addr[22313]= 2146611856;
assign addr[22314]= 2147361045;
assign addr[22315]= 2147429158;
assign addr[22316]= 2146816171;
assign addr[22317]= 2145522281;
assign addr[22318]= 2143547897;
assign addr[22319]= 2140893646;
assign addr[22320]= 2137560369;
assign addr[22321]= 2133549123;
assign addr[22322]= 2128861181;
assign addr[22323]= 2123498030;
assign addr[22324]= 2117461370;
assign addr[22325]= 2110753117;
assign addr[22326]= 2103375398;
assign addr[22327]= 2095330553;
assign addr[22328]= 2086621133;
assign addr[22329]= 2077249901;
assign addr[22330]= 2067219829;
assign addr[22331]= 2056534099;
assign addr[22332]= 2045196100;
assign addr[22333]= 2033209426;
assign addr[22334]= 2020577882;
assign addr[22335]= 2007305472;
assign addr[22336]= 1993396407;
assign addr[22337]= 1978855097;
assign addr[22338]= 1963686155;
assign addr[22339]= 1947894393;
assign addr[22340]= 1931484818;
assign addr[22341]= 1914462636;
assign addr[22342]= 1896833245;
assign addr[22343]= 1878602237;
assign addr[22344]= 1859775393;
assign addr[22345]= 1840358687;
assign addr[22346]= 1820358275;
assign addr[22347]= 1799780501;
assign addr[22348]= 1778631892;
assign addr[22349]= 1756919156;
assign addr[22350]= 1734649179;
assign addr[22351]= 1711829025;
assign addr[22352]= 1688465931;
assign addr[22353]= 1664567307;
assign addr[22354]= 1640140734;
assign addr[22355]= 1615193959;
assign addr[22356]= 1589734894;
assign addr[22357]= 1563771613;
assign addr[22358]= 1537312353;
assign addr[22359]= 1510365504;
assign addr[22360]= 1482939614;
assign addr[22361]= 1455043381;
assign addr[22362]= 1426685652;
assign addr[22363]= 1397875423;
assign addr[22364]= 1368621831;
assign addr[22365]= 1338934154;
assign addr[22366]= 1308821808;
assign addr[22367]= 1278294345;
assign addr[22368]= 1247361445;
assign addr[22369]= 1216032921;
assign addr[22370]= 1184318708;
assign addr[22371]= 1152228866;
assign addr[22372]= 1119773573;
assign addr[22373]= 1086963121;
assign addr[22374]= 1053807919;
assign addr[22375]= 1020318481;
assign addr[22376]= 986505429;
assign addr[22377]= 952379488;
assign addr[22378]= 917951481;
assign addr[22379]= 883232329;
assign addr[22380]= 848233042;
assign addr[22381]= 812964722;
assign addr[22382]= 777438554;
assign addr[22383]= 741665807;
assign addr[22384]= 705657826;
assign addr[22385]= 669426032;
assign addr[22386]= 632981917;
assign addr[22387]= 596337040;
assign addr[22388]= 559503022;
assign addr[22389]= 522491548;
assign addr[22390]= 485314355;
assign addr[22391]= 447983235;
assign addr[22392]= 410510029;
assign addr[22393]= 372906622;
assign addr[22394]= 335184940;
assign addr[22395]= 297356948;
assign addr[22396]= 259434643;
assign addr[22397]= 221430054;
assign addr[22398]= 183355234;
assign addr[22399]= 145222259;
assign addr[22400]= 107043224;
assign addr[22401]= 68830239;
assign addr[22402]= 30595422;
assign addr[22403]= -7649098;
assign addr[22404]= -45891193;
assign addr[22405]= -84118732;
assign addr[22406]= -122319591;
assign addr[22407]= -160481654;
assign addr[22408]= -198592817;
assign addr[22409]= -236640993;
assign addr[22410]= -274614114;
assign addr[22411]= -312500135;
assign addr[22412]= -350287041;
assign addr[22413]= -387962847;
assign addr[22414]= -425515602;
assign addr[22415]= -462933398;
assign addr[22416]= -500204365;
assign addr[22417]= -537316682;
assign addr[22418]= -574258580;
assign addr[22419]= -611018340;
assign addr[22420]= -647584304;
assign addr[22421]= -683944874;
assign addr[22422]= -720088517;
assign addr[22423]= -756003771;
assign addr[22424]= -791679244;
assign addr[22425]= -827103620;
assign addr[22426]= -862265664;
assign addr[22427]= -897154224;
assign addr[22428]= -931758235;
assign addr[22429]= -966066720;
assign addr[22430]= -1000068799;
assign addr[22431]= -1033753687;
assign addr[22432]= -1067110699;
assign addr[22433]= -1100129257;
assign addr[22434]= -1132798888;
assign addr[22435]= -1165109230;
assign addr[22436]= -1197050035;
assign addr[22437]= -1228611172;
assign addr[22438]= -1259782632;
assign addr[22439]= -1290554528;
assign addr[22440]= -1320917099;
assign addr[22441]= -1350860716;
assign addr[22442]= -1380375881;
assign addr[22443]= -1409453233;
assign addr[22444]= -1438083551;
assign addr[22445]= -1466257752;
assign addr[22446]= -1493966902;
assign addr[22447]= -1521202211;
assign addr[22448]= -1547955041;
assign addr[22449]= -1574216908;
assign addr[22450]= -1599979481;
assign addr[22451]= -1625234591;
assign addr[22452]= -1649974225;
assign addr[22453]= -1674190539;
assign addr[22454]= -1697875851;
assign addr[22455]= -1721022648;
assign addr[22456]= -1743623590;
assign addr[22457]= -1765671509;
assign addr[22458]= -1787159411;
assign addr[22459]= -1808080480;
assign addr[22460]= -1828428082;
assign addr[22461]= -1848195763;
assign addr[22462]= -1867377253;
assign addr[22463]= -1885966468;
assign addr[22464]= -1903957513;
assign addr[22465]= -1921344681;
assign addr[22466]= -1938122457;
assign addr[22467]= -1954285520;
assign addr[22468]= -1969828744;
assign addr[22469]= -1984747199;
assign addr[22470]= -1999036154;
assign addr[22471]= -2012691075;
assign addr[22472]= -2025707632;
assign addr[22473]= -2038081698;
assign addr[22474]= -2049809346;
assign addr[22475]= -2060886858;
assign addr[22476]= -2071310720;
assign addr[22477]= -2081077626;
assign addr[22478]= -2090184478;
assign addr[22479]= -2098628387;
assign addr[22480]= -2106406677;
assign addr[22481]= -2113516878;
assign addr[22482]= -2119956737;
assign addr[22483]= -2125724211;
assign addr[22484]= -2130817471;
assign addr[22485]= -2135234901;
assign addr[22486]= -2138975100;
assign addr[22487]= -2142036881;
assign addr[22488]= -2144419275;
assign addr[22489]= -2146121524;
assign addr[22490]= -2147143090;
assign addr[22491]= -2147483648;
assign addr[22492]= -2147143090;
assign addr[22493]= -2146121524;
assign addr[22494]= -2144419275;
assign addr[22495]= -2142036881;
assign addr[22496]= -2138975100;
assign addr[22497]= -2135234901;
assign addr[22498]= -2130817471;
assign addr[22499]= -2125724211;
assign addr[22500]= -2119956737;
assign addr[22501]= -2113516878;
assign addr[22502]= -2106406677;
assign addr[22503]= -2098628387;
assign addr[22504]= -2090184478;
assign addr[22505]= -2081077626;
assign addr[22506]= -2071310720;
assign addr[22507]= -2060886858;
assign addr[22508]= -2049809346;
assign addr[22509]= -2038081698;
assign addr[22510]= -2025707632;
assign addr[22511]= -2012691075;
assign addr[22512]= -1999036154;
assign addr[22513]= -1984747199;
assign addr[22514]= -1969828744;
assign addr[22515]= -1954285520;
assign addr[22516]= -1938122457;
assign addr[22517]= -1921344681;
assign addr[22518]= -1903957513;
assign addr[22519]= -1885966468;
assign addr[22520]= -1867377253;
assign addr[22521]= -1848195763;
assign addr[22522]= -1828428082;
assign addr[22523]= -1808080480;
assign addr[22524]= -1787159411;
assign addr[22525]= -1765671509;
assign addr[22526]= -1743623590;
assign addr[22527]= -1721022648;
assign addr[22528]= -1697875851;
assign addr[22529]= -1674190539;
assign addr[22530]= -1649974225;
assign addr[22531]= -1625234591;
assign addr[22532]= -1599979481;
assign addr[22533]= -1574216908;
assign addr[22534]= -1547955041;
assign addr[22535]= -1521202211;
assign addr[22536]= -1493966902;
assign addr[22537]= -1466257752;
assign addr[22538]= -1438083551;
assign addr[22539]= -1409453233;
assign addr[22540]= -1380375881;
assign addr[22541]= -1350860716;
assign addr[22542]= -1320917099;
assign addr[22543]= -1290554528;
assign addr[22544]= -1259782632;
assign addr[22545]= -1228611172;
assign addr[22546]= -1197050035;
assign addr[22547]= -1165109230;
assign addr[22548]= -1132798888;
assign addr[22549]= -1100129257;
assign addr[22550]= -1067110699;
assign addr[22551]= -1033753687;
assign addr[22552]= -1000068799;
assign addr[22553]= -966066720;
assign addr[22554]= -931758235;
assign addr[22555]= -897154224;
assign addr[22556]= -862265664;
assign addr[22557]= -827103620;
assign addr[22558]= -791679244;
assign addr[22559]= -756003771;
assign addr[22560]= -720088517;
assign addr[22561]= -683944874;
assign addr[22562]= -647584304;
assign addr[22563]= -611018340;
assign addr[22564]= -574258580;
assign addr[22565]= -537316682;
assign addr[22566]= -500204365;
assign addr[22567]= -462933398;
assign addr[22568]= -425515602;
assign addr[22569]= -387962847;
assign addr[22570]= -350287041;
assign addr[22571]= -312500135;
assign addr[22572]= -274614114;
assign addr[22573]= -236640993;
assign addr[22574]= -198592817;
assign addr[22575]= -160481654;
assign addr[22576]= -122319591;
assign addr[22577]= -84118732;
assign addr[22578]= -45891193;
assign addr[22579]= -7649098;
assign addr[22580]= 30595422;
assign addr[22581]= 68830239;
assign addr[22582]= 107043224;
assign addr[22583]= 145222259;
assign addr[22584]= 183355234;
assign addr[22585]= 221430054;
assign addr[22586]= 259434643;
assign addr[22587]= 297356948;
assign addr[22588]= 335184940;
assign addr[22589]= 372906622;
assign addr[22590]= 410510029;
assign addr[22591]= 447983235;
assign addr[22592]= 485314355;
assign addr[22593]= 522491548;
assign addr[22594]= 559503022;
assign addr[22595]= 596337040;
assign addr[22596]= 632981917;
assign addr[22597]= 669426032;
assign addr[22598]= 705657826;
assign addr[22599]= 741665807;
assign addr[22600]= 777438554;
assign addr[22601]= 812964722;
assign addr[22602]= 848233042;
assign addr[22603]= 883232329;
assign addr[22604]= 917951481;
assign addr[22605]= 952379488;
assign addr[22606]= 986505429;
assign addr[22607]= 1020318481;
assign addr[22608]= 1053807919;
assign addr[22609]= 1086963121;
assign addr[22610]= 1119773573;
assign addr[22611]= 1152228866;
assign addr[22612]= 1184318708;
assign addr[22613]= 1216032921;
assign addr[22614]= 1247361445;
assign addr[22615]= 1278294345;
assign addr[22616]= 1308821808;
assign addr[22617]= 1338934154;
assign addr[22618]= 1368621831;
assign addr[22619]= 1397875423;
assign addr[22620]= 1426685652;
assign addr[22621]= 1455043381;
assign addr[22622]= 1482939614;
assign addr[22623]= 1510365504;
assign addr[22624]= 1537312353;
assign addr[22625]= 1563771613;
assign addr[22626]= 1589734894;
assign addr[22627]= 1615193959;
assign addr[22628]= 1640140734;
assign addr[22629]= 1664567307;
assign addr[22630]= 1688465931;
assign addr[22631]= 1711829025;
assign addr[22632]= 1734649179;
assign addr[22633]= 1756919156;
assign addr[22634]= 1778631892;
assign addr[22635]= 1799780501;
assign addr[22636]= 1820358275;
assign addr[22637]= 1840358687;
assign addr[22638]= 1859775393;
assign addr[22639]= 1878602237;
assign addr[22640]= 1896833245;
assign addr[22641]= 1914462636;
assign addr[22642]= 1931484818;
assign addr[22643]= 1947894393;
assign addr[22644]= 1963686155;
assign addr[22645]= 1978855097;
assign addr[22646]= 1993396407;
assign addr[22647]= 2007305472;
assign addr[22648]= 2020577882;
assign addr[22649]= 2033209426;
assign addr[22650]= 2045196100;
assign addr[22651]= 2056534099;
assign addr[22652]= 2067219829;
assign addr[22653]= 2077249901;
assign addr[22654]= 2086621133;
assign addr[22655]= 2095330553;
assign addr[22656]= 2103375398;
assign addr[22657]= 2110753117;
assign addr[22658]= 2117461370;
assign addr[22659]= 2123498030;
assign addr[22660]= 2128861181;
assign addr[22661]= 2133549123;
assign addr[22662]= 2137560369;
assign addr[22663]= 2140893646;
assign addr[22664]= 2143547897;
assign addr[22665]= 2145522281;
assign addr[22666]= 2146816171;
assign addr[22667]= 2147429158;
assign addr[22668]= 2147361045;
assign addr[22669]= 2146611856;
assign addr[22670]= 2145181827;
assign addr[22671]= 2143071413;
assign addr[22672]= 2140281282;
assign addr[22673]= 2136812319;
assign addr[22674]= 2132665626;
assign addr[22675]= 2127842516;
assign addr[22676]= 2122344521;
assign addr[22677]= 2116173382;
assign addr[22678]= 2109331059;
assign addr[22679]= 2101819720;
assign addr[22680]= 2093641749;
assign addr[22681]= 2084799740;
assign addr[22682]= 2075296495;
assign addr[22683]= 2065135031;
assign addr[22684]= 2054318569;
assign addr[22685]= 2042850540;
assign addr[22686]= 2030734582;
assign addr[22687]= 2017974537;
assign addr[22688]= 2004574453;
assign addr[22689]= 1990538579;
assign addr[22690]= 1975871368;
assign addr[22691]= 1960577471;
assign addr[22692]= 1944661739;
assign addr[22693]= 1928129220;
assign addr[22694]= 1910985158;
assign addr[22695]= 1893234990;
assign addr[22696]= 1874884346;
assign addr[22697]= 1855939047;
assign addr[22698]= 1836405100;
assign addr[22699]= 1816288703;
assign addr[22700]= 1795596234;
assign addr[22701]= 1774334257;
assign addr[22702]= 1752509516;
assign addr[22703]= 1730128933;
assign addr[22704]= 1707199606;
assign addr[22705]= 1683728808;
assign addr[22706]= 1659723983;
assign addr[22707]= 1635192744;
assign addr[22708]= 1610142873;
assign addr[22709]= 1584582314;
assign addr[22710]= 1558519173;
assign addr[22711]= 1531961719;
assign addr[22712]= 1504918373;
assign addr[22713]= 1477397714;
assign addr[22714]= 1449408469;
assign addr[22715]= 1420959516;
assign addr[22716]= 1392059879;
assign addr[22717]= 1362718723;
assign addr[22718]= 1332945355;
assign addr[22719]= 1302749217;
assign addr[22720]= 1272139887;
assign addr[22721]= 1241127074;
assign addr[22722]= 1209720613;
assign addr[22723]= 1177930466;
assign addr[22724]= 1145766716;
assign addr[22725]= 1113239564;
assign addr[22726]= 1080359326;
assign addr[22727]= 1047136432;
assign addr[22728]= 1013581418;
assign addr[22729]= 979704927;
assign addr[22730]= 945517704;
assign addr[22731]= 911030591;
assign addr[22732]= 876254528;
assign addr[22733]= 841200544;
assign addr[22734]= 805879757;
assign addr[22735]= 770303369;
assign addr[22736]= 734482665;
assign addr[22737]= 698429006;
assign addr[22738]= 662153826;
assign addr[22739]= 625668632;
assign addr[22740]= 588984994;
assign addr[22741]= 552114549;
assign addr[22742]= 515068990;
assign addr[22743]= 477860067;
assign addr[22744]= 440499581;
assign addr[22745]= 402999383;
assign addr[22746]= 365371365;
assign addr[22747]= 327627463;
assign addr[22748]= 289779648;
assign addr[22749]= 251839923;
assign addr[22750]= 213820322;
assign addr[22751]= 175732905;
assign addr[22752]= 137589750;
assign addr[22753]= 99402956;
assign addr[22754]= 61184634;
assign addr[22755]= 22946906;
assign addr[22756]= -15298099;
assign addr[22757]= -53538253;
assign addr[22758]= -91761426;
assign addr[22759]= -129955495;
assign addr[22760]= -168108346;
assign addr[22761]= -206207878;
assign addr[22762]= -244242007;
assign addr[22763]= -282198671;
assign addr[22764]= -320065829;
assign addr[22765]= -357831473;
assign addr[22766]= -395483624;
assign addr[22767]= -433010339;
assign addr[22768]= -470399716;
assign addr[22769]= -507639898;
assign addr[22770]= -544719071;
assign addr[22771]= -581625477;
assign addr[22772]= -618347408;
assign addr[22773]= -654873219;
assign addr[22774]= -691191324;
assign addr[22775]= -727290205;
assign addr[22776]= -763158411;
assign addr[22777]= -798784567;
assign addr[22778]= -834157373;
assign addr[22779]= -869265610;
assign addr[22780]= -904098143;
assign addr[22781]= -938643924;
assign addr[22782]= -972891995;
assign addr[22783]= -1006831495;
assign addr[22784]= -1040451659;
assign addr[22785]= -1073741824;
assign addr[22786]= -1106691431;
assign addr[22787]= -1139290029;
assign addr[22788]= -1171527280;
assign addr[22789]= -1203392958;
assign addr[22790]= -1234876957;
assign addr[22791]= -1265969291;
assign addr[22792]= -1296660098;
assign addr[22793]= -1326939644;
assign addr[22794]= -1356798326;
assign addr[22795]= -1386226674;
assign addr[22796]= -1415215352;
assign addr[22797]= -1443755168;
assign addr[22798]= -1471837070;
assign addr[22799]= -1499452149;
assign addr[22800]= -1526591649;
assign addr[22801]= -1553246960;
assign addr[22802]= -1579409630;
assign addr[22803]= -1605071359;
assign addr[22804]= -1630224009;
assign addr[22805]= -1654859602;
assign addr[22806]= -1678970324;
assign addr[22807]= -1702548529;
assign addr[22808]= -1725586737;
assign addr[22809]= -1748077642;
assign addr[22810]= -1770014111;
assign addr[22811]= -1791389186;
assign addr[22812]= -1812196087;
assign addr[22813]= -1832428215;
assign addr[22814]= -1852079154;
assign addr[22815]= -1871142669;
assign addr[22816]= -1889612716;
assign addr[22817]= -1907483436;
assign addr[22818]= -1924749160;
assign addr[22819]= -1941404413;
assign addr[22820]= -1957443913;
assign addr[22821]= -1972862571;
assign addr[22822]= -1987655498;
assign addr[22823]= -2001818002;
assign addr[22824]= -2015345591;
assign addr[22825]= -2028233973;
assign addr[22826]= -2040479063;
assign addr[22827]= -2052076975;
assign addr[22828]= -2063024031;
assign addr[22829]= -2073316760;
assign addr[22830]= -2082951896;
assign addr[22831]= -2091926384;
assign addr[22832]= -2100237377;
assign addr[22833]= -2107882239;
assign addr[22834]= -2114858546;
assign addr[22835]= -2121164085;
assign addr[22836]= -2126796855;
assign addr[22837]= -2131755071;
assign addr[22838]= -2136037160;
assign addr[22839]= -2139641764;
assign addr[22840]= -2142567738;
assign addr[22841]= -2144814157;
assign addr[22842]= -2146380306;
assign addr[22843]= -2147265689;
assign addr[22844]= -2147470025;
assign addr[22845]= -2146993250;
assign addr[22846]= -2145835515;
assign addr[22847]= -2143997187;
assign addr[22848]= -2141478848;
assign addr[22849]= -2138281298;
assign addr[22850]= -2134405552;
assign addr[22851]= -2129852837;
assign addr[22852]= -2124624598;
assign addr[22853]= -2118722494;
assign addr[22854]= -2112148396;
assign addr[22855]= -2104904390;
assign addr[22856]= -2096992772;
assign addr[22857]= -2088416053;
assign addr[22858]= -2079176953;
assign addr[22859]= -2069278401;
assign addr[22860]= -2058723538;
assign addr[22861]= -2047515711;
assign addr[22862]= -2035658475;
assign addr[22863]= -2023155591;
assign addr[22864]= -2010011024;
assign addr[22865]= -1996228943;
assign addr[22866]= -1981813720;
assign addr[22867]= -1966769926;
assign addr[22868]= -1951102334;
assign addr[22869]= -1934815911;
assign addr[22870]= -1917915825;
assign addr[22871]= -1900407434;
assign addr[22872]= -1882296293;
assign addr[22873]= -1863588145;
assign addr[22874]= -1844288924;
assign addr[22875]= -1824404752;
assign addr[22876]= -1803941934;
assign addr[22877]= -1782906961;
assign addr[22878]= -1761306505;
assign addr[22879]= -1739147417;
assign addr[22880]= -1716436725;
assign addr[22881]= -1693181631;
assign addr[22882]= -1669389513;
assign addr[22883]= -1645067915;
assign addr[22884]= -1620224553;
assign addr[22885]= -1594867305;
assign addr[22886]= -1569004214;
assign addr[22887]= -1542643483;
assign addr[22888]= -1515793473;
assign addr[22889]= -1488462700;
assign addr[22890]= -1460659832;
assign addr[22891]= -1432393688;
assign addr[22892]= -1403673233;
assign addr[22893]= -1374507575;
assign addr[22894]= -1344905966;
assign addr[22895]= -1314877795;
assign addr[22896]= -1284432584;
assign addr[22897]= -1253579991;
assign addr[22898]= -1222329801;
assign addr[22899]= -1190691925;
assign addr[22900]= -1158676398;
assign addr[22901]= -1126293375;
assign addr[22902]= -1093553126;
assign addr[22903]= -1060466036;
assign addr[22904]= -1027042599;
assign addr[22905]= -993293415;
assign addr[22906]= -959229189;
assign addr[22907]= -924860725;
assign addr[22908]= -890198924;
assign addr[22909]= -855254778;
assign addr[22910]= -820039373;
assign addr[22911]= -784563876;
assign addr[22912]= -748839539;
assign addr[22913]= -712877694;
assign addr[22914]= -676689746;
assign addr[22915]= -640287172;
assign addr[22916]= -603681519;
assign addr[22917]= -566884397;
assign addr[22918]= -529907477;
assign addr[22919]= -492762486;
assign addr[22920]= -455461206;
assign addr[22921]= -418015468;
assign addr[22922]= -380437148;
assign addr[22923]= -342738165;
assign addr[22924]= -304930476;
assign addr[22925]= -267026072;
assign addr[22926]= -229036977;
assign addr[22927]= -190975237;
assign addr[22928]= -152852926;
assign addr[22929]= -114682135;
assign addr[22930]= -76474970;
assign addr[22931]= -38243550;
assign addr[22932]= 0;
assign addr[22933]= 38243550;
assign addr[22934]= 76474970;
assign addr[22935]= 114682135;
assign addr[22936]= 152852926;
assign addr[22937]= 190975237;
assign addr[22938]= 229036977;
assign addr[22939]= 267026072;
assign addr[22940]= 304930476;
assign addr[22941]= 342738165;
assign addr[22942]= 380437148;
assign addr[22943]= 418015468;
assign addr[22944]= 455461206;
assign addr[22945]= 492762486;
assign addr[22946]= 529907477;
assign addr[22947]= 566884397;
assign addr[22948]= 603681519;
assign addr[22949]= 640287172;
assign addr[22950]= 676689746;
assign addr[22951]= 712877694;
assign addr[22952]= 748839539;
assign addr[22953]= 784563876;
assign addr[22954]= 820039373;
assign addr[22955]= 855254778;
assign addr[22956]= 890198924;
assign addr[22957]= 924860725;
assign addr[22958]= 959229189;
assign addr[22959]= 993293415;
assign addr[22960]= 1027042599;
assign addr[22961]= 1060466036;
assign addr[22962]= 1093553126;
assign addr[22963]= 1126293375;
assign addr[22964]= 1158676398;
assign addr[22965]= 1190691925;
assign addr[22966]= 1222329801;
assign addr[22967]= 1253579991;
assign addr[22968]= 1284432584;
assign addr[22969]= 1314877795;
assign addr[22970]= 1344905966;
assign addr[22971]= 1374507575;
assign addr[22972]= 1403673233;
assign addr[22973]= 1432393688;
assign addr[22974]= 1460659832;
assign addr[22975]= 1488462700;
assign addr[22976]= 1515793473;
assign addr[22977]= 1542643483;
assign addr[22978]= 1569004214;
assign addr[22979]= 1594867305;
assign addr[22980]= 1620224553;
assign addr[22981]= 1645067915;
assign addr[22982]= 1669389513;
assign addr[22983]= 1693181631;
assign addr[22984]= 1716436725;
assign addr[22985]= 1739147417;
assign addr[22986]= 1761306505;
assign addr[22987]= 1782906961;
assign addr[22988]= 1803941934;
assign addr[22989]= 1824404752;
assign addr[22990]= 1844288924;
assign addr[22991]= 1863588145;
assign addr[22992]= 1882296293;
assign addr[22993]= 1900407434;
assign addr[22994]= 1917915825;
assign addr[22995]= 1934815911;
assign addr[22996]= 1951102334;
assign addr[22997]= 1966769926;
assign addr[22998]= 1981813720;
assign addr[22999]= 1996228943;
assign addr[23000]= 2010011024;
assign addr[23001]= 2023155591;
assign addr[23002]= 2035658475;
assign addr[23003]= 2047515711;
assign addr[23004]= 2058723538;
assign addr[23005]= 2069278401;
assign addr[23006]= 2079176953;
assign addr[23007]= 2088416053;
assign addr[23008]= 2096992772;
assign addr[23009]= 2104904390;
assign addr[23010]= 2112148396;
assign addr[23011]= 2118722494;
assign addr[23012]= 2124624598;
assign addr[23013]= 2129852837;
assign addr[23014]= 2134405552;
assign addr[23015]= 2138281298;
assign addr[23016]= 2141478848;
assign addr[23017]= 2143997187;
assign addr[23018]= 2145835515;
assign addr[23019]= 2146993250;
assign addr[23020]= 2147470025;
assign addr[23021]= 2147265689;
assign addr[23022]= 2146380306;
assign addr[23023]= 2144814157;
assign addr[23024]= 2142567738;
assign addr[23025]= 2139641764;
assign addr[23026]= 2136037160;
assign addr[23027]= 2131755071;
assign addr[23028]= 2126796855;
assign addr[23029]= 2121164085;
assign addr[23030]= 2114858546;
assign addr[23031]= 2107882239;
assign addr[23032]= 2100237377;
assign addr[23033]= 2091926384;
assign addr[23034]= 2082951896;
assign addr[23035]= 2073316760;
assign addr[23036]= 2063024031;
assign addr[23037]= 2052076975;
assign addr[23038]= 2040479063;
assign addr[23039]= 2028233973;
assign addr[23040]= 2015345591;
assign addr[23041]= 2001818002;
assign addr[23042]= 1987655498;
assign addr[23043]= 1972862571;
assign addr[23044]= 1957443913;
assign addr[23045]= 1941404413;
assign addr[23046]= 1924749160;
assign addr[23047]= 1907483436;
assign addr[23048]= 1889612716;
assign addr[23049]= 1871142669;
assign addr[23050]= 1852079154;
assign addr[23051]= 1832428215;
assign addr[23052]= 1812196087;
assign addr[23053]= 1791389186;
assign addr[23054]= 1770014111;
assign addr[23055]= 1748077642;
assign addr[23056]= 1725586737;
assign addr[23057]= 1702548529;
assign addr[23058]= 1678970324;
assign addr[23059]= 1654859602;
assign addr[23060]= 1630224009;
assign addr[23061]= 1605071359;
assign addr[23062]= 1579409630;
assign addr[23063]= 1553246960;
assign addr[23064]= 1526591649;
assign addr[23065]= 1499452149;
assign addr[23066]= 1471837070;
assign addr[23067]= 1443755168;
assign addr[23068]= 1415215352;
assign addr[23069]= 1386226674;
assign addr[23070]= 1356798326;
assign addr[23071]= 1326939644;
assign addr[23072]= 1296660098;
assign addr[23073]= 1265969291;
assign addr[23074]= 1234876957;
assign addr[23075]= 1203392958;
assign addr[23076]= 1171527280;
assign addr[23077]= 1139290029;
assign addr[23078]= 1106691431;
assign addr[23079]= 1073741824;
assign addr[23080]= 1040451659;
assign addr[23081]= 1006831495;
assign addr[23082]= 972891995;
assign addr[23083]= 938643924;
assign addr[23084]= 904098143;
assign addr[23085]= 869265610;
assign addr[23086]= 834157373;
assign addr[23087]= 798784567;
assign addr[23088]= 763158411;
assign addr[23089]= 727290205;
assign addr[23090]= 691191324;
assign addr[23091]= 654873219;
assign addr[23092]= 618347408;
assign addr[23093]= 581625477;
assign addr[23094]= 544719071;
assign addr[23095]= 507639898;
assign addr[23096]= 470399716;
assign addr[23097]= 433010339;
assign addr[23098]= 395483624;
assign addr[23099]= 357831473;
assign addr[23100]= 320065829;
assign addr[23101]= 282198671;
assign addr[23102]= 244242007;
assign addr[23103]= 206207878;
assign addr[23104]= 168108346;
assign addr[23105]= 129955495;
assign addr[23106]= 91761426;
assign addr[23107]= 53538253;
assign addr[23108]= 15298099;
assign addr[23109]= -22946906;
assign addr[23110]= -61184634;
assign addr[23111]= -99402956;
assign addr[23112]= -137589750;
assign addr[23113]= -175732905;
assign addr[23114]= -213820322;
assign addr[23115]= -251839923;
assign addr[23116]= -289779648;
assign addr[23117]= -327627463;
assign addr[23118]= -365371365;
assign addr[23119]= -402999383;
assign addr[23120]= -440499581;
assign addr[23121]= -477860067;
assign addr[23122]= -515068990;
assign addr[23123]= -552114549;
assign addr[23124]= -588984994;
assign addr[23125]= -625668632;
assign addr[23126]= -662153826;
assign addr[23127]= -698429006;
assign addr[23128]= -734482665;
assign addr[23129]= -770303369;
assign addr[23130]= -805879757;
assign addr[23131]= -841200544;
assign addr[23132]= -876254528;
assign addr[23133]= -911030591;
assign addr[23134]= -945517704;
assign addr[23135]= -979704927;
assign addr[23136]= -1013581418;
assign addr[23137]= -1047136432;
assign addr[23138]= -1080359326;
assign addr[23139]= -1113239564;
assign addr[23140]= -1145766716;
assign addr[23141]= -1177930466;
assign addr[23142]= -1209720613;
assign addr[23143]= -1241127074;
assign addr[23144]= -1272139887;
assign addr[23145]= -1302749217;
assign addr[23146]= -1332945355;
assign addr[23147]= -1362718723;
assign addr[23148]= -1392059879;
assign addr[23149]= -1420959516;
assign addr[23150]= -1449408469;
assign addr[23151]= -1477397714;
assign addr[23152]= -1504918373;
assign addr[23153]= -1531961719;
assign addr[23154]= -1558519173;
assign addr[23155]= -1584582314;
assign addr[23156]= -1610142873;
assign addr[23157]= -1635192744;
assign addr[23158]= -1659723983;
assign addr[23159]= -1683728808;
assign addr[23160]= -1707199606;
assign addr[23161]= -1730128933;
assign addr[23162]= -1752509516;
assign addr[23163]= -1774334257;
assign addr[23164]= -1795596234;
assign addr[23165]= -1816288703;
assign addr[23166]= -1836405100;
assign addr[23167]= -1855939047;
assign addr[23168]= -1874884346;
assign addr[23169]= -1893234990;
assign addr[23170]= -1910985158;
assign addr[23171]= -1928129220;
assign addr[23172]= -1944661739;
assign addr[23173]= -1960577471;
assign addr[23174]= -1975871368;
assign addr[23175]= -1990538579;
assign addr[23176]= -2004574453;
assign addr[23177]= -2017974537;
assign addr[23178]= -2030734582;
assign addr[23179]= -2042850540;
assign addr[23180]= -2054318569;
assign addr[23181]= -2065135031;
assign addr[23182]= -2075296495;
assign addr[23183]= -2084799740;
assign addr[23184]= -2093641749;
assign addr[23185]= -2101819720;
assign addr[23186]= -2109331059;
assign addr[23187]= -2116173382;
assign addr[23188]= -2122344521;
assign addr[23189]= -2127842516;
assign addr[23190]= -2132665626;
assign addr[23191]= -2136812319;
assign addr[23192]= -2140281282;
assign addr[23193]= -2143071413;
assign addr[23194]= -2145181827;
assign addr[23195]= -2146611856;
assign addr[23196]= -2147361045;
assign addr[23197]= -2147429158;
assign addr[23198]= -2146816171;
assign addr[23199]= -2145522281;
assign addr[23200]= -2143547897;
assign addr[23201]= -2140893646;
assign addr[23202]= -2137560369;
assign addr[23203]= -2133549123;
assign addr[23204]= -2128861181;
assign addr[23205]= -2123498030;
assign addr[23206]= -2117461370;
assign addr[23207]= -2110753117;
assign addr[23208]= -2103375398;
assign addr[23209]= -2095330553;
assign addr[23210]= -2086621133;
assign addr[23211]= -2077249901;
assign addr[23212]= -2067219829;
assign addr[23213]= -2056534099;
assign addr[23214]= -2045196100;
assign addr[23215]= -2033209426;
assign addr[23216]= -2020577882;
assign addr[23217]= -2007305472;
assign addr[23218]= -1993396407;
assign addr[23219]= -1978855097;
assign addr[23220]= -1963686155;
assign addr[23221]= -1947894393;
assign addr[23222]= -1931484818;
assign addr[23223]= -1914462636;
assign addr[23224]= -1896833245;
assign addr[23225]= -1878602237;
assign addr[23226]= -1859775393;
assign addr[23227]= -1840358687;
assign addr[23228]= -1820358275;
assign addr[23229]= -1799780501;
assign addr[23230]= -1778631892;
assign addr[23231]= -1756919156;
assign addr[23232]= -1734649179;
assign addr[23233]= -1711829025;
assign addr[23234]= -1688465931;
assign addr[23235]= -1664567307;
assign addr[23236]= -1640140734;
assign addr[23237]= -1615193959;
assign addr[23238]= -1589734894;
assign addr[23239]= -1563771613;
assign addr[23240]= -1537312353;
assign addr[23241]= -1510365504;
assign addr[23242]= -1482939614;
assign addr[23243]= -1455043381;
assign addr[23244]= -1426685652;
assign addr[23245]= -1397875423;
assign addr[23246]= -1368621831;
assign addr[23247]= -1338934154;
assign addr[23248]= -1308821808;
assign addr[23249]= -1278294345;
assign addr[23250]= -1247361445;
assign addr[23251]= -1216032921;
assign addr[23252]= -1184318708;
assign addr[23253]= -1152228866;
assign addr[23254]= -1119773573;
assign addr[23255]= -1086963121;
assign addr[23256]= -1053807919;
assign addr[23257]= -1020318481;
assign addr[23258]= -986505429;
assign addr[23259]= -952379488;
assign addr[23260]= -917951481;
assign addr[23261]= -883232329;
assign addr[23262]= -848233042;
assign addr[23263]= -812964722;
assign addr[23264]= -777438554;
assign addr[23265]= -741665807;
assign addr[23266]= -705657826;
assign addr[23267]= -669426032;
assign addr[23268]= -632981917;
assign addr[23269]= -596337040;
assign addr[23270]= -559503022;
assign addr[23271]= -522491548;
assign addr[23272]= -485314355;
assign addr[23273]= -447983235;
assign addr[23274]= -410510029;
assign addr[23275]= -372906622;
assign addr[23276]= -335184940;
assign addr[23277]= -297356948;
assign addr[23278]= -259434643;
assign addr[23279]= -221430054;
assign addr[23280]= -183355234;
assign addr[23281]= -145222259;
assign addr[23282]= -107043224;
assign addr[23283]= -68830239;
assign addr[23284]= -30595422;
assign addr[23285]= 7649098;
assign addr[23286]= 45891193;
assign addr[23287]= 84118732;
assign addr[23288]= 122319591;
assign addr[23289]= 160481654;
assign addr[23290]= 198592817;
assign addr[23291]= 236640993;
assign addr[23292]= 274614114;
assign addr[23293]= 312500135;
assign addr[23294]= 350287041;
assign addr[23295]= 387962847;
assign addr[23296]= 425515602;
assign addr[23297]= 462933398;
assign addr[23298]= 500204365;
assign addr[23299]= 537316682;
assign addr[23300]= 574258580;
assign addr[23301]= 611018340;
assign addr[23302]= 647584304;
assign addr[23303]= 683944874;
assign addr[23304]= 720088517;
assign addr[23305]= 756003771;
assign addr[23306]= 791679244;
assign addr[23307]= 827103620;
assign addr[23308]= 862265664;
assign addr[23309]= 897154224;
assign addr[23310]= 931758235;
assign addr[23311]= 966066720;
assign addr[23312]= 1000068799;
assign addr[23313]= 1033753687;
assign addr[23314]= 1067110699;
assign addr[23315]= 1100129257;
assign addr[23316]= 1132798888;
assign addr[23317]= 1165109230;
assign addr[23318]= 1197050035;
assign addr[23319]= 1228611172;
assign addr[23320]= 1259782632;
assign addr[23321]= 1290554528;
assign addr[23322]= 1320917099;
assign addr[23323]= 1350860716;
assign addr[23324]= 1380375881;
assign addr[23325]= 1409453233;
assign addr[23326]= 1438083551;
assign addr[23327]= 1466257752;
assign addr[23328]= 1493966902;
assign addr[23329]= 1521202211;
assign addr[23330]= 1547955041;
assign addr[23331]= 1574216908;
assign addr[23332]= 1599979481;
assign addr[23333]= 1625234591;
assign addr[23334]= 1649974225;
assign addr[23335]= 1674190539;
assign addr[23336]= 1697875851;
assign addr[23337]= 1721022648;
assign addr[23338]= 1743623590;
assign addr[23339]= 1765671509;
assign addr[23340]= 1787159411;
assign addr[23341]= 1808080480;
assign addr[23342]= 1828428082;
assign addr[23343]= 1848195763;
assign addr[23344]= 1867377253;
assign addr[23345]= 1885966468;
assign addr[23346]= 1903957513;
assign addr[23347]= 1921344681;
assign addr[23348]= 1938122457;
assign addr[23349]= 1954285520;
assign addr[23350]= 1969828744;
assign addr[23351]= 1984747199;
assign addr[23352]= 1999036154;
assign addr[23353]= 2012691075;
assign addr[23354]= 2025707632;
assign addr[23355]= 2038081698;
assign addr[23356]= 2049809346;
assign addr[23357]= 2060886858;
assign addr[23358]= 2071310720;
assign addr[23359]= 2081077626;
assign addr[23360]= 2090184478;
assign addr[23361]= 2098628387;
assign addr[23362]= 2106406677;
assign addr[23363]= 2113516878;
assign addr[23364]= 2119956737;
assign addr[23365]= 2125724211;
assign addr[23366]= 2130817471;
assign addr[23367]= 2135234901;
assign addr[23368]= 2138975100;
assign addr[23369]= 2142036881;
assign addr[23370]= 2144419275;
assign addr[23371]= 2146121524;
assign addr[23372]= 2147143090;
assign addr[23373]= 2147483648;
assign addr[23374]= 2147143090;
assign addr[23375]= 2146121524;
assign addr[23376]= 2144419275;
assign addr[23377]= 2142036881;
assign addr[23378]= 2138975100;
assign addr[23379]= 2135234901;
assign addr[23380]= 2130817471;
assign addr[23381]= 2125724211;
assign addr[23382]= 2119956737;
assign addr[23383]= 2113516878;
assign addr[23384]= 2106406677;
assign addr[23385]= 2098628387;
assign addr[23386]= 2090184478;
assign addr[23387]= 2081077626;
assign addr[23388]= 2071310720;
assign addr[23389]= 2060886858;
assign addr[23390]= 2049809346;
assign addr[23391]= 2038081698;
assign addr[23392]= 2025707632;
assign addr[23393]= 2012691075;
assign addr[23394]= 1999036154;
assign addr[23395]= 1984747199;
assign addr[23396]= 1969828744;
assign addr[23397]= 1954285520;
assign addr[23398]= 1938122457;
assign addr[23399]= 1921344681;
assign addr[23400]= 1903957513;
assign addr[23401]= 1885966468;
assign addr[23402]= 1867377253;
assign addr[23403]= 1848195763;
assign addr[23404]= 1828428082;
assign addr[23405]= 1808080480;
assign addr[23406]= 1787159411;
assign addr[23407]= 1765671509;
assign addr[23408]= 1743623590;
assign addr[23409]= 1721022648;
assign addr[23410]= 1697875851;
assign addr[23411]= 1674190539;
assign addr[23412]= 1649974225;
assign addr[23413]= 1625234591;
assign addr[23414]= 1599979481;
assign addr[23415]= 1574216908;
assign addr[23416]= 1547955041;
assign addr[23417]= 1521202211;
assign addr[23418]= 1493966902;
assign addr[23419]= 1466257752;
assign addr[23420]= 1438083551;
assign addr[23421]= 1409453233;
assign addr[23422]= 1380375881;
assign addr[23423]= 1350860716;
assign addr[23424]= 1320917099;
assign addr[23425]= 1290554528;
assign addr[23426]= 1259782632;
assign addr[23427]= 1228611172;
assign addr[23428]= 1197050035;
assign addr[23429]= 1165109230;
assign addr[23430]= 1132798888;
assign addr[23431]= 1100129257;
assign addr[23432]= 1067110699;
assign addr[23433]= 1033753687;
assign addr[23434]= 1000068799;
assign addr[23435]= 966066720;
assign addr[23436]= 931758235;
assign addr[23437]= 897154224;
assign addr[23438]= 862265664;
assign addr[23439]= 827103620;
assign addr[23440]= 791679244;
assign addr[23441]= 756003771;
assign addr[23442]= 720088517;
assign addr[23443]= 683944874;
assign addr[23444]= 647584304;
assign addr[23445]= 611018340;
assign addr[23446]= 574258580;
assign addr[23447]= 537316682;
assign addr[23448]= 500204365;
assign addr[23449]= 462933398;
assign addr[23450]= 425515602;
assign addr[23451]= 387962847;
assign addr[23452]= 350287041;
assign addr[23453]= 312500135;
assign addr[23454]= 274614114;
assign addr[23455]= 236640993;
assign addr[23456]= 198592817;
assign addr[23457]= 160481654;
assign addr[23458]= 122319591;
assign addr[23459]= 84118732;
assign addr[23460]= 45891193;
assign addr[23461]= 7649098;
assign addr[23462]= -30595422;
assign addr[23463]= -68830239;
assign addr[23464]= -107043224;
assign addr[23465]= -145222259;
assign addr[23466]= -183355234;
assign addr[23467]= -221430054;
assign addr[23468]= -259434643;
assign addr[23469]= -297356948;
assign addr[23470]= -335184940;
assign addr[23471]= -372906622;
assign addr[23472]= -410510029;
assign addr[23473]= -447983235;
assign addr[23474]= -485314355;
assign addr[23475]= -522491548;
assign addr[23476]= -559503022;
assign addr[23477]= -596337040;
assign addr[23478]= -632981917;
assign addr[23479]= -669426032;
assign addr[23480]= -705657826;
assign addr[23481]= -741665807;
assign addr[23482]= -777438554;
assign addr[23483]= -812964722;
assign addr[23484]= -848233042;
assign addr[23485]= -883232329;
assign addr[23486]= -917951481;
assign addr[23487]= -952379488;
assign addr[23488]= -986505429;
assign addr[23489]= -1020318481;
assign addr[23490]= -1053807919;
assign addr[23491]= -1086963121;
assign addr[23492]= -1119773573;
assign addr[23493]= -1152228866;
assign addr[23494]= -1184318708;
assign addr[23495]= -1216032921;
assign addr[23496]= -1247361445;
assign addr[23497]= -1278294345;
assign addr[23498]= -1308821808;
assign addr[23499]= -1338934154;
assign addr[23500]= -1368621831;
assign addr[23501]= -1397875423;
assign addr[23502]= -1426685652;
assign addr[23503]= -1455043381;
assign addr[23504]= -1482939614;
assign addr[23505]= -1510365504;
assign addr[23506]= -1537312353;
assign addr[23507]= -1563771613;
assign addr[23508]= -1589734894;
assign addr[23509]= -1615193959;
assign addr[23510]= -1640140734;
assign addr[23511]= -1664567307;
assign addr[23512]= -1688465931;
assign addr[23513]= -1711829025;
assign addr[23514]= -1734649179;
assign addr[23515]= -1756919156;
assign addr[23516]= -1778631892;
assign addr[23517]= -1799780501;
assign addr[23518]= -1820358275;
assign addr[23519]= -1840358687;
assign addr[23520]= -1859775393;
assign addr[23521]= -1878602237;
assign addr[23522]= -1896833245;
assign addr[23523]= -1914462636;
assign addr[23524]= -1931484818;
assign addr[23525]= -1947894393;
assign addr[23526]= -1963686155;
assign addr[23527]= -1978855097;
assign addr[23528]= -1993396407;
assign addr[23529]= -2007305472;
assign addr[23530]= -2020577882;
assign addr[23531]= -2033209426;
assign addr[23532]= -2045196100;
assign addr[23533]= -2056534099;
assign addr[23534]= -2067219829;
assign addr[23535]= -2077249901;
assign addr[23536]= -2086621133;
assign addr[23537]= -2095330553;
assign addr[23538]= -2103375398;
assign addr[23539]= -2110753117;
assign addr[23540]= -2117461370;
assign addr[23541]= -2123498030;
assign addr[23542]= -2128861181;
assign addr[23543]= -2133549123;
assign addr[23544]= -2137560369;
assign addr[23545]= -2140893646;
assign addr[23546]= -2143547897;
assign addr[23547]= -2145522281;
assign addr[23548]= -2146816171;
assign addr[23549]= -2147429158;
assign addr[23550]= -2147361045;
assign addr[23551]= -2146611856;
assign addr[23552]= -2145181827;
assign addr[23553]= -2143071413;
assign addr[23554]= -2140281282;
assign addr[23555]= -2136812319;
assign addr[23556]= -2132665626;
assign addr[23557]= -2127842516;
assign addr[23558]= -2122344521;
assign addr[23559]= -2116173382;
assign addr[23560]= -2109331059;
assign addr[23561]= -2101819720;
assign addr[23562]= -2093641749;
assign addr[23563]= -2084799740;
assign addr[23564]= -2075296495;
assign addr[23565]= -2065135031;
assign addr[23566]= -2054318569;
assign addr[23567]= -2042850540;
assign addr[23568]= -2030734582;
assign addr[23569]= -2017974537;
assign addr[23570]= -2004574453;
assign addr[23571]= -1990538579;
assign addr[23572]= -1975871368;
assign addr[23573]= -1960577471;
assign addr[23574]= -1944661739;
assign addr[23575]= -1928129220;
assign addr[23576]= -1910985158;
assign addr[23577]= -1893234990;
assign addr[23578]= -1874884346;
assign addr[23579]= -1855939047;
assign addr[23580]= -1836405100;
assign addr[23581]= -1816288703;
assign addr[23582]= -1795596234;
assign addr[23583]= -1774334257;
assign addr[23584]= -1752509516;
assign addr[23585]= -1730128933;
assign addr[23586]= -1707199606;
assign addr[23587]= -1683728808;
assign addr[23588]= -1659723983;
assign addr[23589]= -1635192744;
assign addr[23590]= -1610142873;
assign addr[23591]= -1584582314;
assign addr[23592]= -1558519173;
assign addr[23593]= -1531961719;
assign addr[23594]= -1504918373;
assign addr[23595]= -1477397714;
assign addr[23596]= -1449408469;
assign addr[23597]= -1420959516;
assign addr[23598]= -1392059879;
assign addr[23599]= -1362718723;
assign addr[23600]= -1332945355;
assign addr[23601]= -1302749217;
assign addr[23602]= -1272139887;
assign addr[23603]= -1241127074;
assign addr[23604]= -1209720613;
assign addr[23605]= -1177930466;
assign addr[23606]= -1145766716;
assign addr[23607]= -1113239564;
assign addr[23608]= -1080359326;
assign addr[23609]= -1047136432;
assign addr[23610]= -1013581418;
assign addr[23611]= -979704927;
assign addr[23612]= -945517704;
assign addr[23613]= -911030591;
assign addr[23614]= -876254528;
assign addr[23615]= -841200544;
assign addr[23616]= -805879757;
assign addr[23617]= -770303369;
assign addr[23618]= -734482665;
assign addr[23619]= -698429006;
assign addr[23620]= -662153826;
assign addr[23621]= -625668632;
assign addr[23622]= -588984994;
assign addr[23623]= -552114549;
assign addr[23624]= -515068990;
assign addr[23625]= -477860067;
assign addr[23626]= -440499581;
assign addr[23627]= -402999383;
assign addr[23628]= -365371365;
assign addr[23629]= -327627463;
assign addr[23630]= -289779648;
assign addr[23631]= -251839923;
assign addr[23632]= -213820322;
assign addr[23633]= -175732905;
assign addr[23634]= -137589750;
assign addr[23635]= -99402956;
assign addr[23636]= -61184634;
assign addr[23637]= -22946906;
assign addr[23638]= 15298099;
assign addr[23639]= 53538253;
assign addr[23640]= 91761426;
assign addr[23641]= 129955495;
assign addr[23642]= 168108346;
assign addr[23643]= 206207878;
assign addr[23644]= 244242007;
assign addr[23645]= 282198671;
assign addr[23646]= 320065829;
assign addr[23647]= 357831473;
assign addr[23648]= 395483624;
assign addr[23649]= 433010339;
assign addr[23650]= 470399716;
assign addr[23651]= 507639898;
assign addr[23652]= 544719071;
assign addr[23653]= 581625477;
assign addr[23654]= 618347408;
assign addr[23655]= 654873219;
assign addr[23656]= 691191324;
assign addr[23657]= 727290205;
assign addr[23658]= 763158411;
assign addr[23659]= 798784567;
assign addr[23660]= 834157373;
assign addr[23661]= 869265610;
assign addr[23662]= 904098143;
assign addr[23663]= 938643924;
assign addr[23664]= 972891995;
assign addr[23665]= 1006831495;
assign addr[23666]= 1040451659;
assign addr[23667]= 1073741824;
assign addr[23668]= 1106691431;
assign addr[23669]= 1139290029;
assign addr[23670]= 1171527280;
assign addr[23671]= 1203392958;
assign addr[23672]= 1234876957;
assign addr[23673]= 1265969291;
assign addr[23674]= 1296660098;
assign addr[23675]= 1326939644;
assign addr[23676]= 1356798326;
assign addr[23677]= 1386226674;
assign addr[23678]= 1415215352;
assign addr[23679]= 1443755168;
assign addr[23680]= 1471837070;
assign addr[23681]= 1499452149;
assign addr[23682]= 1526591649;
assign addr[23683]= 1553246960;
assign addr[23684]= 1579409630;
assign addr[23685]= 1605071359;
assign addr[23686]= 1630224009;
assign addr[23687]= 1654859602;
assign addr[23688]= 1678970324;
assign addr[23689]= 1702548529;
assign addr[23690]= 1725586737;
assign addr[23691]= 1748077642;
assign addr[23692]= 1770014111;
assign addr[23693]= 1791389186;
assign addr[23694]= 1812196087;
assign addr[23695]= 1832428215;
assign addr[23696]= 1852079154;
assign addr[23697]= 1871142669;
assign addr[23698]= 1889612716;
assign addr[23699]= 1907483436;
assign addr[23700]= 1924749160;
assign addr[23701]= 1941404413;
assign addr[23702]= 1957443913;
assign addr[23703]= 1972862571;
assign addr[23704]= 1987655498;
assign addr[23705]= 2001818002;
assign addr[23706]= 2015345591;
assign addr[23707]= 2028233973;
assign addr[23708]= 2040479063;
assign addr[23709]= 2052076975;
assign addr[23710]= 2063024031;
assign addr[23711]= 2073316760;
assign addr[23712]= 2082951896;
assign addr[23713]= 2091926384;
assign addr[23714]= 2100237377;
assign addr[23715]= 2107882239;
assign addr[23716]= 2114858546;
assign addr[23717]= 2121164085;
assign addr[23718]= 2126796855;
assign addr[23719]= 2131755071;
assign addr[23720]= 2136037160;
assign addr[23721]= 2139641764;
assign addr[23722]= 2142567738;
assign addr[23723]= 2144814157;
assign addr[23724]= 2146380306;
assign addr[23725]= 2147265689;
assign addr[23726]= 2147470025;
assign addr[23727]= 2146993250;
assign addr[23728]= 2145835515;
assign addr[23729]= 2143997187;
assign addr[23730]= 2141478848;
assign addr[23731]= 2138281298;
assign addr[23732]= 2134405552;
assign addr[23733]= 2129852837;
assign addr[23734]= 2124624598;
assign addr[23735]= 2118722494;
assign addr[23736]= 2112148396;
assign addr[23737]= 2104904390;
assign addr[23738]= 2096992772;
assign addr[23739]= 2088416053;
assign addr[23740]= 2079176953;
assign addr[23741]= 2069278401;
assign addr[23742]= 2058723538;
assign addr[23743]= 2047515711;
assign addr[23744]= 2035658475;
assign addr[23745]= 2023155591;
assign addr[23746]= 2010011024;
assign addr[23747]= 1996228943;
assign addr[23748]= 1981813720;
assign addr[23749]= 1966769926;
assign addr[23750]= 1951102334;
assign addr[23751]= 1934815911;
assign addr[23752]= 1917915825;
assign addr[23753]= 1900407434;
assign addr[23754]= 1882296293;
assign addr[23755]= 1863588145;
assign addr[23756]= 1844288924;
assign addr[23757]= 1824404752;
assign addr[23758]= 1803941934;
assign addr[23759]= 1782906961;
assign addr[23760]= 1761306505;
assign addr[23761]= 1739147417;
assign addr[23762]= 1716436725;
assign addr[23763]= 1693181631;
assign addr[23764]= 1669389513;
assign addr[23765]= 1645067915;
assign addr[23766]= 1620224553;
assign addr[23767]= 1594867305;
assign addr[23768]= 1569004214;
assign addr[23769]= 1542643483;
assign addr[23770]= 1515793473;
assign addr[23771]= 1488462700;
assign addr[23772]= 1460659832;
assign addr[23773]= 1432393688;
assign addr[23774]= 1403673233;
assign addr[23775]= 1374507575;
assign addr[23776]= 1344905966;
assign addr[23777]= 1314877795;
assign addr[23778]= 1284432584;
assign addr[23779]= 1253579991;
assign addr[23780]= 1222329801;
assign addr[23781]= 1190691925;
assign addr[23782]= 1158676398;
assign addr[23783]= 1126293375;
assign addr[23784]= 1093553126;
assign addr[23785]= 1060466036;
assign addr[23786]= 1027042599;
assign addr[23787]= 993293415;
assign addr[23788]= 959229189;
assign addr[23789]= 924860725;
assign addr[23790]= 890198924;
assign addr[23791]= 855254778;
assign addr[23792]= 820039373;
assign addr[23793]= 784563876;
assign addr[23794]= 748839539;
assign addr[23795]= 712877694;
assign addr[23796]= 676689746;
assign addr[23797]= 640287172;
assign addr[23798]= 603681519;
assign addr[23799]= 566884397;
assign addr[23800]= 529907477;
assign addr[23801]= 492762486;
assign addr[23802]= 455461206;
assign addr[23803]= 418015468;
assign addr[23804]= 380437148;
assign addr[23805]= 342738165;
assign addr[23806]= 304930476;
assign addr[23807]= 267026072;
assign addr[23808]= 229036977;
assign addr[23809]= 190975237;
assign addr[23810]= 152852926;
assign addr[23811]= 114682135;
assign addr[23812]= 76474970;
assign addr[23813]= 38243550;
assign addr[23814]= 0;
assign addr[23815]= -38243550;
assign addr[23816]= -76474970;
assign addr[23817]= -114682135;
assign addr[23818]= -152852926;
assign addr[23819]= -190975237;
assign addr[23820]= -229036977;
assign addr[23821]= -267026072;
assign addr[23822]= -304930476;
assign addr[23823]= -342738165;
assign addr[23824]= -380437148;
assign addr[23825]= -418015468;
assign addr[23826]= -455461206;
assign addr[23827]= -492762486;
assign addr[23828]= -529907477;
assign addr[23829]= -566884397;
assign addr[23830]= -603681519;
assign addr[23831]= -640287172;
assign addr[23832]= -676689746;
assign addr[23833]= -712877694;
assign addr[23834]= -748839539;
assign addr[23835]= -784563876;
assign addr[23836]= -820039373;
assign addr[23837]= -855254778;
assign addr[23838]= -890198924;
assign addr[23839]= -924860725;
assign addr[23840]= -959229189;
assign addr[23841]= -993293415;
assign addr[23842]= -1027042599;
assign addr[23843]= -1060466036;
assign addr[23844]= -1093553126;
assign addr[23845]= -1126293375;
assign addr[23846]= -1158676398;
assign addr[23847]= -1190691925;
assign addr[23848]= -1222329801;
assign addr[23849]= -1253579991;
assign addr[23850]= -1284432584;
assign addr[23851]= -1314877795;
assign addr[23852]= -1344905966;
assign addr[23853]= -1374507575;
assign addr[23854]= -1403673233;
assign addr[23855]= -1432393688;
assign addr[23856]= -1460659832;
assign addr[23857]= -1488462700;
assign addr[23858]= -1515793473;
assign addr[23859]= -1542643483;
assign addr[23860]= -1569004214;
assign addr[23861]= -1594867305;
assign addr[23862]= -1620224553;
assign addr[23863]= -1645067915;
assign addr[23864]= -1669389513;
assign addr[23865]= -1693181631;
assign addr[23866]= -1716436725;
assign addr[23867]= -1739147417;
assign addr[23868]= -1761306505;
assign addr[23869]= -1782906961;
assign addr[23870]= -1803941934;
assign addr[23871]= -1824404752;
assign addr[23872]= -1844288924;
assign addr[23873]= -1863588145;
assign addr[23874]= -1882296293;
assign addr[23875]= -1900407434;
assign addr[23876]= -1917915825;
assign addr[23877]= -1934815911;
assign addr[23878]= -1951102334;
assign addr[23879]= -1966769926;
assign addr[23880]= -1981813720;
assign addr[23881]= -1996228943;
assign addr[23882]= -2010011024;
assign addr[23883]= -2023155591;
assign addr[23884]= -2035658475;
assign addr[23885]= -2047515711;
assign addr[23886]= -2058723538;
assign addr[23887]= -2069278401;
assign addr[23888]= -2079176953;
assign addr[23889]= -2088416053;
assign addr[23890]= -2096992772;
assign addr[23891]= -2104904390;
assign addr[23892]= -2112148396;
assign addr[23893]= -2118722494;
assign addr[23894]= -2124624598;
assign addr[23895]= -2129852837;
assign addr[23896]= -2134405552;
assign addr[23897]= -2138281298;
assign addr[23898]= -2141478848;
assign addr[23899]= -2143997187;
assign addr[23900]= -2145835515;
assign addr[23901]= -2146993250;
assign addr[23902]= -2147470025;
assign addr[23903]= -2147265689;
assign addr[23904]= -2146380306;
assign addr[23905]= -2144814157;
assign addr[23906]= -2142567738;
assign addr[23907]= -2139641764;
assign addr[23908]= -2136037160;
assign addr[23909]= -2131755071;
assign addr[23910]= -2126796855;
assign addr[23911]= -2121164085;
assign addr[23912]= -2114858546;
assign addr[23913]= -2107882239;
assign addr[23914]= -2100237377;
assign addr[23915]= -2091926384;
assign addr[23916]= -2082951896;
assign addr[23917]= -2073316760;
assign addr[23918]= -2063024031;
assign addr[23919]= -2052076975;
assign addr[23920]= -2040479063;
assign addr[23921]= -2028233973;
assign addr[23922]= -2015345591;
assign addr[23923]= -2001818002;
assign addr[23924]= -1987655498;
assign addr[23925]= -1972862571;
assign addr[23926]= -1957443913;
assign addr[23927]= -1941404413;
assign addr[23928]= -1924749160;
assign addr[23929]= -1907483436;
assign addr[23930]= -1889612716;
assign addr[23931]= -1871142669;
assign addr[23932]= -1852079154;
assign addr[23933]= -1832428215;
assign addr[23934]= -1812196087;
assign addr[23935]= -1791389186;
assign addr[23936]= -1770014111;
assign addr[23937]= -1748077642;
assign addr[23938]= -1725586737;
assign addr[23939]= -1702548529;
assign addr[23940]= -1678970324;
assign addr[23941]= -1654859602;
assign addr[23942]= -1630224009;
assign addr[23943]= -1605071359;
assign addr[23944]= -1579409630;
assign addr[23945]= -1553246960;
assign addr[23946]= -1526591649;
assign addr[23947]= -1499452149;
assign addr[23948]= -1471837070;
assign addr[23949]= -1443755168;
assign addr[23950]= -1415215352;
assign addr[23951]= -1386226674;
assign addr[23952]= -1356798326;
assign addr[23953]= -1326939644;
assign addr[23954]= -1296660098;
assign addr[23955]= -1265969291;
assign addr[23956]= -1234876957;
assign addr[23957]= -1203392958;
assign addr[23958]= -1171527280;
assign addr[23959]= -1139290029;
assign addr[23960]= -1106691431;
assign addr[23961]= -1073741824;
assign addr[23962]= -1040451659;
assign addr[23963]= -1006831495;
assign addr[23964]= -972891995;
assign addr[23965]= -938643924;
assign addr[23966]= -904098143;
assign addr[23967]= -869265610;
assign addr[23968]= -834157373;
assign addr[23969]= -798784567;
assign addr[23970]= -763158411;
assign addr[23971]= -727290205;
assign addr[23972]= -691191324;
assign addr[23973]= -654873219;
assign addr[23974]= -618347408;
assign addr[23975]= -581625477;
assign addr[23976]= -544719071;
assign addr[23977]= -507639898;
assign addr[23978]= -470399716;
assign addr[23979]= -433010339;
assign addr[23980]= -395483624;
assign addr[23981]= -357831473;
assign addr[23982]= -320065829;
assign addr[23983]= -282198671;
assign addr[23984]= -244242007;
assign addr[23985]= -206207878;
assign addr[23986]= -168108346;
assign addr[23987]= -129955495;
assign addr[23988]= -91761426;
assign addr[23989]= -53538253;
assign addr[23990]= -15298099;
assign addr[23991]= 22946906;
assign addr[23992]= 61184634;
assign addr[23993]= 99402956;
assign addr[23994]= 137589750;
assign addr[23995]= 175732905;
assign addr[23996]= 213820322;
assign addr[23997]= 251839923;
assign addr[23998]= 289779648;
assign addr[23999]= 327627463;
assign addr[24000]= 365371365;
assign addr[24001]= 402999383;
assign addr[24002]= 440499581;
assign addr[24003]= 477860067;
assign addr[24004]= 515068990;
assign addr[24005]= 552114549;
assign addr[24006]= 588984994;
assign addr[24007]= 625668632;
assign addr[24008]= 662153826;
assign addr[24009]= 698429006;
assign addr[24010]= 734482665;
assign addr[24011]= 770303369;
assign addr[24012]= 805879757;
assign addr[24013]= 841200544;
assign addr[24014]= 876254528;
assign addr[24015]= 911030591;
assign addr[24016]= 945517704;
assign addr[24017]= 979704927;
assign addr[24018]= 1013581418;
assign addr[24019]= 1047136432;
assign addr[24020]= 1080359326;
assign addr[24021]= 1113239564;
assign addr[24022]= 1145766716;
assign addr[24023]= 1177930466;
assign addr[24024]= 1209720613;
assign addr[24025]= 1241127074;
assign addr[24026]= 1272139887;
assign addr[24027]= 1302749217;
assign addr[24028]= 1332945355;
assign addr[24029]= 1362718723;
assign addr[24030]= 1392059879;
assign addr[24031]= 1420959516;
assign addr[24032]= 1449408469;
assign addr[24033]= 1477397714;
assign addr[24034]= 1504918373;
assign addr[24035]= 1531961719;
assign addr[24036]= 1558519173;
assign addr[24037]= 1584582314;
assign addr[24038]= 1610142873;
assign addr[24039]= 1635192744;
assign addr[24040]= 1659723983;
assign addr[24041]= 1683728808;
assign addr[24042]= 1707199606;
assign addr[24043]= 1730128933;
assign addr[24044]= 1752509516;
assign addr[24045]= 1774334257;
assign addr[24046]= 1795596234;
assign addr[24047]= 1816288703;
assign addr[24048]= 1836405100;
assign addr[24049]= 1855939047;
assign addr[24050]= 1874884346;
assign addr[24051]= 1893234990;
assign addr[24052]= 1910985158;
assign addr[24053]= 1928129220;
assign addr[24054]= 1944661739;
assign addr[24055]= 1960577471;
assign addr[24056]= 1975871368;
assign addr[24057]= 1990538579;
assign addr[24058]= 2004574453;
assign addr[24059]= 2017974537;
assign addr[24060]= 2030734582;
assign addr[24061]= 2042850540;
assign addr[24062]= 2054318569;
assign addr[24063]= 2065135031;
assign addr[24064]= 2075296495;
assign addr[24065]= 2084799740;
assign addr[24066]= 2093641749;
assign addr[24067]= 2101819720;
assign addr[24068]= 2109331059;
assign addr[24069]= 2116173382;
assign addr[24070]= 2122344521;
assign addr[24071]= 2127842516;
assign addr[24072]= 2132665626;
assign addr[24073]= 2136812319;
assign addr[24074]= 2140281282;
assign addr[24075]= 2143071413;
assign addr[24076]= 2145181827;
assign addr[24077]= 2146611856;
assign addr[24078]= 2147361045;
assign addr[24079]= 2147429158;
assign addr[24080]= 2146816171;
assign addr[24081]= 2145522281;
assign addr[24082]= 2143547897;
assign addr[24083]= 2140893646;
assign addr[24084]= 2137560369;
assign addr[24085]= 2133549123;
assign addr[24086]= 2128861181;
assign addr[24087]= 2123498030;
assign addr[24088]= 2117461370;
assign addr[24089]= 2110753117;
assign addr[24090]= 2103375398;
assign addr[24091]= 2095330553;
assign addr[24092]= 2086621133;
assign addr[24093]= 2077249901;
assign addr[24094]= 2067219829;
assign addr[24095]= 2056534099;
assign addr[24096]= 2045196100;
assign addr[24097]= 2033209426;
assign addr[24098]= 2020577882;
assign addr[24099]= 2007305472;
assign addr[24100]= 1993396407;
assign addr[24101]= 1978855097;
assign addr[24102]= 1963686155;
assign addr[24103]= 1947894393;
assign addr[24104]= 1931484818;
assign addr[24105]= 1914462636;
assign addr[24106]= 1896833245;
assign addr[24107]= 1878602237;
assign addr[24108]= 1859775393;
assign addr[24109]= 1840358687;
assign addr[24110]= 1820358275;
assign addr[24111]= 1799780501;
assign addr[24112]= 1778631892;
assign addr[24113]= 1756919156;
assign addr[24114]= 1734649179;
assign addr[24115]= 1711829025;
assign addr[24116]= 1688465931;
assign addr[24117]= 1664567307;
assign addr[24118]= 1640140734;
assign addr[24119]= 1615193959;
assign addr[24120]= 1589734894;
assign addr[24121]= 1563771613;
assign addr[24122]= 1537312353;
assign addr[24123]= 1510365504;
assign addr[24124]= 1482939614;
assign addr[24125]= 1455043381;
assign addr[24126]= 1426685652;
assign addr[24127]= 1397875423;
assign addr[24128]= 1368621831;
assign addr[24129]= 1338934154;
assign addr[24130]= 1308821808;
assign addr[24131]= 1278294345;
assign addr[24132]= 1247361445;
assign addr[24133]= 1216032921;
assign addr[24134]= 1184318708;
assign addr[24135]= 1152228866;
assign addr[24136]= 1119773573;
assign addr[24137]= 1086963121;
assign addr[24138]= 1053807919;
assign addr[24139]= 1020318481;
assign addr[24140]= 986505429;
assign addr[24141]= 952379488;
assign addr[24142]= 917951481;
assign addr[24143]= 883232329;
assign addr[24144]= 848233042;
assign addr[24145]= 812964722;
assign addr[24146]= 777438554;
assign addr[24147]= 741665807;
assign addr[24148]= 705657826;
assign addr[24149]= 669426032;
assign addr[24150]= 632981917;
assign addr[24151]= 596337040;
assign addr[24152]= 559503022;
assign addr[24153]= 522491548;
assign addr[24154]= 485314355;
assign addr[24155]= 447983235;
assign addr[24156]= 410510029;
assign addr[24157]= 372906622;
assign addr[24158]= 335184940;
assign addr[24159]= 297356948;
assign addr[24160]= 259434643;
assign addr[24161]= 221430054;
assign addr[24162]= 183355234;
assign addr[24163]= 145222259;
assign addr[24164]= 107043224;
assign addr[24165]= 68830239;
assign addr[24166]= 30595422;
assign addr[24167]= -7649098;
assign addr[24168]= -45891193;
assign addr[24169]= -84118732;
assign addr[24170]= -122319591;
assign addr[24171]= -160481654;
assign addr[24172]= -198592817;
assign addr[24173]= -236640993;
assign addr[24174]= -274614114;
assign addr[24175]= -312500135;
assign addr[24176]= -350287041;
assign addr[24177]= -387962847;
assign addr[24178]= -425515602;
assign addr[24179]= -462933398;
assign addr[24180]= -500204365;
assign addr[24181]= -537316682;
assign addr[24182]= -574258580;
assign addr[24183]= -611018340;
assign addr[24184]= -647584304;
assign addr[24185]= -683944874;
assign addr[24186]= -720088517;
assign addr[24187]= -756003771;
assign addr[24188]= -791679244;
assign addr[24189]= -827103620;
assign addr[24190]= -862265664;
assign addr[24191]= -897154224;
assign addr[24192]= -931758235;
assign addr[24193]= -966066720;
assign addr[24194]= -1000068799;
assign addr[24195]= -1033753687;
assign addr[24196]= -1067110699;
assign addr[24197]= -1100129257;
assign addr[24198]= -1132798888;
assign addr[24199]= -1165109230;
assign addr[24200]= -1197050035;
assign addr[24201]= -1228611172;
assign addr[24202]= -1259782632;
assign addr[24203]= -1290554528;
assign addr[24204]= -1320917099;
assign addr[24205]= -1350860716;
assign addr[24206]= -1380375881;
assign addr[24207]= -1409453233;
assign addr[24208]= -1438083551;
assign addr[24209]= -1466257752;
assign addr[24210]= -1493966902;
assign addr[24211]= -1521202211;
assign addr[24212]= -1547955041;
assign addr[24213]= -1574216908;
assign addr[24214]= -1599979481;
assign addr[24215]= -1625234591;
assign addr[24216]= -1649974225;
assign addr[24217]= -1674190539;
assign addr[24218]= -1697875851;
assign addr[24219]= -1721022648;
assign addr[24220]= -1743623590;
assign addr[24221]= -1765671509;
assign addr[24222]= -1787159411;
assign addr[24223]= -1808080480;
assign addr[24224]= -1828428082;
assign addr[24225]= -1848195763;
assign addr[24226]= -1867377253;
assign addr[24227]= -1885966468;
assign addr[24228]= -1903957513;
assign addr[24229]= -1921344681;
assign addr[24230]= -1938122457;
assign addr[24231]= -1954285520;
assign addr[24232]= -1969828744;
assign addr[24233]= -1984747199;
assign addr[24234]= -1999036154;
assign addr[24235]= -2012691075;
assign addr[24236]= -2025707632;
assign addr[24237]= -2038081698;
assign addr[24238]= -2049809346;
assign addr[24239]= -2060886858;
assign addr[24240]= -2071310720;
assign addr[24241]= -2081077626;
assign addr[24242]= -2090184478;
assign addr[24243]= -2098628387;
assign addr[24244]= -2106406677;
assign addr[24245]= -2113516878;
assign addr[24246]= -2119956737;
assign addr[24247]= -2125724211;
assign addr[24248]= -2130817471;
assign addr[24249]= -2135234901;
assign addr[24250]= -2138975100;
assign addr[24251]= -2142036881;
assign addr[24252]= -2144419275;
assign addr[24253]= -2146121524;
assign addr[24254]= -2147143090;
assign addr[24255]= -2147483648;
assign addr[24256]= -2147143090;
assign addr[24257]= -2146121524;
assign addr[24258]= -2144419275;
assign addr[24259]= -2142036881;
assign addr[24260]= -2138975100;
assign addr[24261]= -2135234901;
assign addr[24262]= -2130817471;
assign addr[24263]= -2125724211;
assign addr[24264]= -2119956737;
assign addr[24265]= -2113516878;
assign addr[24266]= -2106406677;
assign addr[24267]= -2098628387;
assign addr[24268]= -2090184478;
assign addr[24269]= -2081077626;
assign addr[24270]= -2071310720;
assign addr[24271]= -2060886858;
assign addr[24272]= -2049809346;
assign addr[24273]= -2038081698;
assign addr[24274]= -2025707632;
assign addr[24275]= -2012691075;
assign addr[24276]= -1999036154;
assign addr[24277]= -1984747199;
assign addr[24278]= -1969828744;
assign addr[24279]= -1954285520;
assign addr[24280]= -1938122457;
assign addr[24281]= -1921344681;
assign addr[24282]= -1903957513;
assign addr[24283]= -1885966468;
assign addr[24284]= -1867377253;
assign addr[24285]= -1848195763;
assign addr[24286]= -1828428082;
assign addr[24287]= -1808080480;
assign addr[24288]= -1787159411;
assign addr[24289]= -1765671509;
assign addr[24290]= -1743623590;
assign addr[24291]= -1721022648;
assign addr[24292]= -1697875851;
assign addr[24293]= -1674190539;
assign addr[24294]= -1649974225;
assign addr[24295]= -1625234591;
assign addr[24296]= -1599979481;
assign addr[24297]= -1574216908;
assign addr[24298]= -1547955041;
assign addr[24299]= -1521202211;
assign addr[24300]= -1493966902;
assign addr[24301]= -1466257752;
assign addr[24302]= -1438083551;
assign addr[24303]= -1409453233;
assign addr[24304]= -1380375881;
assign addr[24305]= -1350860716;
assign addr[24306]= -1320917099;
assign addr[24307]= -1290554528;
assign addr[24308]= -1259782632;
assign addr[24309]= -1228611172;
assign addr[24310]= -1197050035;
assign addr[24311]= -1165109230;
assign addr[24312]= -1132798888;
assign addr[24313]= -1100129257;
assign addr[24314]= -1067110699;
assign addr[24315]= -1033753687;
assign addr[24316]= -1000068799;
assign addr[24317]= -966066720;
assign addr[24318]= -931758235;
assign addr[24319]= -897154224;
assign addr[24320]= -862265664;
assign addr[24321]= -827103620;
assign addr[24322]= -791679244;
assign addr[24323]= -756003771;
assign addr[24324]= -720088517;
assign addr[24325]= -683944874;
assign addr[24326]= -647584304;
assign addr[24327]= -611018340;
assign addr[24328]= -574258580;
assign addr[24329]= -537316682;
assign addr[24330]= -500204365;
assign addr[24331]= -462933398;
assign addr[24332]= -425515602;
assign addr[24333]= -387962847;
assign addr[24334]= -350287041;
assign addr[24335]= -312500135;
assign addr[24336]= -274614114;
assign addr[24337]= -236640993;
assign addr[24338]= -198592817;
assign addr[24339]= -160481654;
assign addr[24340]= -122319591;
assign addr[24341]= -84118732;
assign addr[24342]= -45891193;
assign addr[24343]= -7649098;
assign addr[24344]= 30595422;
assign addr[24345]= 68830239;
assign addr[24346]= 107043224;
assign addr[24347]= 145222259;
assign addr[24348]= 183355234;
assign addr[24349]= 221430054;
assign addr[24350]= 259434643;
assign addr[24351]= 297356948;
assign addr[24352]= 335184940;
assign addr[24353]= 372906622;
assign addr[24354]= 410510029;
assign addr[24355]= 447983235;
assign addr[24356]= 485314355;
assign addr[24357]= 522491548;
assign addr[24358]= 559503022;
assign addr[24359]= 596337040;
assign addr[24360]= 632981917;
assign addr[24361]= 669426032;
assign addr[24362]= 705657826;
assign addr[24363]= 741665807;
assign addr[24364]= 777438554;
assign addr[24365]= 812964722;
assign addr[24366]= 848233042;
assign addr[24367]= 883232329;
assign addr[24368]= 917951481;
assign addr[24369]= 952379488;
assign addr[24370]= 986505429;
assign addr[24371]= 1020318481;
assign addr[24372]= 1053807919;
assign addr[24373]= 1086963121;
assign addr[24374]= 1119773573;
assign addr[24375]= 1152228866;
assign addr[24376]= 1184318708;
assign addr[24377]= 1216032921;
assign addr[24378]= 1247361445;
assign addr[24379]= 1278294345;
assign addr[24380]= 1308821808;
assign addr[24381]= 1338934154;
assign addr[24382]= 1368621831;
assign addr[24383]= 1397875423;
assign addr[24384]= 1426685652;
assign addr[24385]= 1455043381;
assign addr[24386]= 1482939614;
assign addr[24387]= 1510365504;
assign addr[24388]= 1537312353;
assign addr[24389]= 1563771613;
assign addr[24390]= 1589734894;
assign addr[24391]= 1615193959;
assign addr[24392]= 1640140734;
assign addr[24393]= 1664567307;
assign addr[24394]= 1688465931;
assign addr[24395]= 1711829025;
assign addr[24396]= 1734649179;
assign addr[24397]= 1756919156;
assign addr[24398]= 1778631892;
assign addr[24399]= 1799780501;
assign addr[24400]= 1820358275;
assign addr[24401]= 1840358687;
assign addr[24402]= 1859775393;
assign addr[24403]= 1878602237;
assign addr[24404]= 1896833245;
assign addr[24405]= 1914462636;
assign addr[24406]= 1931484818;
assign addr[24407]= 1947894393;
assign addr[24408]= 1963686155;
assign addr[24409]= 1978855097;
assign addr[24410]= 1993396407;
assign addr[24411]= 2007305472;
assign addr[24412]= 2020577882;
assign addr[24413]= 2033209426;
assign addr[24414]= 2045196100;
assign addr[24415]= 2056534099;
assign addr[24416]= 2067219829;
assign addr[24417]= 2077249901;
assign addr[24418]= 2086621133;
assign addr[24419]= 2095330553;
assign addr[24420]= 2103375398;
assign addr[24421]= 2110753117;
assign addr[24422]= 2117461370;
assign addr[24423]= 2123498030;
assign addr[24424]= 2128861181;
assign addr[24425]= 2133549123;
assign addr[24426]= 2137560369;
assign addr[24427]= 2140893646;
assign addr[24428]= 2143547897;
assign addr[24429]= 2145522281;
assign addr[24430]= 2146816171;
assign addr[24431]= 2147429158;
assign addr[24432]= 2147361045;
assign addr[24433]= 2146611856;
assign addr[24434]= 2145181827;
assign addr[24435]= 2143071413;
assign addr[24436]= 2140281282;
assign addr[24437]= 2136812319;
assign addr[24438]= 2132665626;
assign addr[24439]= 2127842516;
assign addr[24440]= 2122344521;
assign addr[24441]= 2116173382;
assign addr[24442]= 2109331059;
assign addr[24443]= 2101819720;
assign addr[24444]= 2093641749;
assign addr[24445]= 2084799740;
assign addr[24446]= 2075296495;
assign addr[24447]= 2065135031;
assign addr[24448]= 2054318569;
assign addr[24449]= 2042850540;
assign addr[24450]= 2030734582;
assign addr[24451]= 2017974537;
assign addr[24452]= 2004574453;
assign addr[24453]= 1990538579;
assign addr[24454]= 1975871368;
assign addr[24455]= 1960577471;
assign addr[24456]= 1944661739;
assign addr[24457]= 1928129220;
assign addr[24458]= 1910985158;
assign addr[24459]= 1893234990;
assign addr[24460]= 1874884346;
assign addr[24461]= 1855939047;
assign addr[24462]= 1836405100;
assign addr[24463]= 1816288703;
assign addr[24464]= 1795596234;
assign addr[24465]= 1774334257;
assign addr[24466]= 1752509516;
assign addr[24467]= 1730128933;
assign addr[24468]= 1707199606;
assign addr[24469]= 1683728808;
assign addr[24470]= 1659723983;
assign addr[24471]= 1635192744;
assign addr[24472]= 1610142873;
assign addr[24473]= 1584582314;
assign addr[24474]= 1558519173;
assign addr[24475]= 1531961719;
assign addr[24476]= 1504918373;
assign addr[24477]= 1477397714;
assign addr[24478]= 1449408469;
assign addr[24479]= 1420959516;
assign addr[24480]= 1392059879;
assign addr[24481]= 1362718723;
assign addr[24482]= 1332945355;
assign addr[24483]= 1302749217;
assign addr[24484]= 1272139887;
assign addr[24485]= 1241127074;
assign addr[24486]= 1209720613;
assign addr[24487]= 1177930466;
assign addr[24488]= 1145766716;
assign addr[24489]= 1113239564;
assign addr[24490]= 1080359326;
assign addr[24491]= 1047136432;
assign addr[24492]= 1013581418;
assign addr[24493]= 979704927;
assign addr[24494]= 945517704;
assign addr[24495]= 911030591;
assign addr[24496]= 876254528;
assign addr[24497]= 841200544;
assign addr[24498]= 805879757;
assign addr[24499]= 770303369;
assign addr[24500]= 734482665;
assign addr[24501]= 698429006;
assign addr[24502]= 662153826;
assign addr[24503]= 625668632;
assign addr[24504]= 588984994;
assign addr[24505]= 552114549;
assign addr[24506]= 515068990;
assign addr[24507]= 477860067;
assign addr[24508]= 440499581;
assign addr[24509]= 402999383;
assign addr[24510]= 365371365;
assign addr[24511]= 327627463;
assign addr[24512]= 289779648;
assign addr[24513]= 251839923;
assign addr[24514]= 213820322;
assign addr[24515]= 175732905;
assign addr[24516]= 137589750;
assign addr[24517]= 99402956;
assign addr[24518]= 61184634;
assign addr[24519]= 22946906;
assign addr[24520]= -15298099;
assign addr[24521]= -53538253;
assign addr[24522]= -91761426;
assign addr[24523]= -129955495;
assign addr[24524]= -168108346;
assign addr[24525]= -206207878;
assign addr[24526]= -244242007;
assign addr[24527]= -282198671;
assign addr[24528]= -320065829;
assign addr[24529]= -357831473;
assign addr[24530]= -395483624;
assign addr[24531]= -433010339;
assign addr[24532]= -470399716;
assign addr[24533]= -507639898;
assign addr[24534]= -544719071;
assign addr[24535]= -581625477;
assign addr[24536]= -618347408;
assign addr[24537]= -654873219;
assign addr[24538]= -691191324;
assign addr[24539]= -727290205;
assign addr[24540]= -763158411;
assign addr[24541]= -798784567;
assign addr[24542]= -834157373;
assign addr[24543]= -869265610;
assign addr[24544]= -904098143;
assign addr[24545]= -938643924;
assign addr[24546]= -972891995;
assign addr[24547]= -1006831495;
assign addr[24548]= -1040451659;
assign addr[24549]= -1073741824;
assign addr[24550]= -1106691431;
assign addr[24551]= -1139290029;
assign addr[24552]= -1171527280;
assign addr[24553]= -1203392958;
assign addr[24554]= -1234876957;
assign addr[24555]= -1265969291;
assign addr[24556]= -1296660098;
assign addr[24557]= -1326939644;
assign addr[24558]= -1356798326;
assign addr[24559]= -1386226674;
assign addr[24560]= -1415215352;
assign addr[24561]= -1443755168;
assign addr[24562]= -1471837070;
assign addr[24563]= -1499452149;
assign addr[24564]= -1526591649;
assign addr[24565]= -1553246960;
assign addr[24566]= -1579409630;
assign addr[24567]= -1605071359;
assign addr[24568]= -1630224009;
assign addr[24569]= -1654859602;
assign addr[24570]= -1678970324;
assign addr[24571]= -1702548529;
assign addr[24572]= -1725586737;
assign addr[24573]= -1748077642;
assign addr[24574]= -1770014111;
assign addr[24575]= -1791389186;
assign addr[24576]= -1812196087;
assign addr[24577]= -1832428215;
assign addr[24578]= -1852079154;
assign addr[24579]= -1871142669;
assign addr[24580]= -1889612716;
assign addr[24581]= -1907483436;
assign addr[24582]= -1924749160;
assign addr[24583]= -1941404413;
assign addr[24584]= -1957443913;
assign addr[24585]= -1972862571;
assign addr[24586]= -1987655498;
assign addr[24587]= -2001818002;
assign addr[24588]= -2015345591;
assign addr[24589]= -2028233973;
assign addr[24590]= -2040479063;
assign addr[24591]= -2052076975;
assign addr[24592]= -2063024031;
assign addr[24593]= -2073316760;
assign addr[24594]= -2082951896;
assign addr[24595]= -2091926384;
assign addr[24596]= -2100237377;
assign addr[24597]= -2107882239;
assign addr[24598]= -2114858546;
assign addr[24599]= -2121164085;
assign addr[24600]= -2126796855;
assign addr[24601]= -2131755071;
assign addr[24602]= -2136037160;
assign addr[24603]= -2139641764;
assign addr[24604]= -2142567738;
assign addr[24605]= -2144814157;
assign addr[24606]= -2146380306;
assign addr[24607]= -2147265689;
assign addr[24608]= -2147470025;
assign addr[24609]= -2146993250;
assign addr[24610]= -2145835515;
assign addr[24611]= -2143997187;
assign addr[24612]= -2141478848;
assign addr[24613]= -2138281298;
assign addr[24614]= -2134405552;
assign addr[24615]= -2129852837;
assign addr[24616]= -2124624598;
assign addr[24617]= -2118722494;
assign addr[24618]= -2112148396;
assign addr[24619]= -2104904390;
assign addr[24620]= -2096992772;
assign addr[24621]= -2088416053;
assign addr[24622]= -2079176953;
assign addr[24623]= -2069278401;
assign addr[24624]= -2058723538;
assign addr[24625]= -2047515711;
assign addr[24626]= -2035658475;
assign addr[24627]= -2023155591;
assign addr[24628]= -2010011024;
assign addr[24629]= -1996228943;
assign addr[24630]= -1981813720;
assign addr[24631]= -1966769926;
assign addr[24632]= -1951102334;
assign addr[24633]= -1934815911;
assign addr[24634]= -1917915825;
assign addr[24635]= -1900407434;
assign addr[24636]= -1882296293;
assign addr[24637]= -1863588145;
assign addr[24638]= -1844288924;
assign addr[24639]= -1824404752;
assign addr[24640]= -1803941934;
assign addr[24641]= -1782906961;
assign addr[24642]= -1761306505;
assign addr[24643]= -1739147417;
assign addr[24644]= -1716436725;
assign addr[24645]= -1693181631;
assign addr[24646]= -1669389513;
assign addr[24647]= -1645067915;
assign addr[24648]= -1620224553;
assign addr[24649]= -1594867305;
assign addr[24650]= -1569004214;
assign addr[24651]= -1542643483;
assign addr[24652]= -1515793473;
assign addr[24653]= -1488462700;
assign addr[24654]= -1460659832;
assign addr[24655]= -1432393688;
assign addr[24656]= -1403673233;
assign addr[24657]= -1374507575;
assign addr[24658]= -1344905966;
assign addr[24659]= -1314877795;
assign addr[24660]= -1284432584;
assign addr[24661]= -1253579991;
assign addr[24662]= -1222329801;
assign addr[24663]= -1190691925;
assign addr[24664]= -1158676398;
assign addr[24665]= -1126293375;
assign addr[24666]= -1093553126;
assign addr[24667]= -1060466036;
assign addr[24668]= -1027042599;
assign addr[24669]= -993293415;
assign addr[24670]= -959229189;
assign addr[24671]= -924860725;
assign addr[24672]= -890198924;
assign addr[24673]= -855254778;
assign addr[24674]= -820039373;
assign addr[24675]= -784563876;
assign addr[24676]= -748839539;
assign addr[24677]= -712877694;
assign addr[24678]= -676689746;
assign addr[24679]= -640287172;
assign addr[24680]= -603681519;
assign addr[24681]= -566884397;
assign addr[24682]= -529907477;
assign addr[24683]= -492762486;
assign addr[24684]= -455461206;
assign addr[24685]= -418015468;
assign addr[24686]= -380437148;
assign addr[24687]= -342738165;
assign addr[24688]= -304930476;
assign addr[24689]= -267026072;
assign addr[24690]= -229036977;
assign addr[24691]= -190975237;
assign addr[24692]= -152852926;
assign addr[24693]= -114682135;
assign addr[24694]= -76474970;
assign addr[24695]= -38243550;
assign addr[24696]= 0;
assign addr[24697]= 38243550;
assign addr[24698]= 76474970;
assign addr[24699]= 114682135;
assign addr[24700]= 152852926;
assign addr[24701]= 190975237;
assign addr[24702]= 229036977;
assign addr[24703]= 267026072;
assign addr[24704]= 304930476;
assign addr[24705]= 342738165;
assign addr[24706]= 380437148;
assign addr[24707]= 418015468;
assign addr[24708]= 455461206;
assign addr[24709]= 492762486;
assign addr[24710]= 529907477;
assign addr[24711]= 566884397;
assign addr[24712]= 603681519;
assign addr[24713]= 640287172;
assign addr[24714]= 676689746;
assign addr[24715]= 712877694;
assign addr[24716]= 748839539;
assign addr[24717]= 784563876;
assign addr[24718]= 820039373;
assign addr[24719]= 855254778;
assign addr[24720]= 890198924;
assign addr[24721]= 924860725;
assign addr[24722]= 959229189;
assign addr[24723]= 993293415;
assign addr[24724]= 1027042599;
assign addr[24725]= 1060466036;
assign addr[24726]= 1093553126;
assign addr[24727]= 1126293375;
assign addr[24728]= 1158676398;
assign addr[24729]= 1190691925;
assign addr[24730]= 1222329801;
assign addr[24731]= 1253579991;
assign addr[24732]= 1284432584;
assign addr[24733]= 1314877795;
assign addr[24734]= 1344905966;
assign addr[24735]= 1374507575;
assign addr[24736]= 1403673233;
assign addr[24737]= 1432393688;
assign addr[24738]= 1460659832;
assign addr[24739]= 1488462700;
assign addr[24740]= 1515793473;
assign addr[24741]= 1542643483;
assign addr[24742]= 1569004214;
assign addr[24743]= 1594867305;
assign addr[24744]= 1620224553;
assign addr[24745]= 1645067915;
assign addr[24746]= 1669389513;
assign addr[24747]= 1693181631;
assign addr[24748]= 1716436725;
assign addr[24749]= 1739147417;
assign addr[24750]= 1761306505;
assign addr[24751]= 1782906961;
assign addr[24752]= 1803941934;
assign addr[24753]= 1824404752;
assign addr[24754]= 1844288924;
assign addr[24755]= 1863588145;
assign addr[24756]= 1882296293;
assign addr[24757]= 1900407434;
assign addr[24758]= 1917915825;
assign addr[24759]= 1934815911;
assign addr[24760]= 1951102334;
assign addr[24761]= 1966769926;
assign addr[24762]= 1981813720;
assign addr[24763]= 1996228943;
assign addr[24764]= 2010011024;
assign addr[24765]= 2023155591;
assign addr[24766]= 2035658475;
assign addr[24767]= 2047515711;
assign addr[24768]= 2058723538;
assign addr[24769]= 2069278401;
assign addr[24770]= 2079176953;
assign addr[24771]= 2088416053;
assign addr[24772]= 2096992772;
assign addr[24773]= 2104904390;
assign addr[24774]= 2112148396;
assign addr[24775]= 2118722494;
assign addr[24776]= 2124624598;
assign addr[24777]= 2129852837;
assign addr[24778]= 2134405552;
assign addr[24779]= 2138281298;
assign addr[24780]= 2141478848;
assign addr[24781]= 2143997187;
assign addr[24782]= 2145835515;
assign addr[24783]= 2146993250;
assign addr[24784]= 2147470025;
assign addr[24785]= 2147265689;
assign addr[24786]= 2146380306;
assign addr[24787]= 2144814157;
assign addr[24788]= 2142567738;
assign addr[24789]= 2139641764;
assign addr[24790]= 2136037160;
assign addr[24791]= 2131755071;
assign addr[24792]= 2126796855;
assign addr[24793]= 2121164085;
assign addr[24794]= 2114858546;
assign addr[24795]= 2107882239;
assign addr[24796]= 2100237377;
assign addr[24797]= 2091926384;
assign addr[24798]= 2082951896;
assign addr[24799]= 2073316760;
assign addr[24800]= 2063024031;
assign addr[24801]= 2052076975;
assign addr[24802]= 2040479063;
assign addr[24803]= 2028233973;
assign addr[24804]= 2015345591;
assign addr[24805]= 2001818002;
assign addr[24806]= 1987655498;
assign addr[24807]= 1972862571;
assign addr[24808]= 1957443913;
assign addr[24809]= 1941404413;
assign addr[24810]= 1924749160;
assign addr[24811]= 1907483436;
assign addr[24812]= 1889612716;
assign addr[24813]= 1871142669;
assign addr[24814]= 1852079154;
assign addr[24815]= 1832428215;
assign addr[24816]= 1812196087;
assign addr[24817]= 1791389186;
assign addr[24818]= 1770014111;
assign addr[24819]= 1748077642;
assign addr[24820]= 1725586737;
assign addr[24821]= 1702548529;
assign addr[24822]= 1678970324;
assign addr[24823]= 1654859602;
assign addr[24824]= 1630224009;
assign addr[24825]= 1605071359;
assign addr[24826]= 1579409630;
assign addr[24827]= 1553246960;
assign addr[24828]= 1526591649;
assign addr[24829]= 1499452149;
assign addr[24830]= 1471837070;
assign addr[24831]= 1443755168;
assign addr[24832]= 1415215352;
assign addr[24833]= 1386226674;
assign addr[24834]= 1356798326;
assign addr[24835]= 1326939644;
assign addr[24836]= 1296660098;
assign addr[24837]= 1265969291;
assign addr[24838]= 1234876957;
assign addr[24839]= 1203392958;
assign addr[24840]= 1171527280;
assign addr[24841]= 1139290029;
assign addr[24842]= 1106691431;
assign addr[24843]= 1073741824;
assign addr[24844]= 1040451659;
assign addr[24845]= 1006831495;
assign addr[24846]= 972891995;
assign addr[24847]= 938643924;
assign addr[24848]= 904098143;
assign addr[24849]= 869265610;
assign addr[24850]= 834157373;
assign addr[24851]= 798784567;
assign addr[24852]= 763158411;
assign addr[24853]= 727290205;
assign addr[24854]= 691191324;
assign addr[24855]= 654873219;
assign addr[24856]= 618347408;
assign addr[24857]= 581625477;
assign addr[24858]= 544719071;
assign addr[24859]= 507639898;
assign addr[24860]= 470399716;
assign addr[24861]= 433010339;
assign addr[24862]= 395483624;
assign addr[24863]= 357831473;
assign addr[24864]= 320065829;
assign addr[24865]= 282198671;
assign addr[24866]= 244242007;
assign addr[24867]= 206207878;
assign addr[24868]= 168108346;
assign addr[24869]= 129955495;
assign addr[24870]= 91761426;
assign addr[24871]= 53538253;
assign addr[24872]= 15298099;
assign addr[24873]= -22946906;
assign addr[24874]= -61184634;
assign addr[24875]= -99402956;
assign addr[24876]= -137589750;
assign addr[24877]= -175732905;
assign addr[24878]= -213820322;
assign addr[24879]= -251839923;
assign addr[24880]= -289779648;
assign addr[24881]= -327627463;
assign addr[24882]= -365371365;
assign addr[24883]= -402999383;
assign addr[24884]= -440499581;
assign addr[24885]= -477860067;
assign addr[24886]= -515068990;
assign addr[24887]= -552114549;
assign addr[24888]= -588984994;
assign addr[24889]= -625668632;
assign addr[24890]= -662153826;
assign addr[24891]= -698429006;
assign addr[24892]= -734482665;
assign addr[24893]= -770303369;
assign addr[24894]= -805879757;
assign addr[24895]= -841200544;
assign addr[24896]= -876254528;
assign addr[24897]= -911030591;
assign addr[24898]= -945517704;
assign addr[24899]= -979704927;
assign addr[24900]= -1013581418;
assign addr[24901]= -1047136432;
assign addr[24902]= -1080359326;
assign addr[24903]= -1113239564;
assign addr[24904]= -1145766716;
assign addr[24905]= -1177930466;
assign addr[24906]= -1209720613;
assign addr[24907]= -1241127074;
assign addr[24908]= -1272139887;
assign addr[24909]= -1302749217;
assign addr[24910]= -1332945355;
assign addr[24911]= -1362718723;
assign addr[24912]= -1392059879;
assign addr[24913]= -1420959516;
assign addr[24914]= -1449408469;
assign addr[24915]= -1477397714;
assign addr[24916]= -1504918373;
assign addr[24917]= -1531961719;
assign addr[24918]= -1558519173;
assign addr[24919]= -1584582314;
assign addr[24920]= -1610142873;
assign addr[24921]= -1635192744;
assign addr[24922]= -1659723983;
assign addr[24923]= -1683728808;
assign addr[24924]= -1707199606;
assign addr[24925]= -1730128933;
assign addr[24926]= -1752509516;
assign addr[24927]= -1774334257;
assign addr[24928]= -1795596234;
assign addr[24929]= -1816288703;
assign addr[24930]= -1836405100;
assign addr[24931]= -1855939047;
assign addr[24932]= -1874884346;
assign addr[24933]= -1893234990;
assign addr[24934]= -1910985158;
assign addr[24935]= -1928129220;
assign addr[24936]= -1944661739;
assign addr[24937]= -1960577471;
assign addr[24938]= -1975871368;
assign addr[24939]= -1990538579;
assign addr[24940]= -2004574453;
assign addr[24941]= -2017974537;
assign addr[24942]= -2030734582;
assign addr[24943]= -2042850540;
assign addr[24944]= -2054318569;
assign addr[24945]= -2065135031;
assign addr[24946]= -2075296495;
assign addr[24947]= -2084799740;
assign addr[24948]= -2093641749;
assign addr[24949]= -2101819720;
assign addr[24950]= -2109331059;
assign addr[24951]= -2116173382;
assign addr[24952]= -2122344521;
assign addr[24953]= -2127842516;
assign addr[24954]= -2132665626;
assign addr[24955]= -2136812319;
assign addr[24956]= -2140281282;
assign addr[24957]= -2143071413;
assign addr[24958]= -2145181827;
assign addr[24959]= -2146611856;
assign addr[24960]= -2147361045;
assign addr[24961]= -2147429158;
assign addr[24962]= -2146816171;
assign addr[24963]= -2145522281;
assign addr[24964]= -2143547897;
assign addr[24965]= -2140893646;
assign addr[24966]= -2137560369;
assign addr[24967]= -2133549123;
assign addr[24968]= -2128861181;
assign addr[24969]= -2123498030;
assign addr[24970]= -2117461370;
assign addr[24971]= -2110753117;
assign addr[24972]= -2103375398;
assign addr[24973]= -2095330553;
assign addr[24974]= -2086621133;
assign addr[24975]= -2077249901;
assign addr[24976]= -2067219829;
assign addr[24977]= -2056534099;
assign addr[24978]= -2045196100;
assign addr[24979]= -2033209426;
assign addr[24980]= -2020577882;
assign addr[24981]= -2007305472;
assign addr[24982]= -1993396407;
assign addr[24983]= -1978855097;
assign addr[24984]= -1963686155;
assign addr[24985]= -1947894393;
assign addr[24986]= -1931484818;
assign addr[24987]= -1914462636;
assign addr[24988]= -1896833245;
assign addr[24989]= -1878602237;
assign addr[24990]= -1859775393;
assign addr[24991]= -1840358687;
assign addr[24992]= -1820358275;
assign addr[24993]= -1799780501;
assign addr[24994]= -1778631892;
assign addr[24995]= -1756919156;
assign addr[24996]= -1734649179;
assign addr[24997]= -1711829025;
assign addr[24998]= -1688465931;
assign addr[24999]= -1664567307;
assign addr[25000]= -1640140734;
assign addr[25001]= -1615193959;
assign addr[25002]= -1589734894;
assign addr[25003]= -1563771613;
assign addr[25004]= -1537312353;
assign addr[25005]= -1510365504;
assign addr[25006]= -1482939614;
assign addr[25007]= -1455043381;
assign addr[25008]= -1426685652;
assign addr[25009]= -1397875423;
assign addr[25010]= -1368621831;
assign addr[25011]= -1338934154;
assign addr[25012]= -1308821808;
assign addr[25013]= -1278294345;
assign addr[25014]= -1247361445;
assign addr[25015]= -1216032921;
assign addr[25016]= -1184318708;
assign addr[25017]= -1152228866;
assign addr[25018]= -1119773573;
assign addr[25019]= -1086963121;
assign addr[25020]= -1053807919;
assign addr[25021]= -1020318481;
assign addr[25022]= -986505429;
assign addr[25023]= -952379488;
assign addr[25024]= -917951481;
assign addr[25025]= -883232329;
assign addr[25026]= -848233042;
assign addr[25027]= -812964722;
assign addr[25028]= -777438554;
assign addr[25029]= -741665807;
assign addr[25030]= -705657826;
assign addr[25031]= -669426032;
assign addr[25032]= -632981917;
assign addr[25033]= -596337040;
assign addr[25034]= -559503022;
assign addr[25035]= -522491548;
assign addr[25036]= -485314355;
assign addr[25037]= -447983235;
assign addr[25038]= -410510029;
assign addr[25039]= -372906622;
assign addr[25040]= -335184940;
assign addr[25041]= -297356948;
assign addr[25042]= -259434643;
assign addr[25043]= -221430054;
assign addr[25044]= -183355234;
assign addr[25045]= -145222259;
assign addr[25046]= -107043224;
assign addr[25047]= -68830239;
assign addr[25048]= -30595422;
assign addr[25049]= 7649098;
assign addr[25050]= 45891193;
assign addr[25051]= 84118732;
assign addr[25052]= 122319591;
assign addr[25053]= 160481654;
assign addr[25054]= 198592817;
assign addr[25055]= 236640993;
assign addr[25056]= 274614114;
assign addr[25057]= 312500135;
assign addr[25058]= 350287041;
assign addr[25059]= 387962847;
assign addr[25060]= 425515602;
assign addr[25061]= 462933398;
assign addr[25062]= 500204365;
assign addr[25063]= 537316682;
assign addr[25064]= 574258580;
assign addr[25065]= 611018340;
assign addr[25066]= 647584304;
assign addr[25067]= 683944874;
assign addr[25068]= 720088517;
assign addr[25069]= 756003771;
assign addr[25070]= 791679244;
assign addr[25071]= 827103620;
assign addr[25072]= 862265664;
assign addr[25073]= 897154224;
assign addr[25074]= 931758235;
assign addr[25075]= 966066720;
assign addr[25076]= 1000068799;
assign addr[25077]= 1033753687;
assign addr[25078]= 1067110699;
assign addr[25079]= 1100129257;
assign addr[25080]= 1132798888;
assign addr[25081]= 1165109230;
assign addr[25082]= 1197050035;
assign addr[25083]= 1228611172;
assign addr[25084]= 1259782632;
assign addr[25085]= 1290554528;
assign addr[25086]= 1320917099;
assign addr[25087]= 1350860716;
assign addr[25088]= 1380375881;
assign addr[25089]= 1409453233;
assign addr[25090]= 1438083551;
assign addr[25091]= 1466257752;
assign addr[25092]= 1493966902;
assign addr[25093]= 1521202211;
assign addr[25094]= 1547955041;
assign addr[25095]= 1574216908;
assign addr[25096]= 1599979481;
assign addr[25097]= 1625234591;
assign addr[25098]= 1649974225;
assign addr[25099]= 1674190539;
assign addr[25100]= 1697875851;
assign addr[25101]= 1721022648;
assign addr[25102]= 1743623590;
assign addr[25103]= 1765671509;
assign addr[25104]= 1787159411;
assign addr[25105]= 1808080480;
assign addr[25106]= 1828428082;
assign addr[25107]= 1848195763;
assign addr[25108]= 1867377253;
assign addr[25109]= 1885966468;
assign addr[25110]= 1903957513;
assign addr[25111]= 1921344681;
assign addr[25112]= 1938122457;
assign addr[25113]= 1954285520;
assign addr[25114]= 1969828744;
assign addr[25115]= 1984747199;
assign addr[25116]= 1999036154;
assign addr[25117]= 2012691075;
assign addr[25118]= 2025707632;
assign addr[25119]= 2038081698;
assign addr[25120]= 2049809346;
assign addr[25121]= 2060886858;
assign addr[25122]= 2071310720;
assign addr[25123]= 2081077626;
assign addr[25124]= 2090184478;
assign addr[25125]= 2098628387;
assign addr[25126]= 2106406677;
assign addr[25127]= 2113516878;
assign addr[25128]= 2119956737;
assign addr[25129]= 2125724211;
assign addr[25130]= 2130817471;
assign addr[25131]= 2135234901;
assign addr[25132]= 2138975100;
assign addr[25133]= 2142036881;
assign addr[25134]= 2144419275;
assign addr[25135]= 2146121524;
assign addr[25136]= 2147143090;
assign addr[25137]= 2147483648;
assign addr[25138]= 2147143090;
assign addr[25139]= 2146121524;
assign addr[25140]= 2144419275;
assign addr[25141]= 2142036881;
assign addr[25142]= 2138975100;
assign addr[25143]= 2135234901;
assign addr[25144]= 2130817471;
assign addr[25145]= 2125724211;
assign addr[25146]= 2119956737;
assign addr[25147]= 2113516878;
assign addr[25148]= 2106406677;
assign addr[25149]= 2098628387;
assign addr[25150]= 2090184478;
assign addr[25151]= 2081077626;
assign addr[25152]= 2071310720;
assign addr[25153]= 2060886858;
assign addr[25154]= 2049809346;
assign addr[25155]= 2038081698;
assign addr[25156]= 2025707632;
assign addr[25157]= 2012691075;
assign addr[25158]= 1999036154;
assign addr[25159]= 1984747199;
assign addr[25160]= 1969828744;
assign addr[25161]= 1954285520;
assign addr[25162]= 1938122457;
assign addr[25163]= 1921344681;
assign addr[25164]= 1903957513;
assign addr[25165]= 1885966468;
assign addr[25166]= 1867377253;
assign addr[25167]= 1848195763;
assign addr[25168]= 1828428082;
assign addr[25169]= 1808080480;
assign addr[25170]= 1787159411;
assign addr[25171]= 1765671509;
assign addr[25172]= 1743623590;
assign addr[25173]= 1721022648;
assign addr[25174]= 1697875851;
assign addr[25175]= 1674190539;
assign addr[25176]= 1649974225;
assign addr[25177]= 1625234591;
assign addr[25178]= 1599979481;
assign addr[25179]= 1574216908;
assign addr[25180]= 1547955041;
assign addr[25181]= 1521202211;
assign addr[25182]= 1493966902;
assign addr[25183]= 1466257752;
assign addr[25184]= 1438083551;
assign addr[25185]= 1409453233;
assign addr[25186]= 1380375881;
assign addr[25187]= 1350860716;
assign addr[25188]= 1320917099;
assign addr[25189]= 1290554528;
assign addr[25190]= 1259782632;
assign addr[25191]= 1228611172;
assign addr[25192]= 1197050035;
assign addr[25193]= 1165109230;
assign addr[25194]= 1132798888;
assign addr[25195]= 1100129257;
assign addr[25196]= 1067110699;
assign addr[25197]= 1033753687;
assign addr[25198]= 1000068799;
assign addr[25199]= 966066720;
assign addr[25200]= 931758235;
assign addr[25201]= 897154224;
assign addr[25202]= 862265664;
assign addr[25203]= 827103620;
assign addr[25204]= 791679244;
assign addr[25205]= 756003771;
assign addr[25206]= 720088517;
assign addr[25207]= 683944874;
assign addr[25208]= 647584304;
assign addr[25209]= 611018340;
assign addr[25210]= 574258580;
assign addr[25211]= 537316682;
assign addr[25212]= 500204365;
assign addr[25213]= 462933398;
assign addr[25214]= 425515602;
assign addr[25215]= 387962847;
assign addr[25216]= 350287041;
assign addr[25217]= 312500135;
assign addr[25218]= 274614114;
assign addr[25219]= 236640993;
assign addr[25220]= 198592817;
assign addr[25221]= 160481654;
assign addr[25222]= 122319591;
assign addr[25223]= 84118732;
assign addr[25224]= 45891193;
assign addr[25225]= 7649098;
assign addr[25226]= -30595422;
assign addr[25227]= -68830239;
assign addr[25228]= -107043224;
assign addr[25229]= -145222259;
assign addr[25230]= -183355234;
assign addr[25231]= -221430054;
assign addr[25232]= -259434643;
assign addr[25233]= -297356948;
assign addr[25234]= -335184940;
assign addr[25235]= -372906622;
assign addr[25236]= -410510029;
assign addr[25237]= -447983235;
assign addr[25238]= -485314355;
assign addr[25239]= -522491548;
assign addr[25240]= -559503022;
assign addr[25241]= -596337040;
assign addr[25242]= -632981917;
assign addr[25243]= -669426032;
assign addr[25244]= -705657826;
assign addr[25245]= -741665807;
assign addr[25246]= -777438554;
assign addr[25247]= -812964722;
assign addr[25248]= -848233042;
assign addr[25249]= -883232329;
assign addr[25250]= -917951481;
assign addr[25251]= -952379488;
assign addr[25252]= -986505429;
assign addr[25253]= -1020318481;
assign addr[25254]= -1053807919;
assign addr[25255]= -1086963121;
assign addr[25256]= -1119773573;
assign addr[25257]= -1152228866;
assign addr[25258]= -1184318708;
assign addr[25259]= -1216032921;
assign addr[25260]= -1247361445;
assign addr[25261]= -1278294345;
assign addr[25262]= -1308821808;
assign addr[25263]= -1338934154;
assign addr[25264]= -1368621831;
assign addr[25265]= -1397875423;
assign addr[25266]= -1426685652;
assign addr[25267]= -1455043381;
assign addr[25268]= -1482939614;
assign addr[25269]= -1510365504;
assign addr[25270]= -1537312353;
assign addr[25271]= -1563771613;
assign addr[25272]= -1589734894;
assign addr[25273]= -1615193959;
assign addr[25274]= -1640140734;
assign addr[25275]= -1664567307;
assign addr[25276]= -1688465931;
assign addr[25277]= -1711829025;
assign addr[25278]= -1734649179;
assign addr[25279]= -1756919156;
assign addr[25280]= -1778631892;
assign addr[25281]= -1799780501;
assign addr[25282]= -1820358275;
assign addr[25283]= -1840358687;
assign addr[25284]= -1859775393;
assign addr[25285]= -1878602237;
assign addr[25286]= -1896833245;
assign addr[25287]= -1914462636;
assign addr[25288]= -1931484818;
assign addr[25289]= -1947894393;
assign addr[25290]= -1963686155;
assign addr[25291]= -1978855097;
assign addr[25292]= -1993396407;
assign addr[25293]= -2007305472;
assign addr[25294]= -2020577882;
assign addr[25295]= -2033209426;
assign addr[25296]= -2045196100;
assign addr[25297]= -2056534099;
assign addr[25298]= -2067219829;
assign addr[25299]= -2077249901;
assign addr[25300]= -2086621133;
assign addr[25301]= -2095330553;
assign addr[25302]= -2103375398;
assign addr[25303]= -2110753117;
assign addr[25304]= -2117461370;
assign addr[25305]= -2123498030;
assign addr[25306]= -2128861181;
assign addr[25307]= -2133549123;
assign addr[25308]= -2137560369;
assign addr[25309]= -2140893646;
assign addr[25310]= -2143547897;
assign addr[25311]= -2145522281;
assign addr[25312]= -2146816171;
assign addr[25313]= -2147429158;
assign addr[25314]= -2147361045;
assign addr[25315]= -2146611856;
assign addr[25316]= -2145181827;
assign addr[25317]= -2143071413;
assign addr[25318]= -2140281282;
assign addr[25319]= -2136812319;
assign addr[25320]= -2132665626;
assign addr[25321]= -2127842516;
assign addr[25322]= -2122344521;
assign addr[25323]= -2116173382;
assign addr[25324]= -2109331059;
assign addr[25325]= -2101819720;
assign addr[25326]= -2093641749;
assign addr[25327]= -2084799740;
assign addr[25328]= -2075296495;
assign addr[25329]= -2065135031;
assign addr[25330]= -2054318569;
assign addr[25331]= -2042850540;
assign addr[25332]= -2030734582;
assign addr[25333]= -2017974537;
assign addr[25334]= -2004574453;
assign addr[25335]= -1990538579;
assign addr[25336]= -1975871368;
assign addr[25337]= -1960577471;
assign addr[25338]= -1944661739;
assign addr[25339]= -1928129220;
assign addr[25340]= -1910985158;
assign addr[25341]= -1893234990;
assign addr[25342]= -1874884346;
assign addr[25343]= -1855939047;
assign addr[25344]= -1836405100;
assign addr[25345]= -1816288703;
assign addr[25346]= -1795596234;
assign addr[25347]= -1774334257;
assign addr[25348]= -1752509516;
assign addr[25349]= -1730128933;
assign addr[25350]= -1707199606;
assign addr[25351]= -1683728808;
assign addr[25352]= -1659723983;
assign addr[25353]= -1635192744;
assign addr[25354]= -1610142873;
assign addr[25355]= -1584582314;
assign addr[25356]= -1558519173;
assign addr[25357]= -1531961719;
assign addr[25358]= -1504918373;
assign addr[25359]= -1477397714;
assign addr[25360]= -1449408469;
assign addr[25361]= -1420959516;
assign addr[25362]= -1392059879;
assign addr[25363]= -1362718723;
assign addr[25364]= -1332945355;
assign addr[25365]= -1302749217;
assign addr[25366]= -1272139887;
assign addr[25367]= -1241127074;
assign addr[25368]= -1209720613;
assign addr[25369]= -1177930466;
assign addr[25370]= -1145766716;
assign addr[25371]= -1113239564;
assign addr[25372]= -1080359326;
assign addr[25373]= -1047136432;
assign addr[25374]= -1013581418;
assign addr[25375]= -979704927;
assign addr[25376]= -945517704;
assign addr[25377]= -911030591;
assign addr[25378]= -876254528;
assign addr[25379]= -841200544;
assign addr[25380]= -805879757;
assign addr[25381]= -770303369;
assign addr[25382]= -734482665;
assign addr[25383]= -698429006;
assign addr[25384]= -662153826;
assign addr[25385]= -625668632;
assign addr[25386]= -588984994;
assign addr[25387]= -552114549;
assign addr[25388]= -515068990;
assign addr[25389]= -477860067;
assign addr[25390]= -440499581;
assign addr[25391]= -402999383;
assign addr[25392]= -365371365;
assign addr[25393]= -327627463;
assign addr[25394]= -289779648;
assign addr[25395]= -251839923;
assign addr[25396]= -213820322;
assign addr[25397]= -175732905;
assign addr[25398]= -137589750;
assign addr[25399]= -99402956;
assign addr[25400]= -61184634;
assign addr[25401]= -22946906;
assign addr[25402]= 15298099;
assign addr[25403]= 53538253;
assign addr[25404]= 91761426;
assign addr[25405]= 129955495;
assign addr[25406]= 168108346;
assign addr[25407]= 206207878;
assign addr[25408]= 244242007;
assign addr[25409]= 282198671;
assign addr[25410]= 320065829;
assign addr[25411]= 357831473;
assign addr[25412]= 395483624;
assign addr[25413]= 433010339;
assign addr[25414]= 470399716;
assign addr[25415]= 507639898;
assign addr[25416]= 544719071;
assign addr[25417]= 581625477;
assign addr[25418]= 618347408;
assign addr[25419]= 654873219;
assign addr[25420]= 691191324;
assign addr[25421]= 727290205;
assign addr[25422]= 763158411;
assign addr[25423]= 798784567;
assign addr[25424]= 834157373;
assign addr[25425]= 869265610;
assign addr[25426]= 904098143;
assign addr[25427]= 938643924;
assign addr[25428]= 972891995;
assign addr[25429]= 1006831495;
assign addr[25430]= 1040451659;
assign addr[25431]= 1073741824;
assign addr[25432]= 1106691431;
assign addr[25433]= 1139290029;
assign addr[25434]= 1171527280;
assign addr[25435]= 1203392958;
assign addr[25436]= 1234876957;
assign addr[25437]= 1265969291;
assign addr[25438]= 1296660098;
assign addr[25439]= 1326939644;
assign addr[25440]= 1356798326;
assign addr[25441]= 1386226674;
assign addr[25442]= 1415215352;
assign addr[25443]= 1443755168;
assign addr[25444]= 1471837070;
assign addr[25445]= 1499452149;
assign addr[25446]= 1526591649;
assign addr[25447]= 1553246960;
assign addr[25448]= 1579409630;
assign addr[25449]= 1605071359;
assign addr[25450]= 1630224009;
assign addr[25451]= 1654859602;
assign addr[25452]= 1678970324;
assign addr[25453]= 1702548529;
assign addr[25454]= 1725586737;
assign addr[25455]= 1748077642;
assign addr[25456]= 1770014111;
assign addr[25457]= 1791389186;
assign addr[25458]= 1812196087;
assign addr[25459]= 1832428215;
assign addr[25460]= 1852079154;
assign addr[25461]= 1871142669;
assign addr[25462]= 1889612716;
assign addr[25463]= 1907483436;
assign addr[25464]= 1924749160;
assign addr[25465]= 1941404413;
assign addr[25466]= 1957443913;
assign addr[25467]= 1972862571;
assign addr[25468]= 1987655498;
assign addr[25469]= 2001818002;
assign addr[25470]= 2015345591;
assign addr[25471]= 2028233973;
assign addr[25472]= 2040479063;
assign addr[25473]= 2052076975;
assign addr[25474]= 2063024031;
assign addr[25475]= 2073316760;
assign addr[25476]= 2082951896;
assign addr[25477]= 2091926384;
assign addr[25478]= 2100237377;
assign addr[25479]= 2107882239;
assign addr[25480]= 2114858546;
assign addr[25481]= 2121164085;
assign addr[25482]= 2126796855;
assign addr[25483]= 2131755071;
assign addr[25484]= 2136037160;
assign addr[25485]= 2139641764;
assign addr[25486]= 2142567738;
assign addr[25487]= 2144814157;
assign addr[25488]= 2146380306;
assign addr[25489]= 2147265689;
assign addr[25490]= 2147470025;
assign addr[25491]= 2146993250;
assign addr[25492]= 2145835515;
assign addr[25493]= 2143997187;
assign addr[25494]= 2141478848;
assign addr[25495]= 2138281298;
assign addr[25496]= 2134405552;
assign addr[25497]= 2129852837;
assign addr[25498]= 2124624598;
assign addr[25499]= 2118722494;
assign addr[25500]= 2112148396;
assign addr[25501]= 2104904390;
assign addr[25502]= 2096992772;
assign addr[25503]= 2088416053;
assign addr[25504]= 2079176953;
assign addr[25505]= 2069278401;
assign addr[25506]= 2058723538;
assign addr[25507]= 2047515711;
assign addr[25508]= 2035658475;
assign addr[25509]= 2023155591;
assign addr[25510]= 2010011024;
assign addr[25511]= 1996228943;
assign addr[25512]= 1981813720;
assign addr[25513]= 1966769926;
assign addr[25514]= 1951102334;
assign addr[25515]= 1934815911;
assign addr[25516]= 1917915825;
assign addr[25517]= 1900407434;
assign addr[25518]= 1882296293;
assign addr[25519]= 1863588145;
assign addr[25520]= 1844288924;
assign addr[25521]= 1824404752;
assign addr[25522]= 1803941934;
assign addr[25523]= 1782906961;
assign addr[25524]= 1761306505;
assign addr[25525]= 1739147417;
assign addr[25526]= 1716436725;
assign addr[25527]= 1693181631;
assign addr[25528]= 1669389513;
assign addr[25529]= 1645067915;
assign addr[25530]= 1620224553;
assign addr[25531]= 1594867305;
assign addr[25532]= 1569004214;
assign addr[25533]= 1542643483;
assign addr[25534]= 1515793473;
assign addr[25535]= 1488462700;
assign addr[25536]= 1460659832;
assign addr[25537]= 1432393688;
assign addr[25538]= 1403673233;
assign addr[25539]= 1374507575;
assign addr[25540]= 1344905966;
assign addr[25541]= 1314877795;
assign addr[25542]= 1284432584;
assign addr[25543]= 1253579991;
assign addr[25544]= 1222329801;
assign addr[25545]= 1190691925;
assign addr[25546]= 1158676398;
assign addr[25547]= 1126293375;
assign addr[25548]= 1093553126;
assign addr[25549]= 1060466036;
assign addr[25550]= 1027042599;
assign addr[25551]= 993293415;
assign addr[25552]= 959229189;
assign addr[25553]= 924860725;
assign addr[25554]= 890198924;
assign addr[25555]= 855254778;
assign addr[25556]= 820039373;
assign addr[25557]= 784563876;
assign addr[25558]= 748839539;
assign addr[25559]= 712877694;
assign addr[25560]= 676689746;
assign addr[25561]= 640287172;
assign addr[25562]= 603681519;
assign addr[25563]= 566884397;
assign addr[25564]= 529907477;
assign addr[25565]= 492762486;
assign addr[25566]= 455461206;
assign addr[25567]= 418015468;
assign addr[25568]= 380437148;
assign addr[25569]= 342738165;
assign addr[25570]= 304930476;
assign addr[25571]= 267026072;
assign addr[25572]= 229036977;
assign addr[25573]= 190975237;
assign addr[25574]= 152852926;
assign addr[25575]= 114682135;
assign addr[25576]= 76474970;
assign addr[25577]= 38243550;
assign addr[25578]= 0;
assign addr[25579]= -38243550;
assign addr[25580]= -76474970;
assign addr[25581]= -114682135;
assign addr[25582]= -152852926;
assign addr[25583]= -190975237;
assign addr[25584]= -229036977;
assign addr[25585]= -267026072;
assign addr[25586]= -304930476;
assign addr[25587]= -342738165;
assign addr[25588]= -380437148;
assign addr[25589]= -418015468;
assign addr[25590]= -455461206;
assign addr[25591]= -492762486;
assign addr[25592]= -529907477;
assign addr[25593]= -566884397;
assign addr[25594]= -603681519;
assign addr[25595]= -640287172;
assign addr[25596]= -676689746;
assign addr[25597]= -712877694;
assign addr[25598]= -748839539;
assign addr[25599]= -784563876;
assign addr[25600]= -820039373;
assign addr[25601]= -855254778;
assign addr[25602]= -890198924;
assign addr[25603]= -924860725;
assign addr[25604]= -959229189;
assign addr[25605]= -993293415;
assign addr[25606]= -1027042599;
assign addr[25607]= -1060466036;
assign addr[25608]= -1093553126;
assign addr[25609]= -1126293375;
assign addr[25610]= -1158676398;
assign addr[25611]= -1190691925;
assign addr[25612]= -1222329801;
assign addr[25613]= -1253579991;
assign addr[25614]= -1284432584;
assign addr[25615]= -1314877795;
assign addr[25616]= -1344905966;
assign addr[25617]= -1374507575;
assign addr[25618]= -1403673233;
assign addr[25619]= -1432393688;
assign addr[25620]= -1460659832;
assign addr[25621]= -1488462700;
assign addr[25622]= -1515793473;
assign addr[25623]= -1542643483;
assign addr[25624]= -1569004214;
assign addr[25625]= -1594867305;
assign addr[25626]= -1620224553;
assign addr[25627]= -1645067915;
assign addr[25628]= -1669389513;
assign addr[25629]= -1693181631;
assign addr[25630]= -1716436725;
assign addr[25631]= -1739147417;
assign addr[25632]= -1761306505;
assign addr[25633]= -1782906961;
assign addr[25634]= -1803941934;
assign addr[25635]= -1824404752;
assign addr[25636]= -1844288924;
assign addr[25637]= -1863588145;
assign addr[25638]= -1882296293;
assign addr[25639]= -1900407434;
assign addr[25640]= -1917915825;
assign addr[25641]= -1934815911;
assign addr[25642]= -1951102334;
assign addr[25643]= -1966769926;
assign addr[25644]= -1981813720;
assign addr[25645]= -1996228943;
assign addr[25646]= -2010011024;
assign addr[25647]= -2023155591;
assign addr[25648]= -2035658475;
assign addr[25649]= -2047515711;
assign addr[25650]= -2058723538;
assign addr[25651]= -2069278401;
assign addr[25652]= -2079176953;
assign addr[25653]= -2088416053;
assign addr[25654]= -2096992772;
assign addr[25655]= -2104904390;
assign addr[25656]= -2112148396;
assign addr[25657]= -2118722494;
assign addr[25658]= -2124624598;
assign addr[25659]= -2129852837;
assign addr[25660]= -2134405552;
assign addr[25661]= -2138281298;
assign addr[25662]= -2141478848;
assign addr[25663]= -2143997187;
assign addr[25664]= -2145835515;
assign addr[25665]= -2146993250;
assign addr[25666]= -2147470025;
assign addr[25667]= -2147265689;
assign addr[25668]= -2146380306;
assign addr[25669]= -2144814157;
assign addr[25670]= -2142567738;
assign addr[25671]= -2139641764;
assign addr[25672]= -2136037160;
assign addr[25673]= -2131755071;
assign addr[25674]= -2126796855;
assign addr[25675]= -2121164085;
assign addr[25676]= -2114858546;
assign addr[25677]= -2107882239;
assign addr[25678]= -2100237377;
assign addr[25679]= -2091926384;
assign addr[25680]= -2082951896;
assign addr[25681]= -2073316760;
assign addr[25682]= -2063024031;
assign addr[25683]= -2052076975;
assign addr[25684]= -2040479063;
assign addr[25685]= -2028233973;
assign addr[25686]= -2015345591;
assign addr[25687]= -2001818002;
assign addr[25688]= -1987655498;
assign addr[25689]= -1972862571;
assign addr[25690]= -1957443913;
assign addr[25691]= -1941404413;
assign addr[25692]= -1924749160;
assign addr[25693]= -1907483436;
assign addr[25694]= -1889612716;
assign addr[25695]= -1871142669;
assign addr[25696]= -1852079154;
assign addr[25697]= -1832428215;
assign addr[25698]= -1812196087;
assign addr[25699]= -1791389186;
assign addr[25700]= -1770014111;
assign addr[25701]= -1748077642;
assign addr[25702]= -1725586737;
assign addr[25703]= -1702548529;
assign addr[25704]= -1678970324;
assign addr[25705]= -1654859602;
assign addr[25706]= -1630224009;
assign addr[25707]= -1605071359;
assign addr[25708]= -1579409630;
assign addr[25709]= -1553246960;
assign addr[25710]= -1526591649;
assign addr[25711]= -1499452149;
assign addr[25712]= -1471837070;
assign addr[25713]= -1443755168;
assign addr[25714]= -1415215352;
assign addr[25715]= -1386226674;
assign addr[25716]= -1356798326;
assign addr[25717]= -1326939644;
assign addr[25718]= -1296660098;
assign addr[25719]= -1265969291;
assign addr[25720]= -1234876957;
assign addr[25721]= -1203392958;
assign addr[25722]= -1171527280;
assign addr[25723]= -1139290029;
assign addr[25724]= -1106691431;
assign addr[25725]= -1073741824;
assign addr[25726]= -1040451659;
assign addr[25727]= -1006831495;
assign addr[25728]= -972891995;
assign addr[25729]= -938643924;
assign addr[25730]= -904098143;
assign addr[25731]= -869265610;
assign addr[25732]= -834157373;
assign addr[25733]= -798784567;
assign addr[25734]= -763158411;
assign addr[25735]= -727290205;
assign addr[25736]= -691191324;
assign addr[25737]= -654873219;
assign addr[25738]= -618347408;
assign addr[25739]= -581625477;
assign addr[25740]= -544719071;
assign addr[25741]= -507639898;
assign addr[25742]= -470399716;
assign addr[25743]= -433010339;
assign addr[25744]= -395483624;
assign addr[25745]= -357831473;
assign addr[25746]= -320065829;
assign addr[25747]= -282198671;
assign addr[25748]= -244242007;
assign addr[25749]= -206207878;
assign addr[25750]= -168108346;
assign addr[25751]= -129955495;
assign addr[25752]= -91761426;
assign addr[25753]= -53538253;
assign addr[25754]= -15298099;
assign addr[25755]= 22946906;
assign addr[25756]= 61184634;
assign addr[25757]= 99402956;
assign addr[25758]= 137589750;
assign addr[25759]= 175732905;
assign addr[25760]= 213820322;
assign addr[25761]= 251839923;
assign addr[25762]= 289779648;
assign addr[25763]= 327627463;
assign addr[25764]= 365371365;
assign addr[25765]= 402999383;
assign addr[25766]= 440499581;
assign addr[25767]= 477860067;
assign addr[25768]= 515068990;
assign addr[25769]= 552114549;
assign addr[25770]= 588984994;
assign addr[25771]= 625668632;
assign addr[25772]= 662153826;
assign addr[25773]= 698429006;
assign addr[25774]= 734482665;
assign addr[25775]= 770303369;
assign addr[25776]= 805879757;
assign addr[25777]= 841200544;
assign addr[25778]= 876254528;
assign addr[25779]= 911030591;
assign addr[25780]= 945517704;
assign addr[25781]= 979704927;
assign addr[25782]= 1013581418;
assign addr[25783]= 1047136432;
assign addr[25784]= 1080359326;
assign addr[25785]= 1113239564;
assign addr[25786]= 1145766716;
assign addr[25787]= 1177930466;
assign addr[25788]= 1209720613;
assign addr[25789]= 1241127074;
assign addr[25790]= 1272139887;
assign addr[25791]= 1302749217;
assign addr[25792]= 1332945355;
assign addr[25793]= 1362718723;
assign addr[25794]= 1392059879;
assign addr[25795]= 1420959516;
assign addr[25796]= 1449408469;
assign addr[25797]= 1477397714;
assign addr[25798]= 1504918373;
assign addr[25799]= 1531961719;
assign addr[25800]= 1558519173;
assign addr[25801]= 1584582314;
assign addr[25802]= 1610142873;
assign addr[25803]= 1635192744;
assign addr[25804]= 1659723983;
assign addr[25805]= 1683728808;
assign addr[25806]= 1707199606;
assign addr[25807]= 1730128933;
assign addr[25808]= 1752509516;
assign addr[25809]= 1774334257;
assign addr[25810]= 1795596234;
assign addr[25811]= 1816288703;
assign addr[25812]= 1836405100;
assign addr[25813]= 1855939047;
assign addr[25814]= 1874884346;
assign addr[25815]= 1893234990;
assign addr[25816]= 1910985158;
assign addr[25817]= 1928129220;
assign addr[25818]= 1944661739;
assign addr[25819]= 1960577471;
assign addr[25820]= 1975871368;
assign addr[25821]= 1990538579;
assign addr[25822]= 2004574453;
assign addr[25823]= 2017974537;
assign addr[25824]= 2030734582;
assign addr[25825]= 2042850540;
assign addr[25826]= 2054318569;
assign addr[25827]= 2065135031;
assign addr[25828]= 2075296495;
assign addr[25829]= 2084799740;
assign addr[25830]= 2093641749;
assign addr[25831]= 2101819720;
assign addr[25832]= 2109331059;
assign addr[25833]= 2116173382;
assign addr[25834]= 2122344521;
assign addr[25835]= 2127842516;
assign addr[25836]= 2132665626;
assign addr[25837]= 2136812319;
assign addr[25838]= 2140281282;
assign addr[25839]= 2143071413;
assign addr[25840]= 2145181827;
assign addr[25841]= 2146611856;
assign addr[25842]= 2147361045;
assign addr[25843]= 2147429158;
assign addr[25844]= 2146816171;
assign addr[25845]= 2145522281;
assign addr[25846]= 2143547897;
assign addr[25847]= 2140893646;
assign addr[25848]= 2137560369;
assign addr[25849]= 2133549123;
assign addr[25850]= 2128861181;
assign addr[25851]= 2123498030;
assign addr[25852]= 2117461370;
assign addr[25853]= 2110753117;
assign addr[25854]= 2103375398;
assign addr[25855]= 2095330553;
assign addr[25856]= 2086621133;
assign addr[25857]= 2077249901;
assign addr[25858]= 2067219829;
assign addr[25859]= 2056534099;
assign addr[25860]= 2045196100;
assign addr[25861]= 2033209426;
assign addr[25862]= 2020577882;
assign addr[25863]= 2007305472;
assign addr[25864]= 1993396407;
assign addr[25865]= 1978855097;
assign addr[25866]= 1963686155;
assign addr[25867]= 1947894393;
assign addr[25868]= 1931484818;
assign addr[25869]= 1914462636;
assign addr[25870]= 1896833245;
assign addr[25871]= 1878602237;
assign addr[25872]= 1859775393;
assign addr[25873]= 1840358687;
assign addr[25874]= 1820358275;
assign addr[25875]= 1799780501;
assign addr[25876]= 1778631892;
assign addr[25877]= 1756919156;
assign addr[25878]= 1734649179;
assign addr[25879]= 1711829025;
assign addr[25880]= 1688465931;
assign addr[25881]= 1664567307;
assign addr[25882]= 1640140734;
assign addr[25883]= 1615193959;
assign addr[25884]= 1589734894;
assign addr[25885]= 1563771613;
assign addr[25886]= 1537312353;
assign addr[25887]= 1510365504;
assign addr[25888]= 1482939614;
assign addr[25889]= 1455043381;
assign addr[25890]= 1426685652;
assign addr[25891]= 1397875423;
assign addr[25892]= 1368621831;
assign addr[25893]= 1338934154;
assign addr[25894]= 1308821808;
assign addr[25895]= 1278294345;
assign addr[25896]= 1247361445;
assign addr[25897]= 1216032921;
assign addr[25898]= 1184318708;
assign addr[25899]= 1152228866;
assign addr[25900]= 1119773573;
assign addr[25901]= 1086963121;
assign addr[25902]= 1053807919;
assign addr[25903]= 1020318481;
assign addr[25904]= 986505429;
assign addr[25905]= 952379488;
assign addr[25906]= 917951481;
assign addr[25907]= 883232329;
assign addr[25908]= 848233042;
assign addr[25909]= 812964722;
assign addr[25910]= 777438554;
assign addr[25911]= 741665807;
assign addr[25912]= 705657826;
assign addr[25913]= 669426032;
assign addr[25914]= 632981917;
assign addr[25915]= 596337040;
assign addr[25916]= 559503022;
assign addr[25917]= 522491548;
assign addr[25918]= 485314355;
assign addr[25919]= 447983235;
assign addr[25920]= 410510029;
assign addr[25921]= 372906622;
assign addr[25922]= 335184940;
assign addr[25923]= 297356948;
assign addr[25924]= 259434643;
assign addr[25925]= 221430054;
assign addr[25926]= 183355234;
assign addr[25927]= 145222259;
assign addr[25928]= 107043224;
assign addr[25929]= 68830239;
assign addr[25930]= 30595422;
assign addr[25931]= -7649098;
assign addr[25932]= -45891193;
assign addr[25933]= -84118732;
assign addr[25934]= -122319591;
assign addr[25935]= -160481654;
assign addr[25936]= -198592817;
assign addr[25937]= -236640993;
assign addr[25938]= -274614114;
assign addr[25939]= -312500135;
assign addr[25940]= -350287041;
assign addr[25941]= -387962847;
assign addr[25942]= -425515602;
assign addr[25943]= -462933398;
assign addr[25944]= -500204365;
assign addr[25945]= -537316682;
assign addr[25946]= -574258580;
assign addr[25947]= -611018340;
assign addr[25948]= -647584304;
assign addr[25949]= -683944874;
assign addr[25950]= -720088517;
assign addr[25951]= -756003771;
assign addr[25952]= -791679244;
assign addr[25953]= -827103620;
assign addr[25954]= -862265664;
assign addr[25955]= -897154224;
assign addr[25956]= -931758235;
assign addr[25957]= -966066720;
assign addr[25958]= -1000068799;
assign addr[25959]= -1033753687;
assign addr[25960]= -1067110699;
assign addr[25961]= -1100129257;
assign addr[25962]= -1132798888;
assign addr[25963]= -1165109230;
assign addr[25964]= -1197050035;
assign addr[25965]= -1228611172;
assign addr[25966]= -1259782632;
assign addr[25967]= -1290554528;
assign addr[25968]= -1320917099;
assign addr[25969]= -1350860716;
assign addr[25970]= -1380375881;
assign addr[25971]= -1409453233;
assign addr[25972]= -1438083551;
assign addr[25973]= -1466257752;
assign addr[25974]= -1493966902;
assign addr[25975]= -1521202211;
assign addr[25976]= -1547955041;
assign addr[25977]= -1574216908;
assign addr[25978]= -1599979481;
assign addr[25979]= -1625234591;
assign addr[25980]= -1649974225;
assign addr[25981]= -1674190539;
assign addr[25982]= -1697875851;
assign addr[25983]= -1721022648;
assign addr[25984]= -1743623590;
assign addr[25985]= -1765671509;
assign addr[25986]= -1787159411;
assign addr[25987]= -1808080480;
assign addr[25988]= -1828428082;
assign addr[25989]= -1848195763;
assign addr[25990]= -1867377253;
assign addr[25991]= -1885966468;
assign addr[25992]= -1903957513;
assign addr[25993]= -1921344681;
assign addr[25994]= -1938122457;
assign addr[25995]= -1954285520;
assign addr[25996]= -1969828744;
assign addr[25997]= -1984747199;
assign addr[25998]= -1999036154;
assign addr[25999]= -2012691075;
assign addr[26000]= -2025707632;
assign addr[26001]= -2038081698;
assign addr[26002]= -2049809346;
assign addr[26003]= -2060886858;
assign addr[26004]= -2071310720;
assign addr[26005]= -2081077626;
assign addr[26006]= -2090184478;
assign addr[26007]= -2098628387;
assign addr[26008]= -2106406677;
assign addr[26009]= -2113516878;
assign addr[26010]= -2119956737;
assign addr[26011]= -2125724211;
assign addr[26012]= -2130817471;
assign addr[26013]= -2135234901;
assign addr[26014]= -2138975100;
assign addr[26015]= -2142036881;
assign addr[26016]= -2144419275;
assign addr[26017]= -2146121524;
assign addr[26018]= -2147143090;
assign addr[26019]= -2147483648;
assign addr[26020]= -2147143090;
assign addr[26021]= -2146121524;
assign addr[26022]= -2144419275;
assign addr[26023]= -2142036881;
assign addr[26024]= -2138975100;
assign addr[26025]= -2135234901;
assign addr[26026]= -2130817471;
assign addr[26027]= -2125724211;
assign addr[26028]= -2119956737;
assign addr[26029]= -2113516878;
assign addr[26030]= -2106406677;
assign addr[26031]= -2098628387;
assign addr[26032]= -2090184478;
assign addr[26033]= -2081077626;
assign addr[26034]= -2071310720;
assign addr[26035]= -2060886858;
assign addr[26036]= -2049809346;
assign addr[26037]= -2038081698;
assign addr[26038]= -2025707632;
assign addr[26039]= -2012691075;
assign addr[26040]= -1999036154;
assign addr[26041]= -1984747199;
assign addr[26042]= -1969828744;
assign addr[26043]= -1954285520;
assign addr[26044]= -1938122457;
assign addr[26045]= -1921344681;
assign addr[26046]= -1903957513;
assign addr[26047]= -1885966468;
assign addr[26048]= -1867377253;
assign addr[26049]= -1848195763;
assign addr[26050]= -1828428082;
assign addr[26051]= -1808080480;
assign addr[26052]= -1787159411;
assign addr[26053]= -1765671509;
assign addr[26054]= -1743623590;
assign addr[26055]= -1721022648;
assign addr[26056]= -1697875851;
assign addr[26057]= -1674190539;
assign addr[26058]= -1649974225;
assign addr[26059]= -1625234591;
assign addr[26060]= -1599979481;
assign addr[26061]= -1574216908;
assign addr[26062]= -1547955041;
assign addr[26063]= -1521202211;
assign addr[26064]= -1493966902;
assign addr[26065]= -1466257752;
assign addr[26066]= -1438083551;
assign addr[26067]= -1409453233;
assign addr[26068]= -1380375881;
assign addr[26069]= -1350860716;
assign addr[26070]= -1320917099;
assign addr[26071]= -1290554528;
assign addr[26072]= -1259782632;
assign addr[26073]= -1228611172;
assign addr[26074]= -1197050035;
assign addr[26075]= -1165109230;
assign addr[26076]= -1132798888;
assign addr[26077]= -1100129257;
assign addr[26078]= -1067110699;
assign addr[26079]= -1033753687;
assign addr[26080]= -1000068799;
assign addr[26081]= -966066720;
assign addr[26082]= -931758235;
assign addr[26083]= -897154224;
assign addr[26084]= -862265664;
assign addr[26085]= -827103620;
assign addr[26086]= -791679244;
assign addr[26087]= -756003771;
assign addr[26088]= -720088517;
assign addr[26089]= -683944874;
assign addr[26090]= -647584304;
assign addr[26091]= -611018340;
assign addr[26092]= -574258580;
assign addr[26093]= -537316682;
assign addr[26094]= -500204365;
assign addr[26095]= -462933398;
assign addr[26096]= -425515602;
assign addr[26097]= -387962847;
assign addr[26098]= -350287041;
assign addr[26099]= -312500135;
assign addr[26100]= -274614114;
assign addr[26101]= -236640993;
assign addr[26102]= -198592817;
assign addr[26103]= -160481654;
assign addr[26104]= -122319591;
assign addr[26105]= -84118732;
assign addr[26106]= -45891193;
assign addr[26107]= -7649098;
assign addr[26108]= 30595422;
assign addr[26109]= 68830239;
assign addr[26110]= 107043224;
assign addr[26111]= 145222259;
assign addr[26112]= 183355234;
assign addr[26113]= 221430054;
assign addr[26114]= 259434643;
assign addr[26115]= 297356948;
assign addr[26116]= 335184940;
assign addr[26117]= 372906622;
assign addr[26118]= 410510029;
assign addr[26119]= 447983235;
assign addr[26120]= 485314355;
assign addr[26121]= 522491548;
assign addr[26122]= 559503022;
assign addr[26123]= 596337040;
assign addr[26124]= 632981917;
assign addr[26125]= 669426032;
assign addr[26126]= 705657826;
assign addr[26127]= 741665807;
assign addr[26128]= 777438554;
assign addr[26129]= 812964722;
assign addr[26130]= 848233042;
assign addr[26131]= 883232329;
assign addr[26132]= 917951481;
assign addr[26133]= 952379488;
assign addr[26134]= 986505429;
assign addr[26135]= 1020318481;
assign addr[26136]= 1053807919;
assign addr[26137]= 1086963121;
assign addr[26138]= 1119773573;
assign addr[26139]= 1152228866;
assign addr[26140]= 1184318708;
assign addr[26141]= 1216032921;
assign addr[26142]= 1247361445;
assign addr[26143]= 1278294345;
assign addr[26144]= 1308821808;
assign addr[26145]= 1338934154;
assign addr[26146]= 1368621831;
assign addr[26147]= 1397875423;
assign addr[26148]= 1426685652;
assign addr[26149]= 1455043381;
assign addr[26150]= 1482939614;
assign addr[26151]= 1510365504;
assign addr[26152]= 1537312353;
assign addr[26153]= 1563771613;
assign addr[26154]= 1589734894;
assign addr[26155]= 1615193959;
assign addr[26156]= 1640140734;
assign addr[26157]= 1664567307;
assign addr[26158]= 1688465931;
assign addr[26159]= 1711829025;
assign addr[26160]= 1734649179;
assign addr[26161]= 1756919156;
assign addr[26162]= 1778631892;
assign addr[26163]= 1799780501;
assign addr[26164]= 1820358275;
assign addr[26165]= 1840358687;
assign addr[26166]= 1859775393;
assign addr[26167]= 1878602237;
assign addr[26168]= 1896833245;
assign addr[26169]= 1914462636;
assign addr[26170]= 1931484818;
assign addr[26171]= 1947894393;
assign addr[26172]= 1963686155;
assign addr[26173]= 1978855097;
assign addr[26174]= 1993396407;
assign addr[26175]= 2007305472;
assign addr[26176]= 2020577882;
assign addr[26177]= 2033209426;
assign addr[26178]= 2045196100;
assign addr[26179]= 2056534099;
assign addr[26180]= 2067219829;
assign addr[26181]= 2077249901;
assign addr[26182]= 2086621133;
assign addr[26183]= 2095330553;
assign addr[26184]= 2103375398;
assign addr[26185]= 2110753117;
assign addr[26186]= 2117461370;
assign addr[26187]= 2123498030;
assign addr[26188]= 2128861181;
assign addr[26189]= 2133549123;
assign addr[26190]= 2137560369;
assign addr[26191]= 2140893646;
assign addr[26192]= 2143547897;
assign addr[26193]= 2145522281;
assign addr[26194]= 2146816171;
assign addr[26195]= 2147429158;
assign addr[26196]= 2147361045;
assign addr[26197]= 2146611856;
assign addr[26198]= 2145181827;
assign addr[26199]= 2143071413;
assign addr[26200]= 2140281282;
assign addr[26201]= 2136812319;
assign addr[26202]= 2132665626;
assign addr[26203]= 2127842516;
assign addr[26204]= 2122344521;
assign addr[26205]= 2116173382;
assign addr[26206]= 2109331059;
assign addr[26207]= 2101819720;
assign addr[26208]= 2093641749;
assign addr[26209]= 2084799740;
assign addr[26210]= 2075296495;
assign addr[26211]= 2065135031;
assign addr[26212]= 2054318569;
assign addr[26213]= 2042850540;
assign addr[26214]= 2030734582;
assign addr[26215]= 2017974537;
assign addr[26216]= 2004574453;
assign addr[26217]= 1990538579;
assign addr[26218]= 1975871368;
assign addr[26219]= 1960577471;
assign addr[26220]= 1944661739;
assign addr[26221]= 1928129220;
assign addr[26222]= 1910985158;
assign addr[26223]= 1893234990;
assign addr[26224]= 1874884346;
assign addr[26225]= 1855939047;
assign addr[26226]= 1836405100;
assign addr[26227]= 1816288703;
assign addr[26228]= 1795596234;
assign addr[26229]= 1774334257;
assign addr[26230]= 1752509516;
assign addr[26231]= 1730128933;
assign addr[26232]= 1707199606;
assign addr[26233]= 1683728808;
assign addr[26234]= 1659723983;
assign addr[26235]= 1635192744;
assign addr[26236]= 1610142873;
assign addr[26237]= 1584582314;
assign addr[26238]= 1558519173;
assign addr[26239]= 1531961719;
assign addr[26240]= 1504918373;
assign addr[26241]= 1477397714;
assign addr[26242]= 1449408469;
assign addr[26243]= 1420959516;
assign addr[26244]= 1392059879;
assign addr[26245]= 1362718723;
assign addr[26246]= 1332945355;
assign addr[26247]= 1302749217;
assign addr[26248]= 1272139887;
assign addr[26249]= 1241127074;
assign addr[26250]= 1209720613;
assign addr[26251]= 1177930466;
assign addr[26252]= 1145766716;
assign addr[26253]= 1113239564;
assign addr[26254]= 1080359326;
assign addr[26255]= 1047136432;
assign addr[26256]= 1013581418;
assign addr[26257]= 979704927;
assign addr[26258]= 945517704;
assign addr[26259]= 911030591;
assign addr[26260]= 876254528;
assign addr[26261]= 841200544;
assign addr[26262]= 805879757;
assign addr[26263]= 770303369;
assign addr[26264]= 734482665;
assign addr[26265]= 698429006;
assign addr[26266]= 662153826;
assign addr[26267]= 625668632;
assign addr[26268]= 588984994;
assign addr[26269]= 552114549;
assign addr[26270]= 515068990;
assign addr[26271]= 477860067;
assign addr[26272]= 440499581;
assign addr[26273]= 402999383;
assign addr[26274]= 365371365;
assign addr[26275]= 327627463;
assign addr[26276]= 289779648;
assign addr[26277]= 251839923;
assign addr[26278]= 213820322;
assign addr[26279]= 175732905;
assign addr[26280]= 137589750;
assign addr[26281]= 99402956;
assign addr[26282]= 61184634;
assign addr[26283]= 22946906;
assign addr[26284]= -15298099;
assign addr[26285]= -53538253;
assign addr[26286]= -91761426;
assign addr[26287]= -129955495;
assign addr[26288]= -168108346;
assign addr[26289]= -206207878;
assign addr[26290]= -244242007;
assign addr[26291]= -282198671;
assign addr[26292]= -320065829;
assign addr[26293]= -357831473;
assign addr[26294]= -395483624;
assign addr[26295]= -433010339;
assign addr[26296]= -470399716;
assign addr[26297]= -507639898;
assign addr[26298]= -544719071;
assign addr[26299]= -581625477;
assign addr[26300]= -618347408;
assign addr[26301]= -654873219;
assign addr[26302]= -691191324;
assign addr[26303]= -727290205;
assign addr[26304]= -763158411;
assign addr[26305]= -798784567;
assign addr[26306]= -834157373;
assign addr[26307]= -869265610;
assign addr[26308]= -904098143;
assign addr[26309]= -938643924;
assign addr[26310]= -972891995;
assign addr[26311]= -1006831495;
assign addr[26312]= -1040451659;
assign addr[26313]= -1073741824;
assign addr[26314]= -1106691431;
assign addr[26315]= -1139290029;
assign addr[26316]= -1171527280;
assign addr[26317]= -1203392958;
assign addr[26318]= -1234876957;
assign addr[26319]= -1265969291;
assign addr[26320]= -1296660098;
assign addr[26321]= -1326939644;
assign addr[26322]= -1356798326;
assign addr[26323]= -1386226674;
assign addr[26324]= -1415215352;
assign addr[26325]= -1443755168;
assign addr[26326]= -1471837070;
assign addr[26327]= -1499452149;
assign addr[26328]= -1526591649;
assign addr[26329]= -1553246960;
assign addr[26330]= -1579409630;
assign addr[26331]= -1605071359;
assign addr[26332]= -1630224009;
assign addr[26333]= -1654859602;
assign addr[26334]= -1678970324;
assign addr[26335]= -1702548529;
assign addr[26336]= -1725586737;
assign addr[26337]= -1748077642;
assign addr[26338]= -1770014111;
assign addr[26339]= -1791389186;
assign addr[26340]= -1812196087;
assign addr[26341]= -1832428215;
assign addr[26342]= -1852079154;
assign addr[26343]= -1871142669;
assign addr[26344]= -1889612716;
assign addr[26345]= -1907483436;
assign addr[26346]= -1924749160;
assign addr[26347]= -1941404413;
assign addr[26348]= -1957443913;
assign addr[26349]= -1972862571;
assign addr[26350]= -1987655498;
assign addr[26351]= -2001818002;
assign addr[26352]= -2015345591;
assign addr[26353]= -2028233973;
assign addr[26354]= -2040479063;
assign addr[26355]= -2052076975;
assign addr[26356]= -2063024031;
assign addr[26357]= -2073316760;
assign addr[26358]= -2082951896;
assign addr[26359]= -2091926384;
assign addr[26360]= -2100237377;
assign addr[26361]= -2107882239;
assign addr[26362]= -2114858546;
assign addr[26363]= -2121164085;
assign addr[26364]= -2126796855;
assign addr[26365]= -2131755071;
assign addr[26366]= -2136037160;
assign addr[26367]= -2139641764;
assign addr[26368]= -2142567738;
assign addr[26369]= -2144814157;
assign addr[26370]= -2146380306;
assign addr[26371]= -2147265689;
assign addr[26372]= -2147470025;
assign addr[26373]= -2146993250;
assign addr[26374]= -2145835515;
assign addr[26375]= -2143997187;
assign addr[26376]= -2141478848;
assign addr[26377]= -2138281298;
assign addr[26378]= -2134405552;
assign addr[26379]= -2129852837;
assign addr[26380]= -2124624598;
assign addr[26381]= -2118722494;
assign addr[26382]= -2112148396;
assign addr[26383]= -2104904390;
assign addr[26384]= -2096992772;
assign addr[26385]= -2088416053;
assign addr[26386]= -2079176953;
assign addr[26387]= -2069278401;
assign addr[26388]= -2058723538;
assign addr[26389]= -2047515711;
assign addr[26390]= -2035658475;
assign addr[26391]= -2023155591;
assign addr[26392]= -2010011024;
assign addr[26393]= -1996228943;
assign addr[26394]= -1981813720;
assign addr[26395]= -1966769926;
assign addr[26396]= -1951102334;
assign addr[26397]= -1934815911;
assign addr[26398]= -1917915825;
assign addr[26399]= -1900407434;
assign addr[26400]= -1882296293;
assign addr[26401]= -1863588145;
assign addr[26402]= -1844288924;
assign addr[26403]= -1824404752;
assign addr[26404]= -1803941934;
assign addr[26405]= -1782906961;
assign addr[26406]= -1761306505;
assign addr[26407]= -1739147417;
assign addr[26408]= -1716436725;
assign addr[26409]= -1693181631;
assign addr[26410]= -1669389513;
assign addr[26411]= -1645067915;
assign addr[26412]= -1620224553;
assign addr[26413]= -1594867305;
assign addr[26414]= -1569004214;
assign addr[26415]= -1542643483;
assign addr[26416]= -1515793473;
assign addr[26417]= -1488462700;
assign addr[26418]= -1460659832;
assign addr[26419]= -1432393688;
assign addr[26420]= -1403673233;
assign addr[26421]= -1374507575;
assign addr[26422]= -1344905966;
assign addr[26423]= -1314877795;
assign addr[26424]= -1284432584;
assign addr[26425]= -1253579991;
assign addr[26426]= -1222329801;
assign addr[26427]= -1190691925;
assign addr[26428]= -1158676398;
assign addr[26429]= -1126293375;
assign addr[26430]= -1093553126;
assign addr[26431]= -1060466036;
assign addr[26432]= -1027042599;
assign addr[26433]= -993293415;
assign addr[26434]= -959229189;
assign addr[26435]= -924860725;
assign addr[26436]= -890198924;
assign addr[26437]= -855254778;
assign addr[26438]= -820039373;
assign addr[26439]= -784563876;
assign addr[26440]= -748839539;
assign addr[26441]= -712877694;
assign addr[26442]= -676689746;
assign addr[26443]= -640287172;
assign addr[26444]= -603681519;
assign addr[26445]= -566884397;
assign addr[26446]= -529907477;
assign addr[26447]= -492762486;
assign addr[26448]= -455461206;
assign addr[26449]= -418015468;
assign addr[26450]= -380437148;
assign addr[26451]= -342738165;
assign addr[26452]= -304930476;
assign addr[26453]= -267026072;
assign addr[26454]= -229036977;
assign addr[26455]= -190975237;
assign addr[26456]= -152852926;
assign addr[26457]= -114682135;
assign addr[26458]= -76474970;
assign addr[26459]= -38243550;
assign addr[26460]= 0;
assign addr[26461]= 38243550;
assign addr[26462]= 76474970;
assign addr[26463]= 114682135;
assign addr[26464]= 152852926;
assign addr[26465]= 190975237;
assign addr[26466]= 229036977;
assign addr[26467]= 267026072;
assign addr[26468]= 304930476;
assign addr[26469]= 342738165;
assign addr[26470]= 380437148;
assign addr[26471]= 418015468;
assign addr[26472]= 455461206;
assign addr[26473]= 492762486;
assign addr[26474]= 529907477;
assign addr[26475]= 566884397;
assign addr[26476]= 603681519;
assign addr[26477]= 640287172;
assign addr[26478]= 676689746;
assign addr[26479]= 712877694;
assign addr[26480]= 748839539;
assign addr[26481]= 784563876;
assign addr[26482]= 820039373;
assign addr[26483]= 855254778;
assign addr[26484]= 890198924;
assign addr[26485]= 924860725;
assign addr[26486]= 959229189;
assign addr[26487]= 993293415;
assign addr[26488]= 1027042599;
assign addr[26489]= 1060466036;
assign addr[26490]= 1093553126;
assign addr[26491]= 1126293375;
assign addr[26492]= 1158676398;
assign addr[26493]= 1190691925;
assign addr[26494]= 1222329801;
assign addr[26495]= 1253579991;
assign addr[26496]= 1284432584;
assign addr[26497]= 1314877795;
assign addr[26498]= 1344905966;
assign addr[26499]= 1374507575;
assign addr[26500]= 1403673233;
assign addr[26501]= 1432393688;
assign addr[26502]= 1460659832;
assign addr[26503]= 1488462700;
assign addr[26504]= 1515793473;
assign addr[26505]= 1542643483;
assign addr[26506]= 1569004214;
assign addr[26507]= 1594867305;
assign addr[26508]= 1620224553;
assign addr[26509]= 1645067915;
assign addr[26510]= 1669389513;
assign addr[26511]= 1693181631;
assign addr[26512]= 1716436725;
assign addr[26513]= 1739147417;
assign addr[26514]= 1761306505;
assign addr[26515]= 1782906961;
assign addr[26516]= 1803941934;
assign addr[26517]= 1824404752;
assign addr[26518]= 1844288924;
assign addr[26519]= 1863588145;
assign addr[26520]= 1882296293;
assign addr[26521]= 1900407434;
assign addr[26522]= 1917915825;
assign addr[26523]= 1934815911;
assign addr[26524]= 1951102334;
assign addr[26525]= 1966769926;
assign addr[26526]= 1981813720;
assign addr[26527]= 1996228943;
assign addr[26528]= 2010011024;
assign addr[26529]= 2023155591;
assign addr[26530]= 2035658475;
assign addr[26531]= 2047515711;
assign addr[26532]= 2058723538;
assign addr[26533]= 2069278401;
assign addr[26534]= 2079176953;
assign addr[26535]= 2088416053;
assign addr[26536]= 2096992772;
assign addr[26537]= 2104904390;
assign addr[26538]= 2112148396;
assign addr[26539]= 2118722494;
assign addr[26540]= 2124624598;
assign addr[26541]= 2129852837;
assign addr[26542]= 2134405552;
assign addr[26543]= 2138281298;
assign addr[26544]= 2141478848;
assign addr[26545]= 2143997187;
assign addr[26546]= 2145835515;
assign addr[26547]= 2146993250;
assign addr[26548]= 2147470025;
assign addr[26549]= 2147265689;
assign addr[26550]= 2146380306;
assign addr[26551]= 2144814157;
assign addr[26552]= 2142567738;
assign addr[26553]= 2139641764;
assign addr[26554]= 2136037160;
assign addr[26555]= 2131755071;
assign addr[26556]= 2126796855;
assign addr[26557]= 2121164085;
assign addr[26558]= 2114858546;
assign addr[26559]= 2107882239;
assign addr[26560]= 2100237377;
assign addr[26561]= 2091926384;
assign addr[26562]= 2082951896;
assign addr[26563]= 2073316760;
assign addr[26564]= 2063024031;
assign addr[26565]= 2052076975;
assign addr[26566]= 2040479063;
assign addr[26567]= 2028233973;
assign addr[26568]= 2015345591;
assign addr[26569]= 2001818002;
assign addr[26570]= 1987655498;
assign addr[26571]= 1972862571;
assign addr[26572]= 1957443913;
assign addr[26573]= 1941404413;
assign addr[26574]= 1924749160;
assign addr[26575]= 1907483436;
assign addr[26576]= 1889612716;
assign addr[26577]= 1871142669;
assign addr[26578]= 1852079154;
assign addr[26579]= 1832428215;
assign addr[26580]= 1812196087;
assign addr[26581]= 1791389186;
assign addr[26582]= 1770014111;
assign addr[26583]= 1748077642;
assign addr[26584]= 1725586737;
assign addr[26585]= 1702548529;
assign addr[26586]= 1678970324;
assign addr[26587]= 1654859602;
assign addr[26588]= 1630224009;
assign addr[26589]= 1605071359;
assign addr[26590]= 1579409630;
assign addr[26591]= 1553246960;
assign addr[26592]= 1526591649;
assign addr[26593]= 1499452149;
assign addr[26594]= 1471837070;
assign addr[26595]= 1443755168;
assign addr[26596]= 1415215352;
assign addr[26597]= 1386226674;
assign addr[26598]= 1356798326;
assign addr[26599]= 1326939644;
assign addr[26600]= 1296660098;
assign addr[26601]= 1265969291;
assign addr[26602]= 1234876957;
assign addr[26603]= 1203392958;
assign addr[26604]= 1171527280;
assign addr[26605]= 1139290029;
assign addr[26606]= 1106691431;
assign addr[26607]= 1073741824;
assign addr[26608]= 1040451659;
assign addr[26609]= 1006831495;
assign addr[26610]= 972891995;
assign addr[26611]= 938643924;
assign addr[26612]= 904098143;
assign addr[26613]= 869265610;
assign addr[26614]= 834157373;
assign addr[26615]= 798784567;
assign addr[26616]= 763158411;
assign addr[26617]= 727290205;
assign addr[26618]= 691191324;
assign addr[26619]= 654873219;
assign addr[26620]= 618347408;
assign addr[26621]= 581625477;
assign addr[26622]= 544719071;
assign addr[26623]= 507639898;
assign addr[26624]= 470399716;
assign addr[26625]= 433010339;
assign addr[26626]= 395483624;
assign addr[26627]= 357831473;
assign addr[26628]= 320065829;
assign addr[26629]= 282198671;
assign addr[26630]= 244242007;
assign addr[26631]= 206207878;
assign addr[26632]= 168108346;
assign addr[26633]= 129955495;
assign addr[26634]= 91761426;
assign addr[26635]= 53538253;
assign addr[26636]= 15298099;
assign addr[26637]= -22946906;
assign addr[26638]= -61184634;
assign addr[26639]= -99402956;
assign addr[26640]= -137589750;
assign addr[26641]= -175732905;
assign addr[26642]= -213820322;
assign addr[26643]= -251839923;
assign addr[26644]= -289779648;
assign addr[26645]= -327627463;
assign addr[26646]= -365371365;
assign addr[26647]= -402999383;
assign addr[26648]= -440499581;
assign addr[26649]= -477860067;
assign addr[26650]= -515068990;
assign addr[26651]= -552114549;
assign addr[26652]= -588984994;
assign addr[26653]= -625668632;
assign addr[26654]= -662153826;
assign addr[26655]= -698429006;
assign addr[26656]= -734482665;
assign addr[26657]= -770303369;
assign addr[26658]= -805879757;
assign addr[26659]= -841200544;
assign addr[26660]= -876254528;
assign addr[26661]= -911030591;
assign addr[26662]= -945517704;
assign addr[26663]= -979704927;
assign addr[26664]= -1013581418;
assign addr[26665]= -1047136432;
assign addr[26666]= -1080359326;
assign addr[26667]= -1113239564;
assign addr[26668]= -1145766716;
assign addr[26669]= -1177930466;
assign addr[26670]= -1209720613;
assign addr[26671]= -1241127074;
assign addr[26672]= -1272139887;
assign addr[26673]= -1302749217;
assign addr[26674]= -1332945355;
assign addr[26675]= -1362718723;
assign addr[26676]= -1392059879;
assign addr[26677]= -1420959516;
assign addr[26678]= -1449408469;
assign addr[26679]= -1477397714;
assign addr[26680]= -1504918373;
assign addr[26681]= -1531961719;
assign addr[26682]= -1558519173;
assign addr[26683]= -1584582314;
assign addr[26684]= -1610142873;
assign addr[26685]= -1635192744;
assign addr[26686]= -1659723983;
assign addr[26687]= -1683728808;
assign addr[26688]= -1707199606;
assign addr[26689]= -1730128933;
assign addr[26690]= -1752509516;
assign addr[26691]= -1774334257;
assign addr[26692]= -1795596234;
assign addr[26693]= -1816288703;
assign addr[26694]= -1836405100;
assign addr[26695]= -1855939047;
assign addr[26696]= -1874884346;
assign addr[26697]= -1893234990;
assign addr[26698]= -1910985158;
assign addr[26699]= -1928129220;
assign addr[26700]= -1944661739;
assign addr[26701]= -1960577471;
assign addr[26702]= -1975871368;
assign addr[26703]= -1990538579;
assign addr[26704]= -2004574453;
assign addr[26705]= -2017974537;
assign addr[26706]= -2030734582;
assign addr[26707]= -2042850540;
assign addr[26708]= -2054318569;
assign addr[26709]= -2065135031;
assign addr[26710]= -2075296495;
assign addr[26711]= -2084799740;
assign addr[26712]= -2093641749;
assign addr[26713]= -2101819720;
assign addr[26714]= -2109331059;
assign addr[26715]= -2116173382;
assign addr[26716]= -2122344521;
assign addr[26717]= -2127842516;
assign addr[26718]= -2132665626;
assign addr[26719]= -2136812319;
assign addr[26720]= -2140281282;
assign addr[26721]= -2143071413;
assign addr[26722]= -2145181827;
assign addr[26723]= -2146611856;
assign addr[26724]= -2147361045;
assign addr[26725]= -2147429158;
assign addr[26726]= -2146816171;
assign addr[26727]= -2145522281;
assign addr[26728]= -2143547897;
assign addr[26729]= -2140893646;
assign addr[26730]= -2137560369;
assign addr[26731]= -2133549123;
assign addr[26732]= -2128861181;
assign addr[26733]= -2123498030;
assign addr[26734]= -2117461370;
assign addr[26735]= -2110753117;
assign addr[26736]= -2103375398;
assign addr[26737]= -2095330553;
assign addr[26738]= -2086621133;
assign addr[26739]= -2077249901;
assign addr[26740]= -2067219829;
assign addr[26741]= -2056534099;
assign addr[26742]= -2045196100;
assign addr[26743]= -2033209426;
assign addr[26744]= -2020577882;
assign addr[26745]= -2007305472;
assign addr[26746]= -1993396407;
assign addr[26747]= -1978855097;
assign addr[26748]= -1963686155;
assign addr[26749]= -1947894393;
assign addr[26750]= -1931484818;
assign addr[26751]= -1914462636;
assign addr[26752]= -1896833245;
assign addr[26753]= -1878602237;
assign addr[26754]= -1859775393;
assign addr[26755]= -1840358687;
assign addr[26756]= -1820358275;
assign addr[26757]= -1799780501;
assign addr[26758]= -1778631892;
assign addr[26759]= -1756919156;
assign addr[26760]= -1734649179;
assign addr[26761]= -1711829025;
assign addr[26762]= -1688465931;
assign addr[26763]= -1664567307;
assign addr[26764]= -1640140734;
assign addr[26765]= -1615193959;
assign addr[26766]= -1589734894;
assign addr[26767]= -1563771613;
assign addr[26768]= -1537312353;
assign addr[26769]= -1510365504;
assign addr[26770]= -1482939614;
assign addr[26771]= -1455043381;
assign addr[26772]= -1426685652;
assign addr[26773]= -1397875423;
assign addr[26774]= -1368621831;
assign addr[26775]= -1338934154;
assign addr[26776]= -1308821808;
assign addr[26777]= -1278294345;
assign addr[26778]= -1247361445;
assign addr[26779]= -1216032921;
assign addr[26780]= -1184318708;
assign addr[26781]= -1152228866;
assign addr[26782]= -1119773573;
assign addr[26783]= -1086963121;
assign addr[26784]= -1053807919;
assign addr[26785]= -1020318481;
assign addr[26786]= -986505429;
assign addr[26787]= -952379488;
assign addr[26788]= -917951481;
assign addr[26789]= -883232329;
assign addr[26790]= -848233042;
assign addr[26791]= -812964722;
assign addr[26792]= -777438554;
assign addr[26793]= -741665807;
assign addr[26794]= -705657826;
assign addr[26795]= -669426032;
assign addr[26796]= -632981917;
assign addr[26797]= -596337040;
assign addr[26798]= -559503022;
assign addr[26799]= -522491548;
assign addr[26800]= -485314355;
assign addr[26801]= -447983235;
assign addr[26802]= -410510029;
assign addr[26803]= -372906622;
assign addr[26804]= -335184940;
assign addr[26805]= -297356948;
assign addr[26806]= -259434643;
assign addr[26807]= -221430054;
assign addr[26808]= -183355234;
assign addr[26809]= -145222259;
assign addr[26810]= -107043224;
assign addr[26811]= -68830239;
assign addr[26812]= -30595422;
assign addr[26813]= 7649098;
assign addr[26814]= 45891193;
assign addr[26815]= 84118732;
assign addr[26816]= 122319591;
assign addr[26817]= 160481654;
assign addr[26818]= 198592817;
assign addr[26819]= 236640993;
assign addr[26820]= 274614114;
assign addr[26821]= 312500135;
assign addr[26822]= 350287041;
assign addr[26823]= 387962847;
assign addr[26824]= 425515602;
assign addr[26825]= 462933398;
assign addr[26826]= 500204365;
assign addr[26827]= 537316682;
assign addr[26828]= 574258580;
assign addr[26829]= 611018340;
assign addr[26830]= 647584304;
assign addr[26831]= 683944874;
assign addr[26832]= 720088517;
assign addr[26833]= 756003771;
assign addr[26834]= 791679244;
assign addr[26835]= 827103620;
assign addr[26836]= 862265664;
assign addr[26837]= 897154224;
assign addr[26838]= 931758235;
assign addr[26839]= 966066720;
assign addr[26840]= 1000068799;
assign addr[26841]= 1033753687;
assign addr[26842]= 1067110699;
assign addr[26843]= 1100129257;
assign addr[26844]= 1132798888;
assign addr[26845]= 1165109230;
assign addr[26846]= 1197050035;
assign addr[26847]= 1228611172;
assign addr[26848]= 1259782632;
assign addr[26849]= 1290554528;
assign addr[26850]= 1320917099;
assign addr[26851]= 1350860716;
assign addr[26852]= 1380375881;
assign addr[26853]= 1409453233;
assign addr[26854]= 1438083551;
assign addr[26855]= 1466257752;
assign addr[26856]= 1493966902;
assign addr[26857]= 1521202211;
assign addr[26858]= 1547955041;
assign addr[26859]= 1574216908;
assign addr[26860]= 1599979481;
assign addr[26861]= 1625234591;
assign addr[26862]= 1649974225;
assign addr[26863]= 1674190539;
assign addr[26864]= 1697875851;
assign addr[26865]= 1721022648;
assign addr[26866]= 1743623590;
assign addr[26867]= 1765671509;
assign addr[26868]= 1787159411;
assign addr[26869]= 1808080480;
assign addr[26870]= 1828428082;
assign addr[26871]= 1848195763;
assign addr[26872]= 1867377253;
assign addr[26873]= 1885966468;
assign addr[26874]= 1903957513;
assign addr[26875]= 1921344681;
assign addr[26876]= 1938122457;
assign addr[26877]= 1954285520;
assign addr[26878]= 1969828744;
assign addr[26879]= 1984747199;
assign addr[26880]= 1999036154;
assign addr[26881]= 2012691075;
assign addr[26882]= 2025707632;
assign addr[26883]= 2038081698;
assign addr[26884]= 2049809346;
assign addr[26885]= 2060886858;
assign addr[26886]= 2071310720;
assign addr[26887]= 2081077626;
assign addr[26888]= 2090184478;
assign addr[26889]= 2098628387;
assign addr[26890]= 2106406677;
assign addr[26891]= 2113516878;
assign addr[26892]= 2119956737;
assign addr[26893]= 2125724211;
assign addr[26894]= 2130817471;
assign addr[26895]= 2135234901;
assign addr[26896]= 2138975100;
assign addr[26897]= 2142036881;
assign addr[26898]= 2144419275;
assign addr[26899]= 2146121524;
assign addr[26900]= 2147143090;
assign addr[26901]= 2147483648;
assign addr[26902]= 2147143090;
assign addr[26903]= 2146121524;
assign addr[26904]= 2144419275;
assign addr[26905]= 2142036881;
assign addr[26906]= 2138975100;
assign addr[26907]= 2135234901;
assign addr[26908]= 2130817471;
assign addr[26909]= 2125724211;
assign addr[26910]= 2119956737;
assign addr[26911]= 2113516878;
assign addr[26912]= 2106406677;
assign addr[26913]= 2098628387;
assign addr[26914]= 2090184478;
assign addr[26915]= 2081077626;
assign addr[26916]= 2071310720;
assign addr[26917]= 2060886858;
assign addr[26918]= 2049809346;
assign addr[26919]= 2038081698;
assign addr[26920]= 2025707632;
assign addr[26921]= 2012691075;
assign addr[26922]= 1999036154;
assign addr[26923]= 1984747199;
assign addr[26924]= 1969828744;
assign addr[26925]= 1954285520;
assign addr[26926]= 1938122457;
assign addr[26927]= 1921344681;
assign addr[26928]= 1903957513;
assign addr[26929]= 1885966468;
assign addr[26930]= 1867377253;
assign addr[26931]= 1848195763;
assign addr[26932]= 1828428082;
assign addr[26933]= 1808080480;
assign addr[26934]= 1787159411;
assign addr[26935]= 1765671509;
assign addr[26936]= 1743623590;
assign addr[26937]= 1721022648;
assign addr[26938]= 1697875851;
assign addr[26939]= 1674190539;
assign addr[26940]= 1649974225;
assign addr[26941]= 1625234591;
assign addr[26942]= 1599979481;
assign addr[26943]= 1574216908;
assign addr[26944]= 1547955041;
assign addr[26945]= 1521202211;
assign addr[26946]= 1493966902;
assign addr[26947]= 1466257752;
assign addr[26948]= 1438083551;
assign addr[26949]= 1409453233;
assign addr[26950]= 1380375881;
assign addr[26951]= 1350860716;
assign addr[26952]= 1320917099;
assign addr[26953]= 1290554528;
assign addr[26954]= 1259782632;
assign addr[26955]= 1228611172;
assign addr[26956]= 1197050035;
assign addr[26957]= 1165109230;
assign addr[26958]= 1132798888;
assign addr[26959]= 1100129257;
assign addr[26960]= 1067110699;
assign addr[26961]= 1033753687;
assign addr[26962]= 1000068799;
assign addr[26963]= 966066720;
assign addr[26964]= 931758235;
assign addr[26965]= 897154224;
assign addr[26966]= 862265664;
assign addr[26967]= 827103620;
assign addr[26968]= 791679244;
assign addr[26969]= 756003771;
assign addr[26970]= 720088517;
assign addr[26971]= 683944874;
assign addr[26972]= 647584304;
assign addr[26973]= 611018340;
assign addr[26974]= 574258580;
assign addr[26975]= 537316682;
assign addr[26976]= 500204365;
assign addr[26977]= 462933398;
assign addr[26978]= 425515602;
assign addr[26979]= 387962847;
assign addr[26980]= 350287041;
assign addr[26981]= 312500135;
assign addr[26982]= 274614114;
assign addr[26983]= 236640993;
assign addr[26984]= 198592817;
assign addr[26985]= 160481654;
assign addr[26986]= 122319591;
assign addr[26987]= 84118732;
assign addr[26988]= 45891193;
assign addr[26989]= 7649098;
assign addr[26990]= -30595422;
assign addr[26991]= -68830239;
assign addr[26992]= -107043224;
assign addr[26993]= -145222259;
assign addr[26994]= -183355234;
assign addr[26995]= -221430054;
assign addr[26996]= -259434643;
assign addr[26997]= -297356948;
assign addr[26998]= -335184940;
assign addr[26999]= -372906622;
assign addr[27000]= -410510029;
assign addr[27001]= -447983235;
assign addr[27002]= -485314355;
assign addr[27003]= -522491548;
assign addr[27004]= -559503022;
assign addr[27005]= -596337040;
assign addr[27006]= -632981917;
assign addr[27007]= -669426032;
assign addr[27008]= -705657826;
assign addr[27009]= -741665807;
assign addr[27010]= -777438554;
assign addr[27011]= -812964722;
assign addr[27012]= -848233042;
assign addr[27013]= -883232329;
assign addr[27014]= -917951481;
assign addr[27015]= -952379488;
assign addr[27016]= -986505429;
assign addr[27017]= -1020318481;
assign addr[27018]= -1053807919;
assign addr[27019]= -1086963121;
assign addr[27020]= -1119773573;
assign addr[27021]= -1152228866;
assign addr[27022]= -1184318708;
assign addr[27023]= -1216032921;
assign addr[27024]= -1247361445;
assign addr[27025]= -1278294345;
assign addr[27026]= -1308821808;
assign addr[27027]= -1338934154;
assign addr[27028]= -1368621831;
assign addr[27029]= -1397875423;
assign addr[27030]= -1426685652;
assign addr[27031]= -1455043381;
assign addr[27032]= -1482939614;
assign addr[27033]= -1510365504;
assign addr[27034]= -1537312353;
assign addr[27035]= -1563771613;
assign addr[27036]= -1589734894;
assign addr[27037]= -1615193959;
assign addr[27038]= -1640140734;
assign addr[27039]= -1664567307;
assign addr[27040]= -1688465931;
assign addr[27041]= -1711829025;
assign addr[27042]= -1734649179;
assign addr[27043]= -1756919156;
assign addr[27044]= -1778631892;
assign addr[27045]= -1799780501;
assign addr[27046]= -1820358275;
assign addr[27047]= -1840358687;
assign addr[27048]= -1859775393;
assign addr[27049]= -1878602237;
assign addr[27050]= -1896833245;
assign addr[27051]= -1914462636;
assign addr[27052]= -1931484818;
assign addr[27053]= -1947894393;
assign addr[27054]= -1963686155;
assign addr[27055]= -1978855097;
assign addr[27056]= -1993396407;
assign addr[27057]= -2007305472;
assign addr[27058]= -2020577882;
assign addr[27059]= -2033209426;
assign addr[27060]= -2045196100;
assign addr[27061]= -2056534099;
assign addr[27062]= -2067219829;
assign addr[27063]= -2077249901;
assign addr[27064]= -2086621133;
assign addr[27065]= -2095330553;
assign addr[27066]= -2103375398;
assign addr[27067]= -2110753117;
assign addr[27068]= -2117461370;
assign addr[27069]= -2123498030;
assign addr[27070]= -2128861181;
assign addr[27071]= -2133549123;
assign addr[27072]= -2137560369;
assign addr[27073]= -2140893646;
assign addr[27074]= -2143547897;
assign addr[27075]= -2145522281;
assign addr[27076]= -2146816171;
assign addr[27077]= -2147429158;
assign addr[27078]= -2147361045;
assign addr[27079]= -2146611856;
assign addr[27080]= -2145181827;
assign addr[27081]= -2143071413;
assign addr[27082]= -2140281282;
assign addr[27083]= -2136812319;
assign addr[27084]= -2132665626;
assign addr[27085]= -2127842516;
assign addr[27086]= -2122344521;
assign addr[27087]= -2116173382;
assign addr[27088]= -2109331059;
assign addr[27089]= -2101819720;
assign addr[27090]= -2093641749;
assign addr[27091]= -2084799740;
assign addr[27092]= -2075296495;
assign addr[27093]= -2065135031;
assign addr[27094]= -2054318569;
assign addr[27095]= -2042850540;
assign addr[27096]= -2030734582;
assign addr[27097]= -2017974537;
assign addr[27098]= -2004574453;
assign addr[27099]= -1990538579;
assign addr[27100]= -1975871368;
assign addr[27101]= -1960577471;
assign addr[27102]= -1944661739;
assign addr[27103]= -1928129220;
assign addr[27104]= -1910985158;
assign addr[27105]= -1893234990;
assign addr[27106]= -1874884346;
assign addr[27107]= -1855939047;
assign addr[27108]= -1836405100;
assign addr[27109]= -1816288703;
assign addr[27110]= -1795596234;
assign addr[27111]= -1774334257;
assign addr[27112]= -1752509516;
assign addr[27113]= -1730128933;
assign addr[27114]= -1707199606;
assign addr[27115]= -1683728808;
assign addr[27116]= -1659723983;
assign addr[27117]= -1635192744;
assign addr[27118]= -1610142873;
assign addr[27119]= -1584582314;
assign addr[27120]= -1558519173;
assign addr[27121]= -1531961719;
assign addr[27122]= -1504918373;
assign addr[27123]= -1477397714;
assign addr[27124]= -1449408469;
assign addr[27125]= -1420959516;
assign addr[27126]= -1392059879;
assign addr[27127]= -1362718723;
assign addr[27128]= -1332945355;
assign addr[27129]= -1302749217;
assign addr[27130]= -1272139887;
assign addr[27131]= -1241127074;
assign addr[27132]= -1209720613;
assign addr[27133]= -1177930466;
assign addr[27134]= -1145766716;
assign addr[27135]= -1113239564;
assign addr[27136]= -1080359326;
assign addr[27137]= -1047136432;
assign addr[27138]= -1013581418;
assign addr[27139]= -979704927;
assign addr[27140]= -945517704;
assign addr[27141]= -911030591;
assign addr[27142]= -876254528;
assign addr[27143]= -841200544;
assign addr[27144]= -805879757;
assign addr[27145]= -770303369;
assign addr[27146]= -734482665;
assign addr[27147]= -698429006;
assign addr[27148]= -662153826;
assign addr[27149]= -625668632;
assign addr[27150]= -588984994;
assign addr[27151]= -552114549;
assign addr[27152]= -515068990;
assign addr[27153]= -477860067;
assign addr[27154]= -440499581;
assign addr[27155]= -402999383;
assign addr[27156]= -365371365;
assign addr[27157]= -327627463;
assign addr[27158]= -289779648;
assign addr[27159]= -251839923;
assign addr[27160]= -213820322;
assign addr[27161]= -175732905;
assign addr[27162]= -137589750;
assign addr[27163]= -99402956;
assign addr[27164]= -61184634;
assign addr[27165]= -22946906;
assign addr[27166]= 15298099;
assign addr[27167]= 53538253;
assign addr[27168]= 91761426;
assign addr[27169]= 129955495;
assign addr[27170]= 168108346;
assign addr[27171]= 206207878;
assign addr[27172]= 244242007;
assign addr[27173]= 282198671;
assign addr[27174]= 320065829;
assign addr[27175]= 357831473;
assign addr[27176]= 395483624;
assign addr[27177]= 433010339;
assign addr[27178]= 470399716;
assign addr[27179]= 507639898;
assign addr[27180]= 544719071;
assign addr[27181]= 581625477;
assign addr[27182]= 618347408;
assign addr[27183]= 654873219;
assign addr[27184]= 691191324;
assign addr[27185]= 727290205;
assign addr[27186]= 763158411;
assign addr[27187]= 798784567;
assign addr[27188]= 834157373;
assign addr[27189]= 869265610;
assign addr[27190]= 904098143;
assign addr[27191]= 938643924;
assign addr[27192]= 972891995;
assign addr[27193]= 1006831495;
assign addr[27194]= 1040451659;
assign addr[27195]= 1073741824;
assign addr[27196]= 1106691431;
assign addr[27197]= 1139290029;
assign addr[27198]= 1171527280;
assign addr[27199]= 1203392958;
assign addr[27200]= 1234876957;
assign addr[27201]= 1265969291;
assign addr[27202]= 1296660098;
assign addr[27203]= 1326939644;
assign addr[27204]= 1356798326;
assign addr[27205]= 1386226674;
assign addr[27206]= 1415215352;
assign addr[27207]= 1443755168;
assign addr[27208]= 1471837070;
assign addr[27209]= 1499452149;
assign addr[27210]= 1526591649;
assign addr[27211]= 1553246960;
assign addr[27212]= 1579409630;
assign addr[27213]= 1605071359;
assign addr[27214]= 1630224009;
assign addr[27215]= 1654859602;
assign addr[27216]= 1678970324;
assign addr[27217]= 1702548529;
assign addr[27218]= 1725586737;
assign addr[27219]= 1748077642;
assign addr[27220]= 1770014111;
assign addr[27221]= 1791389186;
assign addr[27222]= 1812196087;
assign addr[27223]= 1832428215;
assign addr[27224]= 1852079154;
assign addr[27225]= 1871142669;
assign addr[27226]= 1889612716;
assign addr[27227]= 1907483436;
assign addr[27228]= 1924749160;
assign addr[27229]= 1941404413;
assign addr[27230]= 1957443913;
assign addr[27231]= 1972862571;
assign addr[27232]= 1987655498;
assign addr[27233]= 2001818002;
assign addr[27234]= 2015345591;
assign addr[27235]= 2028233973;
assign addr[27236]= 2040479063;
assign addr[27237]= 2052076975;
assign addr[27238]= 2063024031;
assign addr[27239]= 2073316760;
assign addr[27240]= 2082951896;
assign addr[27241]= 2091926384;
assign addr[27242]= 2100237377;
assign addr[27243]= 2107882239;
assign addr[27244]= 2114858546;
assign addr[27245]= 2121164085;
assign addr[27246]= 2126796855;
assign addr[27247]= 2131755071;
assign addr[27248]= 2136037160;
assign addr[27249]= 2139641764;
assign addr[27250]= 2142567738;
assign addr[27251]= 2144814157;
assign addr[27252]= 2146380306;
assign addr[27253]= 2147265689;
assign addr[27254]= 2147470025;
assign addr[27255]= 2146993250;
assign addr[27256]= 2145835515;
assign addr[27257]= 2143997187;
assign addr[27258]= 2141478848;
assign addr[27259]= 2138281298;
assign addr[27260]= 2134405552;
assign addr[27261]= 2129852837;
assign addr[27262]= 2124624598;
assign addr[27263]= 2118722494;
assign addr[27264]= 2112148396;
assign addr[27265]= 2104904390;
assign addr[27266]= 2096992772;
assign addr[27267]= 2088416053;
assign addr[27268]= 2079176953;
assign addr[27269]= 2069278401;
assign addr[27270]= 2058723538;
assign addr[27271]= 2047515711;
assign addr[27272]= 2035658475;
assign addr[27273]= 2023155591;
assign addr[27274]= 2010011024;
assign addr[27275]= 1996228943;
assign addr[27276]= 1981813720;
assign addr[27277]= 1966769926;
assign addr[27278]= 1951102334;
assign addr[27279]= 1934815911;
assign addr[27280]= 1917915825;
assign addr[27281]= 1900407434;
assign addr[27282]= 1882296293;
assign addr[27283]= 1863588145;
assign addr[27284]= 1844288924;
assign addr[27285]= 1824404752;
assign addr[27286]= 1803941934;
assign addr[27287]= 1782906961;
assign addr[27288]= 1761306505;
assign addr[27289]= 1739147417;
assign addr[27290]= 1716436725;
assign addr[27291]= 1693181631;
assign addr[27292]= 1669389513;
assign addr[27293]= 1645067915;
assign addr[27294]= 1620224553;
assign addr[27295]= 1594867305;
assign addr[27296]= 1569004214;
assign addr[27297]= 1542643483;
assign addr[27298]= 1515793473;
assign addr[27299]= 1488462700;
assign addr[27300]= 1460659832;
assign addr[27301]= 1432393688;
assign addr[27302]= 1403673233;
assign addr[27303]= 1374507575;
assign addr[27304]= 1344905966;
assign addr[27305]= 1314877795;
assign addr[27306]= 1284432584;
assign addr[27307]= 1253579991;
assign addr[27308]= 1222329801;
assign addr[27309]= 1190691925;
assign addr[27310]= 1158676398;
assign addr[27311]= 1126293375;
assign addr[27312]= 1093553126;
assign addr[27313]= 1060466036;
assign addr[27314]= 1027042599;
assign addr[27315]= 993293415;
assign addr[27316]= 959229189;
assign addr[27317]= 924860725;
assign addr[27318]= 890198924;
assign addr[27319]= 855254778;
assign addr[27320]= 820039373;
assign addr[27321]= 784563876;
assign addr[27322]= 748839539;
assign addr[27323]= 712877694;
assign addr[27324]= 676689746;
assign addr[27325]= 640287172;
assign addr[27326]= 603681519;
assign addr[27327]= 566884397;
assign addr[27328]= 529907477;
assign addr[27329]= 492762486;
assign addr[27330]= 455461206;
assign addr[27331]= 418015468;
assign addr[27332]= 380437148;
assign addr[27333]= 342738165;
assign addr[27334]= 304930476;
assign addr[27335]= 267026072;
assign addr[27336]= 229036977;
assign addr[27337]= 190975237;
assign addr[27338]= 152852926;
assign addr[27339]= 114682135;
assign addr[27340]= 76474970;
assign addr[27341]= 38243550;
assign addr[27342]= 0;
assign addr[27343]= -38243550;
assign addr[27344]= -76474970;
assign addr[27345]= -114682135;
assign addr[27346]= -152852926;
assign addr[27347]= -190975237;
assign addr[27348]= -229036977;
assign addr[27349]= -267026072;
assign addr[27350]= -304930476;
assign addr[27351]= -342738165;
assign addr[27352]= -380437148;
assign addr[27353]= -418015468;
assign addr[27354]= -455461206;
assign addr[27355]= -492762486;
assign addr[27356]= -529907477;
assign addr[27357]= -566884397;
assign addr[27358]= -603681519;
assign addr[27359]= -640287172;
assign addr[27360]= -676689746;
assign addr[27361]= -712877694;
assign addr[27362]= -748839539;
assign addr[27363]= -784563876;
assign addr[27364]= -820039373;
assign addr[27365]= -855254778;
assign addr[27366]= -890198924;
assign addr[27367]= -924860725;
assign addr[27368]= -959229189;
assign addr[27369]= -993293415;
assign addr[27370]= -1027042599;
assign addr[27371]= -1060466036;
assign addr[27372]= -1093553126;
assign addr[27373]= -1126293375;
assign addr[27374]= -1158676398;
assign addr[27375]= -1190691925;
assign addr[27376]= -1222329801;
assign addr[27377]= -1253579991;
assign addr[27378]= -1284432584;
assign addr[27379]= -1314877795;
assign addr[27380]= -1344905966;
assign addr[27381]= -1374507575;
assign addr[27382]= -1403673233;
assign addr[27383]= -1432393688;
assign addr[27384]= -1460659832;
assign addr[27385]= -1488462700;
assign addr[27386]= -1515793473;
assign addr[27387]= -1542643483;
assign addr[27388]= -1569004214;
assign addr[27389]= -1594867305;
assign addr[27390]= -1620224553;
assign addr[27391]= -1645067915;
assign addr[27392]= -1669389513;
assign addr[27393]= -1693181631;
assign addr[27394]= -1716436725;
assign addr[27395]= -1739147417;
assign addr[27396]= -1761306505;
assign addr[27397]= -1782906961;
assign addr[27398]= -1803941934;
assign addr[27399]= -1824404752;
assign addr[27400]= -1844288924;
assign addr[27401]= -1863588145;
assign addr[27402]= -1882296293;
assign addr[27403]= -1900407434;
assign addr[27404]= -1917915825;
assign addr[27405]= -1934815911;
assign addr[27406]= -1951102334;
assign addr[27407]= -1966769926;
assign addr[27408]= -1981813720;
assign addr[27409]= -1996228943;
assign addr[27410]= -2010011024;
assign addr[27411]= -2023155591;
assign addr[27412]= -2035658475;
assign addr[27413]= -2047515711;
assign addr[27414]= -2058723538;
assign addr[27415]= -2069278401;
assign addr[27416]= -2079176953;
assign addr[27417]= -2088416053;
assign addr[27418]= -2096992772;
assign addr[27419]= -2104904390;
assign addr[27420]= -2112148396;
assign addr[27421]= -2118722494;
assign addr[27422]= -2124624598;
assign addr[27423]= -2129852837;
assign addr[27424]= -2134405552;
assign addr[27425]= -2138281298;
assign addr[27426]= -2141478848;
assign addr[27427]= -2143997187;
assign addr[27428]= -2145835515;
assign addr[27429]= -2146993250;
assign addr[27430]= -2147470025;
assign addr[27431]= -2147265689;
assign addr[27432]= -2146380306;
assign addr[27433]= -2144814157;
assign addr[27434]= -2142567738;
assign addr[27435]= -2139641764;
assign addr[27436]= -2136037160;
assign addr[27437]= -2131755071;
assign addr[27438]= -2126796855;
assign addr[27439]= -2121164085;
assign addr[27440]= -2114858546;
assign addr[27441]= -2107882239;
assign addr[27442]= -2100237377;
assign addr[27443]= -2091926384;
assign addr[27444]= -2082951896;
assign addr[27445]= -2073316760;
assign addr[27446]= -2063024031;
assign addr[27447]= -2052076975;
assign addr[27448]= -2040479063;
assign addr[27449]= -2028233973;
assign addr[27450]= -2015345591;
assign addr[27451]= -2001818002;
assign addr[27452]= -1987655498;
assign addr[27453]= -1972862571;
assign addr[27454]= -1957443913;
assign addr[27455]= -1941404413;
assign addr[27456]= -1924749160;
assign addr[27457]= -1907483436;
assign addr[27458]= -1889612716;
assign addr[27459]= -1871142669;
assign addr[27460]= -1852079154;
assign addr[27461]= -1832428215;
assign addr[27462]= -1812196087;
assign addr[27463]= -1791389186;
assign addr[27464]= -1770014111;
assign addr[27465]= -1748077642;
assign addr[27466]= -1725586737;
assign addr[27467]= -1702548529;
assign addr[27468]= -1678970324;
assign addr[27469]= -1654859602;
assign addr[27470]= -1630224009;
assign addr[27471]= -1605071359;
assign addr[27472]= -1579409630;
assign addr[27473]= -1553246960;
assign addr[27474]= -1526591649;
assign addr[27475]= -1499452149;
assign addr[27476]= -1471837070;
assign addr[27477]= -1443755168;
assign addr[27478]= -1415215352;
assign addr[27479]= -1386226674;
assign addr[27480]= -1356798326;
assign addr[27481]= -1326939644;
assign addr[27482]= -1296660098;
assign addr[27483]= -1265969291;
assign addr[27484]= -1234876957;
assign addr[27485]= -1203392958;
assign addr[27486]= -1171527280;
assign addr[27487]= -1139290029;
assign addr[27488]= -1106691431;
assign addr[27489]= -1073741824;
assign addr[27490]= -1040451659;
assign addr[27491]= -1006831495;
assign addr[27492]= -972891995;
assign addr[27493]= -938643924;
assign addr[27494]= -904098143;
assign addr[27495]= -869265610;
assign addr[27496]= -834157373;
assign addr[27497]= -798784567;
assign addr[27498]= -763158411;
assign addr[27499]= -727290205;
assign addr[27500]= -691191324;
assign addr[27501]= -654873219;
assign addr[27502]= -618347408;
assign addr[27503]= -581625477;
assign addr[27504]= -544719071;
assign addr[27505]= -507639898;
assign addr[27506]= -470399716;
assign addr[27507]= -433010339;
assign addr[27508]= -395483624;
assign addr[27509]= -357831473;
assign addr[27510]= -320065829;
assign addr[27511]= -282198671;
assign addr[27512]= -244242007;
assign addr[27513]= -206207878;
assign addr[27514]= -168108346;
assign addr[27515]= -129955495;
assign addr[27516]= -91761426;
assign addr[27517]= -53538253;
assign addr[27518]= -15298099;
assign addr[27519]= 22946906;
assign addr[27520]= 61184634;
assign addr[27521]= 99402956;
assign addr[27522]= 137589750;
assign addr[27523]= 175732905;
assign addr[27524]= 213820322;
assign addr[27525]= 251839923;
assign addr[27526]= 289779648;
assign addr[27527]= 327627463;
assign addr[27528]= 365371365;
assign addr[27529]= 402999383;
assign addr[27530]= 440499581;
assign addr[27531]= 477860067;
assign addr[27532]= 515068990;
assign addr[27533]= 552114549;
assign addr[27534]= 588984994;
assign addr[27535]= 625668632;
assign addr[27536]= 662153826;
assign addr[27537]= 698429006;
assign addr[27538]= 734482665;
assign addr[27539]= 770303369;
assign addr[27540]= 805879757;
assign addr[27541]= 841200544;
assign addr[27542]= 876254528;
assign addr[27543]= 911030591;
assign addr[27544]= 945517704;
assign addr[27545]= 979704927;
assign addr[27546]= 1013581418;
assign addr[27547]= 1047136432;
assign addr[27548]= 1080359326;
assign addr[27549]= 1113239564;
assign addr[27550]= 1145766716;
assign addr[27551]= 1177930466;
assign addr[27552]= 1209720613;
assign addr[27553]= 1241127074;
assign addr[27554]= 1272139887;
assign addr[27555]= 1302749217;
assign addr[27556]= 1332945355;
assign addr[27557]= 1362718723;
assign addr[27558]= 1392059879;
assign addr[27559]= 1420959516;
assign addr[27560]= 1449408469;
assign addr[27561]= 1477397714;
assign addr[27562]= 1504918373;
assign addr[27563]= 1531961719;
assign addr[27564]= 1558519173;
assign addr[27565]= 1584582314;
assign addr[27566]= 1610142873;
assign addr[27567]= 1635192744;
assign addr[27568]= 1659723983;
assign addr[27569]= 1683728808;
assign addr[27570]= 1707199606;
assign addr[27571]= 1730128933;
assign addr[27572]= 1752509516;
assign addr[27573]= 1774334257;
assign addr[27574]= 1795596234;
assign addr[27575]= 1816288703;
assign addr[27576]= 1836405100;
assign addr[27577]= 1855939047;
assign addr[27578]= 1874884346;
assign addr[27579]= 1893234990;
assign addr[27580]= 1910985158;
assign addr[27581]= 1928129220;
assign addr[27582]= 1944661739;
assign addr[27583]= 1960577471;
assign addr[27584]= 1975871368;
assign addr[27585]= 1990538579;
assign addr[27586]= 2004574453;
assign addr[27587]= 2017974537;
assign addr[27588]= 2030734582;
assign addr[27589]= 2042850540;
assign addr[27590]= 2054318569;
assign addr[27591]= 2065135031;
assign addr[27592]= 2075296495;
assign addr[27593]= 2084799740;
assign addr[27594]= 2093641749;
assign addr[27595]= 2101819720;
assign addr[27596]= 2109331059;
assign addr[27597]= 2116173382;
assign addr[27598]= 2122344521;
assign addr[27599]= 2127842516;
assign addr[27600]= 2132665626;
assign addr[27601]= 2136812319;
assign addr[27602]= 2140281282;
assign addr[27603]= 2143071413;
assign addr[27604]= 2145181827;
assign addr[27605]= 2146611856;
assign addr[27606]= 2147361045;
assign addr[27607]= 2147429158;
assign addr[27608]= 2146816171;
assign addr[27609]= 2145522281;
assign addr[27610]= 2143547897;
assign addr[27611]= 2140893646;
assign addr[27612]= 2137560369;
assign addr[27613]= 2133549123;
assign addr[27614]= 2128861181;
assign addr[27615]= 2123498030;
assign addr[27616]= 2117461370;
assign addr[27617]= 2110753117;
assign addr[27618]= 2103375398;
assign addr[27619]= 2095330553;
assign addr[27620]= 2086621133;
assign addr[27621]= 2077249901;
assign addr[27622]= 2067219829;
assign addr[27623]= 2056534099;
assign addr[27624]= 2045196100;
assign addr[27625]= 2033209426;
assign addr[27626]= 2020577882;
assign addr[27627]= 2007305472;
assign addr[27628]= 1993396407;
assign addr[27629]= 1978855097;
assign addr[27630]= 1963686155;
assign addr[27631]= 1947894393;
assign addr[27632]= 1931484818;
assign addr[27633]= 1914462636;
assign addr[27634]= 1896833245;
assign addr[27635]= 1878602237;
assign addr[27636]= 1859775393;
assign addr[27637]= 1840358687;
assign addr[27638]= 1820358275;
assign addr[27639]= 1799780501;
assign addr[27640]= 1778631892;
assign addr[27641]= 1756919156;
assign addr[27642]= 1734649179;
assign addr[27643]= 1711829025;
assign addr[27644]= 1688465931;
assign addr[27645]= 1664567307;
assign addr[27646]= 1640140734;
assign addr[27647]= 1615193959;
assign addr[27648]= 1589734894;
assign addr[27649]= 1563771613;
assign addr[27650]= 1537312353;
assign addr[27651]= 1510365504;
assign addr[27652]= 1482939614;
assign addr[27653]= 1455043381;
assign addr[27654]= 1426685652;
assign addr[27655]= 1397875423;
assign addr[27656]= 1368621831;
assign addr[27657]= 1338934154;
assign addr[27658]= 1308821808;
assign addr[27659]= 1278294345;
assign addr[27660]= 1247361445;
assign addr[27661]= 1216032921;
assign addr[27662]= 1184318708;
assign addr[27663]= 1152228866;
assign addr[27664]= 1119773573;
assign addr[27665]= 1086963121;
assign addr[27666]= 1053807919;
assign addr[27667]= 1020318481;
assign addr[27668]= 986505429;
assign addr[27669]= 952379488;
assign addr[27670]= 917951481;
assign addr[27671]= 883232329;
assign addr[27672]= 848233042;
assign addr[27673]= 812964722;
assign addr[27674]= 777438554;
assign addr[27675]= 741665807;
assign addr[27676]= 705657826;
assign addr[27677]= 669426032;
assign addr[27678]= 632981917;
assign addr[27679]= 596337040;
assign addr[27680]= 559503022;
assign addr[27681]= 522491548;
assign addr[27682]= 485314355;
assign addr[27683]= 447983235;
assign addr[27684]= 410510029;
assign addr[27685]= 372906622;
assign addr[27686]= 335184940;
assign addr[27687]= 297356948;
assign addr[27688]= 259434643;
assign addr[27689]= 221430054;
assign addr[27690]= 183355234;
assign addr[27691]= 145222259;
assign addr[27692]= 107043224;
assign addr[27693]= 68830239;
assign addr[27694]= 30595422;
assign addr[27695]= -7649098;
assign addr[27696]= -45891193;
assign addr[27697]= -84118732;
assign addr[27698]= -122319591;
assign addr[27699]= -160481654;
assign addr[27700]= -198592817;
assign addr[27701]= -236640993;
assign addr[27702]= -274614114;
assign addr[27703]= -312500135;
assign addr[27704]= -350287041;
assign addr[27705]= -387962847;
assign addr[27706]= -425515602;
assign addr[27707]= -462933398;
assign addr[27708]= -500204365;
assign addr[27709]= -537316682;
assign addr[27710]= -574258580;
assign addr[27711]= -611018340;
assign addr[27712]= -647584304;
assign addr[27713]= -683944874;
assign addr[27714]= -720088517;
assign addr[27715]= -756003771;
assign addr[27716]= -791679244;
assign addr[27717]= -827103620;
assign addr[27718]= -862265664;
assign addr[27719]= -897154224;
assign addr[27720]= -931758235;
assign addr[27721]= -966066720;
assign addr[27722]= -1000068799;
assign addr[27723]= -1033753687;
assign addr[27724]= -1067110699;
assign addr[27725]= -1100129257;
assign addr[27726]= -1132798888;
assign addr[27727]= -1165109230;
assign addr[27728]= -1197050035;
assign addr[27729]= -1228611172;
assign addr[27730]= -1259782632;
assign addr[27731]= -1290554528;
assign addr[27732]= -1320917099;
assign addr[27733]= -1350860716;
assign addr[27734]= -1380375881;
assign addr[27735]= -1409453233;
assign addr[27736]= -1438083551;
assign addr[27737]= -1466257752;
assign addr[27738]= -1493966902;
assign addr[27739]= -1521202211;
assign addr[27740]= -1547955041;
assign addr[27741]= -1574216908;
assign addr[27742]= -1599979481;
assign addr[27743]= -1625234591;
assign addr[27744]= -1649974225;
assign addr[27745]= -1674190539;
assign addr[27746]= -1697875851;
assign addr[27747]= -1721022648;
assign addr[27748]= -1743623590;
assign addr[27749]= -1765671509;
assign addr[27750]= -1787159411;
assign addr[27751]= -1808080480;
assign addr[27752]= -1828428082;
assign addr[27753]= -1848195763;
assign addr[27754]= -1867377253;
assign addr[27755]= -1885966468;
assign addr[27756]= -1903957513;
assign addr[27757]= -1921344681;
assign addr[27758]= -1938122457;
assign addr[27759]= -1954285520;
assign addr[27760]= -1969828744;
assign addr[27761]= -1984747199;
assign addr[27762]= -1999036154;
assign addr[27763]= -2012691075;
assign addr[27764]= -2025707632;
assign addr[27765]= -2038081698;
assign addr[27766]= -2049809346;
assign addr[27767]= -2060886858;
assign addr[27768]= -2071310720;
assign addr[27769]= -2081077626;
assign addr[27770]= -2090184478;
assign addr[27771]= -2098628387;
assign addr[27772]= -2106406677;
assign addr[27773]= -2113516878;
assign addr[27774]= -2119956737;
assign addr[27775]= -2125724211;
assign addr[27776]= -2130817471;
assign addr[27777]= -2135234901;
assign addr[27778]= -2138975100;
assign addr[27779]= -2142036881;
assign addr[27780]= -2144419275;
assign addr[27781]= -2146121524;
assign addr[27782]= -2147143090;
assign addr[27783]= -2147483648;
assign addr[27784]= -2147143090;
assign addr[27785]= -2146121524;
assign addr[27786]= -2144419275;
assign addr[27787]= -2142036881;
assign addr[27788]= -2138975100;
assign addr[27789]= -2135234901;
assign addr[27790]= -2130817471;
assign addr[27791]= -2125724211;
assign addr[27792]= -2119956737;
assign addr[27793]= -2113516878;
assign addr[27794]= -2106406677;
assign addr[27795]= -2098628387;
assign addr[27796]= -2090184478;
assign addr[27797]= -2081077626;
assign addr[27798]= -2071310720;
assign addr[27799]= -2060886858;
assign addr[27800]= -2049809346;
assign addr[27801]= -2038081698;
assign addr[27802]= -2025707632;
assign addr[27803]= -2012691075;
assign addr[27804]= -1999036154;
assign addr[27805]= -1984747199;
assign addr[27806]= -1969828744;
assign addr[27807]= -1954285520;
assign addr[27808]= -1938122457;
assign addr[27809]= -1921344681;
assign addr[27810]= -1903957513;
assign addr[27811]= -1885966468;
assign addr[27812]= -1867377253;
assign addr[27813]= -1848195763;
assign addr[27814]= -1828428082;
assign addr[27815]= -1808080480;
assign addr[27816]= -1787159411;
assign addr[27817]= -1765671509;
assign addr[27818]= -1743623590;
assign addr[27819]= -1721022648;
assign addr[27820]= -1697875851;
assign addr[27821]= -1674190539;
assign addr[27822]= -1649974225;
assign addr[27823]= -1625234591;
assign addr[27824]= -1599979481;
assign addr[27825]= -1574216908;
assign addr[27826]= -1547955041;
assign addr[27827]= -1521202211;
assign addr[27828]= -1493966902;
assign addr[27829]= -1466257752;
assign addr[27830]= -1438083551;
assign addr[27831]= -1409453233;
assign addr[27832]= -1380375881;
assign addr[27833]= -1350860716;
assign addr[27834]= -1320917099;
assign addr[27835]= -1290554528;
assign addr[27836]= -1259782632;
assign addr[27837]= -1228611172;
assign addr[27838]= -1197050035;
assign addr[27839]= -1165109230;
assign addr[27840]= -1132798888;
assign addr[27841]= -1100129257;
assign addr[27842]= -1067110699;
assign addr[27843]= -1033753687;
assign addr[27844]= -1000068799;
assign addr[27845]= -966066720;
assign addr[27846]= -931758235;
assign addr[27847]= -897154224;
assign addr[27848]= -862265664;
assign addr[27849]= -827103620;
assign addr[27850]= -791679244;
assign addr[27851]= -756003771;
assign addr[27852]= -720088517;
assign addr[27853]= -683944874;
assign addr[27854]= -647584304;
assign addr[27855]= -611018340;
assign addr[27856]= -574258580;
assign addr[27857]= -537316682;
assign addr[27858]= -500204365;
assign addr[27859]= -462933398;
assign addr[27860]= -425515602;
assign addr[27861]= -387962847;
assign addr[27862]= -350287041;
assign addr[27863]= -312500135;
assign addr[27864]= -274614114;
assign addr[27865]= -236640993;
assign addr[27866]= -198592817;
assign addr[27867]= -160481654;
assign addr[27868]= -122319591;
assign addr[27869]= -84118732;
assign addr[27870]= -45891193;
assign addr[27871]= -7649098;
assign addr[27872]= 30595422;
assign addr[27873]= 68830239;
assign addr[27874]= 107043224;
assign addr[27875]= 145222259;
assign addr[27876]= 183355234;
assign addr[27877]= 221430054;
assign addr[27878]= 259434643;
assign addr[27879]= 297356948;
assign addr[27880]= 335184940;
assign addr[27881]= 372906622;
assign addr[27882]= 410510029;
assign addr[27883]= 447983235;
assign addr[27884]= 485314355;
assign addr[27885]= 522491548;
assign addr[27886]= 559503022;
assign addr[27887]= 596337040;
assign addr[27888]= 632981917;
assign addr[27889]= 669426032;
assign addr[27890]= 705657826;
assign addr[27891]= 741665807;
assign addr[27892]= 777438554;
assign addr[27893]= 812964722;
assign addr[27894]= 848233042;
assign addr[27895]= 883232329;
assign addr[27896]= 917951481;
assign addr[27897]= 952379488;
assign addr[27898]= 986505429;
assign addr[27899]= 1020318481;
assign addr[27900]= 1053807919;
assign addr[27901]= 1086963121;
assign addr[27902]= 1119773573;
assign addr[27903]= 1152228866;
assign addr[27904]= 1184318708;
assign addr[27905]= 1216032921;
assign addr[27906]= 1247361445;
assign addr[27907]= 1278294345;
assign addr[27908]= 1308821808;
assign addr[27909]= 1338934154;
assign addr[27910]= 1368621831;
assign addr[27911]= 1397875423;
assign addr[27912]= 1426685652;
assign addr[27913]= 1455043381;
assign addr[27914]= 1482939614;
assign addr[27915]= 1510365504;
assign addr[27916]= 1537312353;
assign addr[27917]= 1563771613;
assign addr[27918]= 1589734894;
assign addr[27919]= 1615193959;
assign addr[27920]= 1640140734;
assign addr[27921]= 1664567307;
assign addr[27922]= 1688465931;
assign addr[27923]= 1711829025;
assign addr[27924]= 1734649179;
assign addr[27925]= 1756919156;
assign addr[27926]= 1778631892;
assign addr[27927]= 1799780501;
assign addr[27928]= 1820358275;
assign addr[27929]= 1840358687;
assign addr[27930]= 1859775393;
assign addr[27931]= 1878602237;
assign addr[27932]= 1896833245;
assign addr[27933]= 1914462636;
assign addr[27934]= 1931484818;
assign addr[27935]= 1947894393;
assign addr[27936]= 1963686155;
assign addr[27937]= 1978855097;
assign addr[27938]= 1993396407;
assign addr[27939]= 2007305472;
assign addr[27940]= 2020577882;
assign addr[27941]= 2033209426;
assign addr[27942]= 2045196100;
assign addr[27943]= 2056534099;
assign addr[27944]= 2067219829;
assign addr[27945]= 2077249901;
assign addr[27946]= 2086621133;
assign addr[27947]= 2095330553;
assign addr[27948]= 2103375398;
assign addr[27949]= 2110753117;
assign addr[27950]= 2117461370;
assign addr[27951]= 2123498030;
assign addr[27952]= 2128861181;
assign addr[27953]= 2133549123;
assign addr[27954]= 2137560369;
assign addr[27955]= 2140893646;
assign addr[27956]= 2143547897;
assign addr[27957]= 2145522281;
assign addr[27958]= 2146816171;
assign addr[27959]= 2147429158;
assign addr[27960]= 2147361045;
assign addr[27961]= 2146611856;
assign addr[27962]= 2145181827;
assign addr[27963]= 2143071413;
assign addr[27964]= 2140281282;
assign addr[27965]= 2136812319;
assign addr[27966]= 2132665626;
assign addr[27967]= 2127842516;
assign addr[27968]= 2122344521;
assign addr[27969]= 2116173382;
assign addr[27970]= 2109331059;
assign addr[27971]= 2101819720;
assign addr[27972]= 2093641749;
assign addr[27973]= 2084799740;
assign addr[27974]= 2075296495;
assign addr[27975]= 2065135031;
assign addr[27976]= 2054318569;
assign addr[27977]= 2042850540;
assign addr[27978]= 2030734582;
assign addr[27979]= 2017974537;
assign addr[27980]= 2004574453;
assign addr[27981]= 1990538579;
assign addr[27982]= 1975871368;
assign addr[27983]= 1960577471;
assign addr[27984]= 1944661739;
assign addr[27985]= 1928129220;
assign addr[27986]= 1910985158;
assign addr[27987]= 1893234990;
assign addr[27988]= 1874884346;
assign addr[27989]= 1855939047;
assign addr[27990]= 1836405100;
assign addr[27991]= 1816288703;
assign addr[27992]= 1795596234;
assign addr[27993]= 1774334257;
assign addr[27994]= 1752509516;
assign addr[27995]= 1730128933;
assign addr[27996]= 1707199606;
assign addr[27997]= 1683728808;
assign addr[27998]= 1659723983;
assign addr[27999]= 1635192744;
assign addr[28000]= 1610142873;
assign addr[28001]= 1584582314;
assign addr[28002]= 1558519173;
assign addr[28003]= 1531961719;
assign addr[28004]= 1504918373;
assign addr[28005]= 1477397714;
assign addr[28006]= 1449408469;
assign addr[28007]= 1420959516;
assign addr[28008]= 1392059879;
assign addr[28009]= 1362718723;
assign addr[28010]= 1332945355;
assign addr[28011]= 1302749217;
assign addr[28012]= 1272139887;
assign addr[28013]= 1241127074;
assign addr[28014]= 1209720613;
assign addr[28015]= 1177930466;
assign addr[28016]= 1145766716;
assign addr[28017]= 1113239564;
assign addr[28018]= 1080359326;
assign addr[28019]= 1047136432;
assign addr[28020]= 1013581418;
assign addr[28021]= 979704927;
assign addr[28022]= 945517704;
assign addr[28023]= 911030591;
assign addr[28024]= 876254528;
assign addr[28025]= 841200544;
assign addr[28026]= 805879757;
assign addr[28027]= 770303369;
assign addr[28028]= 734482665;
assign addr[28029]= 698429006;
assign addr[28030]= 662153826;
assign addr[28031]= 625668632;
assign addr[28032]= 588984994;
assign addr[28033]= 552114549;
assign addr[28034]= 515068990;
assign addr[28035]= 477860067;
assign addr[28036]= 440499581;
assign addr[28037]= 402999383;
assign addr[28038]= 365371365;
assign addr[28039]= 327627463;
assign addr[28040]= 289779648;
assign addr[28041]= 251839923;
assign addr[28042]= 213820322;
assign addr[28043]= 175732905;
assign addr[28044]= 137589750;
assign addr[28045]= 99402956;
assign addr[28046]= 61184634;
assign addr[28047]= 22946906;
assign addr[28048]= -15298099;
assign addr[28049]= -53538253;
assign addr[28050]= -91761426;
assign addr[28051]= -129955495;
assign addr[28052]= -168108346;
assign addr[28053]= -206207878;
assign addr[28054]= -244242007;
assign addr[28055]= -282198671;
assign addr[28056]= -320065829;
assign addr[28057]= -357831473;
assign addr[28058]= -395483624;
assign addr[28059]= -433010339;
assign addr[28060]= -470399716;
assign addr[28061]= -507639898;
assign addr[28062]= -544719071;
assign addr[28063]= -581625477;
assign addr[28064]= -618347408;
assign addr[28065]= -654873219;
assign addr[28066]= -691191324;
assign addr[28067]= -727290205;
assign addr[28068]= -763158411;
assign addr[28069]= -798784567;
assign addr[28070]= -834157373;
assign addr[28071]= -869265610;
assign addr[28072]= -904098143;
assign addr[28073]= -938643924;
assign addr[28074]= -972891995;
assign addr[28075]= -1006831495;
assign addr[28076]= -1040451659;
assign addr[28077]= -1073741824;
assign addr[28078]= -1106691431;
assign addr[28079]= -1139290029;
assign addr[28080]= -1171527280;
assign addr[28081]= -1203392958;
assign addr[28082]= -1234876957;
assign addr[28083]= -1265969291;
assign addr[28084]= -1296660098;
assign addr[28085]= -1326939644;
assign addr[28086]= -1356798326;
assign addr[28087]= -1386226674;
assign addr[28088]= -1415215352;
assign addr[28089]= -1443755168;
assign addr[28090]= -1471837070;
assign addr[28091]= -1499452149;
assign addr[28092]= -1526591649;
assign addr[28093]= -1553246960;
assign addr[28094]= -1579409630;
assign addr[28095]= -1605071359;
assign addr[28096]= -1630224009;
assign addr[28097]= -1654859602;
assign addr[28098]= -1678970324;
assign addr[28099]= -1702548529;
assign addr[28100]= -1725586737;
assign addr[28101]= -1748077642;
assign addr[28102]= -1770014111;
assign addr[28103]= -1791389186;
assign addr[28104]= -1812196087;
assign addr[28105]= -1832428215;
assign addr[28106]= -1852079154;
assign addr[28107]= -1871142669;
assign addr[28108]= -1889612716;
assign addr[28109]= -1907483436;
assign addr[28110]= -1924749160;
assign addr[28111]= -1941404413;
assign addr[28112]= -1957443913;
assign addr[28113]= -1972862571;
assign addr[28114]= -1987655498;
assign addr[28115]= -2001818002;
assign addr[28116]= -2015345591;
assign addr[28117]= -2028233973;
assign addr[28118]= -2040479063;
assign addr[28119]= -2052076975;
assign addr[28120]= -2063024031;
assign addr[28121]= -2073316760;
assign addr[28122]= -2082951896;
assign addr[28123]= -2091926384;
assign addr[28124]= -2100237377;
assign addr[28125]= -2107882239;
assign addr[28126]= -2114858546;
assign addr[28127]= -2121164085;
assign addr[28128]= -2126796855;
assign addr[28129]= -2131755071;
assign addr[28130]= -2136037160;
assign addr[28131]= -2139641764;
assign addr[28132]= -2142567738;
assign addr[28133]= -2144814157;
assign addr[28134]= -2146380306;
assign addr[28135]= -2147265689;
assign addr[28136]= -2147470025;
assign addr[28137]= -2146993250;
assign addr[28138]= -2145835515;
assign addr[28139]= -2143997187;
assign addr[28140]= -2141478848;
assign addr[28141]= -2138281298;
assign addr[28142]= -2134405552;
assign addr[28143]= -2129852837;
assign addr[28144]= -2124624598;
assign addr[28145]= -2118722494;
assign addr[28146]= -2112148396;
assign addr[28147]= -2104904390;
assign addr[28148]= -2096992772;
assign addr[28149]= -2088416053;
assign addr[28150]= -2079176953;
assign addr[28151]= -2069278401;
assign addr[28152]= -2058723538;
assign addr[28153]= -2047515711;
assign addr[28154]= -2035658475;
assign addr[28155]= -2023155591;
assign addr[28156]= -2010011024;
assign addr[28157]= -1996228943;
assign addr[28158]= -1981813720;
assign addr[28159]= -1966769926;
assign addr[28160]= -1951102334;
assign addr[28161]= -1934815911;
assign addr[28162]= -1917915825;
assign addr[28163]= -1900407434;
assign addr[28164]= -1882296293;
assign addr[28165]= -1863588145;
assign addr[28166]= -1844288924;
assign addr[28167]= -1824404752;
assign addr[28168]= -1803941934;
assign addr[28169]= -1782906961;
assign addr[28170]= -1761306505;
assign addr[28171]= -1739147417;
assign addr[28172]= -1716436725;
assign addr[28173]= -1693181631;
assign addr[28174]= -1669389513;
assign addr[28175]= -1645067915;
assign addr[28176]= -1620224553;
assign addr[28177]= -1594867305;
assign addr[28178]= -1569004214;
assign addr[28179]= -1542643483;
assign addr[28180]= -1515793473;
assign addr[28181]= -1488462700;
assign addr[28182]= -1460659832;
assign addr[28183]= -1432393688;
assign addr[28184]= -1403673233;
assign addr[28185]= -1374507575;
assign addr[28186]= -1344905966;
assign addr[28187]= -1314877795;
assign addr[28188]= -1284432584;
assign addr[28189]= -1253579991;
assign addr[28190]= -1222329801;
assign addr[28191]= -1190691925;
assign addr[28192]= -1158676398;
assign addr[28193]= -1126293375;
assign addr[28194]= -1093553126;
assign addr[28195]= -1060466036;
assign addr[28196]= -1027042599;
assign addr[28197]= -993293415;
assign addr[28198]= -959229189;
assign addr[28199]= -924860725;
assign addr[28200]= -890198924;
assign addr[28201]= -855254778;
assign addr[28202]= -820039373;
assign addr[28203]= -784563876;
assign addr[28204]= -748839539;
assign addr[28205]= -712877694;
assign addr[28206]= -676689746;
assign addr[28207]= -640287172;
assign addr[28208]= -603681519;
assign addr[28209]= -566884397;
assign addr[28210]= -529907477;
assign addr[28211]= -492762486;
assign addr[28212]= -455461206;
assign addr[28213]= -418015468;
assign addr[28214]= -380437148;
assign addr[28215]= -342738165;
assign addr[28216]= -304930476;
assign addr[28217]= -267026072;
assign addr[28218]= -229036977;
assign addr[28219]= -190975237;
assign addr[28220]= -152852926;
assign addr[28221]= -114682135;
assign addr[28222]= -76474970;
assign addr[28223]= -38243550;
assign addr[28224]= 0;
assign addr[28225]= 38243550;
assign addr[28226]= 76474970;
assign addr[28227]= 114682135;
assign addr[28228]= 152852926;
assign addr[28229]= 190975237;
assign addr[28230]= 229036977;
assign addr[28231]= 267026072;
assign addr[28232]= 304930476;
assign addr[28233]= 342738165;
assign addr[28234]= 380437148;
assign addr[28235]= 418015468;
assign addr[28236]= 455461206;
assign addr[28237]= 492762486;
assign addr[28238]= 529907477;
assign addr[28239]= 566884397;
assign addr[28240]= 603681519;
assign addr[28241]= 640287172;
assign addr[28242]= 676689746;
assign addr[28243]= 712877694;
assign addr[28244]= 748839539;
assign addr[28245]= 784563876;
assign addr[28246]= 820039373;
assign addr[28247]= 855254778;
assign addr[28248]= 890198924;
assign addr[28249]= 924860725;
assign addr[28250]= 959229189;
assign addr[28251]= 993293415;
assign addr[28252]= 1027042599;
assign addr[28253]= 1060466036;
assign addr[28254]= 1093553126;
assign addr[28255]= 1126293375;
assign addr[28256]= 1158676398;
assign addr[28257]= 1190691925;
assign addr[28258]= 1222329801;
assign addr[28259]= 1253579991;
assign addr[28260]= 1284432584;
assign addr[28261]= 1314877795;
assign addr[28262]= 1344905966;
assign addr[28263]= 1374507575;
assign addr[28264]= 1403673233;
assign addr[28265]= 1432393688;
assign addr[28266]= 1460659832;
assign addr[28267]= 1488462700;
assign addr[28268]= 1515793473;
assign addr[28269]= 1542643483;
assign addr[28270]= 1569004214;
assign addr[28271]= 1594867305;
assign addr[28272]= 1620224553;
assign addr[28273]= 1645067915;
assign addr[28274]= 1669389513;
assign addr[28275]= 1693181631;
assign addr[28276]= 1716436725;
assign addr[28277]= 1739147417;
assign addr[28278]= 1761306505;
assign addr[28279]= 1782906961;
assign addr[28280]= 1803941934;
assign addr[28281]= 1824404752;
assign addr[28282]= 1844288924;
assign addr[28283]= 1863588145;
assign addr[28284]= 1882296293;
assign addr[28285]= 1900407434;
assign addr[28286]= 1917915825;
assign addr[28287]= 1934815911;
assign addr[28288]= 1951102334;
assign addr[28289]= 1966769926;
assign addr[28290]= 1981813720;
assign addr[28291]= 1996228943;
assign addr[28292]= 2010011024;
assign addr[28293]= 2023155591;
assign addr[28294]= 2035658475;
assign addr[28295]= 2047515711;
assign addr[28296]= 2058723538;
assign addr[28297]= 2069278401;
assign addr[28298]= 2079176953;
assign addr[28299]= 2088416053;
assign addr[28300]= 2096992772;
assign addr[28301]= 2104904390;
assign addr[28302]= 2112148396;
assign addr[28303]= 2118722494;
assign addr[28304]= 2124624598;
assign addr[28305]= 2129852837;
assign addr[28306]= 2134405552;
assign addr[28307]= 2138281298;
assign addr[28308]= 2141478848;
assign addr[28309]= 2143997187;
assign addr[28310]= 2145835515;
assign addr[28311]= 2146993250;
assign addr[28312]= 2147470025;
assign addr[28313]= 2147265689;
assign addr[28314]= 2146380306;
assign addr[28315]= 2144814157;
assign addr[28316]= 2142567738;
assign addr[28317]= 2139641764;
assign addr[28318]= 2136037160;
assign addr[28319]= 2131755071;
assign addr[28320]= 2126796855;
assign addr[28321]= 2121164085;
assign addr[28322]= 2114858546;
assign addr[28323]= 2107882239;
assign addr[28324]= 2100237377;
assign addr[28325]= 2091926384;
assign addr[28326]= 2082951896;
assign addr[28327]= 2073316760;
assign addr[28328]= 2063024031;
assign addr[28329]= 2052076975;
assign addr[28330]= 2040479063;
assign addr[28331]= 2028233973;
assign addr[28332]= 2015345591;
assign addr[28333]= 2001818002;
assign addr[28334]= 1987655498;
assign addr[28335]= 1972862571;
assign addr[28336]= 1957443913;
assign addr[28337]= 1941404413;
assign addr[28338]= 1924749160;
assign addr[28339]= 1907483436;
assign addr[28340]= 1889612716;
assign addr[28341]= 1871142669;
assign addr[28342]= 1852079154;
assign addr[28343]= 1832428215;
assign addr[28344]= 1812196087;
assign addr[28345]= 1791389186;
assign addr[28346]= 1770014111;
assign addr[28347]= 1748077642;
assign addr[28348]= 1725586737;
assign addr[28349]= 1702548529;
assign addr[28350]= 1678970324;
assign addr[28351]= 1654859602;
assign addr[28352]= 1630224009;
assign addr[28353]= 1605071359;
assign addr[28354]= 1579409630;
assign addr[28355]= 1553246960;
assign addr[28356]= 1526591649;
assign addr[28357]= 1499452149;
assign addr[28358]= 1471837070;
assign addr[28359]= 1443755168;
assign addr[28360]= 1415215352;
assign addr[28361]= 1386226674;
assign addr[28362]= 1356798326;
assign addr[28363]= 1326939644;
assign addr[28364]= 1296660098;
assign addr[28365]= 1265969291;
assign addr[28366]= 1234876957;
assign addr[28367]= 1203392958;
assign addr[28368]= 1171527280;
assign addr[28369]= 1139290029;
assign addr[28370]= 1106691431;
assign addr[28371]= 1073741824;
assign addr[28372]= 1040451659;
assign addr[28373]= 1006831495;
assign addr[28374]= 972891995;
assign addr[28375]= 938643924;
assign addr[28376]= 904098143;
assign addr[28377]= 869265610;
assign addr[28378]= 834157373;
assign addr[28379]= 798784567;
assign addr[28380]= 763158411;
assign addr[28381]= 727290205;
assign addr[28382]= 691191324;
assign addr[28383]= 654873219;
assign addr[28384]= 618347408;
assign addr[28385]= 581625477;
assign addr[28386]= 544719071;
assign addr[28387]= 507639898;
assign addr[28388]= 470399716;
assign addr[28389]= 433010339;
assign addr[28390]= 395483624;
assign addr[28391]= 357831473;
assign addr[28392]= 320065829;
assign addr[28393]= 282198671;
assign addr[28394]= 244242007;
assign addr[28395]= 206207878;
assign addr[28396]= 168108346;
assign addr[28397]= 129955495;
assign addr[28398]= 91761426;
assign addr[28399]= 53538253;
assign addr[28400]= 15298099;
assign addr[28401]= -22946906;
assign addr[28402]= -61184634;
assign addr[28403]= -99402956;
assign addr[28404]= -137589750;
assign addr[28405]= -175732905;
assign addr[28406]= -213820322;
assign addr[28407]= -251839923;
assign addr[28408]= -289779648;
assign addr[28409]= -327627463;
assign addr[28410]= -365371365;
assign addr[28411]= -402999383;
assign addr[28412]= -440499581;
assign addr[28413]= -477860067;
assign addr[28414]= -515068990;
assign addr[28415]= -552114549;
assign addr[28416]= -588984994;
assign addr[28417]= -625668632;
assign addr[28418]= -662153826;
assign addr[28419]= -698429006;
assign addr[28420]= -734482665;
assign addr[28421]= -770303369;
assign addr[28422]= -805879757;
assign addr[28423]= -841200544;
assign addr[28424]= -876254528;
assign addr[28425]= -911030591;
assign addr[28426]= -945517704;
assign addr[28427]= -979704927;
assign addr[28428]= -1013581418;
assign addr[28429]= -1047136432;
assign addr[28430]= -1080359326;
assign addr[28431]= -1113239564;
assign addr[28432]= -1145766716;
assign addr[28433]= -1177930466;
assign addr[28434]= -1209720613;
assign addr[28435]= -1241127074;
assign addr[28436]= -1272139887;
assign addr[28437]= -1302749217;
assign addr[28438]= -1332945355;
assign addr[28439]= -1362718723;
assign addr[28440]= -1392059879;
assign addr[28441]= -1420959516;
assign addr[28442]= -1449408469;
assign addr[28443]= -1477397714;
assign addr[28444]= -1504918373;
assign addr[28445]= -1531961719;
assign addr[28446]= -1558519173;
assign addr[28447]= -1584582314;
assign addr[28448]= -1610142873;
assign addr[28449]= -1635192744;
assign addr[28450]= -1659723983;
assign addr[28451]= -1683728808;
assign addr[28452]= -1707199606;
assign addr[28453]= -1730128933;
assign addr[28454]= -1752509516;
assign addr[28455]= -1774334257;
assign addr[28456]= -1795596234;
assign addr[28457]= -1816288703;
assign addr[28458]= -1836405100;
assign addr[28459]= -1855939047;
assign addr[28460]= -1874884346;
assign addr[28461]= -1893234990;
assign addr[28462]= -1910985158;
assign addr[28463]= -1928129220;
assign addr[28464]= -1944661739;
assign addr[28465]= -1960577471;
assign addr[28466]= -1975871368;
assign addr[28467]= -1990538579;
assign addr[28468]= -2004574453;
assign addr[28469]= -2017974537;
assign addr[28470]= -2030734582;
assign addr[28471]= -2042850540;
assign addr[28472]= -2054318569;
assign addr[28473]= -2065135031;
assign addr[28474]= -2075296495;
assign addr[28475]= -2084799740;
assign addr[28476]= -2093641749;
assign addr[28477]= -2101819720;
assign addr[28478]= -2109331059;
assign addr[28479]= -2116173382;
assign addr[28480]= -2122344521;
assign addr[28481]= -2127842516;
assign addr[28482]= -2132665626;
assign addr[28483]= -2136812319;
assign addr[28484]= -2140281282;
assign addr[28485]= -2143071413;
assign addr[28486]= -2145181827;
assign addr[28487]= -2146611856;
assign addr[28488]= -2147361045;
assign addr[28489]= -2147429158;
assign addr[28490]= -2146816171;
assign addr[28491]= -2145522281;
assign addr[28492]= -2143547897;
assign addr[28493]= -2140893646;
assign addr[28494]= -2137560369;
assign addr[28495]= -2133549123;
assign addr[28496]= -2128861181;
assign addr[28497]= -2123498030;
assign addr[28498]= -2117461370;
assign addr[28499]= -2110753117;
assign addr[28500]= -2103375398;
assign addr[28501]= -2095330553;
assign addr[28502]= -2086621133;
assign addr[28503]= -2077249901;
assign addr[28504]= -2067219829;
assign addr[28505]= -2056534099;
assign addr[28506]= -2045196100;
assign addr[28507]= -2033209426;
assign addr[28508]= -2020577882;
assign addr[28509]= -2007305472;
assign addr[28510]= -1993396407;
assign addr[28511]= -1978855097;
assign addr[28512]= -1963686155;
assign addr[28513]= -1947894393;
assign addr[28514]= -1931484818;
assign addr[28515]= -1914462636;
assign addr[28516]= -1896833245;
assign addr[28517]= -1878602237;
assign addr[28518]= -1859775393;
assign addr[28519]= -1840358687;
assign addr[28520]= -1820358275;
assign addr[28521]= -1799780501;
assign addr[28522]= -1778631892;
assign addr[28523]= -1756919156;
assign addr[28524]= -1734649179;
assign addr[28525]= -1711829025;
assign addr[28526]= -1688465931;
assign addr[28527]= -1664567307;
assign addr[28528]= -1640140734;
assign addr[28529]= -1615193959;
assign addr[28530]= -1589734894;
assign addr[28531]= -1563771613;
assign addr[28532]= -1537312353;
assign addr[28533]= -1510365504;
assign addr[28534]= -1482939614;
assign addr[28535]= -1455043381;
assign addr[28536]= -1426685652;
assign addr[28537]= -1397875423;
assign addr[28538]= -1368621831;
assign addr[28539]= -1338934154;
assign addr[28540]= -1308821808;
assign addr[28541]= -1278294345;
assign addr[28542]= -1247361445;
assign addr[28543]= -1216032921;
assign addr[28544]= -1184318708;
assign addr[28545]= -1152228866;
assign addr[28546]= -1119773573;
assign addr[28547]= -1086963121;
assign addr[28548]= -1053807919;
assign addr[28549]= -1020318481;
assign addr[28550]= -986505429;
assign addr[28551]= -952379488;
assign addr[28552]= -917951481;
assign addr[28553]= -883232329;
assign addr[28554]= -848233042;
assign addr[28555]= -812964722;
assign addr[28556]= -777438554;
assign addr[28557]= -741665807;
assign addr[28558]= -705657826;
assign addr[28559]= -669426032;
assign addr[28560]= -632981917;
assign addr[28561]= -596337040;
assign addr[28562]= -559503022;
assign addr[28563]= -522491548;
assign addr[28564]= -485314355;
assign addr[28565]= -447983235;
assign addr[28566]= -410510029;
assign addr[28567]= -372906622;
assign addr[28568]= -335184940;
assign addr[28569]= -297356948;
assign addr[28570]= -259434643;
assign addr[28571]= -221430054;
assign addr[28572]= -183355234;
assign addr[28573]= -145222259;
assign addr[28574]= -107043224;
assign addr[28575]= -68830239;
assign addr[28576]= -30595422;
assign addr[28577]= 7649098;
assign addr[28578]= 45891193;
assign addr[28579]= 84118732;
assign addr[28580]= 122319591;
assign addr[28581]= 160481654;
assign addr[28582]= 198592817;
assign addr[28583]= 236640993;
assign addr[28584]= 274614114;
assign addr[28585]= 312500135;
assign addr[28586]= 350287041;
assign addr[28587]= 387962847;
assign addr[28588]= 425515602;
assign addr[28589]= 462933398;
assign addr[28590]= 500204365;
assign addr[28591]= 537316682;
assign addr[28592]= 574258580;
assign addr[28593]= 611018340;
assign addr[28594]= 647584304;
assign addr[28595]= 683944874;
assign addr[28596]= 720088517;
assign addr[28597]= 756003771;
assign addr[28598]= 791679244;
assign addr[28599]= 827103620;
assign addr[28600]= 862265664;
assign addr[28601]= 897154224;
assign addr[28602]= 931758235;
assign addr[28603]= 966066720;
assign addr[28604]= 1000068799;
assign addr[28605]= 1033753687;
assign addr[28606]= 1067110699;
assign addr[28607]= 1100129257;
assign addr[28608]= 1132798888;
assign addr[28609]= 1165109230;
assign addr[28610]= 1197050035;
assign addr[28611]= 1228611172;
assign addr[28612]= 1259782632;
assign addr[28613]= 1290554528;
assign addr[28614]= 1320917099;
assign addr[28615]= 1350860716;
assign addr[28616]= 1380375881;
assign addr[28617]= 1409453233;
assign addr[28618]= 1438083551;
assign addr[28619]= 1466257752;
assign addr[28620]= 1493966902;
assign addr[28621]= 1521202211;
assign addr[28622]= 1547955041;
assign addr[28623]= 1574216908;
assign addr[28624]= 1599979481;
assign addr[28625]= 1625234591;
assign addr[28626]= 1649974225;
assign addr[28627]= 1674190539;
assign addr[28628]= 1697875851;
assign addr[28629]= 1721022648;
assign addr[28630]= 1743623590;
assign addr[28631]= 1765671509;
assign addr[28632]= 1787159411;
assign addr[28633]= 1808080480;
assign addr[28634]= 1828428082;
assign addr[28635]= 1848195763;
assign addr[28636]= 1867377253;
assign addr[28637]= 1885966468;
assign addr[28638]= 1903957513;
assign addr[28639]= 1921344681;
assign addr[28640]= 1938122457;
assign addr[28641]= 1954285520;
assign addr[28642]= 1969828744;
assign addr[28643]= 1984747199;
assign addr[28644]= 1999036154;
assign addr[28645]= 2012691075;
assign addr[28646]= 2025707632;
assign addr[28647]= 2038081698;
assign addr[28648]= 2049809346;
assign addr[28649]= 2060886858;
assign addr[28650]= 2071310720;
assign addr[28651]= 2081077626;
assign addr[28652]= 2090184478;
assign addr[28653]= 2098628387;
assign addr[28654]= 2106406677;
assign addr[28655]= 2113516878;
assign addr[28656]= 2119956737;
assign addr[28657]= 2125724211;
assign addr[28658]= 2130817471;
assign addr[28659]= 2135234901;
assign addr[28660]= 2138975100;
assign addr[28661]= 2142036881;
assign addr[28662]= 2144419275;
assign addr[28663]= 2146121524;
assign addr[28664]= 2147143090;
assign addr[28665]= 2147483648;
assign addr[28666]= 2147143090;
assign addr[28667]= 2146121524;
assign addr[28668]= 2144419275;
assign addr[28669]= 2142036881;
assign addr[28670]= 2138975100;
assign addr[28671]= 2135234901;
assign addr[28672]= 2130817471;
assign addr[28673]= 2125724211;
assign addr[28674]= 2119956737;
assign addr[28675]= 2113516878;
assign addr[28676]= 2106406677;
assign addr[28677]= 2098628387;
assign addr[28678]= 2090184478;
assign addr[28679]= 2081077626;
assign addr[28680]= 2071310720;
assign addr[28681]= 2060886858;
assign addr[28682]= 2049809346;
assign addr[28683]= 2038081698;
assign addr[28684]= 2025707632;
assign addr[28685]= 2012691075;
assign addr[28686]= 1999036154;
assign addr[28687]= 1984747199;
assign addr[28688]= 1969828744;
assign addr[28689]= 1954285520;
assign addr[28690]= 1938122457;
assign addr[28691]= 1921344681;
assign addr[28692]= 1903957513;
assign addr[28693]= 1885966468;
assign addr[28694]= 1867377253;
assign addr[28695]= 1848195763;
assign addr[28696]= 1828428082;
assign addr[28697]= 1808080480;
assign addr[28698]= 1787159411;
assign addr[28699]= 1765671509;
assign addr[28700]= 1743623590;
assign addr[28701]= 1721022648;
assign addr[28702]= 1697875851;
assign addr[28703]= 1674190539;
assign addr[28704]= 1649974225;
assign addr[28705]= 1625234591;
assign addr[28706]= 1599979481;
assign addr[28707]= 1574216908;
assign addr[28708]= 1547955041;
assign addr[28709]= 1521202211;
assign addr[28710]= 1493966902;
assign addr[28711]= 1466257752;
assign addr[28712]= 1438083551;
assign addr[28713]= 1409453233;
assign addr[28714]= 1380375881;
assign addr[28715]= 1350860716;
assign addr[28716]= 1320917099;
assign addr[28717]= 1290554528;
assign addr[28718]= 1259782632;
assign addr[28719]= 1228611172;
assign addr[28720]= 1197050035;
assign addr[28721]= 1165109230;
assign addr[28722]= 1132798888;
assign addr[28723]= 1100129257;
assign addr[28724]= 1067110699;
assign addr[28725]= 1033753687;
assign addr[28726]= 1000068799;
assign addr[28727]= 966066720;
assign addr[28728]= 931758235;
assign addr[28729]= 897154224;
assign addr[28730]= 862265664;
assign addr[28731]= 827103620;
assign addr[28732]= 791679244;
assign addr[28733]= 756003771;
assign addr[28734]= 720088517;
assign addr[28735]= 683944874;
assign addr[28736]= 647584304;
assign addr[28737]= 611018340;
assign addr[28738]= 574258580;
assign addr[28739]= 537316682;
assign addr[28740]= 500204365;
assign addr[28741]= 462933398;
assign addr[28742]= 425515602;
assign addr[28743]= 387962847;
assign addr[28744]= 350287041;
assign addr[28745]= 312500135;
assign addr[28746]= 274614114;
assign addr[28747]= 236640993;
assign addr[28748]= 198592817;
assign addr[28749]= 160481654;
assign addr[28750]= 122319591;
assign addr[28751]= 84118732;
assign addr[28752]= 45891193;
assign addr[28753]= 7649098;
assign addr[28754]= -30595422;
assign addr[28755]= -68830239;
assign addr[28756]= -107043224;
assign addr[28757]= -145222259;
assign addr[28758]= -183355234;
assign addr[28759]= -221430054;
assign addr[28760]= -259434643;
assign addr[28761]= -297356948;
assign addr[28762]= -335184940;
assign addr[28763]= -372906622;
assign addr[28764]= -410510029;
assign addr[28765]= -447983235;
assign addr[28766]= -485314355;
assign addr[28767]= -522491548;
assign addr[28768]= -559503022;
assign addr[28769]= -596337040;
assign addr[28770]= -632981917;
assign addr[28771]= -669426032;
assign addr[28772]= -705657826;
assign addr[28773]= -741665807;
assign addr[28774]= -777438554;
assign addr[28775]= -812964722;
assign addr[28776]= -848233042;
assign addr[28777]= -883232329;
assign addr[28778]= -917951481;
assign addr[28779]= -952379488;
assign addr[28780]= -986505429;
assign addr[28781]= -1020318481;
assign addr[28782]= -1053807919;
assign addr[28783]= -1086963121;
assign addr[28784]= -1119773573;
assign addr[28785]= -1152228866;
assign addr[28786]= -1184318708;
assign addr[28787]= -1216032921;
assign addr[28788]= -1247361445;
assign addr[28789]= -1278294345;
assign addr[28790]= -1308821808;
assign addr[28791]= -1338934154;
assign addr[28792]= -1368621831;
assign addr[28793]= -1397875423;
assign addr[28794]= -1426685652;
assign addr[28795]= -1455043381;
assign addr[28796]= -1482939614;
assign addr[28797]= -1510365504;
assign addr[28798]= -1537312353;
assign addr[28799]= -1563771613;
assign addr[28800]= -1589734894;
assign addr[28801]= -1615193959;
assign addr[28802]= -1640140734;
assign addr[28803]= -1664567307;
assign addr[28804]= -1688465931;
assign addr[28805]= -1711829025;
assign addr[28806]= -1734649179;
assign addr[28807]= -1756919156;
assign addr[28808]= -1778631892;
assign addr[28809]= -1799780501;
assign addr[28810]= -1820358275;
assign addr[28811]= -1840358687;
assign addr[28812]= -1859775393;
assign addr[28813]= -1878602237;
assign addr[28814]= -1896833245;
assign addr[28815]= -1914462636;
assign addr[28816]= -1931484818;
assign addr[28817]= -1947894393;
assign addr[28818]= -1963686155;
assign addr[28819]= -1978855097;
assign addr[28820]= -1993396407;
assign addr[28821]= -2007305472;
assign addr[28822]= -2020577882;
assign addr[28823]= -2033209426;
assign addr[28824]= -2045196100;
assign addr[28825]= -2056534099;
assign addr[28826]= -2067219829;
assign addr[28827]= -2077249901;
assign addr[28828]= -2086621133;
assign addr[28829]= -2095330553;
assign addr[28830]= -2103375398;
assign addr[28831]= -2110753117;
assign addr[28832]= -2117461370;
assign addr[28833]= -2123498030;
assign addr[28834]= -2128861181;
assign addr[28835]= -2133549123;
assign addr[28836]= -2137560369;
assign addr[28837]= -2140893646;
assign addr[28838]= -2143547897;
assign addr[28839]= -2145522281;
assign addr[28840]= -2146816171;
assign addr[28841]= -2147429158;
assign addr[28842]= -2147361045;
assign addr[28843]= -2146611856;
assign addr[28844]= -2145181827;
assign addr[28845]= -2143071413;
assign addr[28846]= -2140281282;
assign addr[28847]= -2136812319;
assign addr[28848]= -2132665626;
assign addr[28849]= -2127842516;
assign addr[28850]= -2122344521;
assign addr[28851]= -2116173382;
assign addr[28852]= -2109331059;
assign addr[28853]= -2101819720;
assign addr[28854]= -2093641749;
assign addr[28855]= -2084799740;
assign addr[28856]= -2075296495;
assign addr[28857]= -2065135031;
assign addr[28858]= -2054318569;
assign addr[28859]= -2042850540;
assign addr[28860]= -2030734582;
assign addr[28861]= -2017974537;
assign addr[28862]= -2004574453;
assign addr[28863]= -1990538579;
assign addr[28864]= -1975871368;
assign addr[28865]= -1960577471;
assign addr[28866]= -1944661739;
assign addr[28867]= -1928129220;
assign addr[28868]= -1910985158;
assign addr[28869]= -1893234990;
assign addr[28870]= -1874884346;
assign addr[28871]= -1855939047;
assign addr[28872]= -1836405100;
assign addr[28873]= -1816288703;
assign addr[28874]= -1795596234;
assign addr[28875]= -1774334257;
assign addr[28876]= -1752509516;
assign addr[28877]= -1730128933;
assign addr[28878]= -1707199606;
assign addr[28879]= -1683728808;
assign addr[28880]= -1659723983;
assign addr[28881]= -1635192744;
assign addr[28882]= -1610142873;
assign addr[28883]= -1584582314;
assign addr[28884]= -1558519173;
assign addr[28885]= -1531961719;
assign addr[28886]= -1504918373;
assign addr[28887]= -1477397714;
assign addr[28888]= -1449408469;
assign addr[28889]= -1420959516;
assign addr[28890]= -1392059879;
assign addr[28891]= -1362718723;
assign addr[28892]= -1332945355;
assign addr[28893]= -1302749217;
assign addr[28894]= -1272139887;
assign addr[28895]= -1241127074;
assign addr[28896]= -1209720613;
assign addr[28897]= -1177930466;
assign addr[28898]= -1145766716;
assign addr[28899]= -1113239564;
assign addr[28900]= -1080359326;
assign addr[28901]= -1047136432;
assign addr[28902]= -1013581418;
assign addr[28903]= -979704927;
assign addr[28904]= -945517704;
assign addr[28905]= -911030591;
assign addr[28906]= -876254528;
assign addr[28907]= -841200544;
assign addr[28908]= -805879757;
assign addr[28909]= -770303369;
assign addr[28910]= -734482665;
assign addr[28911]= -698429006;
assign addr[28912]= -662153826;
assign addr[28913]= -625668632;
assign addr[28914]= -588984994;
assign addr[28915]= -552114549;
assign addr[28916]= -515068990;
assign addr[28917]= -477860067;
assign addr[28918]= -440499581;
assign addr[28919]= -402999383;
assign addr[28920]= -365371365;
assign addr[28921]= -327627463;
assign addr[28922]= -289779648;
assign addr[28923]= -251839923;
assign addr[28924]= -213820322;
assign addr[28925]= -175732905;
assign addr[28926]= -137589750;
assign addr[28927]= -99402956;
assign addr[28928]= -61184634;
assign addr[28929]= -22946906;
assign addr[28930]= 15298099;
assign addr[28931]= 53538253;
assign addr[28932]= 91761426;
assign addr[28933]= 129955495;
assign addr[28934]= 168108346;
assign addr[28935]= 206207878;
assign addr[28936]= 244242007;
assign addr[28937]= 282198671;
assign addr[28938]= 320065829;
assign addr[28939]= 357831473;
assign addr[28940]= 395483624;
assign addr[28941]= 433010339;
assign addr[28942]= 470399716;
assign addr[28943]= 507639898;
assign addr[28944]= 544719071;
assign addr[28945]= 581625477;
assign addr[28946]= 618347408;
assign addr[28947]= 654873219;
assign addr[28948]= 691191324;
assign addr[28949]= 727290205;
assign addr[28950]= 763158411;
assign addr[28951]= 798784567;
assign addr[28952]= 834157373;
assign addr[28953]= 869265610;
assign addr[28954]= 904098143;
assign addr[28955]= 938643924;
assign addr[28956]= 972891995;
assign addr[28957]= 1006831495;
assign addr[28958]= 1040451659;
assign addr[28959]= 1073741824;
assign addr[28960]= 1106691431;
assign addr[28961]= 1139290029;
assign addr[28962]= 1171527280;
assign addr[28963]= 1203392958;
assign addr[28964]= 1234876957;
assign addr[28965]= 1265969291;
assign addr[28966]= 1296660098;
assign addr[28967]= 1326939644;
assign addr[28968]= 1356798326;
assign addr[28969]= 1386226674;
assign addr[28970]= 1415215352;
assign addr[28971]= 1443755168;
assign addr[28972]= 1471837070;
assign addr[28973]= 1499452149;
assign addr[28974]= 1526591649;
assign addr[28975]= 1553246960;
assign addr[28976]= 1579409630;
assign addr[28977]= 1605071359;
assign addr[28978]= 1630224009;
assign addr[28979]= 1654859602;
assign addr[28980]= 1678970324;
assign addr[28981]= 1702548529;
assign addr[28982]= 1725586737;
assign addr[28983]= 1748077642;
assign addr[28984]= 1770014111;
assign addr[28985]= 1791389186;
assign addr[28986]= 1812196087;
assign addr[28987]= 1832428215;
assign addr[28988]= 1852079154;
assign addr[28989]= 1871142669;
assign addr[28990]= 1889612716;
assign addr[28991]= 1907483436;
assign addr[28992]= 1924749160;
assign addr[28993]= 1941404413;
assign addr[28994]= 1957443913;
assign addr[28995]= 1972862571;
assign addr[28996]= 1987655498;
assign addr[28997]= 2001818002;
assign addr[28998]= 2015345591;
assign addr[28999]= 2028233973;
assign addr[29000]= 2040479063;
assign addr[29001]= 2052076975;
assign addr[29002]= 2063024031;
assign addr[29003]= 2073316760;
assign addr[29004]= 2082951896;
assign addr[29005]= 2091926384;
assign addr[29006]= 2100237377;
assign addr[29007]= 2107882239;
assign addr[29008]= 2114858546;
assign addr[29009]= 2121164085;
assign addr[29010]= 2126796855;
assign addr[29011]= 2131755071;
assign addr[29012]= 2136037160;
assign addr[29013]= 2139641764;
assign addr[29014]= 2142567738;
assign addr[29015]= 2144814157;
assign addr[29016]= 2146380306;
assign addr[29017]= 2147265689;
assign addr[29018]= 2147470025;
assign addr[29019]= 2146993250;
assign addr[29020]= 2145835515;
assign addr[29021]= 2143997187;
assign addr[29022]= 2141478848;
assign addr[29023]= 2138281298;
assign addr[29024]= 2134405552;
assign addr[29025]= 2129852837;
assign addr[29026]= 2124624598;
assign addr[29027]= 2118722494;
assign addr[29028]= 2112148396;
assign addr[29029]= 2104904390;
assign addr[29030]= 2096992772;
assign addr[29031]= 2088416053;
assign addr[29032]= 2079176953;
assign addr[29033]= 2069278401;
assign addr[29034]= 2058723538;
assign addr[29035]= 2047515711;
assign addr[29036]= 2035658475;
assign addr[29037]= 2023155591;
assign addr[29038]= 2010011024;
assign addr[29039]= 1996228943;
assign addr[29040]= 1981813720;
assign addr[29041]= 1966769926;
assign addr[29042]= 1951102334;
assign addr[29043]= 1934815911;
assign addr[29044]= 1917915825;
assign addr[29045]= 1900407434;
assign addr[29046]= 1882296293;
assign addr[29047]= 1863588145;
assign addr[29048]= 1844288924;
assign addr[29049]= 1824404752;
assign addr[29050]= 1803941934;
assign addr[29051]= 1782906961;
assign addr[29052]= 1761306505;
assign addr[29053]= 1739147417;
assign addr[29054]= 1716436725;
assign addr[29055]= 1693181631;
assign addr[29056]= 1669389513;
assign addr[29057]= 1645067915;
assign addr[29058]= 1620224553;
assign addr[29059]= 1594867305;
assign addr[29060]= 1569004214;
assign addr[29061]= 1542643483;
assign addr[29062]= 1515793473;
assign addr[29063]= 1488462700;
assign addr[29064]= 1460659832;
assign addr[29065]= 1432393688;
assign addr[29066]= 1403673233;
assign addr[29067]= 1374507575;
assign addr[29068]= 1344905966;
assign addr[29069]= 1314877795;
assign addr[29070]= 1284432584;
assign addr[29071]= 1253579991;
assign addr[29072]= 1222329801;
assign addr[29073]= 1190691925;
assign addr[29074]= 1158676398;
assign addr[29075]= 1126293375;
assign addr[29076]= 1093553126;
assign addr[29077]= 1060466036;
assign addr[29078]= 1027042599;
assign addr[29079]= 993293415;
assign addr[29080]= 959229189;
assign addr[29081]= 924860725;
assign addr[29082]= 890198924;
assign addr[29083]= 855254778;
assign addr[29084]= 820039373;
assign addr[29085]= 784563876;
assign addr[29086]= 748839539;
assign addr[29087]= 712877694;
assign addr[29088]= 676689746;
assign addr[29089]= 640287172;
assign addr[29090]= 603681519;
assign addr[29091]= 566884397;
assign addr[29092]= 529907477;
assign addr[29093]= 492762486;
assign addr[29094]= 455461206;
assign addr[29095]= 418015468;
assign addr[29096]= 380437148;
assign addr[29097]= 342738165;
assign addr[29098]= 304930476;
assign addr[29099]= 267026072;
assign addr[29100]= 229036977;
assign addr[29101]= 190975237;
assign addr[29102]= 152852926;
assign addr[29103]= 114682135;
assign addr[29104]= 76474970;
assign addr[29105]= 38243550;
assign addr[29106]= 0;
assign addr[29107]= -38243550;
assign addr[29108]= -76474970;
assign addr[29109]= -114682135;
assign addr[29110]= -152852926;
assign addr[29111]= -190975237;
assign addr[29112]= -229036977;
assign addr[29113]= -267026072;
assign addr[29114]= -304930476;
assign addr[29115]= -342738165;
assign addr[29116]= -380437148;
assign addr[29117]= -418015468;
assign addr[29118]= -455461206;
assign addr[29119]= -492762486;
assign addr[29120]= -529907477;
assign addr[29121]= -566884397;
assign addr[29122]= -603681519;
assign addr[29123]= -640287172;
assign addr[29124]= -676689746;
assign addr[29125]= -712877694;
assign addr[29126]= -748839539;
assign addr[29127]= -784563876;
assign addr[29128]= -820039373;
assign addr[29129]= -855254778;
assign addr[29130]= -890198924;
assign addr[29131]= -924860725;
assign addr[29132]= -959229189;
assign addr[29133]= -993293415;
assign addr[29134]= -1027042599;
assign addr[29135]= -1060466036;
assign addr[29136]= -1093553126;
assign addr[29137]= -1126293375;
assign addr[29138]= -1158676398;
assign addr[29139]= -1190691925;
assign addr[29140]= -1222329801;
assign addr[29141]= -1253579991;
assign addr[29142]= -1284432584;
assign addr[29143]= -1314877795;
assign addr[29144]= -1344905966;
assign addr[29145]= -1374507575;
assign addr[29146]= -1403673233;
assign addr[29147]= -1432393688;
assign addr[29148]= -1460659832;
assign addr[29149]= -1488462700;
assign addr[29150]= -1515793473;
assign addr[29151]= -1542643483;
assign addr[29152]= -1569004214;
assign addr[29153]= -1594867305;
assign addr[29154]= -1620224553;
assign addr[29155]= -1645067915;
assign addr[29156]= -1669389513;
assign addr[29157]= -1693181631;
assign addr[29158]= -1716436725;
assign addr[29159]= -1739147417;
assign addr[29160]= -1761306505;
assign addr[29161]= -1782906961;
assign addr[29162]= -1803941934;
assign addr[29163]= -1824404752;
assign addr[29164]= -1844288924;
assign addr[29165]= -1863588145;
assign addr[29166]= -1882296293;
assign addr[29167]= -1900407434;
assign addr[29168]= -1917915825;
assign addr[29169]= -1934815911;
assign addr[29170]= -1951102334;
assign addr[29171]= -1966769926;
assign addr[29172]= -1981813720;
assign addr[29173]= -1996228943;
assign addr[29174]= -2010011024;
assign addr[29175]= -2023155591;
assign addr[29176]= -2035658475;
assign addr[29177]= -2047515711;
assign addr[29178]= -2058723538;
assign addr[29179]= -2069278401;
assign addr[29180]= -2079176953;
assign addr[29181]= -2088416053;
assign addr[29182]= -2096992772;
assign addr[29183]= -2104904390;
assign addr[29184]= -2112148396;
assign addr[29185]= -2118722494;
assign addr[29186]= -2124624598;
assign addr[29187]= -2129852837;
assign addr[29188]= -2134405552;
assign addr[29189]= -2138281298;
assign addr[29190]= -2141478848;
assign addr[29191]= -2143997187;
assign addr[29192]= -2145835515;
assign addr[29193]= -2146993250;
assign addr[29194]= -2147470025;
assign addr[29195]= -2147265689;
assign addr[29196]= -2146380306;
assign addr[29197]= -2144814157;
assign addr[29198]= -2142567738;
assign addr[29199]= -2139641764;
assign addr[29200]= -2136037160;
assign addr[29201]= -2131755071;
assign addr[29202]= -2126796855;
assign addr[29203]= -2121164085;
assign addr[29204]= -2114858546;
assign addr[29205]= -2107882239;
assign addr[29206]= -2100237377;
assign addr[29207]= -2091926384;
assign addr[29208]= -2082951896;
assign addr[29209]= -2073316760;
assign addr[29210]= -2063024031;
assign addr[29211]= -2052076975;
assign addr[29212]= -2040479063;
assign addr[29213]= -2028233973;
assign addr[29214]= -2015345591;
assign addr[29215]= -2001818002;
assign addr[29216]= -1987655498;
assign addr[29217]= -1972862571;
assign addr[29218]= -1957443913;
assign addr[29219]= -1941404413;
assign addr[29220]= -1924749160;
assign addr[29221]= -1907483436;
assign addr[29222]= -1889612716;
assign addr[29223]= -1871142669;
assign addr[29224]= -1852079154;
assign addr[29225]= -1832428215;
assign addr[29226]= -1812196087;
assign addr[29227]= -1791389186;
assign addr[29228]= -1770014111;
assign addr[29229]= -1748077642;
assign addr[29230]= -1725586737;
assign addr[29231]= -1702548529;
assign addr[29232]= -1678970324;
assign addr[29233]= -1654859602;
assign addr[29234]= -1630224009;
assign addr[29235]= -1605071359;
assign addr[29236]= -1579409630;
assign addr[29237]= -1553246960;
assign addr[29238]= -1526591649;
assign addr[29239]= -1499452149;
assign addr[29240]= -1471837070;
assign addr[29241]= -1443755168;
assign addr[29242]= -1415215352;
assign addr[29243]= -1386226674;
assign addr[29244]= -1356798326;
assign addr[29245]= -1326939644;
assign addr[29246]= -1296660098;
assign addr[29247]= -1265969291;
assign addr[29248]= -1234876957;
assign addr[29249]= -1203392958;
assign addr[29250]= -1171527280;
assign addr[29251]= -1139290029;
assign addr[29252]= -1106691431;
assign addr[29253]= -1073741824;
assign addr[29254]= -1040451659;
assign addr[29255]= -1006831495;
assign addr[29256]= -972891995;
assign addr[29257]= -938643924;
assign addr[29258]= -904098143;
assign addr[29259]= -869265610;
assign addr[29260]= -834157373;
assign addr[29261]= -798784567;
assign addr[29262]= -763158411;
assign addr[29263]= -727290205;
assign addr[29264]= -691191324;
assign addr[29265]= -654873219;
assign addr[29266]= -618347408;
assign addr[29267]= -581625477;
assign addr[29268]= -544719071;
assign addr[29269]= -507639898;
assign addr[29270]= -470399716;
assign addr[29271]= -433010339;
assign addr[29272]= -395483624;
assign addr[29273]= -357831473;
assign addr[29274]= -320065829;
assign addr[29275]= -282198671;
assign addr[29276]= -244242007;
assign addr[29277]= -206207878;
assign addr[29278]= -168108346;
assign addr[29279]= -129955495;
assign addr[29280]= -91761426;
assign addr[29281]= -53538253;
assign addr[29282]= -15298099;
assign addr[29283]= 22946906;
assign addr[29284]= 61184634;
assign addr[29285]= 99402956;
assign addr[29286]= 137589750;
assign addr[29287]= 175732905;
assign addr[29288]= 213820322;
assign addr[29289]= 251839923;
assign addr[29290]= 289779648;
assign addr[29291]= 327627463;
assign addr[29292]= 365371365;
assign addr[29293]= 402999383;
assign addr[29294]= 440499581;
assign addr[29295]= 477860067;
assign addr[29296]= 515068990;
assign addr[29297]= 552114549;
assign addr[29298]= 588984994;
assign addr[29299]= 625668632;
assign addr[29300]= 662153826;
assign addr[29301]= 698429006;
assign addr[29302]= 734482665;
assign addr[29303]= 770303369;
assign addr[29304]= 805879757;
assign addr[29305]= 841200544;
assign addr[29306]= 876254528;
assign addr[29307]= 911030591;
assign addr[29308]= 945517704;
assign addr[29309]= 979704927;
assign addr[29310]= 1013581418;
assign addr[29311]= 1047136432;
assign addr[29312]= 1080359326;
assign addr[29313]= 1113239564;
assign addr[29314]= 1145766716;
assign addr[29315]= 1177930466;
assign addr[29316]= 1209720613;
assign addr[29317]= 1241127074;
assign addr[29318]= 1272139887;
assign addr[29319]= 1302749217;
assign addr[29320]= 1332945355;
assign addr[29321]= 1362718723;
assign addr[29322]= 1392059879;
assign addr[29323]= 1420959516;
assign addr[29324]= 1449408469;
assign addr[29325]= 1477397714;
assign addr[29326]= 1504918373;
assign addr[29327]= 1531961719;
assign addr[29328]= 1558519173;
assign addr[29329]= 1584582314;
assign addr[29330]= 1610142873;
assign addr[29331]= 1635192744;
assign addr[29332]= 1659723983;
assign addr[29333]= 1683728808;
assign addr[29334]= 1707199606;
assign addr[29335]= 1730128933;
assign addr[29336]= 1752509516;
assign addr[29337]= 1774334257;
assign addr[29338]= 1795596234;
assign addr[29339]= 1816288703;
assign addr[29340]= 1836405100;
assign addr[29341]= 1855939047;
assign addr[29342]= 1874884346;
assign addr[29343]= 1893234990;
assign addr[29344]= 1910985158;
assign addr[29345]= 1928129220;
assign addr[29346]= 1944661739;
assign addr[29347]= 1960577471;
assign addr[29348]= 1975871368;
assign addr[29349]= 1990538579;
assign addr[29350]= 2004574453;
assign addr[29351]= 2017974537;
assign addr[29352]= 2030734582;
assign addr[29353]= 2042850540;
assign addr[29354]= 2054318569;
assign addr[29355]= 2065135031;
assign addr[29356]= 2075296495;
assign addr[29357]= 2084799740;
assign addr[29358]= 2093641749;
assign addr[29359]= 2101819720;
assign addr[29360]= 2109331059;
assign addr[29361]= 2116173382;
assign addr[29362]= 2122344521;
assign addr[29363]= 2127842516;
assign addr[29364]= 2132665626;
assign addr[29365]= 2136812319;
assign addr[29366]= 2140281282;
assign addr[29367]= 2143071413;
assign addr[29368]= 2145181827;
assign addr[29369]= 2146611856;
assign addr[29370]= 2147361045;
assign addr[29371]= 2147429158;
assign addr[29372]= 2146816171;
assign addr[29373]= 2145522281;
assign addr[29374]= 2143547897;
assign addr[29375]= 2140893646;
assign addr[29376]= 2137560369;
assign addr[29377]= 2133549123;
assign addr[29378]= 2128861181;
assign addr[29379]= 2123498030;
assign addr[29380]= 2117461370;
assign addr[29381]= 2110753117;
assign addr[29382]= 2103375398;
assign addr[29383]= 2095330553;
assign addr[29384]= 2086621133;
assign addr[29385]= 2077249901;
assign addr[29386]= 2067219829;
assign addr[29387]= 2056534099;
assign addr[29388]= 2045196100;
assign addr[29389]= 2033209426;
assign addr[29390]= 2020577882;
assign addr[29391]= 2007305472;
assign addr[29392]= 1993396407;
assign addr[29393]= 1978855097;
assign addr[29394]= 1963686155;
assign addr[29395]= 1947894393;
assign addr[29396]= 1931484818;
assign addr[29397]= 1914462636;
assign addr[29398]= 1896833245;
assign addr[29399]= 1878602237;
assign addr[29400]= 1859775393;
assign addr[29401]= 1840358687;
assign addr[29402]= 1820358275;
assign addr[29403]= 1799780501;
assign addr[29404]= 1778631892;
assign addr[29405]= 1756919156;
assign addr[29406]= 1734649179;
assign addr[29407]= 1711829025;
assign addr[29408]= 1688465931;
assign addr[29409]= 1664567307;
assign addr[29410]= 1640140734;
assign addr[29411]= 1615193959;
assign addr[29412]= 1589734894;
assign addr[29413]= 1563771613;
assign addr[29414]= 1537312353;
assign addr[29415]= 1510365504;
assign addr[29416]= 1482939614;
assign addr[29417]= 1455043381;
assign addr[29418]= 1426685652;
assign addr[29419]= 1397875423;
assign addr[29420]= 1368621831;
assign addr[29421]= 1338934154;
assign addr[29422]= 1308821808;
assign addr[29423]= 1278294345;
assign addr[29424]= 1247361445;
assign addr[29425]= 1216032921;
assign addr[29426]= 1184318708;
assign addr[29427]= 1152228866;
assign addr[29428]= 1119773573;
assign addr[29429]= 1086963121;
assign addr[29430]= 1053807919;
assign addr[29431]= 1020318481;
assign addr[29432]= 986505429;
assign addr[29433]= 952379488;
assign addr[29434]= 917951481;
assign addr[29435]= 883232329;
assign addr[29436]= 848233042;
assign addr[29437]= 812964722;
assign addr[29438]= 777438554;
assign addr[29439]= 741665807;
assign addr[29440]= 705657826;
assign addr[29441]= 669426032;
assign addr[29442]= 632981917;
assign addr[29443]= 596337040;
assign addr[29444]= 559503022;
assign addr[29445]= 522491548;
assign addr[29446]= 485314355;
assign addr[29447]= 447983235;
assign addr[29448]= 410510029;
assign addr[29449]= 372906622;
assign addr[29450]= 335184940;
assign addr[29451]= 297356948;
assign addr[29452]= 259434643;
assign addr[29453]= 221430054;
assign addr[29454]= 183355234;
assign addr[29455]= 145222259;
assign addr[29456]= 107043224;
assign addr[29457]= 68830239;
assign addr[29458]= 30595422;
assign addr[29459]= -7649098;
assign addr[29460]= -45891193;
assign addr[29461]= -84118732;
assign addr[29462]= -122319591;
assign addr[29463]= -160481654;
assign addr[29464]= -198592817;
assign addr[29465]= -236640993;
assign addr[29466]= -274614114;
assign addr[29467]= -312500135;
assign addr[29468]= -350287041;
assign addr[29469]= -387962847;
assign addr[29470]= -425515602;
assign addr[29471]= -462933398;
assign addr[29472]= -500204365;
assign addr[29473]= -537316682;
assign addr[29474]= -574258580;
assign addr[29475]= -611018340;
assign addr[29476]= -647584304;
assign addr[29477]= -683944874;
assign addr[29478]= -720088517;
assign addr[29479]= -756003771;
assign addr[29480]= -791679244;
assign addr[29481]= -827103620;
assign addr[29482]= -862265664;
assign addr[29483]= -897154224;
assign addr[29484]= -931758235;
assign addr[29485]= -966066720;
assign addr[29486]= -1000068799;
assign addr[29487]= -1033753687;
assign addr[29488]= -1067110699;
assign addr[29489]= -1100129257;
assign addr[29490]= -1132798888;
assign addr[29491]= -1165109230;
assign addr[29492]= -1197050035;
assign addr[29493]= -1228611172;
assign addr[29494]= -1259782632;
assign addr[29495]= -1290554528;
assign addr[29496]= -1320917099;
assign addr[29497]= -1350860716;
assign addr[29498]= -1380375881;
assign addr[29499]= -1409453233;
assign addr[29500]= -1438083551;
assign addr[29501]= -1466257752;
assign addr[29502]= -1493966902;
assign addr[29503]= -1521202211;
assign addr[29504]= -1547955041;
assign addr[29505]= -1574216908;
assign addr[29506]= -1599979481;
assign addr[29507]= -1625234591;
assign addr[29508]= -1649974225;
assign addr[29509]= -1674190539;
assign addr[29510]= -1697875851;
assign addr[29511]= -1721022648;
assign addr[29512]= -1743623590;
assign addr[29513]= -1765671509;
assign addr[29514]= -1787159411;
assign addr[29515]= -1808080480;
assign addr[29516]= -1828428082;
assign addr[29517]= -1848195763;
assign addr[29518]= -1867377253;
assign addr[29519]= -1885966468;
assign addr[29520]= -1903957513;
assign addr[29521]= -1921344681;
assign addr[29522]= -1938122457;
assign addr[29523]= -1954285520;
assign addr[29524]= -1969828744;
assign addr[29525]= -1984747199;
assign addr[29526]= -1999036154;
assign addr[29527]= -2012691075;
assign addr[29528]= -2025707632;
assign addr[29529]= -2038081698;
assign addr[29530]= -2049809346;
assign addr[29531]= -2060886858;
assign addr[29532]= -2071310720;
assign addr[29533]= -2081077626;
assign addr[29534]= -2090184478;
assign addr[29535]= -2098628387;
assign addr[29536]= -2106406677;
assign addr[29537]= -2113516878;
assign addr[29538]= -2119956737;
assign addr[29539]= -2125724211;
assign addr[29540]= -2130817471;
assign addr[29541]= -2135234901;
assign addr[29542]= -2138975100;
assign addr[29543]= -2142036881;
assign addr[29544]= -2144419275;
assign addr[29545]= -2146121524;
assign addr[29546]= -2147143090;
assign addr[29547]= -2147483648;
assign addr[29548]= -2147143090;
assign addr[29549]= -2146121524;
assign addr[29550]= -2144419275;
assign addr[29551]= -2142036881;
assign addr[29552]= -2138975100;
assign addr[29553]= -2135234901;
assign addr[29554]= -2130817471;
assign addr[29555]= -2125724211;
assign addr[29556]= -2119956737;
assign addr[29557]= -2113516878;
assign addr[29558]= -2106406677;
assign addr[29559]= -2098628387;
assign addr[29560]= -2090184478;
assign addr[29561]= -2081077626;
assign addr[29562]= -2071310720;
assign addr[29563]= -2060886858;
assign addr[29564]= -2049809346;
assign addr[29565]= -2038081698;
assign addr[29566]= -2025707632;
assign addr[29567]= -2012691075;
assign addr[29568]= -1999036154;
assign addr[29569]= -1984747199;
assign addr[29570]= -1969828744;
assign addr[29571]= -1954285520;
assign addr[29572]= -1938122457;
assign addr[29573]= -1921344681;
assign addr[29574]= -1903957513;
assign addr[29575]= -1885966468;
assign addr[29576]= -1867377253;
assign addr[29577]= -1848195763;
assign addr[29578]= -1828428082;
assign addr[29579]= -1808080480;
assign addr[29580]= -1787159411;
assign addr[29581]= -1765671509;
assign addr[29582]= -1743623590;
assign addr[29583]= -1721022648;
assign addr[29584]= -1697875851;
assign addr[29585]= -1674190539;
assign addr[29586]= -1649974225;
assign addr[29587]= -1625234591;
assign addr[29588]= -1599979481;
assign addr[29589]= -1574216908;
assign addr[29590]= -1547955041;
assign addr[29591]= -1521202211;
assign addr[29592]= -1493966902;
assign addr[29593]= -1466257752;
assign addr[29594]= -1438083551;
assign addr[29595]= -1409453233;
assign addr[29596]= -1380375881;
assign addr[29597]= -1350860716;
assign addr[29598]= -1320917099;
assign addr[29599]= -1290554528;
assign addr[29600]= -1259782632;
assign addr[29601]= -1228611172;
assign addr[29602]= -1197050035;
assign addr[29603]= -1165109230;
assign addr[29604]= -1132798888;
assign addr[29605]= -1100129257;
assign addr[29606]= -1067110699;
assign addr[29607]= -1033753687;
assign addr[29608]= -1000068799;
assign addr[29609]= -966066720;
assign addr[29610]= -931758235;
assign addr[29611]= -897154224;
assign addr[29612]= -862265664;
assign addr[29613]= -827103620;
assign addr[29614]= -791679244;
assign addr[29615]= -756003771;
assign addr[29616]= -720088517;
assign addr[29617]= -683944874;
assign addr[29618]= -647584304;
assign addr[29619]= -611018340;
assign addr[29620]= -574258580;
assign addr[29621]= -537316682;
assign addr[29622]= -500204365;
assign addr[29623]= -462933398;
assign addr[29624]= -425515602;
assign addr[29625]= -387962847;
assign addr[29626]= -350287041;
assign addr[29627]= -312500135;
assign addr[29628]= -274614114;
assign addr[29629]= -236640993;
assign addr[29630]= -198592817;
assign addr[29631]= -160481654;
assign addr[29632]= -122319591;
assign addr[29633]= -84118732;
assign addr[29634]= -45891193;
assign addr[29635]= -7649098;
assign addr[29636]= 30595422;
assign addr[29637]= 68830239;
assign addr[29638]= 107043224;
assign addr[29639]= 145222259;
assign addr[29640]= 183355234;
assign addr[29641]= 221430054;
assign addr[29642]= 259434643;
assign addr[29643]= 297356948;
assign addr[29644]= 335184940;
assign addr[29645]= 372906622;
assign addr[29646]= 410510029;
assign addr[29647]= 447983235;
assign addr[29648]= 485314355;
assign addr[29649]= 522491548;
assign addr[29650]= 559503022;
assign addr[29651]= 596337040;
assign addr[29652]= 632981917;
assign addr[29653]= 669426032;
assign addr[29654]= 705657826;
assign addr[29655]= 741665807;
assign addr[29656]= 777438554;
assign addr[29657]= 812964722;
assign addr[29658]= 848233042;
assign addr[29659]= 883232329;
assign addr[29660]= 917951481;
assign addr[29661]= 952379488;
assign addr[29662]= 986505429;
assign addr[29663]= 1020318481;
assign addr[29664]= 1053807919;
assign addr[29665]= 1086963121;
assign addr[29666]= 1119773573;
assign addr[29667]= 1152228866;
assign addr[29668]= 1184318708;
assign addr[29669]= 1216032921;
assign addr[29670]= 1247361445;
assign addr[29671]= 1278294345;
assign addr[29672]= 1308821808;
assign addr[29673]= 1338934154;
assign addr[29674]= 1368621831;
assign addr[29675]= 1397875423;
assign addr[29676]= 1426685652;
assign addr[29677]= 1455043381;
assign addr[29678]= 1482939614;
assign addr[29679]= 1510365504;
assign addr[29680]= 1537312353;
assign addr[29681]= 1563771613;
assign addr[29682]= 1589734894;
assign addr[29683]= 1615193959;
assign addr[29684]= 1640140734;
assign addr[29685]= 1664567307;
assign addr[29686]= 1688465931;
assign addr[29687]= 1711829025;
assign addr[29688]= 1734649179;
assign addr[29689]= 1756919156;
assign addr[29690]= 1778631892;
assign addr[29691]= 1799780501;
assign addr[29692]= 1820358275;
assign addr[29693]= 1840358687;
assign addr[29694]= 1859775393;
assign addr[29695]= 1878602237;
assign addr[29696]= 1896833245;
assign addr[29697]= 1914462636;
assign addr[29698]= 1931484818;
assign addr[29699]= 1947894393;
assign addr[29700]= 1963686155;
assign addr[29701]= 1978855097;
assign addr[29702]= 1993396407;
assign addr[29703]= 2007305472;
assign addr[29704]= 2020577882;
assign addr[29705]= 2033209426;
assign addr[29706]= 2045196100;
assign addr[29707]= 2056534099;
assign addr[29708]= 2067219829;
assign addr[29709]= 2077249901;
assign addr[29710]= 2086621133;
assign addr[29711]= 2095330553;
assign addr[29712]= 2103375398;
assign addr[29713]= 2110753117;
assign addr[29714]= 2117461370;
assign addr[29715]= 2123498030;
assign addr[29716]= 2128861181;
assign addr[29717]= 2133549123;
assign addr[29718]= 2137560369;
assign addr[29719]= 2140893646;
assign addr[29720]= 2143547897;
assign addr[29721]= 2145522281;
assign addr[29722]= 2146816171;
assign addr[29723]= 2147429158;
assign addr[29724]= 2147361045;
assign addr[29725]= 2146611856;
assign addr[29726]= 2145181827;
assign addr[29727]= 2143071413;
assign addr[29728]= 2140281282;
assign addr[29729]= 2136812319;
assign addr[29730]= 2132665626;
assign addr[29731]= 2127842516;
assign addr[29732]= 2122344521;
assign addr[29733]= 2116173382;
assign addr[29734]= 2109331059;
assign addr[29735]= 2101819720;
assign addr[29736]= 2093641749;
assign addr[29737]= 2084799740;
assign addr[29738]= 2075296495;
assign addr[29739]= 2065135031;
assign addr[29740]= 2054318569;
assign addr[29741]= 2042850540;
assign addr[29742]= 2030734582;
assign addr[29743]= 2017974537;
assign addr[29744]= 2004574453;
assign addr[29745]= 1990538579;
assign addr[29746]= 1975871368;
assign addr[29747]= 1960577471;
assign addr[29748]= 1944661739;
assign addr[29749]= 1928129220;
assign addr[29750]= 1910985158;
assign addr[29751]= 1893234990;
assign addr[29752]= 1874884346;
assign addr[29753]= 1855939047;
assign addr[29754]= 1836405100;
assign addr[29755]= 1816288703;
assign addr[29756]= 1795596234;
assign addr[29757]= 1774334257;
assign addr[29758]= 1752509516;
assign addr[29759]= 1730128933;
assign addr[29760]= 1707199606;
assign addr[29761]= 1683728808;
assign addr[29762]= 1659723983;
assign addr[29763]= 1635192744;
assign addr[29764]= 1610142873;
assign addr[29765]= 1584582314;
assign addr[29766]= 1558519173;
assign addr[29767]= 1531961719;
assign addr[29768]= 1504918373;
assign addr[29769]= 1477397714;
assign addr[29770]= 1449408469;
assign addr[29771]= 1420959516;
assign addr[29772]= 1392059879;
assign addr[29773]= 1362718723;
assign addr[29774]= 1332945355;
assign addr[29775]= 1302749217;
assign addr[29776]= 1272139887;
assign addr[29777]= 1241127074;
assign addr[29778]= 1209720613;
assign addr[29779]= 1177930466;
assign addr[29780]= 1145766716;
assign addr[29781]= 1113239564;
assign addr[29782]= 1080359326;
assign addr[29783]= 1047136432;
assign addr[29784]= 1013581418;
assign addr[29785]= 979704927;
assign addr[29786]= 945517704;
assign addr[29787]= 911030591;
assign addr[29788]= 876254528;
assign addr[29789]= 841200544;
assign addr[29790]= 805879757;
assign addr[29791]= 770303369;
assign addr[29792]= 734482665;
assign addr[29793]= 698429006;
assign addr[29794]= 662153826;
assign addr[29795]= 625668632;
assign addr[29796]= 588984994;
assign addr[29797]= 552114549;
assign addr[29798]= 515068990;
assign addr[29799]= 477860067;
assign addr[29800]= 440499581;
assign addr[29801]= 402999383;
assign addr[29802]= 365371365;
assign addr[29803]= 327627463;
assign addr[29804]= 289779648;
assign addr[29805]= 251839923;
assign addr[29806]= 213820322;
assign addr[29807]= 175732905;
assign addr[29808]= 137589750;
assign addr[29809]= 99402956;
assign addr[29810]= 61184634;
assign addr[29811]= 22946906;
assign addr[29812]= -15298099;
assign addr[29813]= -53538253;
assign addr[29814]= -91761426;
assign addr[29815]= -129955495;
assign addr[29816]= -168108346;
assign addr[29817]= -206207878;
assign addr[29818]= -244242007;
assign addr[29819]= -282198671;
assign addr[29820]= -320065829;
assign addr[29821]= -357831473;
assign addr[29822]= -395483624;
assign addr[29823]= -433010339;
assign addr[29824]= -470399716;
assign addr[29825]= -507639898;
assign addr[29826]= -544719071;
assign addr[29827]= -581625477;
assign addr[29828]= -618347408;
assign addr[29829]= -654873219;
assign addr[29830]= -691191324;
assign addr[29831]= -727290205;
assign addr[29832]= -763158411;
assign addr[29833]= -798784567;
assign addr[29834]= -834157373;
assign addr[29835]= -869265610;
assign addr[29836]= -904098143;
assign addr[29837]= -938643924;
assign addr[29838]= -972891995;
assign addr[29839]= -1006831495;
assign addr[29840]= -1040451659;
assign addr[29841]= -1073741824;
assign addr[29842]= -1106691431;
assign addr[29843]= -1139290029;
assign addr[29844]= -1171527280;
assign addr[29845]= -1203392958;
assign addr[29846]= -1234876957;
assign addr[29847]= -1265969291;
assign addr[29848]= -1296660098;
assign addr[29849]= -1326939644;
assign addr[29850]= -1356798326;
assign addr[29851]= -1386226674;
assign addr[29852]= -1415215352;
assign addr[29853]= -1443755168;
assign addr[29854]= -1471837070;
assign addr[29855]= -1499452149;
assign addr[29856]= -1526591649;
assign addr[29857]= -1553246960;
assign addr[29858]= -1579409630;
assign addr[29859]= -1605071359;
assign addr[29860]= -1630224009;
assign addr[29861]= -1654859602;
assign addr[29862]= -1678970324;
assign addr[29863]= -1702548529;
assign addr[29864]= -1725586737;
assign addr[29865]= -1748077642;
assign addr[29866]= -1770014111;
assign addr[29867]= -1791389186;
assign addr[29868]= -1812196087;
assign addr[29869]= -1832428215;
assign addr[29870]= -1852079154;
assign addr[29871]= -1871142669;
assign addr[29872]= -1889612716;
assign addr[29873]= -1907483436;
assign addr[29874]= -1924749160;
assign addr[29875]= -1941404413;
assign addr[29876]= -1957443913;
assign addr[29877]= -1972862571;
assign addr[29878]= -1987655498;
assign addr[29879]= -2001818002;
assign addr[29880]= -2015345591;
assign addr[29881]= -2028233973;
assign addr[29882]= -2040479063;
assign addr[29883]= -2052076975;
assign addr[29884]= -2063024031;
assign addr[29885]= -2073316760;
assign addr[29886]= -2082951896;
assign addr[29887]= -2091926384;
assign addr[29888]= -2100237377;
assign addr[29889]= -2107882239;
assign addr[29890]= -2114858546;
assign addr[29891]= -2121164085;
assign addr[29892]= -2126796855;
assign addr[29893]= -2131755071;
assign addr[29894]= -2136037160;
assign addr[29895]= -2139641764;
assign addr[29896]= -2142567738;
assign addr[29897]= -2144814157;
assign addr[29898]= -2146380306;
assign addr[29899]= -2147265689;
assign addr[29900]= -2147470025;
assign addr[29901]= -2146993250;
assign addr[29902]= -2145835515;
assign addr[29903]= -2143997187;
assign addr[29904]= -2141478848;
assign addr[29905]= -2138281298;
assign addr[29906]= -2134405552;
assign addr[29907]= -2129852837;
assign addr[29908]= -2124624598;
assign addr[29909]= -2118722494;
assign addr[29910]= -2112148396;
assign addr[29911]= -2104904390;
assign addr[29912]= -2096992772;
assign addr[29913]= -2088416053;
assign addr[29914]= -2079176953;
assign addr[29915]= -2069278401;
assign addr[29916]= -2058723538;
assign addr[29917]= -2047515711;
assign addr[29918]= -2035658475;
assign addr[29919]= -2023155591;
assign addr[29920]= -2010011024;
assign addr[29921]= -1996228943;
assign addr[29922]= -1981813720;
assign addr[29923]= -1966769926;
assign addr[29924]= -1951102334;
assign addr[29925]= -1934815911;
assign addr[29926]= -1917915825;
assign addr[29927]= -1900407434;
assign addr[29928]= -1882296293;
assign addr[29929]= -1863588145;
assign addr[29930]= -1844288924;
assign addr[29931]= -1824404752;
assign addr[29932]= -1803941934;
assign addr[29933]= -1782906961;
assign addr[29934]= -1761306505;
assign addr[29935]= -1739147417;
assign addr[29936]= -1716436725;
assign addr[29937]= -1693181631;
assign addr[29938]= -1669389513;
assign addr[29939]= -1645067915;
assign addr[29940]= -1620224553;
assign addr[29941]= -1594867305;
assign addr[29942]= -1569004214;
assign addr[29943]= -1542643483;
assign addr[29944]= -1515793473;
assign addr[29945]= -1488462700;
assign addr[29946]= -1460659832;
assign addr[29947]= -1432393688;
assign addr[29948]= -1403673233;
assign addr[29949]= -1374507575;
assign addr[29950]= -1344905966;
assign addr[29951]= -1314877795;
assign addr[29952]= -1284432584;
assign addr[29953]= -1253579991;
assign addr[29954]= -1222329801;
assign addr[29955]= -1190691925;
assign addr[29956]= -1158676398;
assign addr[29957]= -1126293375;
assign addr[29958]= -1093553126;
assign addr[29959]= -1060466036;
assign addr[29960]= -1027042599;
assign addr[29961]= -993293415;
assign addr[29962]= -959229189;
assign addr[29963]= -924860725;
assign addr[29964]= -890198924;
assign addr[29965]= -855254778;
assign addr[29966]= -820039373;
assign addr[29967]= -784563876;
assign addr[29968]= -748839539;
assign addr[29969]= -712877694;
assign addr[29970]= -676689746;
assign addr[29971]= -640287172;
assign addr[29972]= -603681519;
assign addr[29973]= -566884397;
assign addr[29974]= -529907477;
assign addr[29975]= -492762486;
assign addr[29976]= -455461206;
assign addr[29977]= -418015468;
assign addr[29978]= -380437148;
assign addr[29979]= -342738165;
assign addr[29980]= -304930476;
assign addr[29981]= -267026072;
assign addr[29982]= -229036977;
assign addr[29983]= -190975237;
assign addr[29984]= -152852926;
assign addr[29985]= -114682135;
assign addr[29986]= -76474970;
assign addr[29987]= -38243550;
assign addr[29988]= 0;
assign addr[29989]= 38243550;
assign addr[29990]= 76474970;
assign addr[29991]= 114682135;
assign addr[29992]= 152852926;
assign addr[29993]= 190975237;
assign addr[29994]= 229036977;
assign addr[29995]= 267026072;
assign addr[29996]= 304930476;
assign addr[29997]= 342738165;
assign addr[29998]= 380437148;
assign addr[29999]= 418015468;
assign addr[30000]= 455461206;
assign addr[30001]= 492762486;
assign addr[30002]= 529907477;
assign addr[30003]= 566884397;
assign addr[30004]= 603681519;
assign addr[30005]= 640287172;
assign addr[30006]= 676689746;
assign addr[30007]= 712877694;
assign addr[30008]= 748839539;
assign addr[30009]= 784563876;
assign addr[30010]= 820039373;
assign addr[30011]= 855254778;
assign addr[30012]= 890198924;
assign addr[30013]= 924860725;
assign addr[30014]= 959229189;
assign addr[30015]= 993293415;
assign addr[30016]= 1027042599;
assign addr[30017]= 1060466036;
assign addr[30018]= 1093553126;
assign addr[30019]= 1126293375;
assign addr[30020]= 1158676398;
assign addr[30021]= 1190691925;
assign addr[30022]= 1222329801;
assign addr[30023]= 1253579991;
assign addr[30024]= 1284432584;
assign addr[30025]= 1314877795;
assign addr[30026]= 1344905966;
assign addr[30027]= 1374507575;
assign addr[30028]= 1403673233;
assign addr[30029]= 1432393688;
assign addr[30030]= 1460659832;
assign addr[30031]= 1488462700;
assign addr[30032]= 1515793473;
assign addr[30033]= 1542643483;
assign addr[30034]= 1569004214;
assign addr[30035]= 1594867305;
assign addr[30036]= 1620224553;
assign addr[30037]= 1645067915;
assign addr[30038]= 1669389513;
assign addr[30039]= 1693181631;
assign addr[30040]= 1716436725;
assign addr[30041]= 1739147417;
assign addr[30042]= 1761306505;
assign addr[30043]= 1782906961;
assign addr[30044]= 1803941934;
assign addr[30045]= 1824404752;
assign addr[30046]= 1844288924;
assign addr[30047]= 1863588145;
assign addr[30048]= 1882296293;
assign addr[30049]= 1900407434;
assign addr[30050]= 1917915825;
assign addr[30051]= 1934815911;
assign addr[30052]= 1951102334;
assign addr[30053]= 1966769926;
assign addr[30054]= 1981813720;
assign addr[30055]= 1996228943;
assign addr[30056]= 2010011024;
assign addr[30057]= 2023155591;
assign addr[30058]= 2035658475;
assign addr[30059]= 2047515711;
assign addr[30060]= 2058723538;
assign addr[30061]= 2069278401;
assign addr[30062]= 2079176953;
assign addr[30063]= 2088416053;
assign addr[30064]= 2096992772;
assign addr[30065]= 2104904390;
assign addr[30066]= 2112148396;
assign addr[30067]= 2118722494;
assign addr[30068]= 2124624598;
assign addr[30069]= 2129852837;
assign addr[30070]= 2134405552;
assign addr[30071]= 2138281298;
assign addr[30072]= 2141478848;
assign addr[30073]= 2143997187;
assign addr[30074]= 2145835515;
assign addr[30075]= 2146993250;
assign addr[30076]= 2147470025;
assign addr[30077]= 2147265689;
assign addr[30078]= 2146380306;
assign addr[30079]= 2144814157;
assign addr[30080]= 2142567738;
assign addr[30081]= 2139641764;
assign addr[30082]= 2136037160;
assign addr[30083]= 2131755071;
assign addr[30084]= 2126796855;
assign addr[30085]= 2121164085;
assign addr[30086]= 2114858546;
assign addr[30087]= 2107882239;
assign addr[30088]= 2100237377;
assign addr[30089]= 2091926384;
assign addr[30090]= 2082951896;
assign addr[30091]= 2073316760;
assign addr[30092]= 2063024031;
assign addr[30093]= 2052076975;
assign addr[30094]= 2040479063;
assign addr[30095]= 2028233973;
assign addr[30096]= 2015345591;
assign addr[30097]= 2001818002;
assign addr[30098]= 1987655498;
assign addr[30099]= 1972862571;
assign addr[30100]= 1957443913;
assign addr[30101]= 1941404413;
assign addr[30102]= 1924749160;
assign addr[30103]= 1907483436;
assign addr[30104]= 1889612716;
assign addr[30105]= 1871142669;
assign addr[30106]= 1852079154;
assign addr[30107]= 1832428215;
assign addr[30108]= 1812196087;
assign addr[30109]= 1791389186;
assign addr[30110]= 1770014111;
assign addr[30111]= 1748077642;
assign addr[30112]= 1725586737;
assign addr[30113]= 1702548529;
assign addr[30114]= 1678970324;
assign addr[30115]= 1654859602;
assign addr[30116]= 1630224009;
assign addr[30117]= 1605071359;
assign addr[30118]= 1579409630;
assign addr[30119]= 1553246960;
assign addr[30120]= 1526591649;
assign addr[30121]= 1499452149;
assign addr[30122]= 1471837070;
assign addr[30123]= 1443755168;
assign addr[30124]= 1415215352;
assign addr[30125]= 1386226674;
assign addr[30126]= 1356798326;
assign addr[30127]= 1326939644;
assign addr[30128]= 1296660098;
assign addr[30129]= 1265969291;
assign addr[30130]= 1234876957;
assign addr[30131]= 1203392958;
assign addr[30132]= 1171527280;
assign addr[30133]= 1139290029;
assign addr[30134]= 1106691431;
assign addr[30135]= 1073741824;
assign addr[30136]= 1040451659;
assign addr[30137]= 1006831495;
assign addr[30138]= 972891995;
assign addr[30139]= 938643924;
assign addr[30140]= 904098143;
assign addr[30141]= 869265610;
assign addr[30142]= 834157373;
assign addr[30143]= 798784567;
assign addr[30144]= 763158411;
assign addr[30145]= 727290205;
assign addr[30146]= 691191324;
assign addr[30147]= 654873219;
assign addr[30148]= 618347408;
assign addr[30149]= 581625477;
assign addr[30150]= 544719071;
assign addr[30151]= 507639898;
assign addr[30152]= 470399716;
assign addr[30153]= 433010339;
assign addr[30154]= 395483624;
assign addr[30155]= 357831473;
assign addr[30156]= 320065829;
assign addr[30157]= 282198671;
assign addr[30158]= 244242007;
assign addr[30159]= 206207878;
assign addr[30160]= 168108346;
assign addr[30161]= 129955495;
assign addr[30162]= 91761426;
assign addr[30163]= 53538253;
assign addr[30164]= 15298099;
assign addr[30165]= -22946906;
assign addr[30166]= -61184634;
assign addr[30167]= -99402956;
assign addr[30168]= -137589750;
assign addr[30169]= -175732905;
assign addr[30170]= -213820322;
assign addr[30171]= -251839923;
assign addr[30172]= -289779648;
assign addr[30173]= -327627463;
assign addr[30174]= -365371365;
assign addr[30175]= -402999383;
assign addr[30176]= -440499581;
assign addr[30177]= -477860067;
assign addr[30178]= -515068990;
assign addr[30179]= -552114549;
assign addr[30180]= -588984994;
assign addr[30181]= -625668632;
assign addr[30182]= -662153826;
assign addr[30183]= -698429006;
assign addr[30184]= -734482665;
assign addr[30185]= -770303369;
assign addr[30186]= -805879757;
assign addr[30187]= -841200544;
assign addr[30188]= -876254528;
assign addr[30189]= -911030591;
assign addr[30190]= -945517704;
assign addr[30191]= -979704927;
assign addr[30192]= -1013581418;
assign addr[30193]= -1047136432;
assign addr[30194]= -1080359326;
assign addr[30195]= -1113239564;
assign addr[30196]= -1145766716;
assign addr[30197]= -1177930466;
assign addr[30198]= -1209720613;
assign addr[30199]= -1241127074;
assign addr[30200]= -1272139887;
assign addr[30201]= -1302749217;
assign addr[30202]= -1332945355;
assign addr[30203]= -1362718723;
assign addr[30204]= -1392059879;
assign addr[30205]= -1420959516;
assign addr[30206]= -1449408469;
assign addr[30207]= -1477397714;
assign addr[30208]= -1504918373;
assign addr[30209]= -1531961719;
assign addr[30210]= -1558519173;
assign addr[30211]= -1584582314;
assign addr[30212]= -1610142873;
assign addr[30213]= -1635192744;
assign addr[30214]= -1659723983;
assign addr[30215]= -1683728808;
assign addr[30216]= -1707199606;
assign addr[30217]= -1730128933;
assign addr[30218]= -1752509516;
assign addr[30219]= -1774334257;
assign addr[30220]= -1795596234;
assign addr[30221]= -1816288703;
assign addr[30222]= -1836405100;
assign addr[30223]= -1855939047;
assign addr[30224]= -1874884346;
assign addr[30225]= -1893234990;
assign addr[30226]= -1910985158;
assign addr[30227]= -1928129220;
assign addr[30228]= -1944661739;
assign addr[30229]= -1960577471;
assign addr[30230]= -1975871368;
assign addr[30231]= -1990538579;
assign addr[30232]= -2004574453;
assign addr[30233]= -2017974537;
assign addr[30234]= -2030734582;
assign addr[30235]= -2042850540;
assign addr[30236]= -2054318569;
assign addr[30237]= -2065135031;
assign addr[30238]= -2075296495;
assign addr[30239]= -2084799740;
assign addr[30240]= -2093641749;
assign addr[30241]= -2101819720;
assign addr[30242]= -2109331059;
assign addr[30243]= -2116173382;
assign addr[30244]= -2122344521;
assign addr[30245]= -2127842516;
assign addr[30246]= -2132665626;
assign addr[30247]= -2136812319;
assign addr[30248]= -2140281282;
assign addr[30249]= -2143071413;
assign addr[30250]= -2145181827;
assign addr[30251]= -2146611856;
assign addr[30252]= -2147361045;
assign addr[30253]= -2147429158;
assign addr[30254]= -2146816171;
assign addr[30255]= -2145522281;
assign addr[30256]= -2143547897;
assign addr[30257]= -2140893646;
assign addr[30258]= -2137560369;
assign addr[30259]= -2133549123;
assign addr[30260]= -2128861181;
assign addr[30261]= -2123498030;
assign addr[30262]= -2117461370;
assign addr[30263]= -2110753117;
assign addr[30264]= -2103375398;
assign addr[30265]= -2095330553;
assign addr[30266]= -2086621133;
assign addr[30267]= -2077249901;
assign addr[30268]= -2067219829;
assign addr[30269]= -2056534099;
assign addr[30270]= -2045196100;
assign addr[30271]= -2033209426;
assign addr[30272]= -2020577882;
assign addr[30273]= -2007305472;
assign addr[30274]= -1993396407;
assign addr[30275]= -1978855097;
assign addr[30276]= -1963686155;
assign addr[30277]= -1947894393;
assign addr[30278]= -1931484818;
assign addr[30279]= -1914462636;
assign addr[30280]= -1896833245;
assign addr[30281]= -1878602237;
assign addr[30282]= -1859775393;
assign addr[30283]= -1840358687;
assign addr[30284]= -1820358275;
assign addr[30285]= -1799780501;
assign addr[30286]= -1778631892;
assign addr[30287]= -1756919156;
assign addr[30288]= -1734649179;
assign addr[30289]= -1711829025;
assign addr[30290]= -1688465931;
assign addr[30291]= -1664567307;
assign addr[30292]= -1640140734;
assign addr[30293]= -1615193959;
assign addr[30294]= -1589734894;
assign addr[30295]= -1563771613;
assign addr[30296]= -1537312353;
assign addr[30297]= -1510365504;
assign addr[30298]= -1482939614;
assign addr[30299]= -1455043381;
assign addr[30300]= -1426685652;
assign addr[30301]= -1397875423;
assign addr[30302]= -1368621831;
assign addr[30303]= -1338934154;
assign addr[30304]= -1308821808;
assign addr[30305]= -1278294345;
assign addr[30306]= -1247361445;
assign addr[30307]= -1216032921;
assign addr[30308]= -1184318708;
assign addr[30309]= -1152228866;
assign addr[30310]= -1119773573;
assign addr[30311]= -1086963121;
assign addr[30312]= -1053807919;
assign addr[30313]= -1020318481;
assign addr[30314]= -986505429;
assign addr[30315]= -952379488;
assign addr[30316]= -917951481;
assign addr[30317]= -883232329;
assign addr[30318]= -848233042;
assign addr[30319]= -812964722;
assign addr[30320]= -777438554;
assign addr[30321]= -741665807;
assign addr[30322]= -705657826;
assign addr[30323]= -669426032;
assign addr[30324]= -632981917;
assign addr[30325]= -596337040;
assign addr[30326]= -559503022;
assign addr[30327]= -522491548;
assign addr[30328]= -485314355;
assign addr[30329]= -447983235;
assign addr[30330]= -410510029;
assign addr[30331]= -372906622;
assign addr[30332]= -335184940;
assign addr[30333]= -297356948;
assign addr[30334]= -259434643;
assign addr[30335]= -221430054;
assign addr[30336]= -183355234;
assign addr[30337]= -145222259;
assign addr[30338]= -107043224;
assign addr[30339]= -68830239;
assign addr[30340]= -30595422;
assign addr[30341]= 7649098;
assign addr[30342]= 45891193;
assign addr[30343]= 84118732;
assign addr[30344]= 122319591;
assign addr[30345]= 160481654;
assign addr[30346]= 198592817;
assign addr[30347]= 236640993;
assign addr[30348]= 274614114;
assign addr[30349]= 312500135;
assign addr[30350]= 350287041;
assign addr[30351]= 387962847;
assign addr[30352]= 425515602;
assign addr[30353]= 462933398;
assign addr[30354]= 500204365;
assign addr[30355]= 537316682;
assign addr[30356]= 574258580;
assign addr[30357]= 611018340;
assign addr[30358]= 647584304;
assign addr[30359]= 683944874;
assign addr[30360]= 720088517;
assign addr[30361]= 756003771;
assign addr[30362]= 791679244;
assign addr[30363]= 827103620;
assign addr[30364]= 862265664;
assign addr[30365]= 897154224;
assign addr[30366]= 931758235;
assign addr[30367]= 966066720;
assign addr[30368]= 1000068799;
assign addr[30369]= 1033753687;
assign addr[30370]= 1067110699;
assign addr[30371]= 1100129257;
assign addr[30372]= 1132798888;
assign addr[30373]= 1165109230;
assign addr[30374]= 1197050035;
assign addr[30375]= 1228611172;
assign addr[30376]= 1259782632;
assign addr[30377]= 1290554528;
assign addr[30378]= 1320917099;
assign addr[30379]= 1350860716;
assign addr[30380]= 1380375881;
assign addr[30381]= 1409453233;
assign addr[30382]= 1438083551;
assign addr[30383]= 1466257752;
assign addr[30384]= 1493966902;
assign addr[30385]= 1521202211;
assign addr[30386]= 1547955041;
assign addr[30387]= 1574216908;
assign addr[30388]= 1599979481;
assign addr[30389]= 1625234591;
assign addr[30390]= 1649974225;
assign addr[30391]= 1674190539;
assign addr[30392]= 1697875851;
assign addr[30393]= 1721022648;
assign addr[30394]= 1743623590;
assign addr[30395]= 1765671509;
assign addr[30396]= 1787159411;
assign addr[30397]= 1808080480;
assign addr[30398]= 1828428082;
assign addr[30399]= 1848195763;
assign addr[30400]= 1867377253;
assign addr[30401]= 1885966468;
assign addr[30402]= 1903957513;
assign addr[30403]= 1921344681;
assign addr[30404]= 1938122457;
assign addr[30405]= 1954285520;
assign addr[30406]= 1969828744;
assign addr[30407]= 1984747199;
assign addr[30408]= 1999036154;
assign addr[30409]= 2012691075;
assign addr[30410]= 2025707632;
assign addr[30411]= 2038081698;
assign addr[30412]= 2049809346;
assign addr[30413]= 2060886858;
assign addr[30414]= 2071310720;
assign addr[30415]= 2081077626;
assign addr[30416]= 2090184478;
assign addr[30417]= 2098628387;
assign addr[30418]= 2106406677;
assign addr[30419]= 2113516878;
assign addr[30420]= 2119956737;
assign addr[30421]= 2125724211;
assign addr[30422]= 2130817471;
assign addr[30423]= 2135234901;
assign addr[30424]= 2138975100;
assign addr[30425]= 2142036881;
assign addr[30426]= 2144419275;
assign addr[30427]= 2146121524;
assign addr[30428]= 2147143090;
assign addr[30429]= 2147483648;
assign addr[30430]= 2147143090;
assign addr[30431]= 2146121524;
assign addr[30432]= 2144419275;
assign addr[30433]= 2142036881;
assign addr[30434]= 2138975100;
assign addr[30435]= 2135234901;
assign addr[30436]= 2130817471;
assign addr[30437]= 2125724211;
assign addr[30438]= 2119956737;
assign addr[30439]= 2113516878;
assign addr[30440]= 2106406677;
assign addr[30441]= 2098628387;
assign addr[30442]= 2090184478;
assign addr[30443]= 2081077626;
assign addr[30444]= 2071310720;
assign addr[30445]= 2060886858;
assign addr[30446]= 2049809346;
assign addr[30447]= 2038081698;
assign addr[30448]= 2025707632;
assign addr[30449]= 2012691075;
assign addr[30450]= 1999036154;
assign addr[30451]= 1984747199;
assign addr[30452]= 1969828744;
assign addr[30453]= 1954285520;
assign addr[30454]= 1938122457;
assign addr[30455]= 1921344681;
assign addr[30456]= 1903957513;
assign addr[30457]= 1885966468;
assign addr[30458]= 1867377253;
assign addr[30459]= 1848195763;
assign addr[30460]= 1828428082;
assign addr[30461]= 1808080480;
assign addr[30462]= 1787159411;
assign addr[30463]= 1765671509;
assign addr[30464]= 1743623590;
assign addr[30465]= 1721022648;
assign addr[30466]= 1697875851;
assign addr[30467]= 1674190539;
assign addr[30468]= 1649974225;
assign addr[30469]= 1625234591;
assign addr[30470]= 1599979481;
assign addr[30471]= 1574216908;
assign addr[30472]= 1547955041;
assign addr[30473]= 1521202211;
assign addr[30474]= 1493966902;
assign addr[30475]= 1466257752;
assign addr[30476]= 1438083551;
assign addr[30477]= 1409453233;
assign addr[30478]= 1380375881;
assign addr[30479]= 1350860716;
assign addr[30480]= 1320917099;
assign addr[30481]= 1290554528;
assign addr[30482]= 1259782632;
assign addr[30483]= 1228611172;
assign addr[30484]= 1197050035;
assign addr[30485]= 1165109230;
assign addr[30486]= 1132798888;
assign addr[30487]= 1100129257;
assign addr[30488]= 1067110699;
assign addr[30489]= 1033753687;
assign addr[30490]= 1000068799;
assign addr[30491]= 966066720;
assign addr[30492]= 931758235;
assign addr[30493]= 897154224;
assign addr[30494]= 862265664;
assign addr[30495]= 827103620;
assign addr[30496]= 791679244;
assign addr[30497]= 756003771;
assign addr[30498]= 720088517;
assign addr[30499]= 683944874;
assign addr[30500]= 647584304;
assign addr[30501]= 611018340;
assign addr[30502]= 574258580;
assign addr[30503]= 537316682;
assign addr[30504]= 500204365;
assign addr[30505]= 462933398;
assign addr[30506]= 425515602;
assign addr[30507]= 387962847;
assign addr[30508]= 350287041;
assign addr[30509]= 312500135;
assign addr[30510]= 274614114;
assign addr[30511]= 236640993;
assign addr[30512]= 198592817;
assign addr[30513]= 160481654;
assign addr[30514]= 122319591;
assign addr[30515]= 84118732;
assign addr[30516]= 45891193;
assign addr[30517]= 7649098;
assign addr[30518]= -30595422;
assign addr[30519]= -68830239;
assign addr[30520]= -107043224;
assign addr[30521]= -145222259;
assign addr[30522]= -183355234;
assign addr[30523]= -221430054;
assign addr[30524]= -259434643;
assign addr[30525]= -297356948;
assign addr[30526]= -335184940;
assign addr[30527]= -372906622;
assign addr[30528]= -410510029;
assign addr[30529]= -447983235;
assign addr[30530]= -485314355;
assign addr[30531]= -522491548;
assign addr[30532]= -559503022;
assign addr[30533]= -596337040;
assign addr[30534]= -632981917;
assign addr[30535]= -669426032;
assign addr[30536]= -705657826;
assign addr[30537]= -741665807;
assign addr[30538]= -777438554;
assign addr[30539]= -812964722;
assign addr[30540]= -848233042;
assign addr[30541]= -883232329;
assign addr[30542]= -917951481;
assign addr[30543]= -952379488;
assign addr[30544]= -986505429;
assign addr[30545]= -1020318481;
assign addr[30546]= -1053807919;
assign addr[30547]= -1086963121;
assign addr[30548]= -1119773573;
assign addr[30549]= -1152228866;
assign addr[30550]= -1184318708;
assign addr[30551]= -1216032921;
assign addr[30552]= -1247361445;
assign addr[30553]= -1278294345;
assign addr[30554]= -1308821808;
assign addr[30555]= -1338934154;
assign addr[30556]= -1368621831;
assign addr[30557]= -1397875423;
assign addr[30558]= -1426685652;
assign addr[30559]= -1455043381;
assign addr[30560]= -1482939614;
assign addr[30561]= -1510365504;
assign addr[30562]= -1537312353;
assign addr[30563]= -1563771613;
assign addr[30564]= -1589734894;
assign addr[30565]= -1615193959;
assign addr[30566]= -1640140734;
assign addr[30567]= -1664567307;
assign addr[30568]= -1688465931;
assign addr[30569]= -1711829025;
assign addr[30570]= -1734649179;
assign addr[30571]= -1756919156;
assign addr[30572]= -1778631892;
assign addr[30573]= -1799780501;
assign addr[30574]= -1820358275;
assign addr[30575]= -1840358687;
assign addr[30576]= -1859775393;
assign addr[30577]= -1878602237;
assign addr[30578]= -1896833245;
assign addr[30579]= -1914462636;
assign addr[30580]= -1931484818;
assign addr[30581]= -1947894393;
assign addr[30582]= -1963686155;
assign addr[30583]= -1978855097;
assign addr[30584]= -1993396407;
assign addr[30585]= -2007305472;
assign addr[30586]= -2020577882;
assign addr[30587]= -2033209426;
assign addr[30588]= -2045196100;
assign addr[30589]= -2056534099;
assign addr[30590]= -2067219829;
assign addr[30591]= -2077249901;
assign addr[30592]= -2086621133;
assign addr[30593]= -2095330553;
assign addr[30594]= -2103375398;
assign addr[30595]= -2110753117;
assign addr[30596]= -2117461370;
assign addr[30597]= -2123498030;
assign addr[30598]= -2128861181;
assign addr[30599]= -2133549123;
assign addr[30600]= -2137560369;
assign addr[30601]= -2140893646;
assign addr[30602]= -2143547897;
assign addr[30603]= -2145522281;
assign addr[30604]= -2146816171;
assign addr[30605]= -2147429158;
assign addr[30606]= -2147361045;
assign addr[30607]= -2146611856;
assign addr[30608]= -2145181827;
assign addr[30609]= -2143071413;
assign addr[30610]= -2140281282;
assign addr[30611]= -2136812319;
assign addr[30612]= -2132665626;
assign addr[30613]= -2127842516;
assign addr[30614]= -2122344521;
assign addr[30615]= -2116173382;
assign addr[30616]= -2109331059;
assign addr[30617]= -2101819720;
assign addr[30618]= -2093641749;
assign addr[30619]= -2084799740;
assign addr[30620]= -2075296495;
assign addr[30621]= -2065135031;
assign addr[30622]= -2054318569;
assign addr[30623]= -2042850540;
assign addr[30624]= -2030734582;
assign addr[30625]= -2017974537;
assign addr[30626]= -2004574453;
assign addr[30627]= -1990538579;
assign addr[30628]= -1975871368;
assign addr[30629]= -1960577471;
assign addr[30630]= -1944661739;
assign addr[30631]= -1928129220;
assign addr[30632]= -1910985158;
assign addr[30633]= -1893234990;
assign addr[30634]= -1874884346;
assign addr[30635]= -1855939047;
assign addr[30636]= -1836405100;
assign addr[30637]= -1816288703;
assign addr[30638]= -1795596234;
assign addr[30639]= -1774334257;
assign addr[30640]= -1752509516;
assign addr[30641]= -1730128933;
assign addr[30642]= -1707199606;
assign addr[30643]= -1683728808;
assign addr[30644]= -1659723983;
assign addr[30645]= -1635192744;
assign addr[30646]= -1610142873;
assign addr[30647]= -1584582314;
assign addr[30648]= -1558519173;
assign addr[30649]= -1531961719;
assign addr[30650]= -1504918373;
assign addr[30651]= -1477397714;
assign addr[30652]= -1449408469;
assign addr[30653]= -1420959516;
assign addr[30654]= -1392059879;
assign addr[30655]= -1362718723;
assign addr[30656]= -1332945355;
assign addr[30657]= -1302749217;
assign addr[30658]= -1272139887;
assign addr[30659]= -1241127074;
assign addr[30660]= -1209720613;
assign addr[30661]= -1177930466;
assign addr[30662]= -1145766716;
assign addr[30663]= -1113239564;
assign addr[30664]= -1080359326;
assign addr[30665]= -1047136432;
assign addr[30666]= -1013581418;
assign addr[30667]= -979704927;
assign addr[30668]= -945517704;
assign addr[30669]= -911030591;
assign addr[30670]= -876254528;
assign addr[30671]= -841200544;
assign addr[30672]= -805879757;
assign addr[30673]= -770303369;
assign addr[30674]= -734482665;
assign addr[30675]= -698429006;
assign addr[30676]= -662153826;
assign addr[30677]= -625668632;
assign addr[30678]= -588984994;
assign addr[30679]= -552114549;
assign addr[30680]= -515068990;
assign addr[30681]= -477860067;
assign addr[30682]= -440499581;
assign addr[30683]= -402999383;
assign addr[30684]= -365371365;
assign addr[30685]= -327627463;
assign addr[30686]= -289779648;
assign addr[30687]= -251839923;
assign addr[30688]= -213820322;
assign addr[30689]= -175732905;
assign addr[30690]= -137589750;
assign addr[30691]= -99402956;
assign addr[30692]= -61184634;
assign addr[30693]= -22946906;
assign addr[30694]= 15298099;
assign addr[30695]= 53538253;
assign addr[30696]= 91761426;
assign addr[30697]= 129955495;
assign addr[30698]= 168108346;
assign addr[30699]= 206207878;
assign addr[30700]= 244242007;
assign addr[30701]= 282198671;
assign addr[30702]= 320065829;
assign addr[30703]= 357831473;
assign addr[30704]= 395483624;
assign addr[30705]= 433010339;
assign addr[30706]= 470399716;
assign addr[30707]= 507639898;
assign addr[30708]= 544719071;
assign addr[30709]= 581625477;
assign addr[30710]= 618347408;
assign addr[30711]= 654873219;
assign addr[30712]= 691191324;
assign addr[30713]= 727290205;
assign addr[30714]= 763158411;
assign addr[30715]= 798784567;
assign addr[30716]= 834157373;
assign addr[30717]= 869265610;
assign addr[30718]= 904098143;
assign addr[30719]= 938643924;
assign addr[30720]= 972891995;
assign addr[30721]= 1006831495;
assign addr[30722]= 1040451659;
assign addr[30723]= 1073741824;
assign addr[30724]= 1106691431;
assign addr[30725]= 1139290029;
assign addr[30726]= 1171527280;
assign addr[30727]= 1203392958;
assign addr[30728]= 1234876957;
assign addr[30729]= 1265969291;
assign addr[30730]= 1296660098;
assign addr[30731]= 1326939644;
assign addr[30732]= 1356798326;
assign addr[30733]= 1386226674;
assign addr[30734]= 1415215352;
assign addr[30735]= 1443755168;
assign addr[30736]= 1471837070;
assign addr[30737]= 1499452149;
assign addr[30738]= 1526591649;
assign addr[30739]= 1553246960;
assign addr[30740]= 1579409630;
assign addr[30741]= 1605071359;
assign addr[30742]= 1630224009;
assign addr[30743]= 1654859602;
assign addr[30744]= 1678970324;
assign addr[30745]= 1702548529;
assign addr[30746]= 1725586737;
assign addr[30747]= 1748077642;
assign addr[30748]= 1770014111;
assign addr[30749]= 1791389186;
assign addr[30750]= 1812196087;
assign addr[30751]= 1832428215;
assign addr[30752]= 1852079154;
assign addr[30753]= 1871142669;
assign addr[30754]= 1889612716;
assign addr[30755]= 1907483436;
assign addr[30756]= 1924749160;
assign addr[30757]= 1941404413;
assign addr[30758]= 1957443913;
assign addr[30759]= 1972862571;
assign addr[30760]= 1987655498;
assign addr[30761]= 2001818002;
assign addr[30762]= 2015345591;
assign addr[30763]= 2028233973;
assign addr[30764]= 2040479063;
assign addr[30765]= 2052076975;
assign addr[30766]= 2063024031;
assign addr[30767]= 2073316760;
assign addr[30768]= 2082951896;
assign addr[30769]= 2091926384;
assign addr[30770]= 2100237377;
assign addr[30771]= 2107882239;
assign addr[30772]= 2114858546;
assign addr[30773]= 2121164085;
assign addr[30774]= 2126796855;
assign addr[30775]= 2131755071;
assign addr[30776]= 2136037160;
assign addr[30777]= 2139641764;
assign addr[30778]= 2142567738;
assign addr[30779]= 2144814157;
assign addr[30780]= 2146380306;
assign addr[30781]= 2147265689;
assign addr[30782]= 2147470025;
assign addr[30783]= 2146993250;
assign addr[30784]= 2145835515;
assign addr[30785]= 2143997187;
assign addr[30786]= 2141478848;
assign addr[30787]= 2138281298;
assign addr[30788]= 2134405552;
assign addr[30789]= 2129852837;
assign addr[30790]= 2124624598;
assign addr[30791]= 2118722494;
assign addr[30792]= 2112148396;
assign addr[30793]= 2104904390;
assign addr[30794]= 2096992772;
assign addr[30795]= 2088416053;
assign addr[30796]= 2079176953;
assign addr[30797]= 2069278401;
assign addr[30798]= 2058723538;
assign addr[30799]= 2047515711;
assign addr[30800]= 2035658475;
assign addr[30801]= 2023155591;
assign addr[30802]= 2010011024;
assign addr[30803]= 1996228943;
assign addr[30804]= 1981813720;
assign addr[30805]= 1966769926;
assign addr[30806]= 1951102334;
assign addr[30807]= 1934815911;
assign addr[30808]= 1917915825;
assign addr[30809]= 1900407434;
assign addr[30810]= 1882296293;
assign addr[30811]= 1863588145;
assign addr[30812]= 1844288924;
assign addr[30813]= 1824404752;
assign addr[30814]= 1803941934;
assign addr[30815]= 1782906961;
assign addr[30816]= 1761306505;
assign addr[30817]= 1739147417;
assign addr[30818]= 1716436725;
assign addr[30819]= 1693181631;
assign addr[30820]= 1669389513;
assign addr[30821]= 1645067915;
assign addr[30822]= 1620224553;
assign addr[30823]= 1594867305;
assign addr[30824]= 1569004214;
assign addr[30825]= 1542643483;
assign addr[30826]= 1515793473;
assign addr[30827]= 1488462700;
assign addr[30828]= 1460659832;
assign addr[30829]= 1432393688;
assign addr[30830]= 1403673233;
assign addr[30831]= 1374507575;
assign addr[30832]= 1344905966;
assign addr[30833]= 1314877795;
assign addr[30834]= 1284432584;
assign addr[30835]= 1253579991;
assign addr[30836]= 1222329801;
assign addr[30837]= 1190691925;
assign addr[30838]= 1158676398;
assign addr[30839]= 1126293375;
assign addr[30840]= 1093553126;
assign addr[30841]= 1060466036;
assign addr[30842]= 1027042599;
assign addr[30843]= 993293415;
assign addr[30844]= 959229189;
assign addr[30845]= 924860725;
assign addr[30846]= 890198924;
assign addr[30847]= 855254778;
assign addr[30848]= 820039373;
assign addr[30849]= 784563876;
assign addr[30850]= 748839539;
assign addr[30851]= 712877694;
assign addr[30852]= 676689746;
assign addr[30853]= 640287172;
assign addr[30854]= 603681519;
assign addr[30855]= 566884397;
assign addr[30856]= 529907477;
assign addr[30857]= 492762486;
assign addr[30858]= 455461206;
assign addr[30859]= 418015468;
assign addr[30860]= 380437148;
assign addr[30861]= 342738165;
assign addr[30862]= 304930476;
assign addr[30863]= 267026072;
assign addr[30864]= 229036977;
assign addr[30865]= 190975237;
assign addr[30866]= 152852926;
assign addr[30867]= 114682135;
assign addr[30868]= 76474970;
assign addr[30869]= 38243550;
assign addr[30870]= 0;
assign addr[30871]= -38243550;
assign addr[30872]= -76474970;
assign addr[30873]= -114682135;
assign addr[30874]= -152852926;
assign addr[30875]= -190975237;
assign addr[30876]= -229036977;
assign addr[30877]= -267026072;
assign addr[30878]= -304930476;
assign addr[30879]= -342738165;
assign addr[30880]= -380437148;
assign addr[30881]= -418015468;
assign addr[30882]= -455461206;
assign addr[30883]= -492762486;
assign addr[30884]= -529907477;
assign addr[30885]= -566884397;
assign addr[30886]= -603681519;
assign addr[30887]= -640287172;
assign addr[30888]= -676689746;
assign addr[30889]= -712877694;
assign addr[30890]= -748839539;
assign addr[30891]= -784563876;
assign addr[30892]= -820039373;
assign addr[30893]= -855254778;
assign addr[30894]= -890198924;
assign addr[30895]= -924860725;
assign addr[30896]= -959229189;
assign addr[30897]= -993293415;
assign addr[30898]= -1027042599;
assign addr[30899]= -1060466036;
assign addr[30900]= -1093553126;
assign addr[30901]= -1126293375;
assign addr[30902]= -1158676398;
assign addr[30903]= -1190691925;
assign addr[30904]= -1222329801;
assign addr[30905]= -1253579991;
assign addr[30906]= -1284432584;
assign addr[30907]= -1314877795;
assign addr[30908]= -1344905966;
assign addr[30909]= -1374507575;
assign addr[30910]= -1403673233;
assign addr[30911]= -1432393688;
assign addr[30912]= -1460659832;
assign addr[30913]= -1488462700;
assign addr[30914]= -1515793473;
assign addr[30915]= -1542643483;
assign addr[30916]= -1569004214;
assign addr[30917]= -1594867305;
assign addr[30918]= -1620224553;
assign addr[30919]= -1645067915;
assign addr[30920]= -1669389513;
assign addr[30921]= -1693181631;
assign addr[30922]= -1716436725;
assign addr[30923]= -1739147417;
assign addr[30924]= -1761306505;
assign addr[30925]= -1782906961;
assign addr[30926]= -1803941934;
assign addr[30927]= -1824404752;
assign addr[30928]= -1844288924;
assign addr[30929]= -1863588145;
assign addr[30930]= -1882296293;
assign addr[30931]= -1900407434;
assign addr[30932]= -1917915825;
assign addr[30933]= -1934815911;
assign addr[30934]= -1951102334;
assign addr[30935]= -1966769926;
assign addr[30936]= -1981813720;
assign addr[30937]= -1996228943;
assign addr[30938]= -2010011024;
assign addr[30939]= -2023155591;
assign addr[30940]= -2035658475;
assign addr[30941]= -2047515711;
assign addr[30942]= -2058723538;
assign addr[30943]= -2069278401;
assign addr[30944]= -2079176953;
assign addr[30945]= -2088416053;
assign addr[30946]= -2096992772;
assign addr[30947]= -2104904390;
assign addr[30948]= -2112148396;
assign addr[30949]= -2118722494;
assign addr[30950]= -2124624598;
assign addr[30951]= -2129852837;
assign addr[30952]= -2134405552;
assign addr[30953]= -2138281298;
assign addr[30954]= -2141478848;
assign addr[30955]= -2143997187;
assign addr[30956]= -2145835515;
assign addr[30957]= -2146993250;
assign addr[30958]= -2147470025;
assign addr[30959]= -2147265689;
assign addr[30960]= -2146380306;
assign addr[30961]= -2144814157;
assign addr[30962]= -2142567738;
assign addr[30963]= -2139641764;
assign addr[30964]= -2136037160;
assign addr[30965]= -2131755071;
assign addr[30966]= -2126796855;
assign addr[30967]= -2121164085;
assign addr[30968]= -2114858546;
assign addr[30969]= -2107882239;
assign addr[30970]= -2100237377;
assign addr[30971]= -2091926384;
assign addr[30972]= -2082951896;
assign addr[30973]= -2073316760;
assign addr[30974]= -2063024031;
assign addr[30975]= -2052076975;
assign addr[30976]= -2040479063;
assign addr[30977]= -2028233973;
assign addr[30978]= -2015345591;
assign addr[30979]= -2001818002;
assign addr[30980]= -1987655498;
assign addr[30981]= -1972862571;
assign addr[30982]= -1957443913;
assign addr[30983]= -1941404413;
assign addr[30984]= -1924749160;
assign addr[30985]= -1907483436;
assign addr[30986]= -1889612716;
assign addr[30987]= -1871142669;
assign addr[30988]= -1852079154;
assign addr[30989]= -1832428215;
assign addr[30990]= -1812196087;
assign addr[30991]= -1791389186;
assign addr[30992]= -1770014111;
assign addr[30993]= -1748077642;
assign addr[30994]= -1725586737;
assign addr[30995]= -1702548529;
assign addr[30996]= -1678970324;
assign addr[30997]= -1654859602;
assign addr[30998]= -1630224009;
assign addr[30999]= -1605071359;
assign addr[31000]= -1579409630;
assign addr[31001]= -1553246960;
assign addr[31002]= -1526591649;
assign addr[31003]= -1499452149;
assign addr[31004]= -1471837070;
assign addr[31005]= -1443755168;
assign addr[31006]= -1415215352;
assign addr[31007]= -1386226674;
assign addr[31008]= -1356798326;
assign addr[31009]= -1326939644;
assign addr[31010]= -1296660098;
assign addr[31011]= -1265969291;
assign addr[31012]= -1234876957;
assign addr[31013]= -1203392958;
assign addr[31014]= -1171527280;
assign addr[31015]= -1139290029;
assign addr[31016]= -1106691431;
assign addr[31017]= -1073741824;
assign addr[31018]= -1040451659;
assign addr[31019]= -1006831495;
assign addr[31020]= -972891995;
assign addr[31021]= -938643924;
assign addr[31022]= -904098143;
assign addr[31023]= -869265610;
assign addr[31024]= -834157373;
assign addr[31025]= -798784567;
assign addr[31026]= -763158411;
assign addr[31027]= -727290205;
assign addr[31028]= -691191324;
assign addr[31029]= -654873219;
assign addr[31030]= -618347408;
assign addr[31031]= -581625477;
assign addr[31032]= -544719071;
assign addr[31033]= -507639898;
assign addr[31034]= -470399716;
assign addr[31035]= -433010339;
assign addr[31036]= -395483624;
assign addr[31037]= -357831473;
assign addr[31038]= -320065829;
assign addr[31039]= -282198671;
assign addr[31040]= -244242007;
assign addr[31041]= -206207878;
assign addr[31042]= -168108346;
assign addr[31043]= -129955495;
assign addr[31044]= -91761426;
assign addr[31045]= -53538253;
assign addr[31046]= -15298099;
assign addr[31047]= 22946906;
assign addr[31048]= 61184634;
assign addr[31049]= 99402956;
assign addr[31050]= 137589750;
assign addr[31051]= 175732905;
assign addr[31052]= 213820322;
assign addr[31053]= 251839923;
assign addr[31054]= 289779648;
assign addr[31055]= 327627463;
assign addr[31056]= 365371365;
assign addr[31057]= 402999383;
assign addr[31058]= 440499581;
assign addr[31059]= 477860067;
assign addr[31060]= 515068990;
assign addr[31061]= 552114549;
assign addr[31062]= 588984994;
assign addr[31063]= 625668632;
assign addr[31064]= 662153826;
assign addr[31065]= 698429006;
assign addr[31066]= 734482665;
assign addr[31067]= 770303369;
assign addr[31068]= 805879757;
assign addr[31069]= 841200544;
assign addr[31070]= 876254528;
assign addr[31071]= 911030591;
assign addr[31072]= 945517704;
assign addr[31073]= 979704927;
assign addr[31074]= 1013581418;
assign addr[31075]= 1047136432;
assign addr[31076]= 1080359326;
assign addr[31077]= 1113239564;
assign addr[31078]= 1145766716;
assign addr[31079]= 1177930466;
assign addr[31080]= 1209720613;
assign addr[31081]= 1241127074;
assign addr[31082]= 1272139887;
assign addr[31083]= 1302749217;
assign addr[31084]= 1332945355;
assign addr[31085]= 1362718723;
assign addr[31086]= 1392059879;
assign addr[31087]= 1420959516;
assign addr[31088]= 1449408469;
assign addr[31089]= 1477397714;
assign addr[31090]= 1504918373;
assign addr[31091]= 1531961719;
assign addr[31092]= 1558519173;
assign addr[31093]= 1584582314;
assign addr[31094]= 1610142873;
assign addr[31095]= 1635192744;
assign addr[31096]= 1659723983;
assign addr[31097]= 1683728808;
assign addr[31098]= 1707199606;
assign addr[31099]= 1730128933;
assign addr[31100]= 1752509516;
assign addr[31101]= 1774334257;
assign addr[31102]= 1795596234;
assign addr[31103]= 1816288703;
assign addr[31104]= 1836405100;
assign addr[31105]= 1855939047;
assign addr[31106]= 1874884346;
assign addr[31107]= 1893234990;
assign addr[31108]= 1910985158;
assign addr[31109]= 1928129220;
assign addr[31110]= 1944661739;
assign addr[31111]= 1960577471;
assign addr[31112]= 1975871368;
assign addr[31113]= 1990538579;
assign addr[31114]= 2004574453;
assign addr[31115]= 2017974537;
assign addr[31116]= 2030734582;
assign addr[31117]= 2042850540;
assign addr[31118]= 2054318569;
assign addr[31119]= 2065135031;
assign addr[31120]= 2075296495;
assign addr[31121]= 2084799740;
assign addr[31122]= 2093641749;
assign addr[31123]= 2101819720;
assign addr[31124]= 2109331059;
assign addr[31125]= 2116173382;
assign addr[31126]= 2122344521;
assign addr[31127]= 2127842516;
assign addr[31128]= 2132665626;
assign addr[31129]= 2136812319;
assign addr[31130]= 2140281282;
assign addr[31131]= 2143071413;
assign addr[31132]= 2145181827;
assign addr[31133]= 2146611856;
assign addr[31134]= 2147361045;
assign addr[31135]= 2147429158;
assign addr[31136]= 2146816171;
assign addr[31137]= 2145522281;
assign addr[31138]= 2143547897;
assign addr[31139]= 2140893646;
assign addr[31140]= 2137560369;
assign addr[31141]= 2133549123;
assign addr[31142]= 2128861181;
assign addr[31143]= 2123498030;
assign addr[31144]= 2117461370;
assign addr[31145]= 2110753117;
assign addr[31146]= 2103375398;
assign addr[31147]= 2095330553;
assign addr[31148]= 2086621133;
assign addr[31149]= 2077249901;
assign addr[31150]= 2067219829;
assign addr[31151]= 2056534099;
assign addr[31152]= 2045196100;
assign addr[31153]= 2033209426;
assign addr[31154]= 2020577882;
assign addr[31155]= 2007305472;
assign addr[31156]= 1993396407;
assign addr[31157]= 1978855097;
assign addr[31158]= 1963686155;
assign addr[31159]= 1947894393;
assign addr[31160]= 1931484818;
assign addr[31161]= 1914462636;
assign addr[31162]= 1896833245;
assign addr[31163]= 1878602237;
assign addr[31164]= 1859775393;
assign addr[31165]= 1840358687;
assign addr[31166]= 1820358275;
assign addr[31167]= 1799780501;
assign addr[31168]= 1778631892;
assign addr[31169]= 1756919156;
assign addr[31170]= 1734649179;
assign addr[31171]= 1711829025;
assign addr[31172]= 1688465931;
assign addr[31173]= 1664567307;
assign addr[31174]= 1640140734;
assign addr[31175]= 1615193959;
assign addr[31176]= 1589734894;
assign addr[31177]= 1563771613;
assign addr[31178]= 1537312353;
assign addr[31179]= 1510365504;
assign addr[31180]= 1482939614;
assign addr[31181]= 1455043381;
assign addr[31182]= 1426685652;
assign addr[31183]= 1397875423;
assign addr[31184]= 1368621831;
assign addr[31185]= 1338934154;
assign addr[31186]= 1308821808;
assign addr[31187]= 1278294345;
assign addr[31188]= 1247361445;
assign addr[31189]= 1216032921;
assign addr[31190]= 1184318708;
assign addr[31191]= 1152228866;
assign addr[31192]= 1119773573;
assign addr[31193]= 1086963121;
assign addr[31194]= 1053807919;
assign addr[31195]= 1020318481;
assign addr[31196]= 986505429;
assign addr[31197]= 952379488;
assign addr[31198]= 917951481;
assign addr[31199]= 883232329;
assign addr[31200]= 848233042;
assign addr[31201]= 812964722;
assign addr[31202]= 777438554;
assign addr[31203]= 741665807;
assign addr[31204]= 705657826;
assign addr[31205]= 669426032;
assign addr[31206]= 632981917;
assign addr[31207]= 596337040;
assign addr[31208]= 559503022;
assign addr[31209]= 522491548;
assign addr[31210]= 485314355;
assign addr[31211]= 447983235;
assign addr[31212]= 410510029;
assign addr[31213]= 372906622;
assign addr[31214]= 335184940;
assign addr[31215]= 297356948;
assign addr[31216]= 259434643;
assign addr[31217]= 221430054;
assign addr[31218]= 183355234;
assign addr[31219]= 145222259;
assign addr[31220]= 107043224;
assign addr[31221]= 68830239;
assign addr[31222]= 30595422;
assign addr[31223]= -7649098;
assign addr[31224]= -45891193;
assign addr[31225]= -84118732;
assign addr[31226]= -122319591;
assign addr[31227]= -160481654;
assign addr[31228]= -198592817;
assign addr[31229]= -236640993;
assign addr[31230]= -274614114;
assign addr[31231]= -312500135;
assign addr[31232]= -350287041;
assign addr[31233]= -387962847;
assign addr[31234]= -425515602;
assign addr[31235]= -462933398;
assign addr[31236]= -500204365;
assign addr[31237]= -537316682;
assign addr[31238]= -574258580;
assign addr[31239]= -611018340;
assign addr[31240]= -647584304;
assign addr[31241]= -683944874;
assign addr[31242]= -720088517;
assign addr[31243]= -756003771;
assign addr[31244]= -791679244;
assign addr[31245]= -827103620;
assign addr[31246]= -862265664;
assign addr[31247]= -897154224;
assign addr[31248]= -931758235;
assign addr[31249]= -966066720;
assign addr[31250]= -1000068799;
assign addr[31251]= -1033753687;
assign addr[31252]= -1067110699;
assign addr[31253]= -1100129257;
assign addr[31254]= -1132798888;
assign addr[31255]= -1165109230;
assign addr[31256]= -1197050035;
assign addr[31257]= -1228611172;
assign addr[31258]= -1259782632;
assign addr[31259]= -1290554528;
assign addr[31260]= -1320917099;
assign addr[31261]= -1350860716;
assign addr[31262]= -1380375881;
assign addr[31263]= -1409453233;
assign addr[31264]= -1438083551;
assign addr[31265]= -1466257752;
assign addr[31266]= -1493966902;
assign addr[31267]= -1521202211;
assign addr[31268]= -1547955041;
assign addr[31269]= -1574216908;
assign addr[31270]= -1599979481;
assign addr[31271]= -1625234591;
assign addr[31272]= -1649974225;
assign addr[31273]= -1674190539;
assign addr[31274]= -1697875851;
assign addr[31275]= -1721022648;
assign addr[31276]= -1743623590;
assign addr[31277]= -1765671509;
assign addr[31278]= -1787159411;
assign addr[31279]= -1808080480;
assign addr[31280]= -1828428082;
assign addr[31281]= -1848195763;
assign addr[31282]= -1867377253;
assign addr[31283]= -1885966468;
assign addr[31284]= -1903957513;
assign addr[31285]= -1921344681;
assign addr[31286]= -1938122457;
assign addr[31287]= -1954285520;
assign addr[31288]= -1969828744;
assign addr[31289]= -1984747199;
assign addr[31290]= -1999036154;
assign addr[31291]= -2012691075;
assign addr[31292]= -2025707632;
assign addr[31293]= -2038081698;
assign addr[31294]= -2049809346;
assign addr[31295]= -2060886858;
assign addr[31296]= -2071310720;
assign addr[31297]= -2081077626;
assign addr[31298]= -2090184478;
assign addr[31299]= -2098628387;
assign addr[31300]= -2106406677;
assign addr[31301]= -2113516878;
assign addr[31302]= -2119956737;
assign addr[31303]= -2125724211;
assign addr[31304]= -2130817471;
assign addr[31305]= -2135234901;
assign addr[31306]= -2138975100;
assign addr[31307]= -2142036881;
assign addr[31308]= -2144419275;
assign addr[31309]= -2146121524;
assign addr[31310]= -2147143090;
assign addr[31311]= -2147483648;
assign addr[31312]= -2147143090;
assign addr[31313]= -2146121524;
assign addr[31314]= -2144419275;
assign addr[31315]= -2142036881;
assign addr[31316]= -2138975100;
assign addr[31317]= -2135234901;
assign addr[31318]= -2130817471;
assign addr[31319]= -2125724211;
assign addr[31320]= -2119956737;
assign addr[31321]= -2113516878;
assign addr[31322]= -2106406677;
assign addr[31323]= -2098628387;
assign addr[31324]= -2090184478;
assign addr[31325]= -2081077626;
assign addr[31326]= -2071310720;
assign addr[31327]= -2060886858;
assign addr[31328]= -2049809346;
assign addr[31329]= -2038081698;
assign addr[31330]= -2025707632;
assign addr[31331]= -2012691075;
assign addr[31332]= -1999036154;
assign addr[31333]= -1984747199;
assign addr[31334]= -1969828744;
assign addr[31335]= -1954285520;
assign addr[31336]= -1938122457;
assign addr[31337]= -1921344681;
assign addr[31338]= -1903957513;
assign addr[31339]= -1885966468;
assign addr[31340]= -1867377253;
assign addr[31341]= -1848195763;
assign addr[31342]= -1828428082;
assign addr[31343]= -1808080480;
assign addr[31344]= -1787159411;
assign addr[31345]= -1765671509;
assign addr[31346]= -1743623590;
assign addr[31347]= -1721022648;
assign addr[31348]= -1697875851;
assign addr[31349]= -1674190539;
assign addr[31350]= -1649974225;
assign addr[31351]= -1625234591;
assign addr[31352]= -1599979481;
assign addr[31353]= -1574216908;
assign addr[31354]= -1547955041;
assign addr[31355]= -1521202211;
assign addr[31356]= -1493966902;
assign addr[31357]= -1466257752;
assign addr[31358]= -1438083551;
assign addr[31359]= -1409453233;
assign addr[31360]= -1380375881;
assign addr[31361]= -1350860716;
assign addr[31362]= -1320917099;
assign addr[31363]= -1290554528;
assign addr[31364]= -1259782632;
assign addr[31365]= -1228611172;
assign addr[31366]= -1197050035;
assign addr[31367]= -1165109230;
assign addr[31368]= -1132798888;
assign addr[31369]= -1100129257;
assign addr[31370]= -1067110699;
assign addr[31371]= -1033753687;
assign addr[31372]= -1000068799;
assign addr[31373]= -966066720;
assign addr[31374]= -931758235;
assign addr[31375]= -897154224;
assign addr[31376]= -862265664;
assign addr[31377]= -827103620;
assign addr[31378]= -791679244;
assign addr[31379]= -756003771;
assign addr[31380]= -720088517;
assign addr[31381]= -683944874;
assign addr[31382]= -647584304;
assign addr[31383]= -611018340;
assign addr[31384]= -574258580;
assign addr[31385]= -537316682;
assign addr[31386]= -500204365;
assign addr[31387]= -462933398;
assign addr[31388]= -425515602;
assign addr[31389]= -387962847;
assign addr[31390]= -350287041;
assign addr[31391]= -312500135;
assign addr[31392]= -274614114;
assign addr[31393]= -236640993;
assign addr[31394]= -198592817;
assign addr[31395]= -160481654;
assign addr[31396]= -122319591;
assign addr[31397]= -84118732;
assign addr[31398]= -45891193;
assign addr[31399]= -7649098;
assign addr[31400]= 30595422;
assign addr[31401]= 68830239;
assign addr[31402]= 107043224;
assign addr[31403]= 145222259;
assign addr[31404]= 183355234;
assign addr[31405]= 221430054;
assign addr[31406]= 259434643;
assign addr[31407]= 297356948;
assign addr[31408]= 335184940;
assign addr[31409]= 372906622;
assign addr[31410]= 410510029;
assign addr[31411]= 447983235;
assign addr[31412]= 485314355;
assign addr[31413]= 522491548;
assign addr[31414]= 559503022;
assign addr[31415]= 596337040;
assign addr[31416]= 632981917;
assign addr[31417]= 669426032;
assign addr[31418]= 705657826;
assign addr[31419]= 741665807;
assign addr[31420]= 777438554;
assign addr[31421]= 812964722;
assign addr[31422]= 848233042;
assign addr[31423]= 883232329;
assign addr[31424]= 917951481;
assign addr[31425]= 952379488;
assign addr[31426]= 986505429;
assign addr[31427]= 1020318481;
assign addr[31428]= 1053807919;
assign addr[31429]= 1086963121;
assign addr[31430]= 1119773573;
assign addr[31431]= 1152228866;
assign addr[31432]= 1184318708;
assign addr[31433]= 1216032921;
assign addr[31434]= 1247361445;
assign addr[31435]= 1278294345;
assign addr[31436]= 1308821808;
assign addr[31437]= 1338934154;
assign addr[31438]= 1368621831;
assign addr[31439]= 1397875423;
assign addr[31440]= 1426685652;
assign addr[31441]= 1455043381;
assign addr[31442]= 1482939614;
assign addr[31443]= 1510365504;
assign addr[31444]= 1537312353;
assign addr[31445]= 1563771613;
assign addr[31446]= 1589734894;
assign addr[31447]= 1615193959;
assign addr[31448]= 1640140734;
assign addr[31449]= 1664567307;
assign addr[31450]= 1688465931;
assign addr[31451]= 1711829025;
assign addr[31452]= 1734649179;
assign addr[31453]= 1756919156;
assign addr[31454]= 1778631892;
assign addr[31455]= 1799780501;
assign addr[31456]= 1820358275;
assign addr[31457]= 1840358687;
assign addr[31458]= 1859775393;
assign addr[31459]= 1878602237;
assign addr[31460]= 1896833245;
assign addr[31461]= 1914462636;
assign addr[31462]= 1931484818;
assign addr[31463]= 1947894393;
assign addr[31464]= 1963686155;
assign addr[31465]= 1978855097;
assign addr[31466]= 1993396407;
assign addr[31467]= 2007305472;
assign addr[31468]= 2020577882;
assign addr[31469]= 2033209426;
assign addr[31470]= 2045196100;
assign addr[31471]= 2056534099;
assign addr[31472]= 2067219829;
assign addr[31473]= 2077249901;
assign addr[31474]= 2086621133;
assign addr[31475]= 2095330553;
assign addr[31476]= 2103375398;
assign addr[31477]= 2110753117;
assign addr[31478]= 2117461370;
assign addr[31479]= 2123498030;
assign addr[31480]= 2128861181;
assign addr[31481]= 2133549123;
assign addr[31482]= 2137560369;
assign addr[31483]= 2140893646;
assign addr[31484]= 2143547897;
assign addr[31485]= 2145522281;
assign addr[31486]= 2146816171;
assign addr[31487]= 2147429158;
assign addr[31488]= 2147361045;
assign addr[31489]= 2146611856;
assign addr[31490]= 2145181827;
assign addr[31491]= 2143071413;
assign addr[31492]= 2140281282;
assign addr[31493]= 2136812319;
assign addr[31494]= 2132665626;
assign addr[31495]= 2127842516;
assign addr[31496]= 2122344521;
assign addr[31497]= 2116173382;
assign addr[31498]= 2109331059;
assign addr[31499]= 2101819720;
assign addr[31500]= 2093641749;
assign addr[31501]= 2084799740;
assign addr[31502]= 2075296495;
assign addr[31503]= 2065135031;
assign addr[31504]= 2054318569;
assign addr[31505]= 2042850540;
assign addr[31506]= 2030734582;
assign addr[31507]= 2017974537;
assign addr[31508]= 2004574453;
assign addr[31509]= 1990538579;
assign addr[31510]= 1975871368;
assign addr[31511]= 1960577471;
assign addr[31512]= 1944661739;
assign addr[31513]= 1928129220;
assign addr[31514]= 1910985158;
assign addr[31515]= 1893234990;
assign addr[31516]= 1874884346;
assign addr[31517]= 1855939047;
assign addr[31518]= 1836405100;
assign addr[31519]= 1816288703;
assign addr[31520]= 1795596234;
assign addr[31521]= 1774334257;
assign addr[31522]= 1752509516;
assign addr[31523]= 1730128933;
assign addr[31524]= 1707199606;
assign addr[31525]= 1683728808;
assign addr[31526]= 1659723983;
assign addr[31527]= 1635192744;
assign addr[31528]= 1610142873;
assign addr[31529]= 1584582314;
assign addr[31530]= 1558519173;
assign addr[31531]= 1531961719;
assign addr[31532]= 1504918373;
assign addr[31533]= 1477397714;
assign addr[31534]= 1449408469;
assign addr[31535]= 1420959516;
assign addr[31536]= 1392059879;
assign addr[31537]= 1362718723;
assign addr[31538]= 1332945355;
assign addr[31539]= 1302749217;
assign addr[31540]= 1272139887;
assign addr[31541]= 1241127074;
assign addr[31542]= 1209720613;
assign addr[31543]= 1177930466;
assign addr[31544]= 1145766716;
assign addr[31545]= 1113239564;
assign addr[31546]= 1080359326;
assign addr[31547]= 1047136432;
assign addr[31548]= 1013581418;
assign addr[31549]= 979704927;
assign addr[31550]= 945517704;
assign addr[31551]= 911030591;
assign addr[31552]= 876254528;
assign addr[31553]= 841200544;
assign addr[31554]= 805879757;
assign addr[31555]= 770303369;
assign addr[31556]= 734482665;
assign addr[31557]= 698429006;
assign addr[31558]= 662153826;
assign addr[31559]= 625668632;
assign addr[31560]= 588984994;
assign addr[31561]= 552114549;
assign addr[31562]= 515068990;
assign addr[31563]= 477860067;
assign addr[31564]= 440499581;
assign addr[31565]= 402999383;
assign addr[31566]= 365371365;
assign addr[31567]= 327627463;
assign addr[31568]= 289779648;
assign addr[31569]= 251839923;
assign addr[31570]= 213820322;
assign addr[31571]= 175732905;
assign addr[31572]= 137589750;
assign addr[31573]= 99402956;
assign addr[31574]= 61184634;
assign addr[31575]= 22946906;
assign addr[31576]= -15298099;
assign addr[31577]= -53538253;
assign addr[31578]= -91761426;
assign addr[31579]= -129955495;
assign addr[31580]= -168108346;
assign addr[31581]= -206207878;
assign addr[31582]= -244242007;
assign addr[31583]= -282198671;
assign addr[31584]= -320065829;
assign addr[31585]= -357831473;
assign addr[31586]= -395483624;
assign addr[31587]= -433010339;
assign addr[31588]= -470399716;
assign addr[31589]= -507639898;
assign addr[31590]= -544719071;
assign addr[31591]= -581625477;
assign addr[31592]= -618347408;
assign addr[31593]= -654873219;
assign addr[31594]= -691191324;
assign addr[31595]= -727290205;
assign addr[31596]= -763158411;
assign addr[31597]= -798784567;
assign addr[31598]= -834157373;
assign addr[31599]= -869265610;
assign addr[31600]= -904098143;
assign addr[31601]= -938643924;
assign addr[31602]= -972891995;
assign addr[31603]= -1006831495;
assign addr[31604]= -1040451659;
assign addr[31605]= -1073741824;
assign addr[31606]= -1106691431;
assign addr[31607]= -1139290029;
assign addr[31608]= -1171527280;
assign addr[31609]= -1203392958;
assign addr[31610]= -1234876957;
assign addr[31611]= -1265969291;
assign addr[31612]= -1296660098;
assign addr[31613]= -1326939644;
assign addr[31614]= -1356798326;
assign addr[31615]= -1386226674;
assign addr[31616]= -1415215352;
assign addr[31617]= -1443755168;
assign addr[31618]= -1471837070;
assign addr[31619]= -1499452149;
assign addr[31620]= -1526591649;
assign addr[31621]= -1553246960;
assign addr[31622]= -1579409630;
assign addr[31623]= -1605071359;
assign addr[31624]= -1630224009;
assign addr[31625]= -1654859602;
assign addr[31626]= -1678970324;
assign addr[31627]= -1702548529;
assign addr[31628]= -1725586737;
assign addr[31629]= -1748077642;
assign addr[31630]= -1770014111;
assign addr[31631]= -1791389186;
assign addr[31632]= -1812196087;
assign addr[31633]= -1832428215;
assign addr[31634]= -1852079154;
assign addr[31635]= -1871142669;
assign addr[31636]= -1889612716;
assign addr[31637]= -1907483436;
assign addr[31638]= -1924749160;
assign addr[31639]= -1941404413;
assign addr[31640]= -1957443913;
assign addr[31641]= -1972862571;
assign addr[31642]= -1987655498;
assign addr[31643]= -2001818002;
assign addr[31644]= -2015345591;
assign addr[31645]= -2028233973;
assign addr[31646]= -2040479063;
assign addr[31647]= -2052076975;
assign addr[31648]= -2063024031;
assign addr[31649]= -2073316760;
assign addr[31650]= -2082951896;
assign addr[31651]= -2091926384;
assign addr[31652]= -2100237377;
assign addr[31653]= -2107882239;
assign addr[31654]= -2114858546;
assign addr[31655]= -2121164085;
assign addr[31656]= -2126796855;
assign addr[31657]= -2131755071;
assign addr[31658]= -2136037160;
assign addr[31659]= -2139641764;
assign addr[31660]= -2142567738;
assign addr[31661]= -2144814157;
assign addr[31662]= -2146380306;
assign addr[31663]= -2147265689;
assign addr[31664]= -2147470025;
assign addr[31665]= -2146993250;
assign addr[31666]= -2145835515;
assign addr[31667]= -2143997187;
assign addr[31668]= -2141478848;
assign addr[31669]= -2138281298;
assign addr[31670]= -2134405552;
assign addr[31671]= -2129852837;
assign addr[31672]= -2124624598;
assign addr[31673]= -2118722494;
assign addr[31674]= -2112148396;
assign addr[31675]= -2104904390;
assign addr[31676]= -2096992772;
assign addr[31677]= -2088416053;
assign addr[31678]= -2079176953;
assign addr[31679]= -2069278401;
assign addr[31680]= -2058723538;
assign addr[31681]= -2047515711;
assign addr[31682]= -2035658475;
assign addr[31683]= -2023155591;
assign addr[31684]= -2010011024;
assign addr[31685]= -1996228943;
assign addr[31686]= -1981813720;
assign addr[31687]= -1966769926;
assign addr[31688]= -1951102334;
assign addr[31689]= -1934815911;
assign addr[31690]= -1917915825;
assign addr[31691]= -1900407434;
assign addr[31692]= -1882296293;
assign addr[31693]= -1863588145;
assign addr[31694]= -1844288924;
assign addr[31695]= -1824404752;
assign addr[31696]= -1803941934;
assign addr[31697]= -1782906961;
assign addr[31698]= -1761306505;
assign addr[31699]= -1739147417;
assign addr[31700]= -1716436725;
assign addr[31701]= -1693181631;
assign addr[31702]= -1669389513;
assign addr[31703]= -1645067915;
assign addr[31704]= -1620224553;
assign addr[31705]= -1594867305;
assign addr[31706]= -1569004214;
assign addr[31707]= -1542643483;
assign addr[31708]= -1515793473;
assign addr[31709]= -1488462700;
assign addr[31710]= -1460659832;
assign addr[31711]= -1432393688;
assign addr[31712]= -1403673233;
assign addr[31713]= -1374507575;
assign addr[31714]= -1344905966;
assign addr[31715]= -1314877795;
assign addr[31716]= -1284432584;
assign addr[31717]= -1253579991;
assign addr[31718]= -1222329801;
assign addr[31719]= -1190691925;
assign addr[31720]= -1158676398;
assign addr[31721]= -1126293375;
assign addr[31722]= -1093553126;
assign addr[31723]= -1060466036;
assign addr[31724]= -1027042599;
assign addr[31725]= -993293415;
assign addr[31726]= -959229189;
assign addr[31727]= -924860725;
assign addr[31728]= -890198924;
assign addr[31729]= -855254778;
assign addr[31730]= -820039373;
assign addr[31731]= -784563876;
assign addr[31732]= -748839539;
assign addr[31733]= -712877694;
assign addr[31734]= -676689746;
assign addr[31735]= -640287172;
assign addr[31736]= -603681519;
assign addr[31737]= -566884397;
assign addr[31738]= -529907477;
assign addr[31739]= -492762486;
assign addr[31740]= -455461206;
assign addr[31741]= -418015468;
assign addr[31742]= -380437148;
assign addr[31743]= -342738165;
assign addr[31744]= -304930476;
assign addr[31745]= -267026072;
assign addr[31746]= -229036977;
assign addr[31747]= -190975237;
assign addr[31748]= -152852926;
assign addr[31749]= -114682135;
assign addr[31750]= -76474970;
assign addr[31751]= -38243550;
assign addr[31752]= 0;
assign addr[31753]= 38243550;
assign addr[31754]= 76474970;
assign addr[31755]= 114682135;
assign addr[31756]= 152852926;
assign addr[31757]= 190975237;
assign addr[31758]= 229036977;
assign addr[31759]= 267026072;
assign addr[31760]= 304930476;
assign addr[31761]= 342738165;
assign addr[31762]= 380437148;
assign addr[31763]= 418015468;
assign addr[31764]= 455461206;
assign addr[31765]= 492762486;
assign addr[31766]= 529907477;
assign addr[31767]= 566884397;
assign addr[31768]= 603681519;
assign addr[31769]= 640287172;
assign addr[31770]= 676689746;
assign addr[31771]= 712877694;
assign addr[31772]= 748839539;
assign addr[31773]= 784563876;
assign addr[31774]= 820039373;
assign addr[31775]= 855254778;
assign addr[31776]= 890198924;
assign addr[31777]= 924860725;
assign addr[31778]= 959229189;
assign addr[31779]= 993293415;
assign addr[31780]= 1027042599;
assign addr[31781]= 1060466036;
assign addr[31782]= 1093553126;
assign addr[31783]= 1126293375;
assign addr[31784]= 1158676398;
assign addr[31785]= 1190691925;
assign addr[31786]= 1222329801;
assign addr[31787]= 1253579991;
assign addr[31788]= 1284432584;
assign addr[31789]= 1314877795;
assign addr[31790]= 1344905966;
assign addr[31791]= 1374507575;
assign addr[31792]= 1403673233;
assign addr[31793]= 1432393688;
assign addr[31794]= 1460659832;
assign addr[31795]= 1488462700;
assign addr[31796]= 1515793473;
assign addr[31797]= 1542643483;
assign addr[31798]= 1569004214;
assign addr[31799]= 1594867305;
assign addr[31800]= 1620224553;
assign addr[31801]= 1645067915;
assign addr[31802]= 1669389513;
assign addr[31803]= 1693181631;
assign addr[31804]= 1716436725;
assign addr[31805]= 1739147417;
assign addr[31806]= 1761306505;
assign addr[31807]= 1782906961;
assign addr[31808]= 1803941934;
assign addr[31809]= 1824404752;
assign addr[31810]= 1844288924;
assign addr[31811]= 1863588145;
assign addr[31812]= 1882296293;
assign addr[31813]= 1900407434;
assign addr[31814]= 1917915825;
assign addr[31815]= 1934815911;
assign addr[31816]= 1951102334;
assign addr[31817]= 1966769926;
assign addr[31818]= 1981813720;
assign addr[31819]= 1996228943;
assign addr[31820]= 2010011024;
assign addr[31821]= 2023155591;
assign addr[31822]= 2035658475;
assign addr[31823]= 2047515711;
assign addr[31824]= 2058723538;
assign addr[31825]= 2069278401;
assign addr[31826]= 2079176953;
assign addr[31827]= 2088416053;
assign addr[31828]= 2096992772;
assign addr[31829]= 2104904390;
assign addr[31830]= 2112148396;
assign addr[31831]= 2118722494;
assign addr[31832]= 2124624598;
assign addr[31833]= 2129852837;
assign addr[31834]= 2134405552;
assign addr[31835]= 2138281298;
assign addr[31836]= 2141478848;
assign addr[31837]= 2143997187;
assign addr[31838]= 2145835515;
assign addr[31839]= 2146993250;
assign addr[31840]= 2147470025;
assign addr[31841]= 2147265689;
assign addr[31842]= 2146380306;
assign addr[31843]= 2144814157;
assign addr[31844]= 2142567738;
assign addr[31845]= 2139641764;
assign addr[31846]= 2136037160;
assign addr[31847]= 2131755071;
assign addr[31848]= 2126796855;
assign addr[31849]= 2121164085;
assign addr[31850]= 2114858546;
assign addr[31851]= 2107882239;
assign addr[31852]= 2100237377;
assign addr[31853]= 2091926384;
assign addr[31854]= 2082951896;
assign addr[31855]= 2073316760;
assign addr[31856]= 2063024031;
assign addr[31857]= 2052076975;
assign addr[31858]= 2040479063;
assign addr[31859]= 2028233973;
assign addr[31860]= 2015345591;
assign addr[31861]= 2001818002;
assign addr[31862]= 1987655498;
assign addr[31863]= 1972862571;
assign addr[31864]= 1957443913;
assign addr[31865]= 1941404413;
assign addr[31866]= 1924749160;
assign addr[31867]= 1907483436;
assign addr[31868]= 1889612716;
assign addr[31869]= 1871142669;
assign addr[31870]= 1852079154;
assign addr[31871]= 1832428215;
assign addr[31872]= 1812196087;
assign addr[31873]= 1791389186;
assign addr[31874]= 1770014111;
assign addr[31875]= 1748077642;
assign addr[31876]= 1725586737;
assign addr[31877]= 1702548529;
assign addr[31878]= 1678970324;
assign addr[31879]= 1654859602;
assign addr[31880]= 1630224009;
assign addr[31881]= 1605071359;
assign addr[31882]= 1579409630;
assign addr[31883]= 1553246960;
assign addr[31884]= 1526591649;
assign addr[31885]= 1499452149;
assign addr[31886]= 1471837070;
assign addr[31887]= 1443755168;
assign addr[31888]= 1415215352;
assign addr[31889]= 1386226674;
assign addr[31890]= 1356798326;
assign addr[31891]= 1326939644;
assign addr[31892]= 1296660098;
assign addr[31893]= 1265969291;
assign addr[31894]= 1234876957;
assign addr[31895]= 1203392958;
assign addr[31896]= 1171527280;
assign addr[31897]= 1139290029;
assign addr[31898]= 1106691431;
assign addr[31899]= 1073741824;
assign addr[31900]= 1040451659;
assign addr[31901]= 1006831495;
assign addr[31902]= 972891995;
assign addr[31903]= 938643924;
assign addr[31904]= 904098143;
assign addr[31905]= 869265610;
assign addr[31906]= 834157373;
assign addr[31907]= 798784567;
assign addr[31908]= 763158411;
assign addr[31909]= 727290205;
assign addr[31910]= 691191324;
assign addr[31911]= 654873219;
assign addr[31912]= 618347408;
assign addr[31913]= 581625477;
assign addr[31914]= 544719071;
assign addr[31915]= 507639898;
assign addr[31916]= 470399716;
assign addr[31917]= 433010339;
assign addr[31918]= 395483624;
assign addr[31919]= 357831473;
assign addr[31920]= 320065829;
assign addr[31921]= 282198671;
assign addr[31922]= 244242007;
assign addr[31923]= 206207878;
assign addr[31924]= 168108346;
assign addr[31925]= 129955495;
assign addr[31926]= 91761426;
assign addr[31927]= 53538253;
assign addr[31928]= 15298099;
assign addr[31929]= -22946906;
assign addr[31930]= -61184634;
assign addr[31931]= -99402956;
assign addr[31932]= -137589750;
assign addr[31933]= -175732905;
assign addr[31934]= -213820322;
assign addr[31935]= -251839923;
assign addr[31936]= -289779648;
assign addr[31937]= -327627463;
assign addr[31938]= -365371365;
assign addr[31939]= -402999383;
assign addr[31940]= -440499581;
assign addr[31941]= -477860067;
assign addr[31942]= -515068990;
assign addr[31943]= -552114549;
assign addr[31944]= -588984994;
assign addr[31945]= -625668632;
assign addr[31946]= -662153826;
assign addr[31947]= -698429006;
assign addr[31948]= -734482665;
assign addr[31949]= -770303369;
assign addr[31950]= -805879757;
assign addr[31951]= -841200544;
assign addr[31952]= -876254528;
assign addr[31953]= -911030591;
assign addr[31954]= -945517704;
assign addr[31955]= -979704927;
assign addr[31956]= -1013581418;
assign addr[31957]= -1047136432;
assign addr[31958]= -1080359326;
assign addr[31959]= -1113239564;
assign addr[31960]= -1145766716;
assign addr[31961]= -1177930466;
assign addr[31962]= -1209720613;
assign addr[31963]= -1241127074;
assign addr[31964]= -1272139887;
assign addr[31965]= -1302749217;
assign addr[31966]= -1332945355;
assign addr[31967]= -1362718723;
assign addr[31968]= -1392059879;
assign addr[31969]= -1420959516;
assign addr[31970]= -1449408469;
assign addr[31971]= -1477397714;
assign addr[31972]= -1504918373;
assign addr[31973]= -1531961719;
assign addr[31974]= -1558519173;
assign addr[31975]= -1584582314;
assign addr[31976]= -1610142873;
assign addr[31977]= -1635192744;
assign addr[31978]= -1659723983;
assign addr[31979]= -1683728808;
assign addr[31980]= -1707199606;
assign addr[31981]= -1730128933;
assign addr[31982]= -1752509516;
assign addr[31983]= -1774334257;
assign addr[31984]= -1795596234;
assign addr[31985]= -1816288703;
assign addr[31986]= -1836405100;
assign addr[31987]= -1855939047;
assign addr[31988]= -1874884346;
assign addr[31989]= -1893234990;
assign addr[31990]= -1910985158;
assign addr[31991]= -1928129220;
assign addr[31992]= -1944661739;
assign addr[31993]= -1960577471;
assign addr[31994]= -1975871368;
assign addr[31995]= -1990538579;
assign addr[31996]= -2004574453;
assign addr[31997]= -2017974537;
assign addr[31998]= -2030734582;
assign addr[31999]= -2042850540;
assign addr[32000]= -2054318569;
assign addr[32001]= -2065135031;
assign addr[32002]= -2075296495;
assign addr[32003]= -2084799740;
assign addr[32004]= -2093641749;
assign addr[32005]= -2101819720;
assign addr[32006]= -2109331059;
assign addr[32007]= -2116173382;
assign addr[32008]= -2122344521;
assign addr[32009]= -2127842516;
assign addr[32010]= -2132665626;
assign addr[32011]= -2136812319;
assign addr[32012]= -2140281282;
assign addr[32013]= -2143071413;
assign addr[32014]= -2145181827;
assign addr[32015]= -2146611856;
assign addr[32016]= -2147361045;
assign addr[32017]= -2147429158;
assign addr[32018]= -2146816171;
assign addr[32019]= -2145522281;
assign addr[32020]= -2143547897;
assign addr[32021]= -2140893646;
assign addr[32022]= -2137560369;
assign addr[32023]= -2133549123;
assign addr[32024]= -2128861181;
assign addr[32025]= -2123498030;
assign addr[32026]= -2117461370;
assign addr[32027]= -2110753117;
assign addr[32028]= -2103375398;
assign addr[32029]= -2095330553;
assign addr[32030]= -2086621133;
assign addr[32031]= -2077249901;
assign addr[32032]= -2067219829;
assign addr[32033]= -2056534099;
assign addr[32034]= -2045196100;
assign addr[32035]= -2033209426;
assign addr[32036]= -2020577882;
assign addr[32037]= -2007305472;
assign addr[32038]= -1993396407;
assign addr[32039]= -1978855097;
assign addr[32040]= -1963686155;
assign addr[32041]= -1947894393;
assign addr[32042]= -1931484818;
assign addr[32043]= -1914462636;
assign addr[32044]= -1896833245;
assign addr[32045]= -1878602237;
assign addr[32046]= -1859775393;
assign addr[32047]= -1840358687;
assign addr[32048]= -1820358275;
assign addr[32049]= -1799780501;
assign addr[32050]= -1778631892;
assign addr[32051]= -1756919156;
assign addr[32052]= -1734649179;
assign addr[32053]= -1711829025;
assign addr[32054]= -1688465931;
assign addr[32055]= -1664567307;
assign addr[32056]= -1640140734;
assign addr[32057]= -1615193959;
assign addr[32058]= -1589734894;
assign addr[32059]= -1563771613;
assign addr[32060]= -1537312353;
assign addr[32061]= -1510365504;
assign addr[32062]= -1482939614;
assign addr[32063]= -1455043381;
assign addr[32064]= -1426685652;
assign addr[32065]= -1397875423;
assign addr[32066]= -1368621831;
assign addr[32067]= -1338934154;
assign addr[32068]= -1308821808;
assign addr[32069]= -1278294345;
assign addr[32070]= -1247361445;
assign addr[32071]= -1216032921;
assign addr[32072]= -1184318708;
assign addr[32073]= -1152228866;
assign addr[32074]= -1119773573;
assign addr[32075]= -1086963121;
assign addr[32076]= -1053807919;
assign addr[32077]= -1020318481;
assign addr[32078]= -986505429;
assign addr[32079]= -952379488;
assign addr[32080]= -917951481;
assign addr[32081]= -883232329;
assign addr[32082]= -848233042;
assign addr[32083]= -812964722;
assign addr[32084]= -777438554;
assign addr[32085]= -741665807;
assign addr[32086]= -705657826;
assign addr[32087]= -669426032;
assign addr[32088]= -632981917;
assign addr[32089]= -596337040;
assign addr[32090]= -559503022;
assign addr[32091]= -522491548;
assign addr[32092]= -485314355;
assign addr[32093]= -447983235;
assign addr[32094]= -410510029;
assign addr[32095]= -372906622;
assign addr[32096]= -335184940;
assign addr[32097]= -297356948;
assign addr[32098]= -259434643;
assign addr[32099]= -221430054;
assign addr[32100]= -183355234;
assign addr[32101]= -145222259;
assign addr[32102]= -107043224;
assign addr[32103]= -68830239;
assign addr[32104]= -30595422;
assign addr[32105]= 7649098;
assign addr[32106]= 45891193;
assign addr[32107]= 84118732;
assign addr[32108]= 122319591;
assign addr[32109]= 160481654;
assign addr[32110]= 198592817;
assign addr[32111]= 236640993;
assign addr[32112]= 274614114;
assign addr[32113]= 312500135;
assign addr[32114]= 350287041;
assign addr[32115]= 387962847;
assign addr[32116]= 425515602;
assign addr[32117]= 462933398;
assign addr[32118]= 500204365;
assign addr[32119]= 537316682;
assign addr[32120]= 574258580;
assign addr[32121]= 611018340;
assign addr[32122]= 647584304;
assign addr[32123]= 683944874;
assign addr[32124]= 720088517;
assign addr[32125]= 756003771;
assign addr[32126]= 791679244;
assign addr[32127]= 827103620;
assign addr[32128]= 862265664;
assign addr[32129]= 897154224;
assign addr[32130]= 931758235;
assign addr[32131]= 966066720;
assign addr[32132]= 1000068799;
assign addr[32133]= 1033753687;
assign addr[32134]= 1067110699;
assign addr[32135]= 1100129257;
assign addr[32136]= 1132798888;
assign addr[32137]= 1165109230;
assign addr[32138]= 1197050035;
assign addr[32139]= 1228611172;
assign addr[32140]= 1259782632;
assign addr[32141]= 1290554528;
assign addr[32142]= 1320917099;
assign addr[32143]= 1350860716;
assign addr[32144]= 1380375881;
assign addr[32145]= 1409453233;
assign addr[32146]= 1438083551;
assign addr[32147]= 1466257752;
assign addr[32148]= 1493966902;
assign addr[32149]= 1521202211;
assign addr[32150]= 1547955041;
assign addr[32151]= 1574216908;
assign addr[32152]= 1599979481;
assign addr[32153]= 1625234591;
assign addr[32154]= 1649974225;
assign addr[32155]= 1674190539;
assign addr[32156]= 1697875851;
assign addr[32157]= 1721022648;
assign addr[32158]= 1743623590;
assign addr[32159]= 1765671509;
assign addr[32160]= 1787159411;
assign addr[32161]= 1808080480;
assign addr[32162]= 1828428082;
assign addr[32163]= 1848195763;
assign addr[32164]= 1867377253;
assign addr[32165]= 1885966468;
assign addr[32166]= 1903957513;
assign addr[32167]= 1921344681;
assign addr[32168]= 1938122457;
assign addr[32169]= 1954285520;
assign addr[32170]= 1969828744;
assign addr[32171]= 1984747199;
assign addr[32172]= 1999036154;
assign addr[32173]= 2012691075;
assign addr[32174]= 2025707632;
assign addr[32175]= 2038081698;
assign addr[32176]= 2049809346;
assign addr[32177]= 2060886858;
assign addr[32178]= 2071310720;
assign addr[32179]= 2081077626;
assign addr[32180]= 2090184478;
assign addr[32181]= 2098628387;
assign addr[32182]= 2106406677;
assign addr[32183]= 2113516878;
assign addr[32184]= 2119956737;
assign addr[32185]= 2125724211;
assign addr[32186]= 2130817471;
assign addr[32187]= 2135234901;
assign addr[32188]= 2138975100;
assign addr[32189]= 2142036881;
assign addr[32190]= 2144419275;
assign addr[32191]= 2146121524;
assign addr[32192]= 2147143090;
assign addr[32193]= 2147483648;
assign addr[32194]= 2147143090;
assign addr[32195]= 2146121524;
assign addr[32196]= 2144419275;
assign addr[32197]= 2142036881;
assign addr[32198]= 2138975100;
assign addr[32199]= 2135234901;
assign addr[32200]= 2130817471;
assign addr[32201]= 2125724211;
assign addr[32202]= 2119956737;
assign addr[32203]= 2113516878;
assign addr[32204]= 2106406677;
assign addr[32205]= 2098628387;
assign addr[32206]= 2090184478;
assign addr[32207]= 2081077626;
assign addr[32208]= 2071310720;
assign addr[32209]= 2060886858;
assign addr[32210]= 2049809346;
assign addr[32211]= 2038081698;
assign addr[32212]= 2025707632;
assign addr[32213]= 2012691075;
assign addr[32214]= 1999036154;
assign addr[32215]= 1984747199;
assign addr[32216]= 1969828744;
assign addr[32217]= 1954285520;
assign addr[32218]= 1938122457;
assign addr[32219]= 1921344681;
assign addr[32220]= 1903957513;
assign addr[32221]= 1885966468;
assign addr[32222]= 1867377253;
assign addr[32223]= 1848195763;
assign addr[32224]= 1828428082;
assign addr[32225]= 1808080480;
assign addr[32226]= 1787159411;
assign addr[32227]= 1765671509;
assign addr[32228]= 1743623590;
assign addr[32229]= 1721022648;
assign addr[32230]= 1697875851;
assign addr[32231]= 1674190539;
assign addr[32232]= 1649974225;
assign addr[32233]= 1625234591;
assign addr[32234]= 1599979481;
assign addr[32235]= 1574216908;
assign addr[32236]= 1547955041;
assign addr[32237]= 1521202211;
assign addr[32238]= 1493966902;
assign addr[32239]= 1466257752;
assign addr[32240]= 1438083551;
assign addr[32241]= 1409453233;
assign addr[32242]= 1380375881;
assign addr[32243]= 1350860716;
assign addr[32244]= 1320917099;
assign addr[32245]= 1290554528;
assign addr[32246]= 1259782632;
assign addr[32247]= 1228611172;
assign addr[32248]= 1197050035;
assign addr[32249]= 1165109230;
assign addr[32250]= 1132798888;
assign addr[32251]= 1100129257;
assign addr[32252]= 1067110699;
assign addr[32253]= 1033753687;
assign addr[32254]= 1000068799;
assign addr[32255]= 966066720;
assign addr[32256]= 931758235;
assign addr[32257]= 897154224;
assign addr[32258]= 862265664;
assign addr[32259]= 827103620;
assign addr[32260]= 791679244;
assign addr[32261]= 756003771;
assign addr[32262]= 720088517;
assign addr[32263]= 683944874;
assign addr[32264]= 647584304;
assign addr[32265]= 611018340;
assign addr[32266]= 574258580;
assign addr[32267]= 537316682;
assign addr[32268]= 500204365;
assign addr[32269]= 462933398;
assign addr[32270]= 425515602;
assign addr[32271]= 387962847;
assign addr[32272]= 350287041;
assign addr[32273]= 312500135;
assign addr[32274]= 274614114;
assign addr[32275]= 236640993;
assign addr[32276]= 198592817;
assign addr[32277]= 160481654;
assign addr[32278]= 122319591;
assign addr[32279]= 84118732;
assign addr[32280]= 45891193;
assign addr[32281]= 7649098;
assign addr[32282]= -30595422;
assign addr[32283]= -68830239;
assign addr[32284]= -107043224;
assign addr[32285]= -145222259;
assign addr[32286]= -183355234;
assign addr[32287]= -221430054;
assign addr[32288]= -259434643;
assign addr[32289]= -297356948;
assign addr[32290]= -335184940;
assign addr[32291]= -372906622;
assign addr[32292]= -410510029;
assign addr[32293]= -447983235;
assign addr[32294]= -485314355;
assign addr[32295]= -522491548;
assign addr[32296]= -559503022;
assign addr[32297]= -596337040;
assign addr[32298]= -632981917;
assign addr[32299]= -669426032;
assign addr[32300]= -705657826;
assign addr[32301]= -741665807;
assign addr[32302]= -777438554;
assign addr[32303]= -812964722;
assign addr[32304]= -848233042;
assign addr[32305]= -883232329;
assign addr[32306]= -917951481;
assign addr[32307]= -952379488;
assign addr[32308]= -986505429;
assign addr[32309]= -1020318481;
assign addr[32310]= -1053807919;
assign addr[32311]= -1086963121;
assign addr[32312]= -1119773573;
assign addr[32313]= -1152228866;
assign addr[32314]= -1184318708;
assign addr[32315]= -1216032921;
assign addr[32316]= -1247361445;
assign addr[32317]= -1278294345;
assign addr[32318]= -1308821808;
assign addr[32319]= -1338934154;
assign addr[32320]= -1368621831;
assign addr[32321]= -1397875423;
assign addr[32322]= -1426685652;
assign addr[32323]= -1455043381;
assign addr[32324]= -1482939614;
assign addr[32325]= -1510365504;
assign addr[32326]= -1537312353;
assign addr[32327]= -1563771613;
assign addr[32328]= -1589734894;
assign addr[32329]= -1615193959;
assign addr[32330]= -1640140734;
assign addr[32331]= -1664567307;
assign addr[32332]= -1688465931;
assign addr[32333]= -1711829025;
assign addr[32334]= -1734649179;
assign addr[32335]= -1756919156;
assign addr[32336]= -1778631892;
assign addr[32337]= -1799780501;
assign addr[32338]= -1820358275;
assign addr[32339]= -1840358687;
assign addr[32340]= -1859775393;
assign addr[32341]= -1878602237;
assign addr[32342]= -1896833245;
assign addr[32343]= -1914462636;
assign addr[32344]= -1931484818;
assign addr[32345]= -1947894393;
assign addr[32346]= -1963686155;
assign addr[32347]= -1978855097;
assign addr[32348]= -1993396407;
assign addr[32349]= -2007305472;
assign addr[32350]= -2020577882;
assign addr[32351]= -2033209426;
assign addr[32352]= -2045196100;
assign addr[32353]= -2056534099;
assign addr[32354]= -2067219829;
assign addr[32355]= -2077249901;
assign addr[32356]= -2086621133;
assign addr[32357]= -2095330553;
assign addr[32358]= -2103375398;
assign addr[32359]= -2110753117;
assign addr[32360]= -2117461370;
assign addr[32361]= -2123498030;
assign addr[32362]= -2128861181;
assign addr[32363]= -2133549123;
assign addr[32364]= -2137560369;
assign addr[32365]= -2140893646;
assign addr[32366]= -2143547897;
assign addr[32367]= -2145522281;
assign addr[32368]= -2146816171;
assign addr[32369]= -2147429158;
assign addr[32370]= -2147361045;
assign addr[32371]= -2146611856;
assign addr[32372]= -2145181827;
assign addr[32373]= -2143071413;
assign addr[32374]= -2140281282;
assign addr[32375]= -2136812319;
assign addr[32376]= -2132665626;
assign addr[32377]= -2127842516;
assign addr[32378]= -2122344521;
assign addr[32379]= -2116173382;
assign addr[32380]= -2109331059;
assign addr[32381]= -2101819720;
assign addr[32382]= -2093641749;
assign addr[32383]= -2084799740;
assign addr[32384]= -2075296495;
assign addr[32385]= -2065135031;
assign addr[32386]= -2054318569;
assign addr[32387]= -2042850540;
assign addr[32388]= -2030734582;
assign addr[32389]= -2017974537;
assign addr[32390]= -2004574453;
assign addr[32391]= -1990538579;
assign addr[32392]= -1975871368;
assign addr[32393]= -1960577471;
assign addr[32394]= -1944661739;
assign addr[32395]= -1928129220;
assign addr[32396]= -1910985158;
assign addr[32397]= -1893234990;
assign addr[32398]= -1874884346;
assign addr[32399]= -1855939047;
assign addr[32400]= -1836405100;
assign addr[32401]= -1816288703;
assign addr[32402]= -1795596234;
assign addr[32403]= -1774334257;
assign addr[32404]= -1752509516;
assign addr[32405]= -1730128933;
assign addr[32406]= -1707199606;
assign addr[32407]= -1683728808;
assign addr[32408]= -1659723983;
assign addr[32409]= -1635192744;
assign addr[32410]= -1610142873;
assign addr[32411]= -1584582314;
assign addr[32412]= -1558519173;
assign addr[32413]= -1531961719;
assign addr[32414]= -1504918373;
assign addr[32415]= -1477397714;
assign addr[32416]= -1449408469;
assign addr[32417]= -1420959516;
assign addr[32418]= -1392059879;
assign addr[32419]= -1362718723;
assign addr[32420]= -1332945355;
assign addr[32421]= -1302749217;
assign addr[32422]= -1272139887;
assign addr[32423]= -1241127074;
assign addr[32424]= -1209720613;
assign addr[32425]= -1177930466;
assign addr[32426]= -1145766716;
assign addr[32427]= -1113239564;
assign addr[32428]= -1080359326;
assign addr[32429]= -1047136432;
assign addr[32430]= -1013581418;
assign addr[32431]= -979704927;
assign addr[32432]= -945517704;
assign addr[32433]= -911030591;
assign addr[32434]= -876254528;
assign addr[32435]= -841200544;
assign addr[32436]= -805879757;
assign addr[32437]= -770303369;
assign addr[32438]= -734482665;
assign addr[32439]= -698429006;
assign addr[32440]= -662153826;
assign addr[32441]= -625668632;
assign addr[32442]= -588984994;
assign addr[32443]= -552114549;
assign addr[32444]= -515068990;
assign addr[32445]= -477860067;
assign addr[32446]= -440499581;
assign addr[32447]= -402999383;
assign addr[32448]= -365371365;
assign addr[32449]= -327627463;
assign addr[32450]= -289779648;
assign addr[32451]= -251839923;
assign addr[32452]= -213820322;
assign addr[32453]= -175732905;
assign addr[32454]= -137589750;
assign addr[32455]= -99402956;
assign addr[32456]= -61184634;
assign addr[32457]= -22946906;
assign addr[32458]= 15298099;
assign addr[32459]= 53538253;
assign addr[32460]= 91761426;
assign addr[32461]= 129955495;
assign addr[32462]= 168108346;
assign addr[32463]= 206207878;
assign addr[32464]= 244242007;
assign addr[32465]= 282198671;
assign addr[32466]= 320065829;
assign addr[32467]= 357831473;
assign addr[32468]= 395483624;
assign addr[32469]= 433010339;
assign addr[32470]= 470399716;
assign addr[32471]= 507639898;
assign addr[32472]= 544719071;
assign addr[32473]= 581625477;
assign addr[32474]= 618347408;
assign addr[32475]= 654873219;
assign addr[32476]= 691191324;
assign addr[32477]= 727290205;
assign addr[32478]= 763158411;
assign addr[32479]= 798784567;
assign addr[32480]= 834157373;
assign addr[32481]= 869265610;
assign addr[32482]= 904098143;
assign addr[32483]= 938643924;
assign addr[32484]= 972891995;
assign addr[32485]= 1006831495;
assign addr[32486]= 1040451659;
assign addr[32487]= 1073741824;
assign addr[32488]= 1106691431;
assign addr[32489]= 1139290029;
assign addr[32490]= 1171527280;
assign addr[32491]= 1203392958;
assign addr[32492]= 1234876957;
assign addr[32493]= 1265969291;
assign addr[32494]= 1296660098;
assign addr[32495]= 1326939644;
assign addr[32496]= 1356798326;
assign addr[32497]= 1386226674;
assign addr[32498]= 1415215352;
assign addr[32499]= 1443755168;
assign addr[32500]= 1471837070;
assign addr[32501]= 1499452149;
assign addr[32502]= 1526591649;
assign addr[32503]= 1553246960;
assign addr[32504]= 1579409630;
assign addr[32505]= 1605071359;
assign addr[32506]= 1630224009;
assign addr[32507]= 1654859602;
assign addr[32508]= 1678970324;
assign addr[32509]= 1702548529;
assign addr[32510]= 1725586737;
assign addr[32511]= 1748077642;
assign addr[32512]= 1770014111;
assign addr[32513]= 1791389186;
assign addr[32514]= 1812196087;
assign addr[32515]= 1832428215;
assign addr[32516]= 1852079154;
assign addr[32517]= 1871142669;
assign addr[32518]= 1889612716;
assign addr[32519]= 1907483436;
assign addr[32520]= 1924749160;
assign addr[32521]= 1941404413;
assign addr[32522]= 1957443913;
assign addr[32523]= 1972862571;
assign addr[32524]= 1987655498;
assign addr[32525]= 2001818002;
assign addr[32526]= 2015345591;
assign addr[32527]= 2028233973;
assign addr[32528]= 2040479063;
assign addr[32529]= 2052076975;
assign addr[32530]= 2063024031;
assign addr[32531]= 2073316760;
assign addr[32532]= 2082951896;
assign addr[32533]= 2091926384;
assign addr[32534]= 2100237377;
assign addr[32535]= 2107882239;
assign addr[32536]= 2114858546;
assign addr[32537]= 2121164085;
assign addr[32538]= 2126796855;
assign addr[32539]= 2131755071;
assign addr[32540]= 2136037160;
assign addr[32541]= 2139641764;
assign addr[32542]= 2142567738;
assign addr[32543]= 2144814157;
assign addr[32544]= 2146380306;
assign addr[32545]= 2147265689;
assign addr[32546]= 2147470025;
assign addr[32547]= 2146993250;
assign addr[32548]= 2145835515;
assign addr[32549]= 2143997187;
assign addr[32550]= 2141478848;
assign addr[32551]= 2138281298;
assign addr[32552]= 2134405552;
assign addr[32553]= 2129852837;
assign addr[32554]= 2124624598;
assign addr[32555]= 2118722494;
assign addr[32556]= 2112148396;
assign addr[32557]= 2104904390;
assign addr[32558]= 2096992772;
assign addr[32559]= 2088416053;
assign addr[32560]= 2079176953;
assign addr[32561]= 2069278401;
assign addr[32562]= 2058723538;
assign addr[32563]= 2047515711;
assign addr[32564]= 2035658475;
assign addr[32565]= 2023155591;
assign addr[32566]= 2010011024;
assign addr[32567]= 1996228943;
assign addr[32568]= 1981813720;
assign addr[32569]= 1966769926;
assign addr[32570]= 1951102334;
assign addr[32571]= 1934815911;
assign addr[32572]= 1917915825;
assign addr[32573]= 1900407434;
assign addr[32574]= 1882296293;
assign addr[32575]= 1863588145;
assign addr[32576]= 1844288924;
assign addr[32577]= 1824404752;
assign addr[32578]= 1803941934;
assign addr[32579]= 1782906961;
assign addr[32580]= 1761306505;
assign addr[32581]= 1739147417;
assign addr[32582]= 1716436725;
assign addr[32583]= 1693181631;
assign addr[32584]= 1669389513;
assign addr[32585]= 1645067915;
assign addr[32586]= 1620224553;
assign addr[32587]= 1594867305;
assign addr[32588]= 1569004214;
assign addr[32589]= 1542643483;
assign addr[32590]= 1515793473;
assign addr[32591]= 1488462700;
assign addr[32592]= 1460659832;
assign addr[32593]= 1432393688;
assign addr[32594]= 1403673233;
assign addr[32595]= 1374507575;
assign addr[32596]= 1344905966;
assign addr[32597]= 1314877795;
assign addr[32598]= 1284432584;
assign addr[32599]= 1253579991;
assign addr[32600]= 1222329801;
assign addr[32601]= 1190691925;
assign addr[32602]= 1158676398;
assign addr[32603]= 1126293375;
assign addr[32604]= 1093553126;
assign addr[32605]= 1060466036;
assign addr[32606]= 1027042599;
assign addr[32607]= 993293415;
assign addr[32608]= 959229189;
assign addr[32609]= 924860725;
assign addr[32610]= 890198924;
assign addr[32611]= 855254778;
assign addr[32612]= 820039373;
assign addr[32613]= 784563876;
assign addr[32614]= 748839539;
assign addr[32615]= 712877694;
assign addr[32616]= 676689746;
assign addr[32617]= 640287172;
assign addr[32618]= 603681519;
assign addr[32619]= 566884397;
assign addr[32620]= 529907477;
assign addr[32621]= 492762486;
assign addr[32622]= 455461206;
assign addr[32623]= 418015468;
assign addr[32624]= 380437148;
assign addr[32625]= 342738165;
assign addr[32626]= 304930476;
assign addr[32627]= 267026072;
assign addr[32628]= 229036977;
assign addr[32629]= 190975237;
assign addr[32630]= 152852926;
assign addr[32631]= 114682135;
assign addr[32632]= 76474970;
assign addr[32633]= 38243550;
assign addr[32634]= 0;
assign addr[32635]= -38243550;
assign addr[32636]= -76474970;
assign addr[32637]= -114682135;
assign addr[32638]= -152852926;
assign addr[32639]= -190975237;
assign addr[32640]= -229036977;
assign addr[32641]= -267026072;
assign addr[32642]= -304930476;
assign addr[32643]= -342738165;
assign addr[32644]= -380437148;
assign addr[32645]= -418015468;
assign addr[32646]= -455461206;
assign addr[32647]= -492762486;
assign addr[32648]= -529907477;
assign addr[32649]= -566884397;
assign addr[32650]= -603681519;
assign addr[32651]= -640287172;
assign addr[32652]= -676689746;
assign addr[32653]= -712877694;
assign addr[32654]= -748839539;
assign addr[32655]= -784563876;
assign addr[32656]= -820039373;
assign addr[32657]= -855254778;
assign addr[32658]= -890198924;
assign addr[32659]= -924860725;
assign addr[32660]= -959229189;
assign addr[32661]= -993293415;
assign addr[32662]= -1027042599;
assign addr[32663]= -1060466036;
assign addr[32664]= -1093553126;
assign addr[32665]= -1126293375;
assign addr[32666]= -1158676398;
assign addr[32667]= -1190691925;
assign addr[32668]= -1222329801;
assign addr[32669]= -1253579991;
assign addr[32670]= -1284432584;
assign addr[32671]= -1314877795;
assign addr[32672]= -1344905966;
assign addr[32673]= -1374507575;
assign addr[32674]= -1403673233;
assign addr[32675]= -1432393688;
assign addr[32676]= -1460659832;
assign addr[32677]= -1488462700;
assign addr[32678]= -1515793473;
assign addr[32679]= -1542643483;
assign addr[32680]= -1569004214;
assign addr[32681]= -1594867305;
assign addr[32682]= -1620224553;
assign addr[32683]= -1645067915;
assign addr[32684]= -1669389513;
assign addr[32685]= -1693181631;
assign addr[32686]= -1716436725;
assign addr[32687]= -1739147417;
assign addr[32688]= -1761306505;
assign addr[32689]= -1782906961;
assign addr[32690]= -1803941934;
assign addr[32691]= -1824404752;
assign addr[32692]= -1844288924;
assign addr[32693]= -1863588145;
assign addr[32694]= -1882296293;
assign addr[32695]= -1900407434;
assign addr[32696]= -1917915825;
assign addr[32697]= -1934815911;
assign addr[32698]= -1951102334;
assign addr[32699]= -1966769926;
assign addr[32700]= -1981813720;
assign addr[32701]= -1996228943;
assign addr[32702]= -2010011024;
assign addr[32703]= -2023155591;
assign addr[32704]= -2035658475;
assign addr[32705]= -2047515711;
assign addr[32706]= -2058723538;
assign addr[32707]= -2069278401;
assign addr[32708]= -2079176953;
assign addr[32709]= -2088416053;
assign addr[32710]= -2096992772;
assign addr[32711]= -2104904390;
assign addr[32712]= -2112148396;
assign addr[32713]= -2118722494;
assign addr[32714]= -2124624598;
assign addr[32715]= -2129852837;
assign addr[32716]= -2134405552;
assign addr[32717]= -2138281298;
assign addr[32718]= -2141478848;
assign addr[32719]= -2143997187;
assign addr[32720]= -2145835515;
assign addr[32721]= -2146993250;
assign addr[32722]= -2147470025;
assign addr[32723]= -2147265689;
assign addr[32724]= -2146380306;
assign addr[32725]= -2144814157;
assign addr[32726]= -2142567738;
assign addr[32727]= -2139641764;
assign addr[32728]= -2136037160;
assign addr[32729]= -2131755071;
assign addr[32730]= -2126796855;
assign addr[32731]= -2121164085;
assign addr[32732]= -2114858546;
assign addr[32733]= -2107882239;
assign addr[32734]= -2100237377;
assign addr[32735]= -2091926384;
assign addr[32736]= -2082951896;
assign addr[32737]= -2073316760;
assign addr[32738]= -2063024031;
assign addr[32739]= -2052076975;
assign addr[32740]= -2040479063;
assign addr[32741]= -2028233973;
assign addr[32742]= -2015345591;
assign addr[32743]= -2001818002;
assign addr[32744]= -1987655498;
assign addr[32745]= -1972862571;
assign addr[32746]= -1957443913;
assign addr[32747]= -1941404413;
assign addr[32748]= -1924749160;
assign addr[32749]= -1907483436;
assign addr[32750]= -1889612716;
assign addr[32751]= -1871142669;
assign addr[32752]= -1852079154;
assign addr[32753]= -1832428215;
assign addr[32754]= -1812196087;
assign addr[32755]= -1791389186;
assign addr[32756]= -1770014111;
assign addr[32757]= -1748077642;
assign addr[32758]= -1725586737;
assign addr[32759]= -1702548529;
assign addr[32760]= -1678970324;
assign addr[32761]= -1654859602;
assign addr[32762]= -1630224009;
assign addr[32763]= -1605071359;
assign addr[32764]= -1579409630;
assign addr[32765]= -1553246960;
assign addr[32766]= -1526591649;
assign addr[32767]= -1499452149;
assign addr[32768]= -1471837070;
assign addr[32769]= -1443755168;
assign addr[32770]= -1415215352;
assign addr[32771]= -1386226674;
assign addr[32772]= -1356798326;
assign addr[32773]= -1326939644;
assign addr[32774]= -1296660098;
assign addr[32775]= -1265969291;
assign addr[32776]= -1234876957;
assign addr[32777]= -1203392958;
assign addr[32778]= -1171527280;
assign addr[32779]= -1139290029;
assign addr[32780]= -1106691431;
assign addr[32781]= -1073741824;
assign addr[32782]= -1040451659;
assign addr[32783]= -1006831495;
assign addr[32784]= -972891995;
assign addr[32785]= -938643924;
assign addr[32786]= -904098143;
assign addr[32787]= -869265610;
assign addr[32788]= -834157373;
assign addr[32789]= -798784567;
assign addr[32790]= -763158411;
assign addr[32791]= -727290205;
assign addr[32792]= -691191324;
assign addr[32793]= -654873219;
assign addr[32794]= -618347408;
assign addr[32795]= -581625477;
assign addr[32796]= -544719071;
assign addr[32797]= -507639898;
assign addr[32798]= -470399716;
assign addr[32799]= -433010339;
assign addr[32800]= -395483624;
assign addr[32801]= -357831473;
assign addr[32802]= -320065829;
assign addr[32803]= -282198671;
assign addr[32804]= -244242007;
assign addr[32805]= -206207878;
assign addr[32806]= -168108346;
assign addr[32807]= -129955495;
assign addr[32808]= -91761426;
assign addr[32809]= -53538253;
assign addr[32810]= -15298099;
assign addr[32811]= 22946906;
assign addr[32812]= 61184634;
assign addr[32813]= 99402956;
assign addr[32814]= 137589750;
assign addr[32815]= 175732905;
assign addr[32816]= 213820322;
assign addr[32817]= 251839923;
assign addr[32818]= 289779648;
assign addr[32819]= 327627463;
assign addr[32820]= 365371365;
assign addr[32821]= 402999383;
assign addr[32822]= 440499581;
assign addr[32823]= 477860067;
assign addr[32824]= 515068990;
assign addr[32825]= 552114549;
assign addr[32826]= 588984994;
assign addr[32827]= 625668632;
assign addr[32828]= 662153826;
assign addr[32829]= 698429006;
assign addr[32830]= 734482665;
assign addr[32831]= 770303369;
assign addr[32832]= 805879757;
assign addr[32833]= 841200544;
assign addr[32834]= 876254528;
assign addr[32835]= 911030591;
assign addr[32836]= 945517704;
assign addr[32837]= 979704927;
assign addr[32838]= 1013581418;
assign addr[32839]= 1047136432;
assign addr[32840]= 1080359326;
assign addr[32841]= 1113239564;
assign addr[32842]= 1145766716;
assign addr[32843]= 1177930466;
assign addr[32844]= 1209720613;
assign addr[32845]= 1241127074;
assign addr[32846]= 1272139887;
assign addr[32847]= 1302749217;
assign addr[32848]= 1332945355;
assign addr[32849]= 1362718723;
assign addr[32850]= 1392059879;
assign addr[32851]= 1420959516;
assign addr[32852]= 1449408469;
assign addr[32853]= 1477397714;
assign addr[32854]= 1504918373;
assign addr[32855]= 1531961719;
assign addr[32856]= 1558519173;
assign addr[32857]= 1584582314;
assign addr[32858]= 1610142873;
assign addr[32859]= 1635192744;
assign addr[32860]= 1659723983;
assign addr[32861]= 1683728808;
assign addr[32862]= 1707199606;
assign addr[32863]= 1730128933;
assign addr[32864]= 1752509516;
assign addr[32865]= 1774334257;
assign addr[32866]= 1795596234;
assign addr[32867]= 1816288703;
assign addr[32868]= 1836405100;
assign addr[32869]= 1855939047;
assign addr[32870]= 1874884346;
assign addr[32871]= 1893234990;
assign addr[32872]= 1910985158;
assign addr[32873]= 1928129220;
assign addr[32874]= 1944661739;
assign addr[32875]= 1960577471;
assign addr[32876]= 1975871368;
assign addr[32877]= 1990538579;
assign addr[32878]= 2004574453;
assign addr[32879]= 2017974537;
assign addr[32880]= 2030734582;
assign addr[32881]= 2042850540;
assign addr[32882]= 2054318569;
assign addr[32883]= 2065135031;
assign addr[32884]= 2075296495;
assign addr[32885]= 2084799740;
assign addr[32886]= 2093641749;
assign addr[32887]= 2101819720;
assign addr[32888]= 2109331059;
assign addr[32889]= 2116173382;
assign addr[32890]= 2122344521;
assign addr[32891]= 2127842516;
assign addr[32892]= 2132665626;
assign addr[32893]= 2136812319;
assign addr[32894]= 2140281282;
assign addr[32895]= 2143071413;
assign addr[32896]= 2145181827;
assign addr[32897]= 2146611856;
assign addr[32898]= 2147361045;
assign addr[32899]= 2147429158;
assign addr[32900]= 2146816171;
assign addr[32901]= 2145522281;
assign addr[32902]= 2143547897;
assign addr[32903]= 2140893646;
assign addr[32904]= 2137560369;
assign addr[32905]= 2133549123;
assign addr[32906]= 2128861181;
assign addr[32907]= 2123498030;
assign addr[32908]= 2117461370;
assign addr[32909]= 2110753117;
assign addr[32910]= 2103375398;
assign addr[32911]= 2095330553;
assign addr[32912]= 2086621133;
assign addr[32913]= 2077249901;
assign addr[32914]= 2067219829;
assign addr[32915]= 2056534099;
assign addr[32916]= 2045196100;
assign addr[32917]= 2033209426;
assign addr[32918]= 2020577882;
assign addr[32919]= 2007305472;
assign addr[32920]= 1993396407;
assign addr[32921]= 1978855097;
assign addr[32922]= 1963686155;
assign addr[32923]= 1947894393;
assign addr[32924]= 1931484818;
assign addr[32925]= 1914462636;
assign addr[32926]= 1896833245;
assign addr[32927]= 1878602237;
assign addr[32928]= 1859775393;
assign addr[32929]= 1840358687;
assign addr[32930]= 1820358275;
assign addr[32931]= 1799780501;
assign addr[32932]= 1778631892;
assign addr[32933]= 1756919156;
assign addr[32934]= 1734649179;
assign addr[32935]= 1711829025;
assign addr[32936]= 1688465931;
assign addr[32937]= 1664567307;
assign addr[32938]= 1640140734;
assign addr[32939]= 1615193959;
assign addr[32940]= 1589734894;
assign addr[32941]= 1563771613;
assign addr[32942]= 1537312353;
assign addr[32943]= 1510365504;
assign addr[32944]= 1482939614;
assign addr[32945]= 1455043381;
assign addr[32946]= 1426685652;
assign addr[32947]= 1397875423;
assign addr[32948]= 1368621831;
assign addr[32949]= 1338934154;
assign addr[32950]= 1308821808;
assign addr[32951]= 1278294345;
assign addr[32952]= 1247361445;
assign addr[32953]= 1216032921;
assign addr[32954]= 1184318708;
assign addr[32955]= 1152228866;
assign addr[32956]= 1119773573;
assign addr[32957]= 1086963121;
assign addr[32958]= 1053807919;
assign addr[32959]= 1020318481;
assign addr[32960]= 986505429;
assign addr[32961]= 952379488;
assign addr[32962]= 917951481;
assign addr[32963]= 883232329;
assign addr[32964]= 848233042;
assign addr[32965]= 812964722;
assign addr[32966]= 777438554;
assign addr[32967]= 741665807;
assign addr[32968]= 705657826;
assign addr[32969]= 669426032;
assign addr[32970]= 632981917;
assign addr[32971]= 596337040;
assign addr[32972]= 559503022;
assign addr[32973]= 522491548;
assign addr[32974]= 485314355;
assign addr[32975]= 447983235;
assign addr[32976]= 410510029;
assign addr[32977]= 372906622;
assign addr[32978]= 335184940;
assign addr[32979]= 297356948;
assign addr[32980]= 259434643;
assign addr[32981]= 221430054;
assign addr[32982]= 183355234;
assign addr[32983]= 145222259;
assign addr[32984]= 107043224;
assign addr[32985]= 68830239;
assign addr[32986]= 30595422;
assign addr[32987]= -7649098;
assign addr[32988]= -45891193;
assign addr[32989]= -84118732;
assign addr[32990]= -122319591;
assign addr[32991]= -160481654;
assign addr[32992]= -198592817;
assign addr[32993]= -236640993;
assign addr[32994]= -274614114;
assign addr[32995]= -312500135;
assign addr[32996]= -350287041;
assign addr[32997]= -387962847;
assign addr[32998]= -425515602;
assign addr[32999]= -462933398;
assign addr[33000]= -500204365;
assign addr[33001]= -537316682;
assign addr[33002]= -574258580;
assign addr[33003]= -611018340;
assign addr[33004]= -647584304;
assign addr[33005]= -683944874;
assign addr[33006]= -720088517;
assign addr[33007]= -756003771;
assign addr[33008]= -791679244;
assign addr[33009]= -827103620;
assign addr[33010]= -862265664;
assign addr[33011]= -897154224;
assign addr[33012]= -931758235;
assign addr[33013]= -966066720;
assign addr[33014]= -1000068799;
assign addr[33015]= -1033753687;
assign addr[33016]= -1067110699;
assign addr[33017]= -1100129257;
assign addr[33018]= -1132798888;
assign addr[33019]= -1165109230;
assign addr[33020]= -1197050035;
assign addr[33021]= -1228611172;
assign addr[33022]= -1259782632;
assign addr[33023]= -1290554528;
assign addr[33024]= -1320917099;
assign addr[33025]= -1350860716;
assign addr[33026]= -1380375881;
assign addr[33027]= -1409453233;
assign addr[33028]= -1438083551;
assign addr[33029]= -1466257752;
assign addr[33030]= -1493966902;
assign addr[33031]= -1521202211;
assign addr[33032]= -1547955041;
assign addr[33033]= -1574216908;
assign addr[33034]= -1599979481;
assign addr[33035]= -1625234591;
assign addr[33036]= -1649974225;
assign addr[33037]= -1674190539;
assign addr[33038]= -1697875851;
assign addr[33039]= -1721022648;
assign addr[33040]= -1743623590;
assign addr[33041]= -1765671509;
assign addr[33042]= -1787159411;
assign addr[33043]= -1808080480;
assign addr[33044]= -1828428082;
assign addr[33045]= -1848195763;
assign addr[33046]= -1867377253;
assign addr[33047]= -1885966468;
assign addr[33048]= -1903957513;
assign addr[33049]= -1921344681;
assign addr[33050]= -1938122457;
assign addr[33051]= -1954285520;
assign addr[33052]= -1969828744;
assign addr[33053]= -1984747199;
assign addr[33054]= -1999036154;
assign addr[33055]= -2012691075;
assign addr[33056]= -2025707632;
assign addr[33057]= -2038081698;
assign addr[33058]= -2049809346;
assign addr[33059]= -2060886858;
assign addr[33060]= -2071310720;
assign addr[33061]= -2081077626;
assign addr[33062]= -2090184478;
assign addr[33063]= -2098628387;
assign addr[33064]= -2106406677;
assign addr[33065]= -2113516878;
assign addr[33066]= -2119956737;
assign addr[33067]= -2125724211;
assign addr[33068]= -2130817471;
assign addr[33069]= -2135234901;
assign addr[33070]= -2138975100;
assign addr[33071]= -2142036881;
assign addr[33072]= -2144419275;
assign addr[33073]= -2146121524;
assign addr[33074]= -2147143090;
assign addr[33075]= -2147483648;
assign addr[33076]= -2147143090;
assign addr[33077]= -2146121524;
assign addr[33078]= -2144419275;
assign addr[33079]= -2142036881;
assign addr[33080]= -2138975100;
assign addr[33081]= -2135234901;
assign addr[33082]= -2130817471;
assign addr[33083]= -2125724211;
assign addr[33084]= -2119956737;
assign addr[33085]= -2113516878;
assign addr[33086]= -2106406677;
assign addr[33087]= -2098628387;
assign addr[33088]= -2090184478;
assign addr[33089]= -2081077626;
assign addr[33090]= -2071310720;
assign addr[33091]= -2060886858;
assign addr[33092]= -2049809346;
assign addr[33093]= -2038081698;
assign addr[33094]= -2025707632;
assign addr[33095]= -2012691075;
assign addr[33096]= -1999036154;
assign addr[33097]= -1984747199;
assign addr[33098]= -1969828744;
assign addr[33099]= -1954285520;
assign addr[33100]= -1938122457;
assign addr[33101]= -1921344681;
assign addr[33102]= -1903957513;
assign addr[33103]= -1885966468;
assign addr[33104]= -1867377253;
assign addr[33105]= -1848195763;
assign addr[33106]= -1828428082;
assign addr[33107]= -1808080480;
assign addr[33108]= -1787159411;
assign addr[33109]= -1765671509;
assign addr[33110]= -1743623590;
assign addr[33111]= -1721022648;
assign addr[33112]= -1697875851;
assign addr[33113]= -1674190539;
assign addr[33114]= -1649974225;
assign addr[33115]= -1625234591;
assign addr[33116]= -1599979481;
assign addr[33117]= -1574216908;
assign addr[33118]= -1547955041;
assign addr[33119]= -1521202211;
assign addr[33120]= -1493966902;
assign addr[33121]= -1466257752;
assign addr[33122]= -1438083551;
assign addr[33123]= -1409453233;
assign addr[33124]= -1380375881;
assign addr[33125]= -1350860716;
assign addr[33126]= -1320917099;
assign addr[33127]= -1290554528;
assign addr[33128]= -1259782632;
assign addr[33129]= -1228611172;
assign addr[33130]= -1197050035;
assign addr[33131]= -1165109230;
assign addr[33132]= -1132798888;
assign addr[33133]= -1100129257;
assign addr[33134]= -1067110699;
assign addr[33135]= -1033753687;
assign addr[33136]= -1000068799;
assign addr[33137]= -966066720;
assign addr[33138]= -931758235;
assign addr[33139]= -897154224;
assign addr[33140]= -862265664;
assign addr[33141]= -827103620;
assign addr[33142]= -791679244;
assign addr[33143]= -756003771;
assign addr[33144]= -720088517;
assign addr[33145]= -683944874;
assign addr[33146]= -647584304;
assign addr[33147]= -611018340;
assign addr[33148]= -574258580;
assign addr[33149]= -537316682;
assign addr[33150]= -500204365;
assign addr[33151]= -462933398;
assign addr[33152]= -425515602;
assign addr[33153]= -387962847;
assign addr[33154]= -350287041;
assign addr[33155]= -312500135;
assign addr[33156]= -274614114;
assign addr[33157]= -236640993;
assign addr[33158]= -198592817;
assign addr[33159]= -160481654;
assign addr[33160]= -122319591;
assign addr[33161]= -84118732;
assign addr[33162]= -45891193;
assign addr[33163]= -7649098;
assign addr[33164]= 30595422;
assign addr[33165]= 68830239;
assign addr[33166]= 107043224;
assign addr[33167]= 145222259;
assign addr[33168]= 183355234;
assign addr[33169]= 221430054;
assign addr[33170]= 259434643;
assign addr[33171]= 297356948;
assign addr[33172]= 335184940;
assign addr[33173]= 372906622;
assign addr[33174]= 410510029;
assign addr[33175]= 447983235;
assign addr[33176]= 485314355;
assign addr[33177]= 522491548;
assign addr[33178]= 559503022;
assign addr[33179]= 596337040;
assign addr[33180]= 632981917;
assign addr[33181]= 669426032;
assign addr[33182]= 705657826;
assign addr[33183]= 741665807;
assign addr[33184]= 777438554;
assign addr[33185]= 812964722;
assign addr[33186]= 848233042;
assign addr[33187]= 883232329;
assign addr[33188]= 917951481;
assign addr[33189]= 952379488;
assign addr[33190]= 986505429;
assign addr[33191]= 1020318481;
assign addr[33192]= 1053807919;
assign addr[33193]= 1086963121;
assign addr[33194]= 1119773573;
assign addr[33195]= 1152228866;
assign addr[33196]= 1184318708;
assign addr[33197]= 1216032921;
assign addr[33198]= 1247361445;
assign addr[33199]= 1278294345;
assign addr[33200]= 1308821808;
assign addr[33201]= 1338934154;
assign addr[33202]= 1368621831;
assign addr[33203]= 1397875423;
assign addr[33204]= 1426685652;
assign addr[33205]= 1455043381;
assign addr[33206]= 1482939614;
assign addr[33207]= 1510365504;
assign addr[33208]= 1537312353;
assign addr[33209]= 1563771613;
assign addr[33210]= 1589734894;
assign addr[33211]= 1615193959;
assign addr[33212]= 1640140734;
assign addr[33213]= 1664567307;
assign addr[33214]= 1688465931;
assign addr[33215]= 1711829025;
assign addr[33216]= 1734649179;
assign addr[33217]= 1756919156;
assign addr[33218]= 1778631892;
assign addr[33219]= 1799780501;
assign addr[33220]= 1820358275;
assign addr[33221]= 1840358687;
assign addr[33222]= 1859775393;
assign addr[33223]= 1878602237;
assign addr[33224]= 1896833245;
assign addr[33225]= 1914462636;
assign addr[33226]= 1931484818;
assign addr[33227]= 1947894393;
assign addr[33228]= 1963686155;
assign addr[33229]= 1978855097;
assign addr[33230]= 1993396407;
assign addr[33231]= 2007305472;
assign addr[33232]= 2020577882;
assign addr[33233]= 2033209426;
assign addr[33234]= 2045196100;
assign addr[33235]= 2056534099;
assign addr[33236]= 2067219829;
assign addr[33237]= 2077249901;
assign addr[33238]= 2086621133;
assign addr[33239]= 2095330553;
assign addr[33240]= 2103375398;
assign addr[33241]= 2110753117;
assign addr[33242]= 2117461370;
assign addr[33243]= 2123498030;
assign addr[33244]= 2128861181;
assign addr[33245]= 2133549123;
assign addr[33246]= 2137560369;
assign addr[33247]= 2140893646;
assign addr[33248]= 2143547897;
assign addr[33249]= 2145522281;
assign addr[33250]= 2146816171;
assign addr[33251]= 2147429158;
assign addr[33252]= 2147361045;
assign addr[33253]= 2146611856;
assign addr[33254]= 2145181827;
assign addr[33255]= 2143071413;
assign addr[33256]= 2140281282;
assign addr[33257]= 2136812319;
assign addr[33258]= 2132665626;
assign addr[33259]= 2127842516;
assign addr[33260]= 2122344521;
assign addr[33261]= 2116173382;
assign addr[33262]= 2109331059;
assign addr[33263]= 2101819720;
assign addr[33264]= 2093641749;
assign addr[33265]= 2084799740;
assign addr[33266]= 2075296495;
assign addr[33267]= 2065135031;
assign addr[33268]= 2054318569;
assign addr[33269]= 2042850540;
assign addr[33270]= 2030734582;
assign addr[33271]= 2017974537;
assign addr[33272]= 2004574453;
assign addr[33273]= 1990538579;
assign addr[33274]= 1975871368;
assign addr[33275]= 1960577471;
assign addr[33276]= 1944661739;
assign addr[33277]= 1928129220;
assign addr[33278]= 1910985158;
assign addr[33279]= 1893234990;
assign addr[33280]= 1874884346;
assign addr[33281]= 1855939047;
assign addr[33282]= 1836405100;
assign addr[33283]= 1816288703;
assign addr[33284]= 1795596234;
assign addr[33285]= 1774334257;
assign addr[33286]= 1752509516;
assign addr[33287]= 1730128933;
assign addr[33288]= 1707199606;
assign addr[33289]= 1683728808;
assign addr[33290]= 1659723983;
assign addr[33291]= 1635192744;
assign addr[33292]= 1610142873;
assign addr[33293]= 1584582314;
assign addr[33294]= 1558519173;
assign addr[33295]= 1531961719;
assign addr[33296]= 1504918373;
assign addr[33297]= 1477397714;
assign addr[33298]= 1449408469;
assign addr[33299]= 1420959516;
assign addr[33300]= 1392059879;
assign addr[33301]= 1362718723;
assign addr[33302]= 1332945355;
assign addr[33303]= 1302749217;
assign addr[33304]= 1272139887;
assign addr[33305]= 1241127074;
assign addr[33306]= 1209720613;
assign addr[33307]= 1177930466;
assign addr[33308]= 1145766716;
assign addr[33309]= 1113239564;
assign addr[33310]= 1080359326;
assign addr[33311]= 1047136432;
assign addr[33312]= 1013581418;
assign addr[33313]= 979704927;
assign addr[33314]= 945517704;
assign addr[33315]= 911030591;
assign addr[33316]= 876254528;
assign addr[33317]= 841200544;
assign addr[33318]= 805879757;
assign addr[33319]= 770303369;
assign addr[33320]= 734482665;
assign addr[33321]= 698429006;
assign addr[33322]= 662153826;
assign addr[33323]= 625668632;
assign addr[33324]= 588984994;
assign addr[33325]= 552114549;
assign addr[33326]= 515068990;
assign addr[33327]= 477860067;
assign addr[33328]= 440499581;
assign addr[33329]= 402999383;
assign addr[33330]= 365371365;
assign addr[33331]= 327627463;
assign addr[33332]= 289779648;
assign addr[33333]= 251839923;
assign addr[33334]= 213820322;
assign addr[33335]= 175732905;
assign addr[33336]= 137589750;
assign addr[33337]= 99402956;
assign addr[33338]= 61184634;
assign addr[33339]= 22946906;
assign addr[33340]= -15298099;
assign addr[33341]= -53538253;
assign addr[33342]= -91761426;
assign addr[33343]= -129955495;
assign addr[33344]= -168108346;
assign addr[33345]= -206207878;
assign addr[33346]= -244242007;
assign addr[33347]= -282198671;
assign addr[33348]= -320065829;
assign addr[33349]= -357831473;
assign addr[33350]= -395483624;
assign addr[33351]= -433010339;
assign addr[33352]= -470399716;
assign addr[33353]= -507639898;
assign addr[33354]= -544719071;
assign addr[33355]= -581625477;
assign addr[33356]= -618347408;
assign addr[33357]= -654873219;
assign addr[33358]= -691191324;
assign addr[33359]= -727290205;
assign addr[33360]= -763158411;
assign addr[33361]= -798784567;
assign addr[33362]= -834157373;
assign addr[33363]= -869265610;
assign addr[33364]= -904098143;
assign addr[33365]= -938643924;
assign addr[33366]= -972891995;
assign addr[33367]= -1006831495;
assign addr[33368]= -1040451659;
assign addr[33369]= -1073741824;
assign addr[33370]= -1106691431;
assign addr[33371]= -1139290029;
assign addr[33372]= -1171527280;
assign addr[33373]= -1203392958;
assign addr[33374]= -1234876957;
assign addr[33375]= -1265969291;
assign addr[33376]= -1296660098;
assign addr[33377]= -1326939644;
assign addr[33378]= -1356798326;
assign addr[33379]= -1386226674;
assign addr[33380]= -1415215352;
assign addr[33381]= -1443755168;
assign addr[33382]= -1471837070;
assign addr[33383]= -1499452149;
assign addr[33384]= -1526591649;
assign addr[33385]= -1553246960;
assign addr[33386]= -1579409630;
assign addr[33387]= -1605071359;
assign addr[33388]= -1630224009;
assign addr[33389]= -1654859602;
assign addr[33390]= -1678970324;
assign addr[33391]= -1702548529;
assign addr[33392]= -1725586737;
assign addr[33393]= -1748077642;
assign addr[33394]= -1770014111;
assign addr[33395]= -1791389186;
assign addr[33396]= -1812196087;
assign addr[33397]= -1832428215;
assign addr[33398]= -1852079154;
assign addr[33399]= -1871142669;
assign addr[33400]= -1889612716;
assign addr[33401]= -1907483436;
assign addr[33402]= -1924749160;
assign addr[33403]= -1941404413;
assign addr[33404]= -1957443913;
assign addr[33405]= -1972862571;
assign addr[33406]= -1987655498;
assign addr[33407]= -2001818002;
assign addr[33408]= -2015345591;
assign addr[33409]= -2028233973;
assign addr[33410]= -2040479063;
assign addr[33411]= -2052076975;
assign addr[33412]= -2063024031;
assign addr[33413]= -2073316760;
assign addr[33414]= -2082951896;
assign addr[33415]= -2091926384;
assign addr[33416]= -2100237377;
assign addr[33417]= -2107882239;
assign addr[33418]= -2114858546;
assign addr[33419]= -2121164085;
assign addr[33420]= -2126796855;
assign addr[33421]= -2131755071;
assign addr[33422]= -2136037160;
assign addr[33423]= -2139641764;
assign addr[33424]= -2142567738;
assign addr[33425]= -2144814157;
assign addr[33426]= -2146380306;
assign addr[33427]= -2147265689;
assign addr[33428]= -2147470025;
assign addr[33429]= -2146993250;
assign addr[33430]= -2145835515;
assign addr[33431]= -2143997187;
assign addr[33432]= -2141478848;
assign addr[33433]= -2138281298;
assign addr[33434]= -2134405552;
assign addr[33435]= -2129852837;
assign addr[33436]= -2124624598;
assign addr[33437]= -2118722494;
assign addr[33438]= -2112148396;
assign addr[33439]= -2104904390;
assign addr[33440]= -2096992772;
assign addr[33441]= -2088416053;
assign addr[33442]= -2079176953;
assign addr[33443]= -2069278401;
assign addr[33444]= -2058723538;
assign addr[33445]= -2047515711;
assign addr[33446]= -2035658475;
assign addr[33447]= -2023155591;
assign addr[33448]= -2010011024;
assign addr[33449]= -1996228943;
assign addr[33450]= -1981813720;
assign addr[33451]= -1966769926;
assign addr[33452]= -1951102334;
assign addr[33453]= -1934815911;
assign addr[33454]= -1917915825;
assign addr[33455]= -1900407434;
assign addr[33456]= -1882296293;
assign addr[33457]= -1863588145;
assign addr[33458]= -1844288924;
assign addr[33459]= -1824404752;
assign addr[33460]= -1803941934;
assign addr[33461]= -1782906961;
assign addr[33462]= -1761306505;
assign addr[33463]= -1739147417;
assign addr[33464]= -1716436725;
assign addr[33465]= -1693181631;
assign addr[33466]= -1669389513;
assign addr[33467]= -1645067915;
assign addr[33468]= -1620224553;
assign addr[33469]= -1594867305;
assign addr[33470]= -1569004214;
assign addr[33471]= -1542643483;
assign addr[33472]= -1515793473;
assign addr[33473]= -1488462700;
assign addr[33474]= -1460659832;
assign addr[33475]= -1432393688;
assign addr[33476]= -1403673233;
assign addr[33477]= -1374507575;
assign addr[33478]= -1344905966;
assign addr[33479]= -1314877795;
assign addr[33480]= -1284432584;
assign addr[33481]= -1253579991;
assign addr[33482]= -1222329801;
assign addr[33483]= -1190691925;
assign addr[33484]= -1158676398;
assign addr[33485]= -1126293375;
assign addr[33486]= -1093553126;
assign addr[33487]= -1060466036;
assign addr[33488]= -1027042599;
assign addr[33489]= -993293415;
assign addr[33490]= -959229189;
assign addr[33491]= -924860725;
assign addr[33492]= -890198924;
assign addr[33493]= -855254778;
assign addr[33494]= -820039373;
assign addr[33495]= -784563876;
assign addr[33496]= -748839539;
assign addr[33497]= -712877694;
assign addr[33498]= -676689746;
assign addr[33499]= -640287172;
assign addr[33500]= -603681519;
assign addr[33501]= -566884397;
assign addr[33502]= -529907477;
assign addr[33503]= -492762486;
assign addr[33504]= -455461206;
assign addr[33505]= -418015468;
assign addr[33506]= -380437148;
assign addr[33507]= -342738165;
assign addr[33508]= -304930476;
assign addr[33509]= -267026072;
assign addr[33510]= -229036977;
assign addr[33511]= -190975237;
assign addr[33512]= -152852926;
assign addr[33513]= -114682135;
assign addr[33514]= -76474970;
assign addr[33515]= -38243550;
assign addr[33516]= 0;
assign addr[33517]= 38243550;
assign addr[33518]= 76474970;
assign addr[33519]= 114682135;
assign addr[33520]= 152852926;
assign addr[33521]= 190975237;
assign addr[33522]= 229036977;
assign addr[33523]= 267026072;
assign addr[33524]= 304930476;
assign addr[33525]= 342738165;
assign addr[33526]= 380437148;
assign addr[33527]= 418015468;
assign addr[33528]= 455461206;
assign addr[33529]= 492762486;
assign addr[33530]= 529907477;
assign addr[33531]= 566884397;
assign addr[33532]= 603681519;
assign addr[33533]= 640287172;
assign addr[33534]= 676689746;
assign addr[33535]= 712877694;
assign addr[33536]= 748839539;
assign addr[33537]= 784563876;
assign addr[33538]= 820039373;
assign addr[33539]= 855254778;
assign addr[33540]= 890198924;
assign addr[33541]= 924860725;
assign addr[33542]= 959229189;
assign addr[33543]= 993293415;
assign addr[33544]= 1027042599;
assign addr[33545]= 1060466036;
assign addr[33546]= 1093553126;
assign addr[33547]= 1126293375;
assign addr[33548]= 1158676398;
assign addr[33549]= 1190691925;
assign addr[33550]= 1222329801;
assign addr[33551]= 1253579991;
assign addr[33552]= 1284432584;
assign addr[33553]= 1314877795;
assign addr[33554]= 1344905966;
assign addr[33555]= 1374507575;
assign addr[33556]= 1403673233;
assign addr[33557]= 1432393688;
assign addr[33558]= 1460659832;
assign addr[33559]= 1488462700;
assign addr[33560]= 1515793473;
assign addr[33561]= 1542643483;
assign addr[33562]= 1569004214;
assign addr[33563]= 1594867305;
assign addr[33564]= 1620224553;
assign addr[33565]= 1645067915;
assign addr[33566]= 1669389513;
assign addr[33567]= 1693181631;
assign addr[33568]= 1716436725;
assign addr[33569]= 1739147417;
assign addr[33570]= 1761306505;
assign addr[33571]= 1782906961;
assign addr[33572]= 1803941934;
assign addr[33573]= 1824404752;
assign addr[33574]= 1844288924;
assign addr[33575]= 1863588145;
assign addr[33576]= 1882296293;
assign addr[33577]= 1900407434;
assign addr[33578]= 1917915825;
assign addr[33579]= 1934815911;
assign addr[33580]= 1951102334;
assign addr[33581]= 1966769926;
assign addr[33582]= 1981813720;
assign addr[33583]= 1996228943;
assign addr[33584]= 2010011024;
assign addr[33585]= 2023155591;
assign addr[33586]= 2035658475;
assign addr[33587]= 2047515711;
assign addr[33588]= 2058723538;
assign addr[33589]= 2069278401;
assign addr[33590]= 2079176953;
assign addr[33591]= 2088416053;
assign addr[33592]= 2096992772;
assign addr[33593]= 2104904390;
assign addr[33594]= 2112148396;
assign addr[33595]= 2118722494;
assign addr[33596]= 2124624598;
assign addr[33597]= 2129852837;
assign addr[33598]= 2134405552;
assign addr[33599]= 2138281298;
assign addr[33600]= 2141478848;
assign addr[33601]= 2143997187;
assign addr[33602]= 2145835515;
assign addr[33603]= 2146993250;
assign addr[33604]= 2147470025;
assign addr[33605]= 2147265689;
assign addr[33606]= 2146380306;
assign addr[33607]= 2144814157;
assign addr[33608]= 2142567738;
assign addr[33609]= 2139641764;
assign addr[33610]= 2136037160;
assign addr[33611]= 2131755071;
assign addr[33612]= 2126796855;
assign addr[33613]= 2121164085;
assign addr[33614]= 2114858546;
assign addr[33615]= 2107882239;
assign addr[33616]= 2100237377;
assign addr[33617]= 2091926384;
assign addr[33618]= 2082951896;
assign addr[33619]= 2073316760;
assign addr[33620]= 2063024031;
assign addr[33621]= 2052076975;
assign addr[33622]= 2040479063;
assign addr[33623]= 2028233973;
assign addr[33624]= 2015345591;
assign addr[33625]= 2001818002;
assign addr[33626]= 1987655498;
assign addr[33627]= 1972862571;
assign addr[33628]= 1957443913;
assign addr[33629]= 1941404413;
assign addr[33630]= 1924749160;
assign addr[33631]= 1907483436;
assign addr[33632]= 1889612716;
assign addr[33633]= 1871142669;
assign addr[33634]= 1852079154;
assign addr[33635]= 1832428215;
assign addr[33636]= 1812196087;
assign addr[33637]= 1791389186;
assign addr[33638]= 1770014111;
assign addr[33639]= 1748077642;
assign addr[33640]= 1725586737;
assign addr[33641]= 1702548529;
assign addr[33642]= 1678970324;
assign addr[33643]= 1654859602;
assign addr[33644]= 1630224009;
assign addr[33645]= 1605071359;
assign addr[33646]= 1579409630;
assign addr[33647]= 1553246960;
assign addr[33648]= 1526591649;
assign addr[33649]= 1499452149;
assign addr[33650]= 1471837070;
assign addr[33651]= 1443755168;
assign addr[33652]= 1415215352;
assign addr[33653]= 1386226674;
assign addr[33654]= 1356798326;
assign addr[33655]= 1326939644;
assign addr[33656]= 1296660098;
assign addr[33657]= 1265969291;
assign addr[33658]= 1234876957;
assign addr[33659]= 1203392958;
assign addr[33660]= 1171527280;
assign addr[33661]= 1139290029;
assign addr[33662]= 1106691431;
assign addr[33663]= 1073741824;
assign addr[33664]= 1040451659;
assign addr[33665]= 1006831495;
assign addr[33666]= 972891995;
assign addr[33667]= 938643924;
assign addr[33668]= 904098143;
assign addr[33669]= 869265610;
assign addr[33670]= 834157373;
assign addr[33671]= 798784567;
assign addr[33672]= 763158411;
assign addr[33673]= 727290205;
assign addr[33674]= 691191324;
assign addr[33675]= 654873219;
assign addr[33676]= 618347408;
assign addr[33677]= 581625477;
assign addr[33678]= 544719071;
assign addr[33679]= 507639898;
assign addr[33680]= 470399716;
assign addr[33681]= 433010339;
assign addr[33682]= 395483624;
assign addr[33683]= 357831473;
assign addr[33684]= 320065829;
assign addr[33685]= 282198671;
assign addr[33686]= 244242007;
assign addr[33687]= 206207878;
assign addr[33688]= 168108346;
assign addr[33689]= 129955495;
assign addr[33690]= 91761426;
assign addr[33691]= 53538253;
assign addr[33692]= 15298099;
assign addr[33693]= -22946906;
assign addr[33694]= -61184634;
assign addr[33695]= -99402956;
assign addr[33696]= -137589750;
assign addr[33697]= -175732905;
assign addr[33698]= -213820322;
assign addr[33699]= -251839923;
assign addr[33700]= -289779648;
assign addr[33701]= -327627463;
assign addr[33702]= -365371365;
assign addr[33703]= -402999383;
assign addr[33704]= -440499581;
assign addr[33705]= -477860067;
assign addr[33706]= -515068990;
assign addr[33707]= -552114549;
assign addr[33708]= -588984994;
assign addr[33709]= -625668632;
assign addr[33710]= -662153826;
assign addr[33711]= -698429006;
assign addr[33712]= -734482665;
assign addr[33713]= -770303369;
assign addr[33714]= -805879757;
assign addr[33715]= -841200544;
assign addr[33716]= -876254528;
assign addr[33717]= -911030591;
assign addr[33718]= -945517704;
assign addr[33719]= -979704927;
assign addr[33720]= -1013581418;
assign addr[33721]= -1047136432;
assign addr[33722]= -1080359326;
assign addr[33723]= -1113239564;
assign addr[33724]= -1145766716;
assign addr[33725]= -1177930466;
assign addr[33726]= -1209720613;
assign addr[33727]= -1241127074;
assign addr[33728]= -1272139887;
assign addr[33729]= -1302749217;
assign addr[33730]= -1332945355;
assign addr[33731]= -1362718723;
assign addr[33732]= -1392059879;
assign addr[33733]= -1420959516;
assign addr[33734]= -1449408469;
assign addr[33735]= -1477397714;
assign addr[33736]= -1504918373;
assign addr[33737]= -1531961719;
assign addr[33738]= -1558519173;
assign addr[33739]= -1584582314;
assign addr[33740]= -1610142873;
assign addr[33741]= -1635192744;
assign addr[33742]= -1659723983;
assign addr[33743]= -1683728808;
assign addr[33744]= -1707199606;
assign addr[33745]= -1730128933;
assign addr[33746]= -1752509516;
assign addr[33747]= -1774334257;
assign addr[33748]= -1795596234;
assign addr[33749]= -1816288703;
assign addr[33750]= -1836405100;
assign addr[33751]= -1855939047;
assign addr[33752]= -1874884346;
assign addr[33753]= -1893234990;
assign addr[33754]= -1910985158;
assign addr[33755]= -1928129220;
assign addr[33756]= -1944661739;
assign addr[33757]= -1960577471;
assign addr[33758]= -1975871368;
assign addr[33759]= -1990538579;
assign addr[33760]= -2004574453;
assign addr[33761]= -2017974537;
assign addr[33762]= -2030734582;
assign addr[33763]= -2042850540;
assign addr[33764]= -2054318569;
assign addr[33765]= -2065135031;
assign addr[33766]= -2075296495;
assign addr[33767]= -2084799740;
assign addr[33768]= -2093641749;
assign addr[33769]= -2101819720;
assign addr[33770]= -2109331059;
assign addr[33771]= -2116173382;
assign addr[33772]= -2122344521;
assign addr[33773]= -2127842516;
assign addr[33774]= -2132665626;
assign addr[33775]= -2136812319;
assign addr[33776]= -2140281282;
assign addr[33777]= -2143071413;
assign addr[33778]= -2145181827;
assign addr[33779]= -2146611856;
assign addr[33780]= -2147361045;
assign addr[33781]= -2147429158;
assign addr[33782]= -2146816171;
assign addr[33783]= -2145522281;
assign addr[33784]= -2143547897;
assign addr[33785]= -2140893646;
assign addr[33786]= -2137560369;
assign addr[33787]= -2133549123;
assign addr[33788]= -2128861181;
assign addr[33789]= -2123498030;
assign addr[33790]= -2117461370;
assign addr[33791]= -2110753117;
assign addr[33792]= -2103375398;
assign addr[33793]= -2095330553;
assign addr[33794]= -2086621133;
assign addr[33795]= -2077249901;
assign addr[33796]= -2067219829;
assign addr[33797]= -2056534099;
assign addr[33798]= -2045196100;
assign addr[33799]= -2033209426;
assign addr[33800]= -2020577882;
assign addr[33801]= -2007305472;
assign addr[33802]= -1993396407;
assign addr[33803]= -1978855097;
assign addr[33804]= -1963686155;
assign addr[33805]= -1947894393;
assign addr[33806]= -1931484818;
assign addr[33807]= -1914462636;
assign addr[33808]= -1896833245;
assign addr[33809]= -1878602237;
assign addr[33810]= -1859775393;
assign addr[33811]= -1840358687;
assign addr[33812]= -1820358275;
assign addr[33813]= -1799780501;
assign addr[33814]= -1778631892;
assign addr[33815]= -1756919156;
assign addr[33816]= -1734649179;
assign addr[33817]= -1711829025;
assign addr[33818]= -1688465931;
assign addr[33819]= -1664567307;
assign addr[33820]= -1640140734;
assign addr[33821]= -1615193959;
assign addr[33822]= -1589734894;
assign addr[33823]= -1563771613;
assign addr[33824]= -1537312353;
assign addr[33825]= -1510365504;
assign addr[33826]= -1482939614;
assign addr[33827]= -1455043381;
assign addr[33828]= -1426685652;
assign addr[33829]= -1397875423;
assign addr[33830]= -1368621831;
assign addr[33831]= -1338934154;
assign addr[33832]= -1308821808;
assign addr[33833]= -1278294345;
assign addr[33834]= -1247361445;
assign addr[33835]= -1216032921;
assign addr[33836]= -1184318708;
assign addr[33837]= -1152228866;
assign addr[33838]= -1119773573;
assign addr[33839]= -1086963121;
assign addr[33840]= -1053807919;
assign addr[33841]= -1020318481;
assign addr[33842]= -986505429;
assign addr[33843]= -952379488;
assign addr[33844]= -917951481;
assign addr[33845]= -883232329;
assign addr[33846]= -848233042;
assign addr[33847]= -812964722;
assign addr[33848]= -777438554;
assign addr[33849]= -741665807;
assign addr[33850]= -705657826;
assign addr[33851]= -669426032;
assign addr[33852]= -632981917;
assign addr[33853]= -596337040;
assign addr[33854]= -559503022;
assign addr[33855]= -522491548;
assign addr[33856]= -485314355;
assign addr[33857]= -447983235;
assign addr[33858]= -410510029;
assign addr[33859]= -372906622;
assign addr[33860]= -335184940;
assign addr[33861]= -297356948;
assign addr[33862]= -259434643;
assign addr[33863]= -221430054;
assign addr[33864]= -183355234;
assign addr[33865]= -145222259;
assign addr[33866]= -107043224;
assign addr[33867]= -68830239;
assign addr[33868]= -30595422;
assign addr[33869]= 7649098;
assign addr[33870]= 45891193;
assign addr[33871]= 84118732;
assign addr[33872]= 122319591;
assign addr[33873]= 160481654;
assign addr[33874]= 198592817;
assign addr[33875]= 236640993;
assign addr[33876]= 274614114;
assign addr[33877]= 312500135;
assign addr[33878]= 350287041;
assign addr[33879]= 387962847;
assign addr[33880]= 425515602;
assign addr[33881]= 462933398;
assign addr[33882]= 500204365;
assign addr[33883]= 537316682;
assign addr[33884]= 574258580;
assign addr[33885]= 611018340;
assign addr[33886]= 647584304;
assign addr[33887]= 683944874;
assign addr[33888]= 720088517;
assign addr[33889]= 756003771;
assign addr[33890]= 791679244;
assign addr[33891]= 827103620;
assign addr[33892]= 862265664;
assign addr[33893]= 897154224;
assign addr[33894]= 931758235;
assign addr[33895]= 966066720;
assign addr[33896]= 1000068799;
assign addr[33897]= 1033753687;
assign addr[33898]= 1067110699;
assign addr[33899]= 1100129257;
assign addr[33900]= 1132798888;
assign addr[33901]= 1165109230;
assign addr[33902]= 1197050035;
assign addr[33903]= 1228611172;
assign addr[33904]= 1259782632;
assign addr[33905]= 1290554528;
assign addr[33906]= 1320917099;
assign addr[33907]= 1350860716;
assign addr[33908]= 1380375881;
assign addr[33909]= 1409453233;
assign addr[33910]= 1438083551;
assign addr[33911]= 1466257752;
assign addr[33912]= 1493966902;
assign addr[33913]= 1521202211;
assign addr[33914]= 1547955041;
assign addr[33915]= 1574216908;
assign addr[33916]= 1599979481;
assign addr[33917]= 1625234591;
assign addr[33918]= 1649974225;
assign addr[33919]= 1674190539;
assign addr[33920]= 1697875851;
assign addr[33921]= 1721022648;
assign addr[33922]= 1743623590;
assign addr[33923]= 1765671509;
assign addr[33924]= 1787159411;
assign addr[33925]= 1808080480;
assign addr[33926]= 1828428082;
assign addr[33927]= 1848195763;
assign addr[33928]= 1867377253;
assign addr[33929]= 1885966468;
assign addr[33930]= 1903957513;
assign addr[33931]= 1921344681;
assign addr[33932]= 1938122457;
assign addr[33933]= 1954285520;
assign addr[33934]= 1969828744;
assign addr[33935]= 1984747199;
assign addr[33936]= 1999036154;
assign addr[33937]= 2012691075;
assign addr[33938]= 2025707632;
assign addr[33939]= 2038081698;
assign addr[33940]= 2049809346;
assign addr[33941]= 2060886858;
assign addr[33942]= 2071310720;
assign addr[33943]= 2081077626;
assign addr[33944]= 2090184478;
assign addr[33945]= 2098628387;
assign addr[33946]= 2106406677;
assign addr[33947]= 2113516878;
assign addr[33948]= 2119956737;
assign addr[33949]= 2125724211;
assign addr[33950]= 2130817471;
assign addr[33951]= 2135234901;
assign addr[33952]= 2138975100;
assign addr[33953]= 2142036881;
assign addr[33954]= 2144419275;
assign addr[33955]= 2146121524;
assign addr[33956]= 2147143090;
assign addr[33957]= 2147483648;
assign addr[33958]= 2147143090;
assign addr[33959]= 2146121524;
assign addr[33960]= 2144419275;
assign addr[33961]= 2142036881;
assign addr[33962]= 2138975100;
assign addr[33963]= 2135234901;
assign addr[33964]= 2130817471;
assign addr[33965]= 2125724211;
assign addr[33966]= 2119956737;
assign addr[33967]= 2113516878;
assign addr[33968]= 2106406677;
assign addr[33969]= 2098628387;
assign addr[33970]= 2090184478;
assign addr[33971]= 2081077626;
assign addr[33972]= 2071310720;
assign addr[33973]= 2060886858;
assign addr[33974]= 2049809346;
assign addr[33975]= 2038081698;
assign addr[33976]= 2025707632;
assign addr[33977]= 2012691075;
assign addr[33978]= 1999036154;
assign addr[33979]= 1984747199;
assign addr[33980]= 1969828744;
assign addr[33981]= 1954285520;
assign addr[33982]= 1938122457;
assign addr[33983]= 1921344681;
assign addr[33984]= 1903957513;
assign addr[33985]= 1885966468;
assign addr[33986]= 1867377253;
assign addr[33987]= 1848195763;
assign addr[33988]= 1828428082;
assign addr[33989]= 1808080480;
assign addr[33990]= 1787159411;
assign addr[33991]= 1765671509;
assign addr[33992]= 1743623590;
assign addr[33993]= 1721022648;
assign addr[33994]= 1697875851;
assign addr[33995]= 1674190539;
assign addr[33996]= 1649974225;
assign addr[33997]= 1625234591;
assign addr[33998]= 1599979481;
assign addr[33999]= 1574216908;
assign addr[34000]= 1547955041;
assign addr[34001]= 1521202211;
assign addr[34002]= 1493966902;
assign addr[34003]= 1466257752;
assign addr[34004]= 1438083551;
assign addr[34005]= 1409453233;
assign addr[34006]= 1380375881;
assign addr[34007]= 1350860716;
assign addr[34008]= 1320917099;
assign addr[34009]= 1290554528;
assign addr[34010]= 1259782632;
assign addr[34011]= 1228611172;
assign addr[34012]= 1197050035;
assign addr[34013]= 1165109230;
assign addr[34014]= 1132798888;
assign addr[34015]= 1100129257;
assign addr[34016]= 1067110699;
assign addr[34017]= 1033753687;
assign addr[34018]= 1000068799;
assign addr[34019]= 966066720;
assign addr[34020]= 931758235;
assign addr[34021]= 897154224;
assign addr[34022]= 862265664;
assign addr[34023]= 827103620;
assign addr[34024]= 791679244;
assign addr[34025]= 756003771;
assign addr[34026]= 720088517;
assign addr[34027]= 683944874;
assign addr[34028]= 647584304;
assign addr[34029]= 611018340;
assign addr[34030]= 574258580;
assign addr[34031]= 537316682;
assign addr[34032]= 500204365;
assign addr[34033]= 462933398;
assign addr[34034]= 425515602;
assign addr[34035]= 387962847;
assign addr[34036]= 350287041;
assign addr[34037]= 312500135;
assign addr[34038]= 274614114;
assign addr[34039]= 236640993;
assign addr[34040]= 198592817;
assign addr[34041]= 160481654;
assign addr[34042]= 122319591;
assign addr[34043]= 84118732;
assign addr[34044]= 45891193;
assign addr[34045]= 7649098;
assign addr[34046]= -30595422;
assign addr[34047]= -68830239;
assign addr[34048]= -107043224;
assign addr[34049]= -145222259;
assign addr[34050]= -183355234;
assign addr[34051]= -221430054;
assign addr[34052]= -259434643;
assign addr[34053]= -297356948;
assign addr[34054]= -335184940;
assign addr[34055]= -372906622;
assign addr[34056]= -410510029;
assign addr[34057]= -447983235;
assign addr[34058]= -485314355;
assign addr[34059]= -522491548;
assign addr[34060]= -559503022;
assign addr[34061]= -596337040;
assign addr[34062]= -632981917;
assign addr[34063]= -669426032;
assign addr[34064]= -705657826;
assign addr[34065]= -741665807;
assign addr[34066]= -777438554;
assign addr[34067]= -812964722;
assign addr[34068]= -848233042;
assign addr[34069]= -883232329;
assign addr[34070]= -917951481;
assign addr[34071]= -952379488;
assign addr[34072]= -986505429;
assign addr[34073]= -1020318481;
assign addr[34074]= -1053807919;
assign addr[34075]= -1086963121;
assign addr[34076]= -1119773573;
assign addr[34077]= -1152228866;
assign addr[34078]= -1184318708;
assign addr[34079]= -1216032921;
assign addr[34080]= -1247361445;
assign addr[34081]= -1278294345;
assign addr[34082]= -1308821808;
assign addr[34083]= -1338934154;
assign addr[34084]= -1368621831;
assign addr[34085]= -1397875423;
assign addr[34086]= -1426685652;
assign addr[34087]= -1455043381;
assign addr[34088]= -1482939614;
assign addr[34089]= -1510365504;
assign addr[34090]= -1537312353;
assign addr[34091]= -1563771613;
assign addr[34092]= -1589734894;
assign addr[34093]= -1615193959;
assign addr[34094]= -1640140734;
assign addr[34095]= -1664567307;
assign addr[34096]= -1688465931;
assign addr[34097]= -1711829025;
assign addr[34098]= -1734649179;
assign addr[34099]= -1756919156;
assign addr[34100]= -1778631892;
assign addr[34101]= -1799780501;
assign addr[34102]= -1820358275;
assign addr[34103]= -1840358687;
assign addr[34104]= -1859775393;
assign addr[34105]= -1878602237;
assign addr[34106]= -1896833245;
assign addr[34107]= -1914462636;
assign addr[34108]= -1931484818;
assign addr[34109]= -1947894393;
assign addr[34110]= -1963686155;
assign addr[34111]= -1978855097;
assign addr[34112]= -1993396407;
assign addr[34113]= -2007305472;
assign addr[34114]= -2020577882;
assign addr[34115]= -2033209426;
assign addr[34116]= -2045196100;
assign addr[34117]= -2056534099;
assign addr[34118]= -2067219829;
assign addr[34119]= -2077249901;
assign addr[34120]= -2086621133;
assign addr[34121]= -2095330553;
assign addr[34122]= -2103375398;
assign addr[34123]= -2110753117;
assign addr[34124]= -2117461370;
assign addr[34125]= -2123498030;
assign addr[34126]= -2128861181;
assign addr[34127]= -2133549123;
assign addr[34128]= -2137560369;
assign addr[34129]= -2140893646;
assign addr[34130]= -2143547897;
assign addr[34131]= -2145522281;
assign addr[34132]= -2146816171;
assign addr[34133]= -2147429158;
assign addr[34134]= -2147361045;
assign addr[34135]= -2146611856;
assign addr[34136]= -2145181827;
assign addr[34137]= -2143071413;
assign addr[34138]= -2140281282;
assign addr[34139]= -2136812319;
assign addr[34140]= -2132665626;
assign addr[34141]= -2127842516;
assign addr[34142]= -2122344521;
assign addr[34143]= -2116173382;
assign addr[34144]= -2109331059;
assign addr[34145]= -2101819720;
assign addr[34146]= -2093641749;
assign addr[34147]= -2084799740;
assign addr[34148]= -2075296495;
assign addr[34149]= -2065135031;
assign addr[34150]= -2054318569;
assign addr[34151]= -2042850540;
assign addr[34152]= -2030734582;
assign addr[34153]= -2017974537;
assign addr[34154]= -2004574453;
assign addr[34155]= -1990538579;
assign addr[34156]= -1975871368;
assign addr[34157]= -1960577471;
assign addr[34158]= -1944661739;
assign addr[34159]= -1928129220;
assign addr[34160]= -1910985158;
assign addr[34161]= -1893234990;
assign addr[34162]= -1874884346;
assign addr[34163]= -1855939047;
assign addr[34164]= -1836405100;
assign addr[34165]= -1816288703;
assign addr[34166]= -1795596234;
assign addr[34167]= -1774334257;
assign addr[34168]= -1752509516;
assign addr[34169]= -1730128933;
assign addr[34170]= -1707199606;
assign addr[34171]= -1683728808;
assign addr[34172]= -1659723983;
assign addr[34173]= -1635192744;
assign addr[34174]= -1610142873;
assign addr[34175]= -1584582314;
assign addr[34176]= -1558519173;
assign addr[34177]= -1531961719;
assign addr[34178]= -1504918373;
assign addr[34179]= -1477397714;
assign addr[34180]= -1449408469;
assign addr[34181]= -1420959516;
assign addr[34182]= -1392059879;
assign addr[34183]= -1362718723;
assign addr[34184]= -1332945355;
assign addr[34185]= -1302749217;
assign addr[34186]= -1272139887;
assign addr[34187]= -1241127074;
assign addr[34188]= -1209720613;
assign addr[34189]= -1177930466;
assign addr[34190]= -1145766716;
assign addr[34191]= -1113239564;
assign addr[34192]= -1080359326;
assign addr[34193]= -1047136432;
assign addr[34194]= -1013581418;
assign addr[34195]= -979704927;
assign addr[34196]= -945517704;
assign addr[34197]= -911030591;
assign addr[34198]= -876254528;
assign addr[34199]= -841200544;
assign addr[34200]= -805879757;
assign addr[34201]= -770303369;
assign addr[34202]= -734482665;
assign addr[34203]= -698429006;
assign addr[34204]= -662153826;
assign addr[34205]= -625668632;
assign addr[34206]= -588984994;
assign addr[34207]= -552114549;
assign addr[34208]= -515068990;
assign addr[34209]= -477860067;
assign addr[34210]= -440499581;
assign addr[34211]= -402999383;
assign addr[34212]= -365371365;
assign addr[34213]= -327627463;
assign addr[34214]= -289779648;
assign addr[34215]= -251839923;
assign addr[34216]= -213820322;
assign addr[34217]= -175732905;
assign addr[34218]= -137589750;
assign addr[34219]= -99402956;
assign addr[34220]= -61184634;
assign addr[34221]= -22946906;
assign addr[34222]= 15298099;
assign addr[34223]= 53538253;
assign addr[34224]= 91761426;
assign addr[34225]= 129955495;
assign addr[34226]= 168108346;
assign addr[34227]= 206207878;
assign addr[34228]= 244242007;
assign addr[34229]= 282198671;
assign addr[34230]= 320065829;
assign addr[34231]= 357831473;
assign addr[34232]= 395483624;
assign addr[34233]= 433010339;
assign addr[34234]= 470399716;
assign addr[34235]= 507639898;
assign addr[34236]= 544719071;
assign addr[34237]= 581625477;
assign addr[34238]= 618347408;
assign addr[34239]= 654873219;
assign addr[34240]= 691191324;
assign addr[34241]= 727290205;
assign addr[34242]= 763158411;
assign addr[34243]= 798784567;
assign addr[34244]= 834157373;
assign addr[34245]= 869265610;
assign addr[34246]= 904098143;
assign addr[34247]= 938643924;
assign addr[34248]= 972891995;
assign addr[34249]= 1006831495;
assign addr[34250]= 1040451659;
assign addr[34251]= 1073741824;
assign addr[34252]= 1106691431;
assign addr[34253]= 1139290029;
assign addr[34254]= 1171527280;
assign addr[34255]= 1203392958;
assign addr[34256]= 1234876957;
assign addr[34257]= 1265969291;
assign addr[34258]= 1296660098;
assign addr[34259]= 1326939644;
assign addr[34260]= 1356798326;
assign addr[34261]= 1386226674;
assign addr[34262]= 1415215352;
assign addr[34263]= 1443755168;
assign addr[34264]= 1471837070;
assign addr[34265]= 1499452149;
assign addr[34266]= 1526591649;
assign addr[34267]= 1553246960;
assign addr[34268]= 1579409630;
assign addr[34269]= 1605071359;
assign addr[34270]= 1630224009;
assign addr[34271]= 1654859602;
assign addr[34272]= 1678970324;
assign addr[34273]= 1702548529;
assign addr[34274]= 1725586737;
assign addr[34275]= 1748077642;
assign addr[34276]= 1770014111;
assign addr[34277]= 1791389186;
assign addr[34278]= 1812196087;
assign addr[34279]= 1832428215;
assign addr[34280]= 1852079154;
assign addr[34281]= 1871142669;
assign addr[34282]= 1889612716;
assign addr[34283]= 1907483436;
assign addr[34284]= 1924749160;
assign addr[34285]= 1941404413;
assign addr[34286]= 1957443913;
assign addr[34287]= 1972862571;
assign addr[34288]= 1987655498;
assign addr[34289]= 2001818002;
assign addr[34290]= 2015345591;
assign addr[34291]= 2028233973;
assign addr[34292]= 2040479063;
assign addr[34293]= 2052076975;
assign addr[34294]= 2063024031;
assign addr[34295]= 2073316760;
assign addr[34296]= 2082951896;
assign addr[34297]= 2091926384;
assign addr[34298]= 2100237377;
assign addr[34299]= 2107882239;
assign addr[34300]= 2114858546;
assign addr[34301]= 2121164085;
assign addr[34302]= 2126796855;
assign addr[34303]= 2131755071;
assign addr[34304]= 2136037160;
assign addr[34305]= 2139641764;
assign addr[34306]= 2142567738;
assign addr[34307]= 2144814157;
assign addr[34308]= 2146380306;
assign addr[34309]= 2147265689;
assign addr[34310]= 2147470025;
assign addr[34311]= 2146993250;
assign addr[34312]= 2145835515;
assign addr[34313]= 2143997187;
assign addr[34314]= 2141478848;
assign addr[34315]= 2138281298;
assign addr[34316]= 2134405552;
assign addr[34317]= 2129852837;
assign addr[34318]= 2124624598;
assign addr[34319]= 2118722494;
assign addr[34320]= 2112148396;
assign addr[34321]= 2104904390;
assign addr[34322]= 2096992772;
assign addr[34323]= 2088416053;
assign addr[34324]= 2079176953;
assign addr[34325]= 2069278401;
assign addr[34326]= 2058723538;
assign addr[34327]= 2047515711;
assign addr[34328]= 2035658475;
assign addr[34329]= 2023155591;
assign addr[34330]= 2010011024;
assign addr[34331]= 1996228943;
assign addr[34332]= 1981813720;
assign addr[34333]= 1966769926;
assign addr[34334]= 1951102334;
assign addr[34335]= 1934815911;
assign addr[34336]= 1917915825;
assign addr[34337]= 1900407434;
assign addr[34338]= 1882296293;
assign addr[34339]= 1863588145;
assign addr[34340]= 1844288924;
assign addr[34341]= 1824404752;
assign addr[34342]= 1803941934;
assign addr[34343]= 1782906961;
assign addr[34344]= 1761306505;
assign addr[34345]= 1739147417;
assign addr[34346]= 1716436725;
assign addr[34347]= 1693181631;
assign addr[34348]= 1669389513;
assign addr[34349]= 1645067915;
assign addr[34350]= 1620224553;
assign addr[34351]= 1594867305;
assign addr[34352]= 1569004214;
assign addr[34353]= 1542643483;
assign addr[34354]= 1515793473;
assign addr[34355]= 1488462700;
assign addr[34356]= 1460659832;
assign addr[34357]= 1432393688;
assign addr[34358]= 1403673233;
assign addr[34359]= 1374507575;
assign addr[34360]= 1344905966;
assign addr[34361]= 1314877795;
assign addr[34362]= 1284432584;
assign addr[34363]= 1253579991;
assign addr[34364]= 1222329801;
assign addr[34365]= 1190691925;
assign addr[34366]= 1158676398;
assign addr[34367]= 1126293375;
assign addr[34368]= 1093553126;
assign addr[34369]= 1060466036;
assign addr[34370]= 1027042599;
assign addr[34371]= 993293415;
assign addr[34372]= 959229189;
assign addr[34373]= 924860725;
assign addr[34374]= 890198924;
assign addr[34375]= 855254778;
assign addr[34376]= 820039373;
assign addr[34377]= 784563876;
assign addr[34378]= 748839539;
assign addr[34379]= 712877694;
assign addr[34380]= 676689746;
assign addr[34381]= 640287172;
assign addr[34382]= 603681519;
assign addr[34383]= 566884397;
assign addr[34384]= 529907477;
assign addr[34385]= 492762486;
assign addr[34386]= 455461206;
assign addr[34387]= 418015468;
assign addr[34388]= 380437148;
assign addr[34389]= 342738165;
assign addr[34390]= 304930476;
assign addr[34391]= 267026072;
assign addr[34392]= 229036977;
assign addr[34393]= 190975237;
assign addr[34394]= 152852926;
assign addr[34395]= 114682135;
assign addr[34396]= 76474970;
assign addr[34397]= 38243550;
assign addr[34398]= 0;
assign addr[34399]= -38243550;
assign addr[34400]= -76474970;
assign addr[34401]= -114682135;
assign addr[34402]= -152852926;
assign addr[34403]= -190975237;
assign addr[34404]= -229036977;
assign addr[34405]= -267026072;
assign addr[34406]= -304930476;
assign addr[34407]= -342738165;
assign addr[34408]= -380437148;
assign addr[34409]= -418015468;
assign addr[34410]= -455461206;
assign addr[34411]= -492762486;
assign addr[34412]= -529907477;
assign addr[34413]= -566884397;
assign addr[34414]= -603681519;
assign addr[34415]= -640287172;
assign addr[34416]= -676689746;
assign addr[34417]= -712877694;
assign addr[34418]= -748839539;
assign addr[34419]= -784563876;
assign addr[34420]= -820039373;
assign addr[34421]= -855254778;
assign addr[34422]= -890198924;
assign addr[34423]= -924860725;
assign addr[34424]= -959229189;
assign addr[34425]= -993293415;
assign addr[34426]= -1027042599;
assign addr[34427]= -1060466036;
assign addr[34428]= -1093553126;
assign addr[34429]= -1126293375;
assign addr[34430]= -1158676398;
assign addr[34431]= -1190691925;
assign addr[34432]= -1222329801;
assign addr[34433]= -1253579991;
assign addr[34434]= -1284432584;
assign addr[34435]= -1314877795;
assign addr[34436]= -1344905966;
assign addr[34437]= -1374507575;
assign addr[34438]= -1403673233;
assign addr[34439]= -1432393688;
assign addr[34440]= -1460659832;
assign addr[34441]= -1488462700;
assign addr[34442]= -1515793473;
assign addr[34443]= -1542643483;
assign addr[34444]= -1569004214;
assign addr[34445]= -1594867305;
assign addr[34446]= -1620224553;
assign addr[34447]= -1645067915;
assign addr[34448]= -1669389513;
assign addr[34449]= -1693181631;
assign addr[34450]= -1716436725;
assign addr[34451]= -1739147417;
assign addr[34452]= -1761306505;
assign addr[34453]= -1782906961;
assign addr[34454]= -1803941934;
assign addr[34455]= -1824404752;
assign addr[34456]= -1844288924;
assign addr[34457]= -1863588145;
assign addr[34458]= -1882296293;
assign addr[34459]= -1900407434;
assign addr[34460]= -1917915825;
assign addr[34461]= -1934815911;
assign addr[34462]= -1951102334;
assign addr[34463]= -1966769926;
assign addr[34464]= -1981813720;
assign addr[34465]= -1996228943;
assign addr[34466]= -2010011024;
assign addr[34467]= -2023155591;
assign addr[34468]= -2035658475;
assign addr[34469]= -2047515711;
assign addr[34470]= -2058723538;
assign addr[34471]= -2069278401;
assign addr[34472]= -2079176953;
assign addr[34473]= -2088416053;
assign addr[34474]= -2096992772;
assign addr[34475]= -2104904390;
assign addr[34476]= -2112148396;
assign addr[34477]= -2118722494;
assign addr[34478]= -2124624598;
assign addr[34479]= -2129852837;
assign addr[34480]= -2134405552;
assign addr[34481]= -2138281298;
assign addr[34482]= -2141478848;
assign addr[34483]= -2143997187;
assign addr[34484]= -2145835515;
assign addr[34485]= -2146993250;
assign addr[34486]= -2147470025;
assign addr[34487]= -2147265689;
assign addr[34488]= -2146380306;
assign addr[34489]= -2144814157;
assign addr[34490]= -2142567738;
assign addr[34491]= -2139641764;
assign addr[34492]= -2136037160;
assign addr[34493]= -2131755071;
assign addr[34494]= -2126796855;
assign addr[34495]= -2121164085;
assign addr[34496]= -2114858546;
assign addr[34497]= -2107882239;
assign addr[34498]= -2100237377;
assign addr[34499]= -2091926384;
assign addr[34500]= -2082951896;
assign addr[34501]= -2073316760;
assign addr[34502]= -2063024031;
assign addr[34503]= -2052076975;
assign addr[34504]= -2040479063;
assign addr[34505]= -2028233973;
assign addr[34506]= -2015345591;
assign addr[34507]= -2001818002;
assign addr[34508]= -1987655498;
assign addr[34509]= -1972862571;
assign addr[34510]= -1957443913;
assign addr[34511]= -1941404413;
assign addr[34512]= -1924749160;
assign addr[34513]= -1907483436;
assign addr[34514]= -1889612716;
assign addr[34515]= -1871142669;
assign addr[34516]= -1852079154;
assign addr[34517]= -1832428215;
assign addr[34518]= -1812196087;
assign addr[34519]= -1791389186;
assign addr[34520]= -1770014111;
assign addr[34521]= -1748077642;
assign addr[34522]= -1725586737;
assign addr[34523]= -1702548529;
assign addr[34524]= -1678970324;
assign addr[34525]= -1654859602;
assign addr[34526]= -1630224009;
assign addr[34527]= -1605071359;
assign addr[34528]= -1579409630;
assign addr[34529]= -1553246960;
assign addr[34530]= -1526591649;
assign addr[34531]= -1499452149;
assign addr[34532]= -1471837070;
assign addr[34533]= -1443755168;
assign addr[34534]= -1415215352;
assign addr[34535]= -1386226674;
assign addr[34536]= -1356798326;
assign addr[34537]= -1326939644;
assign addr[34538]= -1296660098;
assign addr[34539]= -1265969291;
assign addr[34540]= -1234876957;
assign addr[34541]= -1203392958;
assign addr[34542]= -1171527280;
assign addr[34543]= -1139290029;
assign addr[34544]= -1106691431;
assign addr[34545]= -1073741824;
assign addr[34546]= -1040451659;
assign addr[34547]= -1006831495;
assign addr[34548]= -972891995;
assign addr[34549]= -938643924;
assign addr[34550]= -904098143;
assign addr[34551]= -869265610;
assign addr[34552]= -834157373;
assign addr[34553]= -798784567;
assign addr[34554]= -763158411;
assign addr[34555]= -727290205;
assign addr[34556]= -691191324;
assign addr[34557]= -654873219;
assign addr[34558]= -618347408;
assign addr[34559]= -581625477;
assign addr[34560]= -544719071;
assign addr[34561]= -507639898;
assign addr[34562]= -470399716;
assign addr[34563]= -433010339;
assign addr[34564]= -395483624;
assign addr[34565]= -357831473;
assign addr[34566]= -320065829;
assign addr[34567]= -282198671;
assign addr[34568]= -244242007;
assign addr[34569]= -206207878;
assign addr[34570]= -168108346;
assign addr[34571]= -129955495;
assign addr[34572]= -91761426;
assign addr[34573]= -53538253;
assign addr[34574]= -15298099;
assign addr[34575]= 22946906;
assign addr[34576]= 61184634;
assign addr[34577]= 99402956;
assign addr[34578]= 137589750;
assign addr[34579]= 175732905;
assign addr[34580]= 213820322;
assign addr[34581]= 251839923;
assign addr[34582]= 289779648;
assign addr[34583]= 327627463;
assign addr[34584]= 365371365;
assign addr[34585]= 402999383;
assign addr[34586]= 440499581;
assign addr[34587]= 477860067;
assign addr[34588]= 515068990;
assign addr[34589]= 552114549;
assign addr[34590]= 588984994;
assign addr[34591]= 625668632;
assign addr[34592]= 662153826;
assign addr[34593]= 698429006;
assign addr[34594]= 734482665;
assign addr[34595]= 770303369;
assign addr[34596]= 805879757;
assign addr[34597]= 841200544;
assign addr[34598]= 876254528;
assign addr[34599]= 911030591;
assign addr[34600]= 945517704;
assign addr[34601]= 979704927;
assign addr[34602]= 1013581418;
assign addr[34603]= 1047136432;
assign addr[34604]= 1080359326;
assign addr[34605]= 1113239564;
assign addr[34606]= 1145766716;
assign addr[34607]= 1177930466;
assign addr[34608]= 1209720613;
assign addr[34609]= 1241127074;
assign addr[34610]= 1272139887;
assign addr[34611]= 1302749217;
assign addr[34612]= 1332945355;
assign addr[34613]= 1362718723;
assign addr[34614]= 1392059879;
assign addr[34615]= 1420959516;
assign addr[34616]= 1449408469;
assign addr[34617]= 1477397714;
assign addr[34618]= 1504918373;
assign addr[34619]= 1531961719;
assign addr[34620]= 1558519173;
assign addr[34621]= 1584582314;
assign addr[34622]= 1610142873;
assign addr[34623]= 1635192744;
assign addr[34624]= 1659723983;
assign addr[34625]= 1683728808;
assign addr[34626]= 1707199606;
assign addr[34627]= 1730128933;
assign addr[34628]= 1752509516;
assign addr[34629]= 1774334257;
assign addr[34630]= 1795596234;
assign addr[34631]= 1816288703;
assign addr[34632]= 1836405100;
assign addr[34633]= 1855939047;
assign addr[34634]= 1874884346;
assign addr[34635]= 1893234990;
assign addr[34636]= 1910985158;
assign addr[34637]= 1928129220;
assign addr[34638]= 1944661739;
assign addr[34639]= 1960577471;
assign addr[34640]= 1975871368;
assign addr[34641]= 1990538579;
assign addr[34642]= 2004574453;
assign addr[34643]= 2017974537;
assign addr[34644]= 2030734582;
assign addr[34645]= 2042850540;
assign addr[34646]= 2054318569;
assign addr[34647]= 2065135031;
assign addr[34648]= 2075296495;
assign addr[34649]= 2084799740;
assign addr[34650]= 2093641749;
assign addr[34651]= 2101819720;
assign addr[34652]= 2109331059;
assign addr[34653]= 2116173382;
assign addr[34654]= 2122344521;
assign addr[34655]= 2127842516;
assign addr[34656]= 2132665626;
assign addr[34657]= 2136812319;
assign addr[34658]= 2140281282;
assign addr[34659]= 2143071413;
assign addr[34660]= 2145181827;
assign addr[34661]= 2146611856;
assign addr[34662]= 2147361045;
assign addr[34663]= 2147429158;
assign addr[34664]= 2146816171;
assign addr[34665]= 2145522281;
assign addr[34666]= 2143547897;
assign addr[34667]= 2140893646;
assign addr[34668]= 2137560369;
assign addr[34669]= 2133549123;
assign addr[34670]= 2128861181;
assign addr[34671]= 2123498030;
assign addr[34672]= 2117461370;
assign addr[34673]= 2110753117;
assign addr[34674]= 2103375398;
assign addr[34675]= 2095330553;
assign addr[34676]= 2086621133;
assign addr[34677]= 2077249901;
assign addr[34678]= 2067219829;
assign addr[34679]= 2056534099;
assign addr[34680]= 2045196100;
assign addr[34681]= 2033209426;
assign addr[34682]= 2020577882;
assign addr[34683]= 2007305472;
assign addr[34684]= 1993396407;
assign addr[34685]= 1978855097;
assign addr[34686]= 1963686155;
assign addr[34687]= 1947894393;
assign addr[34688]= 1931484818;
assign addr[34689]= 1914462636;
assign addr[34690]= 1896833245;
assign addr[34691]= 1878602237;
assign addr[34692]= 1859775393;
assign addr[34693]= 1840358687;
assign addr[34694]= 1820358275;
assign addr[34695]= 1799780501;
assign addr[34696]= 1778631892;
assign addr[34697]= 1756919156;
assign addr[34698]= 1734649179;
assign addr[34699]= 1711829025;
assign addr[34700]= 1688465931;
assign addr[34701]= 1664567307;
assign addr[34702]= 1640140734;
assign addr[34703]= 1615193959;
assign addr[34704]= 1589734894;
assign addr[34705]= 1563771613;
assign addr[34706]= 1537312353;
assign addr[34707]= 1510365504;
assign addr[34708]= 1482939614;
assign addr[34709]= 1455043381;
assign addr[34710]= 1426685652;
assign addr[34711]= 1397875423;
assign addr[34712]= 1368621831;
assign addr[34713]= 1338934154;
assign addr[34714]= 1308821808;
assign addr[34715]= 1278294345;
assign addr[34716]= 1247361445;
assign addr[34717]= 1216032921;
assign addr[34718]= 1184318708;
assign addr[34719]= 1152228866;
assign addr[34720]= 1119773573;
assign addr[34721]= 1086963121;
assign addr[34722]= 1053807919;
assign addr[34723]= 1020318481;
assign addr[34724]= 986505429;
assign addr[34725]= 952379488;
assign addr[34726]= 917951481;
assign addr[34727]= 883232329;
assign addr[34728]= 848233042;
assign addr[34729]= 812964722;
assign addr[34730]= 777438554;
assign addr[34731]= 741665807;
assign addr[34732]= 705657826;
assign addr[34733]= 669426032;
assign addr[34734]= 632981917;
assign addr[34735]= 596337040;
assign addr[34736]= 559503022;
assign addr[34737]= 522491548;
assign addr[34738]= 485314355;
assign addr[34739]= 447983235;
assign addr[34740]= 410510029;
assign addr[34741]= 372906622;
assign addr[34742]= 335184940;
assign addr[34743]= 297356948;
assign addr[34744]= 259434643;
assign addr[34745]= 221430054;
assign addr[34746]= 183355234;
assign addr[34747]= 145222259;
assign addr[34748]= 107043224;
assign addr[34749]= 68830239;
assign addr[34750]= 30595422;
assign addr[34751]= -7649098;
assign addr[34752]= -45891193;
assign addr[34753]= -84118732;
assign addr[34754]= -122319591;
assign addr[34755]= -160481654;
assign addr[34756]= -198592817;
assign addr[34757]= -236640993;
assign addr[34758]= -274614114;
assign addr[34759]= -312500135;
assign addr[34760]= -350287041;
assign addr[34761]= -387962847;
assign addr[34762]= -425515602;
assign addr[34763]= -462933398;
assign addr[34764]= -500204365;
assign addr[34765]= -537316682;
assign addr[34766]= -574258580;
assign addr[34767]= -611018340;
assign addr[34768]= -647584304;
assign addr[34769]= -683944874;
assign addr[34770]= -720088517;
assign addr[34771]= -756003771;
assign addr[34772]= -791679244;
assign addr[34773]= -827103620;
assign addr[34774]= -862265664;
assign addr[34775]= -897154224;
assign addr[34776]= -931758235;
assign addr[34777]= -966066720;
assign addr[34778]= -1000068799;
assign addr[34779]= -1033753687;
assign addr[34780]= -1067110699;
assign addr[34781]= -1100129257;
assign addr[34782]= -1132798888;
assign addr[34783]= -1165109230;
assign addr[34784]= -1197050035;
assign addr[34785]= -1228611172;
assign addr[34786]= -1259782632;
assign addr[34787]= -1290554528;
assign addr[34788]= -1320917099;
assign addr[34789]= -1350860716;
assign addr[34790]= -1380375881;
assign addr[34791]= -1409453233;
assign addr[34792]= -1438083551;
assign addr[34793]= -1466257752;
assign addr[34794]= -1493966902;
assign addr[34795]= -1521202211;
assign addr[34796]= -1547955041;
assign addr[34797]= -1574216908;
assign addr[34798]= -1599979481;
assign addr[34799]= -1625234591;
assign addr[34800]= -1649974225;
assign addr[34801]= -1674190539;
assign addr[34802]= -1697875851;
assign addr[34803]= -1721022648;
assign addr[34804]= -1743623590;
assign addr[34805]= -1765671509;
assign addr[34806]= -1787159411;
assign addr[34807]= -1808080480;
assign addr[34808]= -1828428082;
assign addr[34809]= -1848195763;
assign addr[34810]= -1867377253;
assign addr[34811]= -1885966468;
assign addr[34812]= -1903957513;
assign addr[34813]= -1921344681;
assign addr[34814]= -1938122457;
assign addr[34815]= -1954285520;
assign addr[34816]= -1969828744;
assign addr[34817]= -1984747199;
assign addr[34818]= -1999036154;
assign addr[34819]= -2012691075;
assign addr[34820]= -2025707632;
assign addr[34821]= -2038081698;
assign addr[34822]= -2049809346;
assign addr[34823]= -2060886858;
assign addr[34824]= -2071310720;
assign addr[34825]= -2081077626;
assign addr[34826]= -2090184478;
assign addr[34827]= -2098628387;
assign addr[34828]= -2106406677;
assign addr[34829]= -2113516878;
assign addr[34830]= -2119956737;
assign addr[34831]= -2125724211;
assign addr[34832]= -2130817471;
assign addr[34833]= -2135234901;
assign addr[34834]= -2138975100;
assign addr[34835]= -2142036881;
assign addr[34836]= -2144419275;
assign addr[34837]= -2146121524;
assign addr[34838]= -2147143090;
assign addr[34839]= -2147483648;
assign addr[34840]= -2147143090;
assign addr[34841]= -2146121524;
assign addr[34842]= -2144419275;
assign addr[34843]= -2142036881;
assign addr[34844]= -2138975100;
assign addr[34845]= -2135234901;
assign addr[34846]= -2130817471;
assign addr[34847]= -2125724211;
assign addr[34848]= -2119956737;
assign addr[34849]= -2113516878;
assign addr[34850]= -2106406677;
assign addr[34851]= -2098628387;
assign addr[34852]= -2090184478;
assign addr[34853]= -2081077626;
assign addr[34854]= -2071310720;
assign addr[34855]= -2060886858;
assign addr[34856]= -2049809346;
assign addr[34857]= -2038081698;
assign addr[34858]= -2025707632;
assign addr[34859]= -2012691075;
assign addr[34860]= -1999036154;
assign addr[34861]= -1984747199;
assign addr[34862]= -1969828744;
assign addr[34863]= -1954285520;
assign addr[34864]= -1938122457;
assign addr[34865]= -1921344681;
assign addr[34866]= -1903957513;
assign addr[34867]= -1885966468;
assign addr[34868]= -1867377253;
assign addr[34869]= -1848195763;
assign addr[34870]= -1828428082;
assign addr[34871]= -1808080480;
assign addr[34872]= -1787159411;
assign addr[34873]= -1765671509;
assign addr[34874]= -1743623590;
assign addr[34875]= -1721022648;
assign addr[34876]= -1697875851;
assign addr[34877]= -1674190539;
assign addr[34878]= -1649974225;
assign addr[34879]= -1625234591;
assign addr[34880]= -1599979481;
assign addr[34881]= -1574216908;
assign addr[34882]= -1547955041;
assign addr[34883]= -1521202211;
assign addr[34884]= -1493966902;
assign addr[34885]= -1466257752;
assign addr[34886]= -1438083551;
assign addr[34887]= -1409453233;
assign addr[34888]= -1380375881;
assign addr[34889]= -1350860716;
assign addr[34890]= -1320917099;
assign addr[34891]= -1290554528;
assign addr[34892]= -1259782632;
assign addr[34893]= -1228611172;
assign addr[34894]= -1197050035;
assign addr[34895]= -1165109230;
assign addr[34896]= -1132798888;
assign addr[34897]= -1100129257;
assign addr[34898]= -1067110699;
assign addr[34899]= -1033753687;
assign addr[34900]= -1000068799;
assign addr[34901]= -966066720;
assign addr[34902]= -931758235;
assign addr[34903]= -897154224;
assign addr[34904]= -862265664;
assign addr[34905]= -827103620;
assign addr[34906]= -791679244;
assign addr[34907]= -756003771;
assign addr[34908]= -720088517;
assign addr[34909]= -683944874;
assign addr[34910]= -647584304;
assign addr[34911]= -611018340;
assign addr[34912]= -574258580;
assign addr[34913]= -537316682;
assign addr[34914]= -500204365;
assign addr[34915]= -462933398;
assign addr[34916]= -425515602;
assign addr[34917]= -387962847;
assign addr[34918]= -350287041;
assign addr[34919]= -312500135;
assign addr[34920]= -274614114;
assign addr[34921]= -236640993;
assign addr[34922]= -198592817;
assign addr[34923]= -160481654;
assign addr[34924]= -122319591;
assign addr[34925]= -84118732;
assign addr[34926]= -45891193;
assign addr[34927]= -7649098;
assign addr[34928]= 30595422;
assign addr[34929]= 68830239;
assign addr[34930]= 107043224;
assign addr[34931]= 145222259;
assign addr[34932]= 183355234;
assign addr[34933]= 221430054;
assign addr[34934]= 259434643;
assign addr[34935]= 297356948;
assign addr[34936]= 335184940;
assign addr[34937]= 372906622;
assign addr[34938]= 410510029;
assign addr[34939]= 447983235;
assign addr[34940]= 485314355;
assign addr[34941]= 522491548;
assign addr[34942]= 559503022;
assign addr[34943]= 596337040;
assign addr[34944]= 632981917;
assign addr[34945]= 669426032;
assign addr[34946]= 705657826;
assign addr[34947]= 741665807;
assign addr[34948]= 777438554;
assign addr[34949]= 812964722;
assign addr[34950]= 848233042;
assign addr[34951]= 883232329;
assign addr[34952]= 917951481;
assign addr[34953]= 952379488;
assign addr[34954]= 986505429;
assign addr[34955]= 1020318481;
assign addr[34956]= 1053807919;
assign addr[34957]= 1086963121;
assign addr[34958]= 1119773573;
assign addr[34959]= 1152228866;
assign addr[34960]= 1184318708;
assign addr[34961]= 1216032921;
assign addr[34962]= 1247361445;
assign addr[34963]= 1278294345;
assign addr[34964]= 1308821808;
assign addr[34965]= 1338934154;
assign addr[34966]= 1368621831;
assign addr[34967]= 1397875423;
assign addr[34968]= 1426685652;
assign addr[34969]= 1455043381;
assign addr[34970]= 1482939614;
assign addr[34971]= 1510365504;
assign addr[34972]= 1537312353;
assign addr[34973]= 1563771613;
assign addr[34974]= 1589734894;
assign addr[34975]= 1615193959;
assign addr[34976]= 1640140734;
assign addr[34977]= 1664567307;
assign addr[34978]= 1688465931;
assign addr[34979]= 1711829025;
assign addr[34980]= 1734649179;
assign addr[34981]= 1756919156;
assign addr[34982]= 1778631892;
assign addr[34983]= 1799780501;
assign addr[34984]= 1820358275;
assign addr[34985]= 1840358687;
assign addr[34986]= 1859775393;
assign addr[34987]= 1878602237;
assign addr[34988]= 1896833245;
assign addr[34989]= 1914462636;
assign addr[34990]= 1931484818;
assign addr[34991]= 1947894393;
assign addr[34992]= 1963686155;
assign addr[34993]= 1978855097;
assign addr[34994]= 1993396407;
assign addr[34995]= 2007305472;
assign addr[34996]= 2020577882;
assign addr[34997]= 2033209426;
assign addr[34998]= 2045196100;
assign addr[34999]= 2056534099;
assign addr[35000]= 2067219829;
assign addr[35001]= 2077249901;
assign addr[35002]= 2086621133;
assign addr[35003]= 2095330553;
assign addr[35004]= 2103375398;
assign addr[35005]= 2110753117;
assign addr[35006]= 2117461370;
assign addr[35007]= 2123498030;
assign addr[35008]= 2128861181;
assign addr[35009]= 2133549123;
assign addr[35010]= 2137560369;
assign addr[35011]= 2140893646;
assign addr[35012]= 2143547897;
assign addr[35013]= 2145522281;
assign addr[35014]= 2146816171;
assign addr[35015]= 2147429158;
assign addr[35016]= 2147361045;
assign addr[35017]= 2146611856;
assign addr[35018]= 2145181827;
assign addr[35019]= 2143071413;
assign addr[35020]= 2140281282;
assign addr[35021]= 2136812319;
assign addr[35022]= 2132665626;
assign addr[35023]= 2127842516;
assign addr[35024]= 2122344521;
assign addr[35025]= 2116173382;
assign addr[35026]= 2109331059;
assign addr[35027]= 2101819720;
assign addr[35028]= 2093641749;
assign addr[35029]= 2084799740;
assign addr[35030]= 2075296495;
assign addr[35031]= 2065135031;
assign addr[35032]= 2054318569;
assign addr[35033]= 2042850540;
assign addr[35034]= 2030734582;
assign addr[35035]= 2017974537;
assign addr[35036]= 2004574453;
assign addr[35037]= 1990538579;
assign addr[35038]= 1975871368;
assign addr[35039]= 1960577471;
assign addr[35040]= 1944661739;
assign addr[35041]= 1928129220;
assign addr[35042]= 1910985158;
assign addr[35043]= 1893234990;
assign addr[35044]= 1874884346;
assign addr[35045]= 1855939047;
assign addr[35046]= 1836405100;
assign addr[35047]= 1816288703;
assign addr[35048]= 1795596234;
assign addr[35049]= 1774334257;
assign addr[35050]= 1752509516;
assign addr[35051]= 1730128933;
assign addr[35052]= 1707199606;
assign addr[35053]= 1683728808;
assign addr[35054]= 1659723983;
assign addr[35055]= 1635192744;
assign addr[35056]= 1610142873;
assign addr[35057]= 1584582314;
assign addr[35058]= 1558519173;
assign addr[35059]= 1531961719;
assign addr[35060]= 1504918373;
assign addr[35061]= 1477397714;
assign addr[35062]= 1449408469;
assign addr[35063]= 1420959516;
assign addr[35064]= 1392059879;
assign addr[35065]= 1362718723;
assign addr[35066]= 1332945355;
assign addr[35067]= 1302749217;
assign addr[35068]= 1272139887;
assign addr[35069]= 1241127074;
assign addr[35070]= 1209720613;
assign addr[35071]= 1177930466;
assign addr[35072]= 1145766716;
assign addr[35073]= 1113239564;
assign addr[35074]= 1080359326;
assign addr[35075]= 1047136432;
assign addr[35076]= 1013581418;
assign addr[35077]= 979704927;
assign addr[35078]= 945517704;
assign addr[35079]= 911030591;
assign addr[35080]= 876254528;
assign addr[35081]= 841200544;
assign addr[35082]= 805879757;
assign addr[35083]= 770303369;
assign addr[35084]= 734482665;
assign addr[35085]= 698429006;
assign addr[35086]= 662153826;
assign addr[35087]= 625668632;
assign addr[35088]= 588984994;
assign addr[35089]= 552114549;
assign addr[35090]= 515068990;
assign addr[35091]= 477860067;
assign addr[35092]= 440499581;
assign addr[35093]= 402999383;
assign addr[35094]= 365371365;
assign addr[35095]= 327627463;
assign addr[35096]= 289779648;
assign addr[35097]= 251839923;
assign addr[35098]= 213820322;
assign addr[35099]= 175732905;
assign addr[35100]= 137589750;
assign addr[35101]= 99402956;
assign addr[35102]= 61184634;
assign addr[35103]= 22946906;
assign addr[35104]= -15298099;
assign addr[35105]= -53538253;
assign addr[35106]= -91761426;
assign addr[35107]= -129955495;
assign addr[35108]= -168108346;
assign addr[35109]= -206207878;
assign addr[35110]= -244242007;
assign addr[35111]= -282198671;
assign addr[35112]= -320065829;
assign addr[35113]= -357831473;
assign addr[35114]= -395483624;
assign addr[35115]= -433010339;
assign addr[35116]= -470399716;
assign addr[35117]= -507639898;
assign addr[35118]= -544719071;
assign addr[35119]= -581625477;
assign addr[35120]= -618347408;
assign addr[35121]= -654873219;
assign addr[35122]= -691191324;
assign addr[35123]= -727290205;
assign addr[35124]= -763158411;
assign addr[35125]= -798784567;
assign addr[35126]= -834157373;
assign addr[35127]= -869265610;
assign addr[35128]= -904098143;
assign addr[35129]= -938643924;
assign addr[35130]= -972891995;
assign addr[35131]= -1006831495;
assign addr[35132]= -1040451659;
assign addr[35133]= -1073741824;
assign addr[35134]= -1106691431;
assign addr[35135]= -1139290029;
assign addr[35136]= -1171527280;
assign addr[35137]= -1203392958;
assign addr[35138]= -1234876957;
assign addr[35139]= -1265969291;
assign addr[35140]= -1296660098;
assign addr[35141]= -1326939644;
assign addr[35142]= -1356798326;
assign addr[35143]= -1386226674;
assign addr[35144]= -1415215352;
assign addr[35145]= -1443755168;
assign addr[35146]= -1471837070;
assign addr[35147]= -1499452149;
assign addr[35148]= -1526591649;
assign addr[35149]= -1553246960;
assign addr[35150]= -1579409630;
assign addr[35151]= -1605071359;
assign addr[35152]= -1630224009;
assign addr[35153]= -1654859602;
assign addr[35154]= -1678970324;
assign addr[35155]= -1702548529;
assign addr[35156]= -1725586737;
assign addr[35157]= -1748077642;
assign addr[35158]= -1770014111;
assign addr[35159]= -1791389186;
assign addr[35160]= -1812196087;
assign addr[35161]= -1832428215;
assign addr[35162]= -1852079154;
assign addr[35163]= -1871142669;
assign addr[35164]= -1889612716;
assign addr[35165]= -1907483436;
assign addr[35166]= -1924749160;
assign addr[35167]= -1941404413;
assign addr[35168]= -1957443913;
assign addr[35169]= -1972862571;
assign addr[35170]= -1987655498;
assign addr[35171]= -2001818002;
assign addr[35172]= -2015345591;
assign addr[35173]= -2028233973;
assign addr[35174]= -2040479063;
assign addr[35175]= -2052076975;
assign addr[35176]= -2063024031;
assign addr[35177]= -2073316760;
assign addr[35178]= -2082951896;
assign addr[35179]= -2091926384;
assign addr[35180]= -2100237377;
assign addr[35181]= -2107882239;
assign addr[35182]= -2114858546;
assign addr[35183]= -2121164085;
assign addr[35184]= -2126796855;
assign addr[35185]= -2131755071;
assign addr[35186]= -2136037160;
assign addr[35187]= -2139641764;
assign addr[35188]= -2142567738;
assign addr[35189]= -2144814157;
assign addr[35190]= -2146380306;
assign addr[35191]= -2147265689;
assign addr[35192]= -2147470025;
assign addr[35193]= -2146993250;
assign addr[35194]= -2145835515;
assign addr[35195]= -2143997187;
assign addr[35196]= -2141478848;
assign addr[35197]= -2138281298;
assign addr[35198]= -2134405552;
assign addr[35199]= -2129852837;
assign addr[35200]= -2124624598;
assign addr[35201]= -2118722494;
assign addr[35202]= -2112148396;
assign addr[35203]= -2104904390;
assign addr[35204]= -2096992772;
assign addr[35205]= -2088416053;
assign addr[35206]= -2079176953;
assign addr[35207]= -2069278401;
assign addr[35208]= -2058723538;
assign addr[35209]= -2047515711;
assign addr[35210]= -2035658475;
assign addr[35211]= -2023155591;
assign addr[35212]= -2010011024;
assign addr[35213]= -1996228943;
assign addr[35214]= -1981813720;
assign addr[35215]= -1966769926;
assign addr[35216]= -1951102334;
assign addr[35217]= -1934815911;
assign addr[35218]= -1917915825;
assign addr[35219]= -1900407434;
assign addr[35220]= -1882296293;
assign addr[35221]= -1863588145;
assign addr[35222]= -1844288924;
assign addr[35223]= -1824404752;
assign addr[35224]= -1803941934;
assign addr[35225]= -1782906961;
assign addr[35226]= -1761306505;
assign addr[35227]= -1739147417;
assign addr[35228]= -1716436725;
assign addr[35229]= -1693181631;
assign addr[35230]= -1669389513;
assign addr[35231]= -1645067915;
assign addr[35232]= -1620224553;
assign addr[35233]= -1594867305;
assign addr[35234]= -1569004214;
assign addr[35235]= -1542643483;
assign addr[35236]= -1515793473;
assign addr[35237]= -1488462700;
assign addr[35238]= -1460659832;
assign addr[35239]= -1432393688;
assign addr[35240]= -1403673233;
assign addr[35241]= -1374507575;
assign addr[35242]= -1344905966;
assign addr[35243]= -1314877795;
assign addr[35244]= -1284432584;
assign addr[35245]= -1253579991;
assign addr[35246]= -1222329801;
assign addr[35247]= -1190691925;
assign addr[35248]= -1158676398;
assign addr[35249]= -1126293375;
assign addr[35250]= -1093553126;
assign addr[35251]= -1060466036;
assign addr[35252]= -1027042599;
assign addr[35253]= -993293415;
assign addr[35254]= -959229189;
assign addr[35255]= -924860725;
assign addr[35256]= -890198924;
assign addr[35257]= -855254778;
assign addr[35258]= -820039373;
assign addr[35259]= -784563876;
assign addr[35260]= -748839539;
assign addr[35261]= -712877694;
assign addr[35262]= -676689746;
assign addr[35263]= -640287172;
assign addr[35264]= -603681519;
assign addr[35265]= -566884397;
assign addr[35266]= -529907477;
assign addr[35267]= -492762486;
assign addr[35268]= -455461206;
assign addr[35269]= -418015468;
assign addr[35270]= -380437148;
assign addr[35271]= -342738165;
assign addr[35272]= -304930476;
assign addr[35273]= -267026072;
assign addr[35274]= -229036977;
assign addr[35275]= -190975237;
assign addr[35276]= -152852926;
assign addr[35277]= -114682135;
assign addr[35278]= -76474970;
assign addr[35279]= -38243550;
assign addr[35280]= 0;
assign addr[35281]= 38243550;
assign addr[35282]= 76474970;
assign addr[35283]= 114682135;
assign addr[35284]= 152852926;
assign addr[35285]= 190975237;
assign addr[35286]= 229036977;
assign addr[35287]= 267026072;
assign addr[35288]= 304930476;
assign addr[35289]= 342738165;
assign addr[35290]= 380437148;
assign addr[35291]= 418015468;
assign addr[35292]= 455461206;
assign addr[35293]= 492762486;
assign addr[35294]= 529907477;
assign addr[35295]= 566884397;
assign addr[35296]= 603681519;
assign addr[35297]= 640287172;
assign addr[35298]= 676689746;
assign addr[35299]= 712877694;
assign addr[35300]= 748839539;
assign addr[35301]= 784563876;
assign addr[35302]= 820039373;
assign addr[35303]= 855254778;
assign addr[35304]= 890198924;
assign addr[35305]= 924860725;
assign addr[35306]= 959229189;
assign addr[35307]= 993293415;
assign addr[35308]= 1027042599;
assign addr[35309]= 1060466036;
assign addr[35310]= 1093553126;
assign addr[35311]= 1126293375;
assign addr[35312]= 1158676398;
assign addr[35313]= 1190691925;
assign addr[35314]= 1222329801;
assign addr[35315]= 1253579991;
assign addr[35316]= 1284432584;
assign addr[35317]= 1314877795;
assign addr[35318]= 1344905966;
assign addr[35319]= 1374507575;
assign addr[35320]= 1403673233;
assign addr[35321]= 1432393688;
assign addr[35322]= 1460659832;
assign addr[35323]= 1488462700;
assign addr[35324]= 1515793473;
assign addr[35325]= 1542643483;
assign addr[35326]= 1569004214;
assign addr[35327]= 1594867305;
assign addr[35328]= 1620224553;
assign addr[35329]= 1645067915;
assign addr[35330]= 1669389513;
assign addr[35331]= 1693181631;
assign addr[35332]= 1716436725;
assign addr[35333]= 1739147417;
assign addr[35334]= 1761306505;
assign addr[35335]= 1782906961;
assign addr[35336]= 1803941934;
assign addr[35337]= 1824404752;
assign addr[35338]= 1844288924;
assign addr[35339]= 1863588145;
assign addr[35340]= 1882296293;
assign addr[35341]= 1900407434;
assign addr[35342]= 1917915825;
assign addr[35343]= 1934815911;
assign addr[35344]= 1951102334;
assign addr[35345]= 1966769926;
assign addr[35346]= 1981813720;
assign addr[35347]= 1996228943;
assign addr[35348]= 2010011024;
assign addr[35349]= 2023155591;
assign addr[35350]= 2035658475;
assign addr[35351]= 2047515711;
assign addr[35352]= 2058723538;
assign addr[35353]= 2069278401;
assign addr[35354]= 2079176953;
assign addr[35355]= 2088416053;
assign addr[35356]= 2096992772;
assign addr[35357]= 2104904390;
assign addr[35358]= 2112148396;
assign addr[35359]= 2118722494;
assign addr[35360]= 2124624598;
assign addr[35361]= 2129852837;
assign addr[35362]= 2134405552;
assign addr[35363]= 2138281298;
assign addr[35364]= 2141478848;
assign addr[35365]= 2143997187;
assign addr[35366]= 2145835515;
assign addr[35367]= 2146993250;
assign addr[35368]= 2147470025;
assign addr[35369]= 2147265689;
assign addr[35370]= 2146380306;
assign addr[35371]= 2144814157;
assign addr[35372]= 2142567738;
assign addr[35373]= 2139641764;
assign addr[35374]= 2136037160;
assign addr[35375]= 2131755071;
assign addr[35376]= 2126796855;
assign addr[35377]= 2121164085;
assign addr[35378]= 2114858546;
assign addr[35379]= 2107882239;
assign addr[35380]= 2100237377;
assign addr[35381]= 2091926384;
assign addr[35382]= 2082951896;
assign addr[35383]= 2073316760;
assign addr[35384]= 2063024031;
assign addr[35385]= 2052076975;
assign addr[35386]= 2040479063;
assign addr[35387]= 2028233973;
assign addr[35388]= 2015345591;
assign addr[35389]= 2001818002;
assign addr[35390]= 1987655498;
assign addr[35391]= 1972862571;
assign addr[35392]= 1957443913;
assign addr[35393]= 1941404413;
assign addr[35394]= 1924749160;
assign addr[35395]= 1907483436;
assign addr[35396]= 1889612716;
assign addr[35397]= 1871142669;
assign addr[35398]= 1852079154;
assign addr[35399]= 1832428215;
assign addr[35400]= 1812196087;
assign addr[35401]= 1791389186;
assign addr[35402]= 1770014111;
assign addr[35403]= 1748077642;
assign addr[35404]= 1725586737;
assign addr[35405]= 1702548529;
assign addr[35406]= 1678970324;
assign addr[35407]= 1654859602;
assign addr[35408]= 1630224009;
assign addr[35409]= 1605071359;
assign addr[35410]= 1579409630;
assign addr[35411]= 1553246960;
assign addr[35412]= 1526591649;
assign addr[35413]= 1499452149;
assign addr[35414]= 1471837070;
assign addr[35415]= 1443755168;
assign addr[35416]= 1415215352;
assign addr[35417]= 1386226674;
assign addr[35418]= 1356798326;
assign addr[35419]= 1326939644;
assign addr[35420]= 1296660098;
assign addr[35421]= 1265969291;
assign addr[35422]= 1234876957;
assign addr[35423]= 1203392958;
assign addr[35424]= 1171527280;
assign addr[35425]= 1139290029;
assign addr[35426]= 1106691431;
assign addr[35427]= 1073741824;
assign addr[35428]= 1040451659;
assign addr[35429]= 1006831495;
assign addr[35430]= 972891995;
assign addr[35431]= 938643924;
assign addr[35432]= 904098143;
assign addr[35433]= 869265610;
assign addr[35434]= 834157373;
assign addr[35435]= 798784567;
assign addr[35436]= 763158411;
assign addr[35437]= 727290205;
assign addr[35438]= 691191324;
assign addr[35439]= 654873219;
assign addr[35440]= 618347408;
assign addr[35441]= 581625477;
assign addr[35442]= 544719071;
assign addr[35443]= 507639898;
assign addr[35444]= 470399716;
assign addr[35445]= 433010339;
assign addr[35446]= 395483624;
assign addr[35447]= 357831473;
assign addr[35448]= 320065829;
assign addr[35449]= 282198671;
assign addr[35450]= 244242007;
assign addr[35451]= 206207878;
assign addr[35452]= 168108346;
assign addr[35453]= 129955495;
assign addr[35454]= 91761426;
assign addr[35455]= 53538253;
assign addr[35456]= 15298099;
assign addr[35457]= -22946906;
assign addr[35458]= -61184634;
assign addr[35459]= -99402956;
assign addr[35460]= -137589750;
assign addr[35461]= -175732905;
assign addr[35462]= -213820322;
assign addr[35463]= -251839923;
assign addr[35464]= -289779648;
assign addr[35465]= -327627463;
assign addr[35466]= -365371365;
assign addr[35467]= -402999383;
assign addr[35468]= -440499581;
assign addr[35469]= -477860067;
assign addr[35470]= -515068990;
assign addr[35471]= -552114549;
assign addr[35472]= -588984994;
assign addr[35473]= -625668632;
assign addr[35474]= -662153826;
assign addr[35475]= -698429006;
assign addr[35476]= -734482665;
assign addr[35477]= -770303369;
assign addr[35478]= -805879757;
assign addr[35479]= -841200544;
assign addr[35480]= -876254528;
assign addr[35481]= -911030591;
assign addr[35482]= -945517704;
assign addr[35483]= -979704927;
assign addr[35484]= -1013581418;
assign addr[35485]= -1047136432;
assign addr[35486]= -1080359326;
assign addr[35487]= -1113239564;
assign addr[35488]= -1145766716;
assign addr[35489]= -1177930466;
assign addr[35490]= -1209720613;
assign addr[35491]= -1241127074;
assign addr[35492]= -1272139887;
assign addr[35493]= -1302749217;
assign addr[35494]= -1332945355;
assign addr[35495]= -1362718723;
assign addr[35496]= -1392059879;
assign addr[35497]= -1420959516;
assign addr[35498]= -1449408469;
assign addr[35499]= -1477397714;
assign addr[35500]= -1504918373;
assign addr[35501]= -1531961719;
assign addr[35502]= -1558519173;
assign addr[35503]= -1584582314;
assign addr[35504]= -1610142873;
assign addr[35505]= -1635192744;
assign addr[35506]= -1659723983;
assign addr[35507]= -1683728808;
assign addr[35508]= -1707199606;
assign addr[35509]= -1730128933;
assign addr[35510]= -1752509516;
assign addr[35511]= -1774334257;
assign addr[35512]= -1795596234;
assign addr[35513]= -1816288703;
assign addr[35514]= -1836405100;
assign addr[35515]= -1855939047;
assign addr[35516]= -1874884346;
assign addr[35517]= -1893234990;
assign addr[35518]= -1910985158;
assign addr[35519]= -1928129220;
assign addr[35520]= -1944661739;
assign addr[35521]= -1960577471;
assign addr[35522]= -1975871368;
assign addr[35523]= -1990538579;
assign addr[35524]= -2004574453;
assign addr[35525]= -2017974537;
assign addr[35526]= -2030734582;
assign addr[35527]= -2042850540;
assign addr[35528]= -2054318569;
assign addr[35529]= -2065135031;
assign addr[35530]= -2075296495;
assign addr[35531]= -2084799740;
assign addr[35532]= -2093641749;
assign addr[35533]= -2101819720;
assign addr[35534]= -2109331059;
assign addr[35535]= -2116173382;
assign addr[35536]= -2122344521;
assign addr[35537]= -2127842516;
assign addr[35538]= -2132665626;
assign addr[35539]= -2136812319;
assign addr[35540]= -2140281282;
assign addr[35541]= -2143071413;
assign addr[35542]= -2145181827;
assign addr[35543]= -2146611856;
assign addr[35544]= -2147361045;
assign addr[35545]= -2147429158;
assign addr[35546]= -2146816171;
assign addr[35547]= -2145522281;
assign addr[35548]= -2143547897;
assign addr[35549]= -2140893646;
assign addr[35550]= -2137560369;
assign addr[35551]= -2133549123;
assign addr[35552]= -2128861181;
assign addr[35553]= -2123498030;
assign addr[35554]= -2117461370;
assign addr[35555]= -2110753117;
assign addr[35556]= -2103375398;
assign addr[35557]= -2095330553;
assign addr[35558]= -2086621133;
assign addr[35559]= -2077249901;
assign addr[35560]= -2067219829;
assign addr[35561]= -2056534099;
assign addr[35562]= -2045196100;
assign addr[35563]= -2033209426;
assign addr[35564]= -2020577882;
assign addr[35565]= -2007305472;
assign addr[35566]= -1993396407;
assign addr[35567]= -1978855097;
assign addr[35568]= -1963686155;
assign addr[35569]= -1947894393;
assign addr[35570]= -1931484818;
assign addr[35571]= -1914462636;
assign addr[35572]= -1896833245;
assign addr[35573]= -1878602237;
assign addr[35574]= -1859775393;
assign addr[35575]= -1840358687;
assign addr[35576]= -1820358275;
assign addr[35577]= -1799780501;
assign addr[35578]= -1778631892;
assign addr[35579]= -1756919156;
assign addr[35580]= -1734649179;
assign addr[35581]= -1711829025;
assign addr[35582]= -1688465931;
assign addr[35583]= -1664567307;
assign addr[35584]= -1640140734;
assign addr[35585]= -1615193959;
assign addr[35586]= -1589734894;
assign addr[35587]= -1563771613;
assign addr[35588]= -1537312353;
assign addr[35589]= -1510365504;
assign addr[35590]= -1482939614;
assign addr[35591]= -1455043381;
assign addr[35592]= -1426685652;
assign addr[35593]= -1397875423;
assign addr[35594]= -1368621831;
assign addr[35595]= -1338934154;
assign addr[35596]= -1308821808;
assign addr[35597]= -1278294345;
assign addr[35598]= -1247361445;
assign addr[35599]= -1216032921;
assign addr[35600]= -1184318708;
assign addr[35601]= -1152228866;
assign addr[35602]= -1119773573;
assign addr[35603]= -1086963121;
assign addr[35604]= -1053807919;
assign addr[35605]= -1020318481;
assign addr[35606]= -986505429;
assign addr[35607]= -952379488;
assign addr[35608]= -917951481;
assign addr[35609]= -883232329;
assign addr[35610]= -848233042;
assign addr[35611]= -812964722;
assign addr[35612]= -777438554;
assign addr[35613]= -741665807;
assign addr[35614]= -705657826;
assign addr[35615]= -669426032;
assign addr[35616]= -632981917;
assign addr[35617]= -596337040;
assign addr[35618]= -559503022;
assign addr[35619]= -522491548;
assign addr[35620]= -485314355;
assign addr[35621]= -447983235;
assign addr[35622]= -410510029;
assign addr[35623]= -372906622;
assign addr[35624]= -335184940;
assign addr[35625]= -297356948;
assign addr[35626]= -259434643;
assign addr[35627]= -221430054;
assign addr[35628]= -183355234;
assign addr[35629]= -145222259;
assign addr[35630]= -107043224;
assign addr[35631]= -68830239;
assign addr[35632]= -30595422;
assign addr[35633]= 7649098;
assign addr[35634]= 45891193;
assign addr[35635]= 84118732;
assign addr[35636]= 122319591;
assign addr[35637]= 160481654;
assign addr[35638]= 198592817;
assign addr[35639]= 236640993;
assign addr[35640]= 274614114;
assign addr[35641]= 312500135;
assign addr[35642]= 350287041;
assign addr[35643]= 387962847;
assign addr[35644]= 425515602;
assign addr[35645]= 462933398;
assign addr[35646]= 500204365;
assign addr[35647]= 537316682;
assign addr[35648]= 574258580;
assign addr[35649]= 611018340;
assign addr[35650]= 647584304;
assign addr[35651]= 683944874;
assign addr[35652]= 720088517;
assign addr[35653]= 756003771;
assign addr[35654]= 791679244;
assign addr[35655]= 827103620;
assign addr[35656]= 862265664;
assign addr[35657]= 897154224;
assign addr[35658]= 931758235;
assign addr[35659]= 966066720;
assign addr[35660]= 1000068799;
assign addr[35661]= 1033753687;
assign addr[35662]= 1067110699;
assign addr[35663]= 1100129257;
assign addr[35664]= 1132798888;
assign addr[35665]= 1165109230;
assign addr[35666]= 1197050035;
assign addr[35667]= 1228611172;
assign addr[35668]= 1259782632;
assign addr[35669]= 1290554528;
assign addr[35670]= 1320917099;
assign addr[35671]= 1350860716;
assign addr[35672]= 1380375881;
assign addr[35673]= 1409453233;
assign addr[35674]= 1438083551;
assign addr[35675]= 1466257752;
assign addr[35676]= 1493966902;
assign addr[35677]= 1521202211;
assign addr[35678]= 1547955041;
assign addr[35679]= 1574216908;
assign addr[35680]= 1599979481;
assign addr[35681]= 1625234591;
assign addr[35682]= 1649974225;
assign addr[35683]= 1674190539;
assign addr[35684]= 1697875851;
assign addr[35685]= 1721022648;
assign addr[35686]= 1743623590;
assign addr[35687]= 1765671509;
assign addr[35688]= 1787159411;
assign addr[35689]= 1808080480;
assign addr[35690]= 1828428082;
assign addr[35691]= 1848195763;
assign addr[35692]= 1867377253;
assign addr[35693]= 1885966468;
assign addr[35694]= 1903957513;
assign addr[35695]= 1921344681;
assign addr[35696]= 1938122457;
assign addr[35697]= 1954285520;
assign addr[35698]= 1969828744;
assign addr[35699]= 1984747199;
assign addr[35700]= 1999036154;
assign addr[35701]= 2012691075;
assign addr[35702]= 2025707632;
assign addr[35703]= 2038081698;
assign addr[35704]= 2049809346;
assign addr[35705]= 2060886858;
assign addr[35706]= 2071310720;
assign addr[35707]= 2081077626;
assign addr[35708]= 2090184478;
assign addr[35709]= 2098628387;
assign addr[35710]= 2106406677;
assign addr[35711]= 2113516878;
assign addr[35712]= 2119956737;
assign addr[35713]= 2125724211;
assign addr[35714]= 2130817471;
assign addr[35715]= 2135234901;
assign addr[35716]= 2138975100;
assign addr[35717]= 2142036881;
assign addr[35718]= 2144419275;
assign addr[35719]= 2146121524;
assign addr[35720]= 2147143090;
assign addr[35721]= 2147483648;
assign addr[35722]= 2147143090;
assign addr[35723]= 2146121524;
assign addr[35724]= 2144419275;
assign addr[35725]= 2142036881;
assign addr[35726]= 2138975100;
assign addr[35727]= 2135234901;
assign addr[35728]= 2130817471;
assign addr[35729]= 2125724211;
assign addr[35730]= 2119956737;
assign addr[35731]= 2113516878;
assign addr[35732]= 2106406677;
assign addr[35733]= 2098628387;
assign addr[35734]= 2090184478;
assign addr[35735]= 2081077626;
assign addr[35736]= 2071310720;
assign addr[35737]= 2060886858;
assign addr[35738]= 2049809346;
assign addr[35739]= 2038081698;
assign addr[35740]= 2025707632;
assign addr[35741]= 2012691075;
assign addr[35742]= 1999036154;
assign addr[35743]= 1984747199;
assign addr[35744]= 1969828744;
assign addr[35745]= 1954285520;
assign addr[35746]= 1938122457;
assign addr[35747]= 1921344681;
assign addr[35748]= 1903957513;
assign addr[35749]= 1885966468;
assign addr[35750]= 1867377253;
assign addr[35751]= 1848195763;
assign addr[35752]= 1828428082;
assign addr[35753]= 1808080480;
assign addr[35754]= 1787159411;
assign addr[35755]= 1765671509;
assign addr[35756]= 1743623590;
assign addr[35757]= 1721022648;
assign addr[35758]= 1697875851;
assign addr[35759]= 1674190539;
assign addr[35760]= 1649974225;
assign addr[35761]= 1625234591;
assign addr[35762]= 1599979481;
assign addr[35763]= 1574216908;
assign addr[35764]= 1547955041;
assign addr[35765]= 1521202211;
assign addr[35766]= 1493966902;
assign addr[35767]= 1466257752;
assign addr[35768]= 1438083551;
assign addr[35769]= 1409453233;
assign addr[35770]= 1380375881;
assign addr[35771]= 1350860716;
assign addr[35772]= 1320917099;
assign addr[35773]= 1290554528;
assign addr[35774]= 1259782632;
assign addr[35775]= 1228611172;
assign addr[35776]= 1197050035;
assign addr[35777]= 1165109230;
assign addr[35778]= 1132798888;
assign addr[35779]= 1100129257;
assign addr[35780]= 1067110699;
assign addr[35781]= 1033753687;
assign addr[35782]= 1000068799;
assign addr[35783]= 966066720;
assign addr[35784]= 931758235;
assign addr[35785]= 897154224;
assign addr[35786]= 862265664;
assign addr[35787]= 827103620;
assign addr[35788]= 791679244;
assign addr[35789]= 756003771;
assign addr[35790]= 720088517;
assign addr[35791]= 683944874;
assign addr[35792]= 647584304;
assign addr[35793]= 611018340;
assign addr[35794]= 574258580;
assign addr[35795]= 537316682;
assign addr[35796]= 500204365;
assign addr[35797]= 462933398;
assign addr[35798]= 425515602;
assign addr[35799]= 387962847;
assign addr[35800]= 350287041;
assign addr[35801]= 312500135;
assign addr[35802]= 274614114;
assign addr[35803]= 236640993;
assign addr[35804]= 198592817;
assign addr[35805]= 160481654;
assign addr[35806]= 122319591;
assign addr[35807]= 84118732;
assign addr[35808]= 45891193;
assign addr[35809]= 7649098;
assign addr[35810]= -30595422;
assign addr[35811]= -68830239;
assign addr[35812]= -107043224;
assign addr[35813]= -145222259;
assign addr[35814]= -183355234;
assign addr[35815]= -221430054;
assign addr[35816]= -259434643;
assign addr[35817]= -297356948;
assign addr[35818]= -335184940;
assign addr[35819]= -372906622;
assign addr[35820]= -410510029;
assign addr[35821]= -447983235;
assign addr[35822]= -485314355;
assign addr[35823]= -522491548;
assign addr[35824]= -559503022;
assign addr[35825]= -596337040;
assign addr[35826]= -632981917;
assign addr[35827]= -669426032;
assign addr[35828]= -705657826;
assign addr[35829]= -741665807;
assign addr[35830]= -777438554;
assign addr[35831]= -812964722;
assign addr[35832]= -848233042;
assign addr[35833]= -883232329;
assign addr[35834]= -917951481;
assign addr[35835]= -952379488;
assign addr[35836]= -986505429;
assign addr[35837]= -1020318481;
assign addr[35838]= -1053807919;
assign addr[35839]= -1086963121;
assign addr[35840]= -1119773573;
assign addr[35841]= -1152228866;
assign addr[35842]= -1184318708;
assign addr[35843]= -1216032921;
assign addr[35844]= -1247361445;
assign addr[35845]= -1278294345;
assign addr[35846]= -1308821808;
assign addr[35847]= -1338934154;
assign addr[35848]= -1368621831;
assign addr[35849]= -1397875423;
assign addr[35850]= -1426685652;
assign addr[35851]= -1455043381;
assign addr[35852]= -1482939614;
assign addr[35853]= -1510365504;
assign addr[35854]= -1537312353;
assign addr[35855]= -1563771613;
assign addr[35856]= -1589734894;
assign addr[35857]= -1615193959;
assign addr[35858]= -1640140734;
assign addr[35859]= -1664567307;
assign addr[35860]= -1688465931;
assign addr[35861]= -1711829025;
assign addr[35862]= -1734649179;
assign addr[35863]= -1756919156;
assign addr[35864]= -1778631892;
assign addr[35865]= -1799780501;
assign addr[35866]= -1820358275;
assign addr[35867]= -1840358687;
assign addr[35868]= -1859775393;
assign addr[35869]= -1878602237;
assign addr[35870]= -1896833245;
assign addr[35871]= -1914462636;
assign addr[35872]= -1931484818;
assign addr[35873]= -1947894393;
assign addr[35874]= -1963686155;
assign addr[35875]= -1978855097;
assign addr[35876]= -1993396407;
assign addr[35877]= -2007305472;
assign addr[35878]= -2020577882;
assign addr[35879]= -2033209426;
assign addr[35880]= -2045196100;
assign addr[35881]= -2056534099;
assign addr[35882]= -2067219829;
assign addr[35883]= -2077249901;
assign addr[35884]= -2086621133;
assign addr[35885]= -2095330553;
assign addr[35886]= -2103375398;
assign addr[35887]= -2110753117;
assign addr[35888]= -2117461370;
assign addr[35889]= -2123498030;
assign addr[35890]= -2128861181;
assign addr[35891]= -2133549123;
assign addr[35892]= -2137560369;
assign addr[35893]= -2140893646;
assign addr[35894]= -2143547897;
assign addr[35895]= -2145522281;
assign addr[35896]= -2146816171;
assign addr[35897]= -2147429158;
assign addr[35898]= -2147361045;
assign addr[35899]= -2146611856;
assign addr[35900]= -2145181827;
assign addr[35901]= -2143071413;
assign addr[35902]= -2140281282;
assign addr[35903]= -2136812319;
assign addr[35904]= -2132665626;
assign addr[35905]= -2127842516;
assign addr[35906]= -2122344521;
assign addr[35907]= -2116173382;
assign addr[35908]= -2109331059;
assign addr[35909]= -2101819720;
assign addr[35910]= -2093641749;
assign addr[35911]= -2084799740;
assign addr[35912]= -2075296495;
assign addr[35913]= -2065135031;
assign addr[35914]= -2054318569;
assign addr[35915]= -2042850540;
assign addr[35916]= -2030734582;
assign addr[35917]= -2017974537;
assign addr[35918]= -2004574453;
assign addr[35919]= -1990538579;
assign addr[35920]= -1975871368;
assign addr[35921]= -1960577471;
assign addr[35922]= -1944661739;
assign addr[35923]= -1928129220;
assign addr[35924]= -1910985158;
assign addr[35925]= -1893234990;
assign addr[35926]= -1874884346;
assign addr[35927]= -1855939047;
assign addr[35928]= -1836405100;
assign addr[35929]= -1816288703;
assign addr[35930]= -1795596234;
assign addr[35931]= -1774334257;
assign addr[35932]= -1752509516;
assign addr[35933]= -1730128933;
assign addr[35934]= -1707199606;
assign addr[35935]= -1683728808;
assign addr[35936]= -1659723983;
assign addr[35937]= -1635192744;
assign addr[35938]= -1610142873;
assign addr[35939]= -1584582314;
assign addr[35940]= -1558519173;
assign addr[35941]= -1531961719;
assign addr[35942]= -1504918373;
assign addr[35943]= -1477397714;
assign addr[35944]= -1449408469;
assign addr[35945]= -1420959516;
assign addr[35946]= -1392059879;
assign addr[35947]= -1362718723;
assign addr[35948]= -1332945355;
assign addr[35949]= -1302749217;
assign addr[35950]= -1272139887;
assign addr[35951]= -1241127074;
assign addr[35952]= -1209720613;
assign addr[35953]= -1177930466;
assign addr[35954]= -1145766716;
assign addr[35955]= -1113239564;
assign addr[35956]= -1080359326;
assign addr[35957]= -1047136432;
assign addr[35958]= -1013581418;
assign addr[35959]= -979704927;
assign addr[35960]= -945517704;
assign addr[35961]= -911030591;
assign addr[35962]= -876254528;
assign addr[35963]= -841200544;
assign addr[35964]= -805879757;
assign addr[35965]= -770303369;
assign addr[35966]= -734482665;
assign addr[35967]= -698429006;
assign addr[35968]= -662153826;
assign addr[35969]= -625668632;
assign addr[35970]= -588984994;
assign addr[35971]= -552114549;
assign addr[35972]= -515068990;
assign addr[35973]= -477860067;
assign addr[35974]= -440499581;
assign addr[35975]= -402999383;
assign addr[35976]= -365371365;
assign addr[35977]= -327627463;
assign addr[35978]= -289779648;
assign addr[35979]= -251839923;
assign addr[35980]= -213820322;
assign addr[35981]= -175732905;
assign addr[35982]= -137589750;
assign addr[35983]= -99402956;
assign addr[35984]= -61184634;
assign addr[35985]= -22946906;
assign addr[35986]= 15298099;
assign addr[35987]= 53538253;
assign addr[35988]= 91761426;
assign addr[35989]= 129955495;
assign addr[35990]= 168108346;
assign addr[35991]= 206207878;
assign addr[35992]= 244242007;
assign addr[35993]= 282198671;
assign addr[35994]= 320065829;
assign addr[35995]= 357831473;
assign addr[35996]= 395483624;
assign addr[35997]= 433010339;
assign addr[35998]= 470399716;
assign addr[35999]= 507639898;
assign addr[36000]= 544719071;
assign addr[36001]= 581625477;
assign addr[36002]= 618347408;
assign addr[36003]= 654873219;
assign addr[36004]= 691191324;
assign addr[36005]= 727290205;
assign addr[36006]= 763158411;
assign addr[36007]= 798784567;
assign addr[36008]= 834157373;
assign addr[36009]= 869265610;
assign addr[36010]= 904098143;
assign addr[36011]= 938643924;
assign addr[36012]= 972891995;
assign addr[36013]= 1006831495;
assign addr[36014]= 1040451659;
assign addr[36015]= 1073741824;
assign addr[36016]= 1106691431;
assign addr[36017]= 1139290029;
assign addr[36018]= 1171527280;
assign addr[36019]= 1203392958;
assign addr[36020]= 1234876957;
assign addr[36021]= 1265969291;
assign addr[36022]= 1296660098;
assign addr[36023]= 1326939644;
assign addr[36024]= 1356798326;
assign addr[36025]= 1386226674;
assign addr[36026]= 1415215352;
assign addr[36027]= 1443755168;
assign addr[36028]= 1471837070;
assign addr[36029]= 1499452149;
assign addr[36030]= 1526591649;
assign addr[36031]= 1553246960;
assign addr[36032]= 1579409630;
assign addr[36033]= 1605071359;
assign addr[36034]= 1630224009;
assign addr[36035]= 1654859602;
assign addr[36036]= 1678970324;
assign addr[36037]= 1702548529;
assign addr[36038]= 1725586737;
assign addr[36039]= 1748077642;
assign addr[36040]= 1770014111;
assign addr[36041]= 1791389186;
assign addr[36042]= 1812196087;
assign addr[36043]= 1832428215;
assign addr[36044]= 1852079154;
assign addr[36045]= 1871142669;
assign addr[36046]= 1889612716;
assign addr[36047]= 1907483436;
assign addr[36048]= 1924749160;
assign addr[36049]= 1941404413;
assign addr[36050]= 1957443913;
assign addr[36051]= 1972862571;
assign addr[36052]= 1987655498;
assign addr[36053]= 2001818002;
assign addr[36054]= 2015345591;
assign addr[36055]= 2028233973;
assign addr[36056]= 2040479063;
assign addr[36057]= 2052076975;
assign addr[36058]= 2063024031;
assign addr[36059]= 2073316760;
assign addr[36060]= 2082951896;
assign addr[36061]= 2091926384;
assign addr[36062]= 2100237377;
assign addr[36063]= 2107882239;
assign addr[36064]= 2114858546;
assign addr[36065]= 2121164085;
assign addr[36066]= 2126796855;
assign addr[36067]= 2131755071;
assign addr[36068]= 2136037160;
assign addr[36069]= 2139641764;
assign addr[36070]= 2142567738;
assign addr[36071]= 2144814157;
assign addr[36072]= 2146380306;
assign addr[36073]= 2147265689;
assign addr[36074]= 2147470025;
assign addr[36075]= 2146993250;
assign addr[36076]= 2145835515;
assign addr[36077]= 2143997187;
assign addr[36078]= 2141478848;
assign addr[36079]= 2138281298;
assign addr[36080]= 2134405552;
assign addr[36081]= 2129852837;
assign addr[36082]= 2124624598;
assign addr[36083]= 2118722494;
assign addr[36084]= 2112148396;
assign addr[36085]= 2104904390;
assign addr[36086]= 2096992772;
assign addr[36087]= 2088416053;
assign addr[36088]= 2079176953;
assign addr[36089]= 2069278401;
assign addr[36090]= 2058723538;
assign addr[36091]= 2047515711;
assign addr[36092]= 2035658475;
assign addr[36093]= 2023155591;
assign addr[36094]= 2010011024;
assign addr[36095]= 1996228943;
assign addr[36096]= 1981813720;
assign addr[36097]= 1966769926;
assign addr[36098]= 1951102334;
assign addr[36099]= 1934815911;
assign addr[36100]= 1917915825;
assign addr[36101]= 1900407434;
assign addr[36102]= 1882296293;
assign addr[36103]= 1863588145;
assign addr[36104]= 1844288924;
assign addr[36105]= 1824404752;
assign addr[36106]= 1803941934;
assign addr[36107]= 1782906961;
assign addr[36108]= 1761306505;
assign addr[36109]= 1739147417;
assign addr[36110]= 1716436725;
assign addr[36111]= 1693181631;
assign addr[36112]= 1669389513;
assign addr[36113]= 1645067915;
assign addr[36114]= 1620224553;
assign addr[36115]= 1594867305;
assign addr[36116]= 1569004214;
assign addr[36117]= 1542643483;
assign addr[36118]= 1515793473;
assign addr[36119]= 1488462700;
assign addr[36120]= 1460659832;
assign addr[36121]= 1432393688;
assign addr[36122]= 1403673233;
assign addr[36123]= 1374507575;
assign addr[36124]= 1344905966;
assign addr[36125]= 1314877795;
assign addr[36126]= 1284432584;
assign addr[36127]= 1253579991;
assign addr[36128]= 1222329801;
assign addr[36129]= 1190691925;
assign addr[36130]= 1158676398;
assign addr[36131]= 1126293375;
assign addr[36132]= 1093553126;
assign addr[36133]= 1060466036;
assign addr[36134]= 1027042599;
assign addr[36135]= 993293415;
assign addr[36136]= 959229189;
assign addr[36137]= 924860725;
assign addr[36138]= 890198924;
assign addr[36139]= 855254778;
assign addr[36140]= 820039373;
assign addr[36141]= 784563876;
assign addr[36142]= 748839539;
assign addr[36143]= 712877694;
assign addr[36144]= 676689746;
assign addr[36145]= 640287172;
assign addr[36146]= 603681519;
assign addr[36147]= 566884397;
assign addr[36148]= 529907477;
assign addr[36149]= 492762486;
assign addr[36150]= 455461206;
assign addr[36151]= 418015468;
assign addr[36152]= 380437148;
assign addr[36153]= 342738165;
assign addr[36154]= 304930476;
assign addr[36155]= 267026072;
assign addr[36156]= 229036977;
assign addr[36157]= 190975237;
assign addr[36158]= 152852926;
assign addr[36159]= 114682135;
assign addr[36160]= 76474970;
assign addr[36161]= 38243550;
assign addr[36162]= 0;
assign addr[36163]= -38243550;
assign addr[36164]= -76474970;
assign addr[36165]= -114682135;
assign addr[36166]= -152852926;
assign addr[36167]= -190975237;
assign addr[36168]= -229036977;
assign addr[36169]= -267026072;
assign addr[36170]= -304930476;
assign addr[36171]= -342738165;
assign addr[36172]= -380437148;
assign addr[36173]= -418015468;
assign addr[36174]= -455461206;
assign addr[36175]= -492762486;
assign addr[36176]= -529907477;
assign addr[36177]= -566884397;
assign addr[36178]= -603681519;
assign addr[36179]= -640287172;
assign addr[36180]= -676689746;
assign addr[36181]= -712877694;
assign addr[36182]= -748839539;
assign addr[36183]= -784563876;
assign addr[36184]= -820039373;
assign addr[36185]= -855254778;
assign addr[36186]= -890198924;
assign addr[36187]= -924860725;
assign addr[36188]= -959229189;
assign addr[36189]= -993293415;
assign addr[36190]= -1027042599;
assign addr[36191]= -1060466036;
assign addr[36192]= -1093553126;
assign addr[36193]= -1126293375;
assign addr[36194]= -1158676398;
assign addr[36195]= -1190691925;
assign addr[36196]= -1222329801;
assign addr[36197]= -1253579991;
assign addr[36198]= -1284432584;
assign addr[36199]= -1314877795;
assign addr[36200]= -1344905966;
assign addr[36201]= -1374507575;
assign addr[36202]= -1403673233;
assign addr[36203]= -1432393688;
assign addr[36204]= -1460659832;
assign addr[36205]= -1488462700;
assign addr[36206]= -1515793473;
assign addr[36207]= -1542643483;
assign addr[36208]= -1569004214;
assign addr[36209]= -1594867305;
assign addr[36210]= -1620224553;
assign addr[36211]= -1645067915;
assign addr[36212]= -1669389513;
assign addr[36213]= -1693181631;
assign addr[36214]= -1716436725;
assign addr[36215]= -1739147417;
assign addr[36216]= -1761306505;
assign addr[36217]= -1782906961;
assign addr[36218]= -1803941934;
assign addr[36219]= -1824404752;
assign addr[36220]= -1844288924;
assign addr[36221]= -1863588145;
assign addr[36222]= -1882296293;
assign addr[36223]= -1900407434;
assign addr[36224]= -1917915825;
assign addr[36225]= -1934815911;
assign addr[36226]= -1951102334;
assign addr[36227]= -1966769926;
assign addr[36228]= -1981813720;
assign addr[36229]= -1996228943;
assign addr[36230]= -2010011024;
assign addr[36231]= -2023155591;
assign addr[36232]= -2035658475;
assign addr[36233]= -2047515711;
assign addr[36234]= -2058723538;
assign addr[36235]= -2069278401;
assign addr[36236]= -2079176953;
assign addr[36237]= -2088416053;
assign addr[36238]= -2096992772;
assign addr[36239]= -2104904390;
assign addr[36240]= -2112148396;
assign addr[36241]= -2118722494;
assign addr[36242]= -2124624598;
assign addr[36243]= -2129852837;
assign addr[36244]= -2134405552;
assign addr[36245]= -2138281298;
assign addr[36246]= -2141478848;
assign addr[36247]= -2143997187;
assign addr[36248]= -2145835515;
assign addr[36249]= -2146993250;
assign addr[36250]= -2147470025;
assign addr[36251]= -2147265689;
assign addr[36252]= -2146380306;
assign addr[36253]= -2144814157;
assign addr[36254]= -2142567738;
assign addr[36255]= -2139641764;
assign addr[36256]= -2136037160;
assign addr[36257]= -2131755071;
assign addr[36258]= -2126796855;
assign addr[36259]= -2121164085;
assign addr[36260]= -2114858546;
assign addr[36261]= -2107882239;
assign addr[36262]= -2100237377;
assign addr[36263]= -2091926384;
assign addr[36264]= -2082951896;
assign addr[36265]= -2073316760;
assign addr[36266]= -2063024031;
assign addr[36267]= -2052076975;
assign addr[36268]= -2040479063;
assign addr[36269]= -2028233973;
assign addr[36270]= -2015345591;
assign addr[36271]= -2001818002;
assign addr[36272]= -1987655498;
assign addr[36273]= -1972862571;
assign addr[36274]= -1957443913;
assign addr[36275]= -1941404413;
assign addr[36276]= -1924749160;
assign addr[36277]= -1907483436;
assign addr[36278]= -1889612716;
assign addr[36279]= -1871142669;
assign addr[36280]= -1852079154;
assign addr[36281]= -1832428215;
assign addr[36282]= -1812196087;
assign addr[36283]= -1791389186;
assign addr[36284]= -1770014111;
assign addr[36285]= -1748077642;
assign addr[36286]= -1725586737;
assign addr[36287]= -1702548529;
assign addr[36288]= -1678970324;
assign addr[36289]= -1654859602;
assign addr[36290]= -1630224009;
assign addr[36291]= -1605071359;
assign addr[36292]= -1579409630;
assign addr[36293]= -1553246960;
assign addr[36294]= -1526591649;
assign addr[36295]= -1499452149;
assign addr[36296]= -1471837070;
assign addr[36297]= -1443755168;
assign addr[36298]= -1415215352;
assign addr[36299]= -1386226674;
assign addr[36300]= -1356798326;
assign addr[36301]= -1326939644;
assign addr[36302]= -1296660098;
assign addr[36303]= -1265969291;
assign addr[36304]= -1234876957;
assign addr[36305]= -1203392958;
assign addr[36306]= -1171527280;
assign addr[36307]= -1139290029;
assign addr[36308]= -1106691431;
assign addr[36309]= -1073741824;
assign addr[36310]= -1040451659;
assign addr[36311]= -1006831495;
assign addr[36312]= -972891995;
assign addr[36313]= -938643924;
assign addr[36314]= -904098143;
assign addr[36315]= -869265610;
assign addr[36316]= -834157373;
assign addr[36317]= -798784567;
assign addr[36318]= -763158411;
assign addr[36319]= -727290205;
assign addr[36320]= -691191324;
assign addr[36321]= -654873219;
assign addr[36322]= -618347408;
assign addr[36323]= -581625477;
assign addr[36324]= -544719071;
assign addr[36325]= -507639898;
assign addr[36326]= -470399716;
assign addr[36327]= -433010339;
assign addr[36328]= -395483624;
assign addr[36329]= -357831473;
assign addr[36330]= -320065829;
assign addr[36331]= -282198671;
assign addr[36332]= -244242007;
assign addr[36333]= -206207878;
assign addr[36334]= -168108346;
assign addr[36335]= -129955495;
assign addr[36336]= -91761426;
assign addr[36337]= -53538253;
assign addr[36338]= -15298099;
assign addr[36339]= 22946906;
assign addr[36340]= 61184634;
assign addr[36341]= 99402956;
assign addr[36342]= 137589750;
assign addr[36343]= 175732905;
assign addr[36344]= 213820322;
assign addr[36345]= 251839923;
assign addr[36346]= 289779648;
assign addr[36347]= 327627463;
assign addr[36348]= 365371365;
assign addr[36349]= 402999383;
assign addr[36350]= 440499581;
assign addr[36351]= 477860067;
assign addr[36352]= 515068990;
assign addr[36353]= 552114549;
assign addr[36354]= 588984994;
assign addr[36355]= 625668632;
assign addr[36356]= 662153826;
assign addr[36357]= 698429006;
assign addr[36358]= 734482665;
assign addr[36359]= 770303369;
assign addr[36360]= 805879757;
assign addr[36361]= 841200544;
assign addr[36362]= 876254528;
assign addr[36363]= 911030591;
assign addr[36364]= 945517704;
assign addr[36365]= 979704927;
assign addr[36366]= 1013581418;
assign addr[36367]= 1047136432;
assign addr[36368]= 1080359326;
assign addr[36369]= 1113239564;
assign addr[36370]= 1145766716;
assign addr[36371]= 1177930466;
assign addr[36372]= 1209720613;
assign addr[36373]= 1241127074;
assign addr[36374]= 1272139887;
assign addr[36375]= 1302749217;
assign addr[36376]= 1332945355;
assign addr[36377]= 1362718723;
assign addr[36378]= 1392059879;
assign addr[36379]= 1420959516;
assign addr[36380]= 1449408469;
assign addr[36381]= 1477397714;
assign addr[36382]= 1504918373;
assign addr[36383]= 1531961719;
assign addr[36384]= 1558519173;
assign addr[36385]= 1584582314;
assign addr[36386]= 1610142873;
assign addr[36387]= 1635192744;
assign addr[36388]= 1659723983;
assign addr[36389]= 1683728808;
assign addr[36390]= 1707199606;
assign addr[36391]= 1730128933;
assign addr[36392]= 1752509516;
assign addr[36393]= 1774334257;
assign addr[36394]= 1795596234;
assign addr[36395]= 1816288703;
assign addr[36396]= 1836405100;
assign addr[36397]= 1855939047;
assign addr[36398]= 1874884346;
assign addr[36399]= 1893234990;
assign addr[36400]= 1910985158;
assign addr[36401]= 1928129220;
assign addr[36402]= 1944661739;
assign addr[36403]= 1960577471;
assign addr[36404]= 1975871368;
assign addr[36405]= 1990538579;
assign addr[36406]= 2004574453;
assign addr[36407]= 2017974537;
assign addr[36408]= 2030734582;
assign addr[36409]= 2042850540;
assign addr[36410]= 2054318569;
assign addr[36411]= 2065135031;
assign addr[36412]= 2075296495;
assign addr[36413]= 2084799740;
assign addr[36414]= 2093641749;
assign addr[36415]= 2101819720;
assign addr[36416]= 2109331059;
assign addr[36417]= 2116173382;
assign addr[36418]= 2122344521;
assign addr[36419]= 2127842516;
assign addr[36420]= 2132665626;
assign addr[36421]= 2136812319;
assign addr[36422]= 2140281282;
assign addr[36423]= 2143071413;
assign addr[36424]= 2145181827;
assign addr[36425]= 2146611856;
assign addr[36426]= 2147361045;
assign addr[36427]= 2147429158;
assign addr[36428]= 2146816171;
assign addr[36429]= 2145522281;
assign addr[36430]= 2143547897;
assign addr[36431]= 2140893646;
assign addr[36432]= 2137560369;
assign addr[36433]= 2133549123;
assign addr[36434]= 2128861181;
assign addr[36435]= 2123498030;
assign addr[36436]= 2117461370;
assign addr[36437]= 2110753117;
assign addr[36438]= 2103375398;
assign addr[36439]= 2095330553;
assign addr[36440]= 2086621133;
assign addr[36441]= 2077249901;
assign addr[36442]= 2067219829;
assign addr[36443]= 2056534099;
assign addr[36444]= 2045196100;
assign addr[36445]= 2033209426;
assign addr[36446]= 2020577882;
assign addr[36447]= 2007305472;
assign addr[36448]= 1993396407;
assign addr[36449]= 1978855097;
assign addr[36450]= 1963686155;
assign addr[36451]= 1947894393;
assign addr[36452]= 1931484818;
assign addr[36453]= 1914462636;
assign addr[36454]= 1896833245;
assign addr[36455]= 1878602237;
assign addr[36456]= 1859775393;
assign addr[36457]= 1840358687;
assign addr[36458]= 1820358275;
assign addr[36459]= 1799780501;
assign addr[36460]= 1778631892;
assign addr[36461]= 1756919156;
assign addr[36462]= 1734649179;
assign addr[36463]= 1711829025;
assign addr[36464]= 1688465931;
assign addr[36465]= 1664567307;
assign addr[36466]= 1640140734;
assign addr[36467]= 1615193959;
assign addr[36468]= 1589734894;
assign addr[36469]= 1563771613;
assign addr[36470]= 1537312353;
assign addr[36471]= 1510365504;
assign addr[36472]= 1482939614;
assign addr[36473]= 1455043381;
assign addr[36474]= 1426685652;
assign addr[36475]= 1397875423;
assign addr[36476]= 1368621831;
assign addr[36477]= 1338934154;
assign addr[36478]= 1308821808;
assign addr[36479]= 1278294345;
assign addr[36480]= 1247361445;
assign addr[36481]= 1216032921;
assign addr[36482]= 1184318708;
assign addr[36483]= 1152228866;
assign addr[36484]= 1119773573;
assign addr[36485]= 1086963121;
assign addr[36486]= 1053807919;
assign addr[36487]= 1020318481;
assign addr[36488]= 986505429;
assign addr[36489]= 952379488;
assign addr[36490]= 917951481;
assign addr[36491]= 883232329;
assign addr[36492]= 848233042;
assign addr[36493]= 812964722;
assign addr[36494]= 777438554;
assign addr[36495]= 741665807;
assign addr[36496]= 705657826;
assign addr[36497]= 669426032;
assign addr[36498]= 632981917;
assign addr[36499]= 596337040;
assign addr[36500]= 559503022;
assign addr[36501]= 522491548;
assign addr[36502]= 485314355;
assign addr[36503]= 447983235;
assign addr[36504]= 410510029;
assign addr[36505]= 372906622;
assign addr[36506]= 335184940;
assign addr[36507]= 297356948;
assign addr[36508]= 259434643;
assign addr[36509]= 221430054;
assign addr[36510]= 183355234;
assign addr[36511]= 145222259;
assign addr[36512]= 107043224;
assign addr[36513]= 68830239;
assign addr[36514]= 30595422;
assign addr[36515]= -7649098;
assign addr[36516]= -45891193;
assign addr[36517]= -84118732;
assign addr[36518]= -122319591;
assign addr[36519]= -160481654;
assign addr[36520]= -198592817;
assign addr[36521]= -236640993;
assign addr[36522]= -274614114;
assign addr[36523]= -312500135;
assign addr[36524]= -350287041;
assign addr[36525]= -387962847;
assign addr[36526]= -425515602;
assign addr[36527]= -462933398;
assign addr[36528]= -500204365;
assign addr[36529]= -537316682;
assign addr[36530]= -574258580;
assign addr[36531]= -611018340;
assign addr[36532]= -647584304;
assign addr[36533]= -683944874;
assign addr[36534]= -720088517;
assign addr[36535]= -756003771;
assign addr[36536]= -791679244;
assign addr[36537]= -827103620;
assign addr[36538]= -862265664;
assign addr[36539]= -897154224;
assign addr[36540]= -931758235;
assign addr[36541]= -966066720;
assign addr[36542]= -1000068799;
assign addr[36543]= -1033753687;
assign addr[36544]= -1067110699;
assign addr[36545]= -1100129257;
assign addr[36546]= -1132798888;
assign addr[36547]= -1165109230;
assign addr[36548]= -1197050035;
assign addr[36549]= -1228611172;
assign addr[36550]= -1259782632;
assign addr[36551]= -1290554528;
assign addr[36552]= -1320917099;
assign addr[36553]= -1350860716;
assign addr[36554]= -1380375881;
assign addr[36555]= -1409453233;
assign addr[36556]= -1438083551;
assign addr[36557]= -1466257752;
assign addr[36558]= -1493966902;
assign addr[36559]= -1521202211;
assign addr[36560]= -1547955041;
assign addr[36561]= -1574216908;
assign addr[36562]= -1599979481;
assign addr[36563]= -1625234591;
assign addr[36564]= -1649974225;
assign addr[36565]= -1674190539;
assign addr[36566]= -1697875851;
assign addr[36567]= -1721022648;
assign addr[36568]= -1743623590;
assign addr[36569]= -1765671509;
assign addr[36570]= -1787159411;
assign addr[36571]= -1808080480;
assign addr[36572]= -1828428082;
assign addr[36573]= -1848195763;
assign addr[36574]= -1867377253;
assign addr[36575]= -1885966468;
assign addr[36576]= -1903957513;
assign addr[36577]= -1921344681;
assign addr[36578]= -1938122457;
assign addr[36579]= -1954285520;
assign addr[36580]= -1969828744;
assign addr[36581]= -1984747199;
assign addr[36582]= -1999036154;
assign addr[36583]= -2012691075;
assign addr[36584]= -2025707632;
assign addr[36585]= -2038081698;
assign addr[36586]= -2049809346;
assign addr[36587]= -2060886858;
assign addr[36588]= -2071310720;
assign addr[36589]= -2081077626;
assign addr[36590]= -2090184478;
assign addr[36591]= -2098628387;
assign addr[36592]= -2106406677;
assign addr[36593]= -2113516878;
assign addr[36594]= -2119956737;
assign addr[36595]= -2125724211;
assign addr[36596]= -2130817471;
assign addr[36597]= -2135234901;
assign addr[36598]= -2138975100;
assign addr[36599]= -2142036881;
assign addr[36600]= -2144419275;
assign addr[36601]= -2146121524;
assign addr[36602]= -2147143090;
assign addr[36603]= -2147483648;
assign addr[36604]= -2147143090;
assign addr[36605]= -2146121524;
assign addr[36606]= -2144419275;
assign addr[36607]= -2142036881;
assign addr[36608]= -2138975100;
assign addr[36609]= -2135234901;
assign addr[36610]= -2130817471;
assign addr[36611]= -2125724211;
assign addr[36612]= -2119956737;
assign addr[36613]= -2113516878;
assign addr[36614]= -2106406677;
assign addr[36615]= -2098628387;
assign addr[36616]= -2090184478;
assign addr[36617]= -2081077626;
assign addr[36618]= -2071310720;
assign addr[36619]= -2060886858;
assign addr[36620]= -2049809346;
assign addr[36621]= -2038081698;
assign addr[36622]= -2025707632;
assign addr[36623]= -2012691075;
assign addr[36624]= -1999036154;
assign addr[36625]= -1984747199;
assign addr[36626]= -1969828744;
assign addr[36627]= -1954285520;
assign addr[36628]= -1938122457;
assign addr[36629]= -1921344681;
assign addr[36630]= -1903957513;
assign addr[36631]= -1885966468;
assign addr[36632]= -1867377253;
assign addr[36633]= -1848195763;
assign addr[36634]= -1828428082;
assign addr[36635]= -1808080480;
assign addr[36636]= -1787159411;
assign addr[36637]= -1765671509;
assign addr[36638]= -1743623590;
assign addr[36639]= -1721022648;
assign addr[36640]= -1697875851;
assign addr[36641]= -1674190539;
assign addr[36642]= -1649974225;
assign addr[36643]= -1625234591;
assign addr[36644]= -1599979481;
assign addr[36645]= -1574216908;
assign addr[36646]= -1547955041;
assign addr[36647]= -1521202211;
assign addr[36648]= -1493966902;
assign addr[36649]= -1466257752;
assign addr[36650]= -1438083551;
assign addr[36651]= -1409453233;
assign addr[36652]= -1380375881;
assign addr[36653]= -1350860716;
assign addr[36654]= -1320917099;
assign addr[36655]= -1290554528;
assign addr[36656]= -1259782632;
assign addr[36657]= -1228611172;
assign addr[36658]= -1197050035;
assign addr[36659]= -1165109230;
assign addr[36660]= -1132798888;
assign addr[36661]= -1100129257;
assign addr[36662]= -1067110699;
assign addr[36663]= -1033753687;
assign addr[36664]= -1000068799;
assign addr[36665]= -966066720;
assign addr[36666]= -931758235;
assign addr[36667]= -897154224;
assign addr[36668]= -862265664;
assign addr[36669]= -827103620;
assign addr[36670]= -791679244;
assign addr[36671]= -756003771;
assign addr[36672]= -720088517;
assign addr[36673]= -683944874;
assign addr[36674]= -647584304;
assign addr[36675]= -611018340;
assign addr[36676]= -574258580;
assign addr[36677]= -537316682;
assign addr[36678]= -500204365;
assign addr[36679]= -462933398;
assign addr[36680]= -425515602;
assign addr[36681]= -387962847;
assign addr[36682]= -350287041;
assign addr[36683]= -312500135;
assign addr[36684]= -274614114;
assign addr[36685]= -236640993;
assign addr[36686]= -198592817;
assign addr[36687]= -160481654;
assign addr[36688]= -122319591;
assign addr[36689]= -84118732;
assign addr[36690]= -45891193;
assign addr[36691]= -7649098;
assign addr[36692]= 30595422;
assign addr[36693]= 68830239;
assign addr[36694]= 107043224;
assign addr[36695]= 145222259;
assign addr[36696]= 183355234;
assign addr[36697]= 221430054;
assign addr[36698]= 259434643;
assign addr[36699]= 297356948;
assign addr[36700]= 335184940;
assign addr[36701]= 372906622;
assign addr[36702]= 410510029;
assign addr[36703]= 447983235;
assign addr[36704]= 485314355;
assign addr[36705]= 522491548;
assign addr[36706]= 559503022;
assign addr[36707]= 596337040;
assign addr[36708]= 632981917;
assign addr[36709]= 669426032;
assign addr[36710]= 705657826;
assign addr[36711]= 741665807;
assign addr[36712]= 777438554;
assign addr[36713]= 812964722;
assign addr[36714]= 848233042;
assign addr[36715]= 883232329;
assign addr[36716]= 917951481;
assign addr[36717]= 952379488;
assign addr[36718]= 986505429;
assign addr[36719]= 1020318481;
assign addr[36720]= 1053807919;
assign addr[36721]= 1086963121;
assign addr[36722]= 1119773573;
assign addr[36723]= 1152228866;
assign addr[36724]= 1184318708;
assign addr[36725]= 1216032921;
assign addr[36726]= 1247361445;
assign addr[36727]= 1278294345;
assign addr[36728]= 1308821808;
assign addr[36729]= 1338934154;
assign addr[36730]= 1368621831;
assign addr[36731]= 1397875423;
assign addr[36732]= 1426685652;
assign addr[36733]= 1455043381;
assign addr[36734]= 1482939614;
assign addr[36735]= 1510365504;
assign addr[36736]= 1537312353;
assign addr[36737]= 1563771613;
assign addr[36738]= 1589734894;
assign addr[36739]= 1615193959;
assign addr[36740]= 1640140734;
assign addr[36741]= 1664567307;
assign addr[36742]= 1688465931;
assign addr[36743]= 1711829025;
assign addr[36744]= 1734649179;
assign addr[36745]= 1756919156;
assign addr[36746]= 1778631892;
assign addr[36747]= 1799780501;
assign addr[36748]= 1820358275;
assign addr[36749]= 1840358687;
assign addr[36750]= 1859775393;
assign addr[36751]= 1878602237;
assign addr[36752]= 1896833245;
assign addr[36753]= 1914462636;
assign addr[36754]= 1931484818;
assign addr[36755]= 1947894393;
assign addr[36756]= 1963686155;
assign addr[36757]= 1978855097;
assign addr[36758]= 1993396407;
assign addr[36759]= 2007305472;
assign addr[36760]= 2020577882;
assign addr[36761]= 2033209426;
assign addr[36762]= 2045196100;
assign addr[36763]= 2056534099;
assign addr[36764]= 2067219829;
assign addr[36765]= 2077249901;
assign addr[36766]= 2086621133;
assign addr[36767]= 2095330553;
assign addr[36768]= 2103375398;
assign addr[36769]= 2110753117;
assign addr[36770]= 2117461370;
assign addr[36771]= 2123498030;
assign addr[36772]= 2128861181;
assign addr[36773]= 2133549123;
assign addr[36774]= 2137560369;
assign addr[36775]= 2140893646;
assign addr[36776]= 2143547897;
assign addr[36777]= 2145522281;
assign addr[36778]= 2146816171;
assign addr[36779]= 2147429158;
assign addr[36780]= 2147361045;
assign addr[36781]= 2146611856;
assign addr[36782]= 2145181827;
assign addr[36783]= 2143071413;
assign addr[36784]= 2140281282;
assign addr[36785]= 2136812319;
assign addr[36786]= 2132665626;
assign addr[36787]= 2127842516;
assign addr[36788]= 2122344521;
assign addr[36789]= 2116173382;
assign addr[36790]= 2109331059;
assign addr[36791]= 2101819720;
assign addr[36792]= 2093641749;
assign addr[36793]= 2084799740;
assign addr[36794]= 2075296495;
assign addr[36795]= 2065135031;
assign addr[36796]= 2054318569;
assign addr[36797]= 2042850540;
assign addr[36798]= 2030734582;
assign addr[36799]= 2017974537;
assign addr[36800]= 2004574453;
assign addr[36801]= 1990538579;
assign addr[36802]= 1975871368;
assign addr[36803]= 1960577471;
assign addr[36804]= 1944661739;
assign addr[36805]= 1928129220;
assign addr[36806]= 1910985158;
assign addr[36807]= 1893234990;
assign addr[36808]= 1874884346;
assign addr[36809]= 1855939047;
assign addr[36810]= 1836405100;
assign addr[36811]= 1816288703;
assign addr[36812]= 1795596234;
assign addr[36813]= 1774334257;
assign addr[36814]= 1752509516;
assign addr[36815]= 1730128933;
assign addr[36816]= 1707199606;
assign addr[36817]= 1683728808;
assign addr[36818]= 1659723983;
assign addr[36819]= 1635192744;
assign addr[36820]= 1610142873;
assign addr[36821]= 1584582314;
assign addr[36822]= 1558519173;
assign addr[36823]= 1531961719;
assign addr[36824]= 1504918373;
assign addr[36825]= 1477397714;
assign addr[36826]= 1449408469;
assign addr[36827]= 1420959516;
assign addr[36828]= 1392059879;
assign addr[36829]= 1362718723;
assign addr[36830]= 1332945355;
assign addr[36831]= 1302749217;
assign addr[36832]= 1272139887;
assign addr[36833]= 1241127074;
assign addr[36834]= 1209720613;
assign addr[36835]= 1177930466;
assign addr[36836]= 1145766716;
assign addr[36837]= 1113239564;
assign addr[36838]= 1080359326;
assign addr[36839]= 1047136432;
assign addr[36840]= 1013581418;
assign addr[36841]= 979704927;
assign addr[36842]= 945517704;
assign addr[36843]= 911030591;
assign addr[36844]= 876254528;
assign addr[36845]= 841200544;
assign addr[36846]= 805879757;
assign addr[36847]= 770303369;
assign addr[36848]= 734482665;
assign addr[36849]= 698429006;
assign addr[36850]= 662153826;
assign addr[36851]= 625668632;
assign addr[36852]= 588984994;
assign addr[36853]= 552114549;
assign addr[36854]= 515068990;
assign addr[36855]= 477860067;
assign addr[36856]= 440499581;
assign addr[36857]= 402999383;
assign addr[36858]= 365371365;
assign addr[36859]= 327627463;
assign addr[36860]= 289779648;
assign addr[36861]= 251839923;
assign addr[36862]= 213820322;
assign addr[36863]= 175732905;
assign addr[36864]= 137589750;
assign addr[36865]= 99402956;
assign addr[36866]= 61184634;
assign addr[36867]= 22946906;
assign addr[36868]= -15298099;
assign addr[36869]= -53538253;
assign addr[36870]= -91761426;
assign addr[36871]= -129955495;
assign addr[36872]= -168108346;
assign addr[36873]= -206207878;
assign addr[36874]= -244242007;
assign addr[36875]= -282198671;
assign addr[36876]= -320065829;
assign addr[36877]= -357831473;
assign addr[36878]= -395483624;
assign addr[36879]= -433010339;
assign addr[36880]= -470399716;
assign addr[36881]= -507639898;
assign addr[36882]= -544719071;
assign addr[36883]= -581625477;
assign addr[36884]= -618347408;
assign addr[36885]= -654873219;
assign addr[36886]= -691191324;
assign addr[36887]= -727290205;
assign addr[36888]= -763158411;
assign addr[36889]= -798784567;
assign addr[36890]= -834157373;
assign addr[36891]= -869265610;
assign addr[36892]= -904098143;
assign addr[36893]= -938643924;
assign addr[36894]= -972891995;
assign addr[36895]= -1006831495;
assign addr[36896]= -1040451659;
assign addr[36897]= -1073741824;
assign addr[36898]= -1106691431;
assign addr[36899]= -1139290029;
assign addr[36900]= -1171527280;
assign addr[36901]= -1203392958;
assign addr[36902]= -1234876957;
assign addr[36903]= -1265969291;
assign addr[36904]= -1296660098;
assign addr[36905]= -1326939644;
assign addr[36906]= -1356798326;
assign addr[36907]= -1386226674;
assign addr[36908]= -1415215352;
assign addr[36909]= -1443755168;
assign addr[36910]= -1471837070;
assign addr[36911]= -1499452149;
assign addr[36912]= -1526591649;
assign addr[36913]= -1553246960;
assign addr[36914]= -1579409630;
assign addr[36915]= -1605071359;
assign addr[36916]= -1630224009;
assign addr[36917]= -1654859602;
assign addr[36918]= -1678970324;
assign addr[36919]= -1702548529;
assign addr[36920]= -1725586737;
assign addr[36921]= -1748077642;
assign addr[36922]= -1770014111;
assign addr[36923]= -1791389186;
assign addr[36924]= -1812196087;
assign addr[36925]= -1832428215;
assign addr[36926]= -1852079154;
assign addr[36927]= -1871142669;
assign addr[36928]= -1889612716;
assign addr[36929]= -1907483436;
assign addr[36930]= -1924749160;
assign addr[36931]= -1941404413;
assign addr[36932]= -1957443913;
assign addr[36933]= -1972862571;
assign addr[36934]= -1987655498;
assign addr[36935]= -2001818002;
assign addr[36936]= -2015345591;
assign addr[36937]= -2028233973;
assign addr[36938]= -2040479063;
assign addr[36939]= -2052076975;
assign addr[36940]= -2063024031;
assign addr[36941]= -2073316760;
assign addr[36942]= -2082951896;
assign addr[36943]= -2091926384;
assign addr[36944]= -2100237377;
assign addr[36945]= -2107882239;
assign addr[36946]= -2114858546;
assign addr[36947]= -2121164085;
assign addr[36948]= -2126796855;
assign addr[36949]= -2131755071;
assign addr[36950]= -2136037160;
assign addr[36951]= -2139641764;
assign addr[36952]= -2142567738;
assign addr[36953]= -2144814157;
assign addr[36954]= -2146380306;
assign addr[36955]= -2147265689;
assign addr[36956]= -2147470025;
assign addr[36957]= -2146993250;
assign addr[36958]= -2145835515;
assign addr[36959]= -2143997187;
assign addr[36960]= -2141478848;
assign addr[36961]= -2138281298;
assign addr[36962]= -2134405552;
assign addr[36963]= -2129852837;
assign addr[36964]= -2124624598;
assign addr[36965]= -2118722494;
assign addr[36966]= -2112148396;
assign addr[36967]= -2104904390;
assign addr[36968]= -2096992772;
assign addr[36969]= -2088416053;
assign addr[36970]= -2079176953;
assign addr[36971]= -2069278401;
assign addr[36972]= -2058723538;
assign addr[36973]= -2047515711;
assign addr[36974]= -2035658475;
assign addr[36975]= -2023155591;
assign addr[36976]= -2010011024;
assign addr[36977]= -1996228943;
assign addr[36978]= -1981813720;
assign addr[36979]= -1966769926;
assign addr[36980]= -1951102334;
assign addr[36981]= -1934815911;
assign addr[36982]= -1917915825;
assign addr[36983]= -1900407434;
assign addr[36984]= -1882296293;
assign addr[36985]= -1863588145;
assign addr[36986]= -1844288924;
assign addr[36987]= -1824404752;
assign addr[36988]= -1803941934;
assign addr[36989]= -1782906961;
assign addr[36990]= -1761306505;
assign addr[36991]= -1739147417;
assign addr[36992]= -1716436725;
assign addr[36993]= -1693181631;
assign addr[36994]= -1669389513;
assign addr[36995]= -1645067915;
assign addr[36996]= -1620224553;
assign addr[36997]= -1594867305;
assign addr[36998]= -1569004214;
assign addr[36999]= -1542643483;
assign addr[37000]= -1515793473;
assign addr[37001]= -1488462700;
assign addr[37002]= -1460659832;
assign addr[37003]= -1432393688;
assign addr[37004]= -1403673233;
assign addr[37005]= -1374507575;
assign addr[37006]= -1344905966;
assign addr[37007]= -1314877795;
assign addr[37008]= -1284432584;
assign addr[37009]= -1253579991;
assign addr[37010]= -1222329801;
assign addr[37011]= -1190691925;
assign addr[37012]= -1158676398;
assign addr[37013]= -1126293375;
assign addr[37014]= -1093553126;
assign addr[37015]= -1060466036;
assign addr[37016]= -1027042599;
assign addr[37017]= -993293415;
assign addr[37018]= -959229189;
assign addr[37019]= -924860725;
assign addr[37020]= -890198924;
assign addr[37021]= -855254778;
assign addr[37022]= -820039373;
assign addr[37023]= -784563876;
assign addr[37024]= -748839539;
assign addr[37025]= -712877694;
assign addr[37026]= -676689746;
assign addr[37027]= -640287172;
assign addr[37028]= -603681519;
assign addr[37029]= -566884397;
assign addr[37030]= -529907477;
assign addr[37031]= -492762486;
assign addr[37032]= -455461206;
assign addr[37033]= -418015468;
assign addr[37034]= -380437148;
assign addr[37035]= -342738165;
assign addr[37036]= -304930476;
assign addr[37037]= -267026072;
assign addr[37038]= -229036977;
assign addr[37039]= -190975237;
assign addr[37040]= -152852926;
assign addr[37041]= -114682135;
assign addr[37042]= -76474970;
assign addr[37043]= -38243550;
assign addr[37044]= 0;
assign addr[37045]= 38243550;
assign addr[37046]= 76474970;
assign addr[37047]= 114682135;
assign addr[37048]= 152852926;
assign addr[37049]= 190975237;
assign addr[37050]= 229036977;
assign addr[37051]= 267026072;
assign addr[37052]= 304930476;
assign addr[37053]= 342738165;
assign addr[37054]= 380437148;
assign addr[37055]= 418015468;
assign addr[37056]= 455461206;
assign addr[37057]= 492762486;
assign addr[37058]= 529907477;
assign addr[37059]= 566884397;
assign addr[37060]= 603681519;
assign addr[37061]= 640287172;
assign addr[37062]= 676689746;
assign addr[37063]= 712877694;
assign addr[37064]= 748839539;
assign addr[37065]= 784563876;
assign addr[37066]= 820039373;
assign addr[37067]= 855254778;
assign addr[37068]= 890198924;
assign addr[37069]= 924860725;
assign addr[37070]= 959229189;
assign addr[37071]= 993293415;
assign addr[37072]= 1027042599;
assign addr[37073]= 1060466036;
assign addr[37074]= 1093553126;
assign addr[37075]= 1126293375;
assign addr[37076]= 1158676398;
assign addr[37077]= 1190691925;
assign addr[37078]= 1222329801;
assign addr[37079]= 1253579991;
assign addr[37080]= 1284432584;
assign addr[37081]= 1314877795;
assign addr[37082]= 1344905966;
assign addr[37083]= 1374507575;
assign addr[37084]= 1403673233;
assign addr[37085]= 1432393688;
assign addr[37086]= 1460659832;
assign addr[37087]= 1488462700;
assign addr[37088]= 1515793473;
assign addr[37089]= 1542643483;
assign addr[37090]= 1569004214;
assign addr[37091]= 1594867305;
assign addr[37092]= 1620224553;
assign addr[37093]= 1645067915;
assign addr[37094]= 1669389513;
assign addr[37095]= 1693181631;
assign addr[37096]= 1716436725;
assign addr[37097]= 1739147417;
assign addr[37098]= 1761306505;
assign addr[37099]= 1782906961;
assign addr[37100]= 1803941934;
assign addr[37101]= 1824404752;
assign addr[37102]= 1844288924;
assign addr[37103]= 1863588145;
assign addr[37104]= 1882296293;
assign addr[37105]= 1900407434;
assign addr[37106]= 1917915825;
assign addr[37107]= 1934815911;
assign addr[37108]= 1951102334;
assign addr[37109]= 1966769926;
assign addr[37110]= 1981813720;
assign addr[37111]= 1996228943;
assign addr[37112]= 2010011024;
assign addr[37113]= 2023155591;
assign addr[37114]= 2035658475;
assign addr[37115]= 2047515711;
assign addr[37116]= 2058723538;
assign addr[37117]= 2069278401;
assign addr[37118]= 2079176953;
assign addr[37119]= 2088416053;
assign addr[37120]= 2096992772;
assign addr[37121]= 2104904390;
assign addr[37122]= 2112148396;
assign addr[37123]= 2118722494;
assign addr[37124]= 2124624598;
assign addr[37125]= 2129852837;
assign addr[37126]= 2134405552;
assign addr[37127]= 2138281298;
assign addr[37128]= 2141478848;
assign addr[37129]= 2143997187;
assign addr[37130]= 2145835515;
assign addr[37131]= 2146993250;
assign addr[37132]= 2147470025;
assign addr[37133]= 2147265689;
assign addr[37134]= 2146380306;
assign addr[37135]= 2144814157;
assign addr[37136]= 2142567738;
assign addr[37137]= 2139641764;
assign addr[37138]= 2136037160;
assign addr[37139]= 2131755071;
assign addr[37140]= 2126796855;
assign addr[37141]= 2121164085;
assign addr[37142]= 2114858546;
assign addr[37143]= 2107882239;
assign addr[37144]= 2100237377;
assign addr[37145]= 2091926384;
assign addr[37146]= 2082951896;
assign addr[37147]= 2073316760;
assign addr[37148]= 2063024031;
assign addr[37149]= 2052076975;
assign addr[37150]= 2040479063;
assign addr[37151]= 2028233973;
assign addr[37152]= 2015345591;
assign addr[37153]= 2001818002;
assign addr[37154]= 1987655498;
assign addr[37155]= 1972862571;
assign addr[37156]= 1957443913;
assign addr[37157]= 1941404413;
assign addr[37158]= 1924749160;
assign addr[37159]= 1907483436;
assign addr[37160]= 1889612716;
assign addr[37161]= 1871142669;
assign addr[37162]= 1852079154;
assign addr[37163]= 1832428215;
assign addr[37164]= 1812196087;
assign addr[37165]= 1791389186;
assign addr[37166]= 1770014111;
assign addr[37167]= 1748077642;
assign addr[37168]= 1725586737;
assign addr[37169]= 1702548529;
assign addr[37170]= 1678970324;
assign addr[37171]= 1654859602;
assign addr[37172]= 1630224009;
assign addr[37173]= 1605071359;
assign addr[37174]= 1579409630;
assign addr[37175]= 1553246960;
assign addr[37176]= 1526591649;
assign addr[37177]= 1499452149;
assign addr[37178]= 1471837070;
assign addr[37179]= 1443755168;
assign addr[37180]= 1415215352;
assign addr[37181]= 1386226674;
assign addr[37182]= 1356798326;
assign addr[37183]= 1326939644;
assign addr[37184]= 1296660098;
assign addr[37185]= 1265969291;
assign addr[37186]= 1234876957;
assign addr[37187]= 1203392958;
assign addr[37188]= 1171527280;
assign addr[37189]= 1139290029;
assign addr[37190]= 1106691431;
assign addr[37191]= 1073741824;
assign addr[37192]= 1040451659;
assign addr[37193]= 1006831495;
assign addr[37194]= 972891995;
assign addr[37195]= 938643924;
assign addr[37196]= 904098143;
assign addr[37197]= 869265610;
assign addr[37198]= 834157373;
assign addr[37199]= 798784567;
assign addr[37200]= 763158411;
assign addr[37201]= 727290205;
assign addr[37202]= 691191324;
assign addr[37203]= 654873219;
assign addr[37204]= 618347408;
assign addr[37205]= 581625477;
assign addr[37206]= 544719071;
assign addr[37207]= 507639898;
assign addr[37208]= 470399716;
assign addr[37209]= 433010339;
assign addr[37210]= 395483624;
assign addr[37211]= 357831473;
assign addr[37212]= 320065829;
assign addr[37213]= 282198671;
assign addr[37214]= 244242007;
assign addr[37215]= 206207878;
assign addr[37216]= 168108346;
assign addr[37217]= 129955495;
assign addr[37218]= 91761426;
assign addr[37219]= 53538253;
assign addr[37220]= 15298099;
assign addr[37221]= -22946906;
assign addr[37222]= -61184634;
assign addr[37223]= -99402956;
assign addr[37224]= -137589750;
assign addr[37225]= -175732905;
assign addr[37226]= -213820322;
assign addr[37227]= -251839923;
assign addr[37228]= -289779648;
assign addr[37229]= -327627463;
assign addr[37230]= -365371365;
assign addr[37231]= -402999383;
assign addr[37232]= -440499581;
assign addr[37233]= -477860067;
assign addr[37234]= -515068990;
assign addr[37235]= -552114549;
assign addr[37236]= -588984994;
assign addr[37237]= -625668632;
assign addr[37238]= -662153826;
assign addr[37239]= -698429006;
assign addr[37240]= -734482665;
assign addr[37241]= -770303369;
assign addr[37242]= -805879757;
assign addr[37243]= -841200544;
assign addr[37244]= -876254528;
assign addr[37245]= -911030591;
assign addr[37246]= -945517704;
assign addr[37247]= -979704927;
assign addr[37248]= -1013581418;
assign addr[37249]= -1047136432;
assign addr[37250]= -1080359326;
assign addr[37251]= -1113239564;
assign addr[37252]= -1145766716;
assign addr[37253]= -1177930466;
assign addr[37254]= -1209720613;
assign addr[37255]= -1241127074;
assign addr[37256]= -1272139887;
assign addr[37257]= -1302749217;
assign addr[37258]= -1332945355;
assign addr[37259]= -1362718723;
assign addr[37260]= -1392059879;
assign addr[37261]= -1420959516;
assign addr[37262]= -1449408469;
assign addr[37263]= -1477397714;
assign addr[37264]= -1504918373;
assign addr[37265]= -1531961719;
assign addr[37266]= -1558519173;
assign addr[37267]= -1584582314;
assign addr[37268]= -1610142873;
assign addr[37269]= -1635192744;
assign addr[37270]= -1659723983;
assign addr[37271]= -1683728808;
assign addr[37272]= -1707199606;
assign addr[37273]= -1730128933;
assign addr[37274]= -1752509516;
assign addr[37275]= -1774334257;
assign addr[37276]= -1795596234;
assign addr[37277]= -1816288703;
assign addr[37278]= -1836405100;
assign addr[37279]= -1855939047;
assign addr[37280]= -1874884346;
assign addr[37281]= -1893234990;
assign addr[37282]= -1910985158;
assign addr[37283]= -1928129220;
assign addr[37284]= -1944661739;
assign addr[37285]= -1960577471;
assign addr[37286]= -1975871368;
assign addr[37287]= -1990538579;
assign addr[37288]= -2004574453;
assign addr[37289]= -2017974537;
assign addr[37290]= -2030734582;
assign addr[37291]= -2042850540;
assign addr[37292]= -2054318569;
assign addr[37293]= -2065135031;
assign addr[37294]= -2075296495;
assign addr[37295]= -2084799740;
assign addr[37296]= -2093641749;
assign addr[37297]= -2101819720;
assign addr[37298]= -2109331059;
assign addr[37299]= -2116173382;
assign addr[37300]= -2122344521;
assign addr[37301]= -2127842516;
assign addr[37302]= -2132665626;
assign addr[37303]= -2136812319;
assign addr[37304]= -2140281282;
assign addr[37305]= -2143071413;
assign addr[37306]= -2145181827;
assign addr[37307]= -2146611856;
assign addr[37308]= -2147361045;
assign addr[37309]= -2147429158;
assign addr[37310]= -2146816171;
assign addr[37311]= -2145522281;
assign addr[37312]= -2143547897;
assign addr[37313]= -2140893646;
assign addr[37314]= -2137560369;
assign addr[37315]= -2133549123;
assign addr[37316]= -2128861181;
assign addr[37317]= -2123498030;
assign addr[37318]= -2117461370;
assign addr[37319]= -2110753117;
assign addr[37320]= -2103375398;
assign addr[37321]= -2095330553;
assign addr[37322]= -2086621133;
assign addr[37323]= -2077249901;
assign addr[37324]= -2067219829;
assign addr[37325]= -2056534099;
assign addr[37326]= -2045196100;
assign addr[37327]= -2033209426;
assign addr[37328]= -2020577882;
assign addr[37329]= -2007305472;
assign addr[37330]= -1993396407;
assign addr[37331]= -1978855097;
assign addr[37332]= -1963686155;
assign addr[37333]= -1947894393;
assign addr[37334]= -1931484818;
assign addr[37335]= -1914462636;
assign addr[37336]= -1896833245;
assign addr[37337]= -1878602237;
assign addr[37338]= -1859775393;
assign addr[37339]= -1840358687;
assign addr[37340]= -1820358275;
assign addr[37341]= -1799780501;
assign addr[37342]= -1778631892;
assign addr[37343]= -1756919156;
assign addr[37344]= -1734649179;
assign addr[37345]= -1711829025;
assign addr[37346]= -1688465931;
assign addr[37347]= -1664567307;
assign addr[37348]= -1640140734;
assign addr[37349]= -1615193959;
assign addr[37350]= -1589734894;
assign addr[37351]= -1563771613;
assign addr[37352]= -1537312353;
assign addr[37353]= -1510365504;
assign addr[37354]= -1482939614;
assign addr[37355]= -1455043381;
assign addr[37356]= -1426685652;
assign addr[37357]= -1397875423;
assign addr[37358]= -1368621831;
assign addr[37359]= -1338934154;
assign addr[37360]= -1308821808;
assign addr[37361]= -1278294345;
assign addr[37362]= -1247361445;
assign addr[37363]= -1216032921;
assign addr[37364]= -1184318708;
assign addr[37365]= -1152228866;
assign addr[37366]= -1119773573;
assign addr[37367]= -1086963121;
assign addr[37368]= -1053807919;
assign addr[37369]= -1020318481;
assign addr[37370]= -986505429;
assign addr[37371]= -952379488;
assign addr[37372]= -917951481;
assign addr[37373]= -883232329;
assign addr[37374]= -848233042;
assign addr[37375]= -812964722;
assign addr[37376]= -777438554;
assign addr[37377]= -741665807;
assign addr[37378]= -705657826;
assign addr[37379]= -669426032;
assign addr[37380]= -632981917;
assign addr[37381]= -596337040;
assign addr[37382]= -559503022;
assign addr[37383]= -522491548;
assign addr[37384]= -485314355;
assign addr[37385]= -447983235;
assign addr[37386]= -410510029;
assign addr[37387]= -372906622;
assign addr[37388]= -335184940;
assign addr[37389]= -297356948;
assign addr[37390]= -259434643;
assign addr[37391]= -221430054;
assign addr[37392]= -183355234;
assign addr[37393]= -145222259;
assign addr[37394]= -107043224;
assign addr[37395]= -68830239;
assign addr[37396]= -30595422;
assign addr[37397]= 7649098;
assign addr[37398]= 45891193;
assign addr[37399]= 84118732;
assign addr[37400]= 122319591;
assign addr[37401]= 160481654;
assign addr[37402]= 198592817;
assign addr[37403]= 236640993;
assign addr[37404]= 274614114;
assign addr[37405]= 312500135;
assign addr[37406]= 350287041;
assign addr[37407]= 387962847;
assign addr[37408]= 425515602;
assign addr[37409]= 462933398;
assign addr[37410]= 500204365;
assign addr[37411]= 537316682;
assign addr[37412]= 574258580;
assign addr[37413]= 611018340;
assign addr[37414]= 647584304;
assign addr[37415]= 683944874;
assign addr[37416]= 720088517;
assign addr[37417]= 756003771;
assign addr[37418]= 791679244;
assign addr[37419]= 827103620;
assign addr[37420]= 862265664;
assign addr[37421]= 897154224;
assign addr[37422]= 931758235;
assign addr[37423]= 966066720;
assign addr[37424]= 1000068799;
assign addr[37425]= 1033753687;
assign addr[37426]= 1067110699;
assign addr[37427]= 1100129257;
assign addr[37428]= 1132798888;
assign addr[37429]= 1165109230;
assign addr[37430]= 1197050035;
assign addr[37431]= 1228611172;
assign addr[37432]= 1259782632;
assign addr[37433]= 1290554528;
assign addr[37434]= 1320917099;
assign addr[37435]= 1350860716;
assign addr[37436]= 1380375881;
assign addr[37437]= 1409453233;
assign addr[37438]= 1438083551;
assign addr[37439]= 1466257752;
assign addr[37440]= 1493966902;
assign addr[37441]= 1521202211;
assign addr[37442]= 1547955041;
assign addr[37443]= 1574216908;
assign addr[37444]= 1599979481;
assign addr[37445]= 1625234591;
assign addr[37446]= 1649974225;
assign addr[37447]= 1674190539;
assign addr[37448]= 1697875851;
assign addr[37449]= 1721022648;
assign addr[37450]= 1743623590;
assign addr[37451]= 1765671509;
assign addr[37452]= 1787159411;
assign addr[37453]= 1808080480;
assign addr[37454]= 1828428082;
assign addr[37455]= 1848195763;
assign addr[37456]= 1867377253;
assign addr[37457]= 1885966468;
assign addr[37458]= 1903957513;
assign addr[37459]= 1921344681;
assign addr[37460]= 1938122457;
assign addr[37461]= 1954285520;
assign addr[37462]= 1969828744;
assign addr[37463]= 1984747199;
assign addr[37464]= 1999036154;
assign addr[37465]= 2012691075;
assign addr[37466]= 2025707632;
assign addr[37467]= 2038081698;
assign addr[37468]= 2049809346;
assign addr[37469]= 2060886858;
assign addr[37470]= 2071310720;
assign addr[37471]= 2081077626;
assign addr[37472]= 2090184478;
assign addr[37473]= 2098628387;
assign addr[37474]= 2106406677;
assign addr[37475]= 2113516878;
assign addr[37476]= 2119956737;
assign addr[37477]= 2125724211;
assign addr[37478]= 2130817471;
assign addr[37479]= 2135234901;
assign addr[37480]= 2138975100;
assign addr[37481]= 2142036881;
assign addr[37482]= 2144419275;
assign addr[37483]= 2146121524;
assign addr[37484]= 2147143090;
assign addr[37485]= 2147483648;
assign addr[37486]= 2147143090;
assign addr[37487]= 2146121524;
assign addr[37488]= 2144419275;
assign addr[37489]= 2142036881;
assign addr[37490]= 2138975100;
assign addr[37491]= 2135234901;
assign addr[37492]= 2130817471;
assign addr[37493]= 2125724211;
assign addr[37494]= 2119956737;
assign addr[37495]= 2113516878;
assign addr[37496]= 2106406677;
assign addr[37497]= 2098628387;
assign addr[37498]= 2090184478;
assign addr[37499]= 2081077626;
assign addr[37500]= 2071310720;
assign addr[37501]= 2060886858;
assign addr[37502]= 2049809346;
assign addr[37503]= 2038081698;
assign addr[37504]= 2025707632;
assign addr[37505]= 2012691075;
assign addr[37506]= 1999036154;
assign addr[37507]= 1984747199;
assign addr[37508]= 1969828744;
assign addr[37509]= 1954285520;
assign addr[37510]= 1938122457;
assign addr[37511]= 1921344681;
assign addr[37512]= 1903957513;
assign addr[37513]= 1885966468;
assign addr[37514]= 1867377253;
assign addr[37515]= 1848195763;
assign addr[37516]= 1828428082;
assign addr[37517]= 1808080480;
assign addr[37518]= 1787159411;
assign addr[37519]= 1765671509;
assign addr[37520]= 1743623590;
assign addr[37521]= 1721022648;
assign addr[37522]= 1697875851;
assign addr[37523]= 1674190539;
assign addr[37524]= 1649974225;
assign addr[37525]= 1625234591;
assign addr[37526]= 1599979481;
assign addr[37527]= 1574216908;
assign addr[37528]= 1547955041;
assign addr[37529]= 1521202211;
assign addr[37530]= 1493966902;
assign addr[37531]= 1466257752;
assign addr[37532]= 1438083551;
assign addr[37533]= 1409453233;
assign addr[37534]= 1380375881;
assign addr[37535]= 1350860716;
assign addr[37536]= 1320917099;
assign addr[37537]= 1290554528;
assign addr[37538]= 1259782632;
assign addr[37539]= 1228611172;
assign addr[37540]= 1197050035;
assign addr[37541]= 1165109230;
assign addr[37542]= 1132798888;
assign addr[37543]= 1100129257;
assign addr[37544]= 1067110699;
assign addr[37545]= 1033753687;
assign addr[37546]= 1000068799;
assign addr[37547]= 966066720;
assign addr[37548]= 931758235;
assign addr[37549]= 897154224;
assign addr[37550]= 862265664;
assign addr[37551]= 827103620;
assign addr[37552]= 791679244;
assign addr[37553]= 756003771;
assign addr[37554]= 720088517;
assign addr[37555]= 683944874;
assign addr[37556]= 647584304;
assign addr[37557]= 611018340;
assign addr[37558]= 574258580;
assign addr[37559]= 537316682;
assign addr[37560]= 500204365;
assign addr[37561]= 462933398;
assign addr[37562]= 425515602;
assign addr[37563]= 387962847;
assign addr[37564]= 350287041;
assign addr[37565]= 312500135;
assign addr[37566]= 274614114;
assign addr[37567]= 236640993;
assign addr[37568]= 198592817;
assign addr[37569]= 160481654;
assign addr[37570]= 122319591;
assign addr[37571]= 84118732;
assign addr[37572]= 45891193;
assign addr[37573]= 7649098;
assign addr[37574]= -30595422;
assign addr[37575]= -68830239;
assign addr[37576]= -107043224;
assign addr[37577]= -145222259;
assign addr[37578]= -183355234;
assign addr[37579]= -221430054;
assign addr[37580]= -259434643;
assign addr[37581]= -297356948;
assign addr[37582]= -335184940;
assign addr[37583]= -372906622;
assign addr[37584]= -410510029;
assign addr[37585]= -447983235;
assign addr[37586]= -485314355;
assign addr[37587]= -522491548;
assign addr[37588]= -559503022;
assign addr[37589]= -596337040;
assign addr[37590]= -632981917;
assign addr[37591]= -669426032;
assign addr[37592]= -705657826;
assign addr[37593]= -741665807;
assign addr[37594]= -777438554;
assign addr[37595]= -812964722;
assign addr[37596]= -848233042;
assign addr[37597]= -883232329;
assign addr[37598]= -917951481;
assign addr[37599]= -952379488;
assign addr[37600]= -986505429;
assign addr[37601]= -1020318481;
assign addr[37602]= -1053807919;
assign addr[37603]= -1086963121;
assign addr[37604]= -1119773573;
assign addr[37605]= -1152228866;
assign addr[37606]= -1184318708;
assign addr[37607]= -1216032921;
assign addr[37608]= -1247361445;
assign addr[37609]= -1278294345;
assign addr[37610]= -1308821808;
assign addr[37611]= -1338934154;
assign addr[37612]= -1368621831;
assign addr[37613]= -1397875423;
assign addr[37614]= -1426685652;
assign addr[37615]= -1455043381;
assign addr[37616]= -1482939614;
assign addr[37617]= -1510365504;
assign addr[37618]= -1537312353;
assign addr[37619]= -1563771613;
assign addr[37620]= -1589734894;
assign addr[37621]= -1615193959;
assign addr[37622]= -1640140734;
assign addr[37623]= -1664567307;
assign addr[37624]= -1688465931;
assign addr[37625]= -1711829025;
assign addr[37626]= -1734649179;
assign addr[37627]= -1756919156;
assign addr[37628]= -1778631892;
assign addr[37629]= -1799780501;
assign addr[37630]= -1820358275;
assign addr[37631]= -1840358687;
assign addr[37632]= -1859775393;
assign addr[37633]= -1878602237;
assign addr[37634]= -1896833245;
assign addr[37635]= -1914462636;
assign addr[37636]= -1931484818;
assign addr[37637]= -1947894393;
assign addr[37638]= -1963686155;
assign addr[37639]= -1978855097;
assign addr[37640]= -1993396407;
assign addr[37641]= -2007305472;
assign addr[37642]= -2020577882;
assign addr[37643]= -2033209426;
assign addr[37644]= -2045196100;
assign addr[37645]= -2056534099;
assign addr[37646]= -2067219829;
assign addr[37647]= -2077249901;
assign addr[37648]= -2086621133;
assign addr[37649]= -2095330553;
assign addr[37650]= -2103375398;
assign addr[37651]= -2110753117;
assign addr[37652]= -2117461370;
assign addr[37653]= -2123498030;
assign addr[37654]= -2128861181;
assign addr[37655]= -2133549123;
assign addr[37656]= -2137560369;
assign addr[37657]= -2140893646;
assign addr[37658]= -2143547897;
assign addr[37659]= -2145522281;
assign addr[37660]= -2146816171;
assign addr[37661]= -2147429158;
assign addr[37662]= -2147361045;
assign addr[37663]= -2146611856;
assign addr[37664]= -2145181827;
assign addr[37665]= -2143071413;
assign addr[37666]= -2140281282;
assign addr[37667]= -2136812319;
assign addr[37668]= -2132665626;
assign addr[37669]= -2127842516;
assign addr[37670]= -2122344521;
assign addr[37671]= -2116173382;
assign addr[37672]= -2109331059;
assign addr[37673]= -2101819720;
assign addr[37674]= -2093641749;
assign addr[37675]= -2084799740;
assign addr[37676]= -2075296495;
assign addr[37677]= -2065135031;
assign addr[37678]= -2054318569;
assign addr[37679]= -2042850540;
assign addr[37680]= -2030734582;
assign addr[37681]= -2017974537;
assign addr[37682]= -2004574453;
assign addr[37683]= -1990538579;
assign addr[37684]= -1975871368;
assign addr[37685]= -1960577471;
assign addr[37686]= -1944661739;
assign addr[37687]= -1928129220;
assign addr[37688]= -1910985158;
assign addr[37689]= -1893234990;
assign addr[37690]= -1874884346;
assign addr[37691]= -1855939047;
assign addr[37692]= -1836405100;
assign addr[37693]= -1816288703;
assign addr[37694]= -1795596234;
assign addr[37695]= -1774334257;
assign addr[37696]= -1752509516;
assign addr[37697]= -1730128933;
assign addr[37698]= -1707199606;
assign addr[37699]= -1683728808;
assign addr[37700]= -1659723983;
assign addr[37701]= -1635192744;
assign addr[37702]= -1610142873;
assign addr[37703]= -1584582314;
assign addr[37704]= -1558519173;
assign addr[37705]= -1531961719;
assign addr[37706]= -1504918373;
assign addr[37707]= -1477397714;
assign addr[37708]= -1449408469;
assign addr[37709]= -1420959516;
assign addr[37710]= -1392059879;
assign addr[37711]= -1362718723;
assign addr[37712]= -1332945355;
assign addr[37713]= -1302749217;
assign addr[37714]= -1272139887;
assign addr[37715]= -1241127074;
assign addr[37716]= -1209720613;
assign addr[37717]= -1177930466;
assign addr[37718]= -1145766716;
assign addr[37719]= -1113239564;
assign addr[37720]= -1080359326;
assign addr[37721]= -1047136432;
assign addr[37722]= -1013581418;
assign addr[37723]= -979704927;
assign addr[37724]= -945517704;
assign addr[37725]= -911030591;
assign addr[37726]= -876254528;
assign addr[37727]= -841200544;
assign addr[37728]= -805879757;
assign addr[37729]= -770303369;
assign addr[37730]= -734482665;
assign addr[37731]= -698429006;
assign addr[37732]= -662153826;
assign addr[37733]= -625668632;
assign addr[37734]= -588984994;
assign addr[37735]= -552114549;
assign addr[37736]= -515068990;
assign addr[37737]= -477860067;
assign addr[37738]= -440499581;
assign addr[37739]= -402999383;
assign addr[37740]= -365371365;
assign addr[37741]= -327627463;
assign addr[37742]= -289779648;
assign addr[37743]= -251839923;
assign addr[37744]= -213820322;
assign addr[37745]= -175732905;
assign addr[37746]= -137589750;
assign addr[37747]= -99402956;
assign addr[37748]= -61184634;
assign addr[37749]= -22946906;
assign addr[37750]= 15298099;
assign addr[37751]= 53538253;
assign addr[37752]= 91761426;
assign addr[37753]= 129955495;
assign addr[37754]= 168108346;
assign addr[37755]= 206207878;
assign addr[37756]= 244242007;
assign addr[37757]= 282198671;
assign addr[37758]= 320065829;
assign addr[37759]= 357831473;
assign addr[37760]= 395483624;
assign addr[37761]= 433010339;
assign addr[37762]= 470399716;
assign addr[37763]= 507639898;
assign addr[37764]= 544719071;
assign addr[37765]= 581625477;
assign addr[37766]= 618347408;
assign addr[37767]= 654873219;
assign addr[37768]= 691191324;
assign addr[37769]= 727290205;
assign addr[37770]= 763158411;
assign addr[37771]= 798784567;
assign addr[37772]= 834157373;
assign addr[37773]= 869265610;
assign addr[37774]= 904098143;
assign addr[37775]= 938643924;
assign addr[37776]= 972891995;
assign addr[37777]= 1006831495;
assign addr[37778]= 1040451659;
assign addr[37779]= 1073741824;
assign addr[37780]= 1106691431;
assign addr[37781]= 1139290029;
assign addr[37782]= 1171527280;
assign addr[37783]= 1203392958;
assign addr[37784]= 1234876957;
assign addr[37785]= 1265969291;
assign addr[37786]= 1296660098;
assign addr[37787]= 1326939644;
assign addr[37788]= 1356798326;
assign addr[37789]= 1386226674;
assign addr[37790]= 1415215352;
assign addr[37791]= 1443755168;
assign addr[37792]= 1471837070;
assign addr[37793]= 1499452149;
assign addr[37794]= 1526591649;
assign addr[37795]= 1553246960;
assign addr[37796]= 1579409630;
assign addr[37797]= 1605071359;
assign addr[37798]= 1630224009;
assign addr[37799]= 1654859602;
assign addr[37800]= 1678970324;
assign addr[37801]= 1702548529;
assign addr[37802]= 1725586737;
assign addr[37803]= 1748077642;
assign addr[37804]= 1770014111;
assign addr[37805]= 1791389186;
assign addr[37806]= 1812196087;
assign addr[37807]= 1832428215;
assign addr[37808]= 1852079154;
assign addr[37809]= 1871142669;
assign addr[37810]= 1889612716;
assign addr[37811]= 1907483436;
assign addr[37812]= 1924749160;
assign addr[37813]= 1941404413;
assign addr[37814]= 1957443913;
assign addr[37815]= 1972862571;
assign addr[37816]= 1987655498;
assign addr[37817]= 2001818002;
assign addr[37818]= 2015345591;
assign addr[37819]= 2028233973;
assign addr[37820]= 2040479063;
assign addr[37821]= 2052076975;
assign addr[37822]= 2063024031;
assign addr[37823]= 2073316760;
assign addr[37824]= 2082951896;
assign addr[37825]= 2091926384;
assign addr[37826]= 2100237377;
assign addr[37827]= 2107882239;
assign addr[37828]= 2114858546;
assign addr[37829]= 2121164085;
assign addr[37830]= 2126796855;
assign addr[37831]= 2131755071;
assign addr[37832]= 2136037160;
assign addr[37833]= 2139641764;
assign addr[37834]= 2142567738;
assign addr[37835]= 2144814157;
assign addr[37836]= 2146380306;
assign addr[37837]= 2147265689;
assign addr[37838]= 2147470025;
assign addr[37839]= 2146993250;
assign addr[37840]= 2145835515;
assign addr[37841]= 2143997187;
assign addr[37842]= 2141478848;
assign addr[37843]= 2138281298;
assign addr[37844]= 2134405552;
assign addr[37845]= 2129852837;
assign addr[37846]= 2124624598;
assign addr[37847]= 2118722494;
assign addr[37848]= 2112148396;
assign addr[37849]= 2104904390;
assign addr[37850]= 2096992772;
assign addr[37851]= 2088416053;
assign addr[37852]= 2079176953;
assign addr[37853]= 2069278401;
assign addr[37854]= 2058723538;
assign addr[37855]= 2047515711;
assign addr[37856]= 2035658475;
assign addr[37857]= 2023155591;
assign addr[37858]= 2010011024;
assign addr[37859]= 1996228943;
assign addr[37860]= 1981813720;
assign addr[37861]= 1966769926;
assign addr[37862]= 1951102334;
assign addr[37863]= 1934815911;
assign addr[37864]= 1917915825;
assign addr[37865]= 1900407434;
assign addr[37866]= 1882296293;
assign addr[37867]= 1863588145;
assign addr[37868]= 1844288924;
assign addr[37869]= 1824404752;
assign addr[37870]= 1803941934;
assign addr[37871]= 1782906961;
assign addr[37872]= 1761306505;
assign addr[37873]= 1739147417;
assign addr[37874]= 1716436725;
assign addr[37875]= 1693181631;
assign addr[37876]= 1669389513;
assign addr[37877]= 1645067915;
assign addr[37878]= 1620224553;
assign addr[37879]= 1594867305;
assign addr[37880]= 1569004214;
assign addr[37881]= 1542643483;
assign addr[37882]= 1515793473;
assign addr[37883]= 1488462700;
assign addr[37884]= 1460659832;
assign addr[37885]= 1432393688;
assign addr[37886]= 1403673233;
assign addr[37887]= 1374507575;
assign addr[37888]= 1344905966;
assign addr[37889]= 1314877795;
assign addr[37890]= 1284432584;
assign addr[37891]= 1253579991;
assign addr[37892]= 1222329801;
assign addr[37893]= 1190691925;
assign addr[37894]= 1158676398;
assign addr[37895]= 1126293375;
assign addr[37896]= 1093553126;
assign addr[37897]= 1060466036;
assign addr[37898]= 1027042599;
assign addr[37899]= 993293415;
assign addr[37900]= 959229189;
assign addr[37901]= 924860725;
assign addr[37902]= 890198924;
assign addr[37903]= 855254778;
assign addr[37904]= 820039373;
assign addr[37905]= 784563876;
assign addr[37906]= 748839539;
assign addr[37907]= 712877694;
assign addr[37908]= 676689746;
assign addr[37909]= 640287172;
assign addr[37910]= 603681519;
assign addr[37911]= 566884397;
assign addr[37912]= 529907477;
assign addr[37913]= 492762486;
assign addr[37914]= 455461206;
assign addr[37915]= 418015468;
assign addr[37916]= 380437148;
assign addr[37917]= 342738165;
assign addr[37918]= 304930476;
assign addr[37919]= 267026072;
assign addr[37920]= 229036977;
assign addr[37921]= 190975237;
assign addr[37922]= 152852926;
assign addr[37923]= 114682135;
assign addr[37924]= 76474970;
assign addr[37925]= 38243550;
assign addr[37926]= 0;
assign addr[37927]= -38243550;
assign addr[37928]= -76474970;
assign addr[37929]= -114682135;
assign addr[37930]= -152852926;
assign addr[37931]= -190975237;
assign addr[37932]= -229036977;
assign addr[37933]= -267026072;
assign addr[37934]= -304930476;
assign addr[37935]= -342738165;
assign addr[37936]= -380437148;
assign addr[37937]= -418015468;
assign addr[37938]= -455461206;
assign addr[37939]= -492762486;
assign addr[37940]= -529907477;
assign addr[37941]= -566884397;
assign addr[37942]= -603681519;
assign addr[37943]= -640287172;
assign addr[37944]= -676689746;
assign addr[37945]= -712877694;
assign addr[37946]= -748839539;
assign addr[37947]= -784563876;
assign addr[37948]= -820039373;
assign addr[37949]= -855254778;
assign addr[37950]= -890198924;
assign addr[37951]= -924860725;
assign addr[37952]= -959229189;
assign addr[37953]= -993293415;
assign addr[37954]= -1027042599;
assign addr[37955]= -1060466036;
assign addr[37956]= -1093553126;
assign addr[37957]= -1126293375;
assign addr[37958]= -1158676398;
assign addr[37959]= -1190691925;
assign addr[37960]= -1222329801;
assign addr[37961]= -1253579991;
assign addr[37962]= -1284432584;
assign addr[37963]= -1314877795;
assign addr[37964]= -1344905966;
assign addr[37965]= -1374507575;
assign addr[37966]= -1403673233;
assign addr[37967]= -1432393688;
assign addr[37968]= -1460659832;
assign addr[37969]= -1488462700;
assign addr[37970]= -1515793473;
assign addr[37971]= -1542643483;
assign addr[37972]= -1569004214;
assign addr[37973]= -1594867305;
assign addr[37974]= -1620224553;
assign addr[37975]= -1645067915;
assign addr[37976]= -1669389513;
assign addr[37977]= -1693181631;
assign addr[37978]= -1716436725;
assign addr[37979]= -1739147417;
assign addr[37980]= -1761306505;
assign addr[37981]= -1782906961;
assign addr[37982]= -1803941934;
assign addr[37983]= -1824404752;
assign addr[37984]= -1844288924;
assign addr[37985]= -1863588145;
assign addr[37986]= -1882296293;
assign addr[37987]= -1900407434;
assign addr[37988]= -1917915825;
assign addr[37989]= -1934815911;
assign addr[37990]= -1951102334;
assign addr[37991]= -1966769926;
assign addr[37992]= -1981813720;
assign addr[37993]= -1996228943;
assign addr[37994]= -2010011024;
assign addr[37995]= -2023155591;
assign addr[37996]= -2035658475;
assign addr[37997]= -2047515711;
assign addr[37998]= -2058723538;
assign addr[37999]= -2069278401;
assign addr[38000]= -2079176953;
assign addr[38001]= -2088416053;
assign addr[38002]= -2096992772;
assign addr[38003]= -2104904390;
assign addr[38004]= -2112148396;
assign addr[38005]= -2118722494;
assign addr[38006]= -2124624598;
assign addr[38007]= -2129852837;
assign addr[38008]= -2134405552;
assign addr[38009]= -2138281298;
assign addr[38010]= -2141478848;
assign addr[38011]= -2143997187;
assign addr[38012]= -2145835515;
assign addr[38013]= -2146993250;
assign addr[38014]= -2147470025;
assign addr[38015]= -2147265689;
assign addr[38016]= -2146380306;
assign addr[38017]= -2144814157;
assign addr[38018]= -2142567738;
assign addr[38019]= -2139641764;
assign addr[38020]= -2136037160;
assign addr[38021]= -2131755071;
assign addr[38022]= -2126796855;
assign addr[38023]= -2121164085;
assign addr[38024]= -2114858546;
assign addr[38025]= -2107882239;
assign addr[38026]= -2100237377;
assign addr[38027]= -2091926384;
assign addr[38028]= -2082951896;
assign addr[38029]= -2073316760;
assign addr[38030]= -2063024031;
assign addr[38031]= -2052076975;
assign addr[38032]= -2040479063;
assign addr[38033]= -2028233973;
assign addr[38034]= -2015345591;
assign addr[38035]= -2001818002;
assign addr[38036]= -1987655498;
assign addr[38037]= -1972862571;
assign addr[38038]= -1957443913;
assign addr[38039]= -1941404413;
assign addr[38040]= -1924749160;
assign addr[38041]= -1907483436;
assign addr[38042]= -1889612716;
assign addr[38043]= -1871142669;
assign addr[38044]= -1852079154;
assign addr[38045]= -1832428215;
assign addr[38046]= -1812196087;
assign addr[38047]= -1791389186;
assign addr[38048]= -1770014111;
assign addr[38049]= -1748077642;
assign addr[38050]= -1725586737;
assign addr[38051]= -1702548529;
assign addr[38052]= -1678970324;
assign addr[38053]= -1654859602;
assign addr[38054]= -1630224009;
assign addr[38055]= -1605071359;
assign addr[38056]= -1579409630;
assign addr[38057]= -1553246960;
assign addr[38058]= -1526591649;
assign addr[38059]= -1499452149;
assign addr[38060]= -1471837070;
assign addr[38061]= -1443755168;
assign addr[38062]= -1415215352;
assign addr[38063]= -1386226674;
assign addr[38064]= -1356798326;
assign addr[38065]= -1326939644;
assign addr[38066]= -1296660098;
assign addr[38067]= -1265969291;
assign addr[38068]= -1234876957;
assign addr[38069]= -1203392958;
assign addr[38070]= -1171527280;
assign addr[38071]= -1139290029;
assign addr[38072]= -1106691431;
assign addr[38073]= -1073741824;
assign addr[38074]= -1040451659;
assign addr[38075]= -1006831495;
assign addr[38076]= -972891995;
assign addr[38077]= -938643924;
assign addr[38078]= -904098143;
assign addr[38079]= -869265610;
assign addr[38080]= -834157373;
assign addr[38081]= -798784567;
assign addr[38082]= -763158411;
assign addr[38083]= -727290205;
assign addr[38084]= -691191324;
assign addr[38085]= -654873219;
assign addr[38086]= -618347408;
assign addr[38087]= -581625477;
assign addr[38088]= -544719071;
assign addr[38089]= -507639898;
assign addr[38090]= -470399716;
assign addr[38091]= -433010339;
assign addr[38092]= -395483624;
assign addr[38093]= -357831473;
assign addr[38094]= -320065829;
assign addr[38095]= -282198671;
assign addr[38096]= -244242007;
assign addr[38097]= -206207878;
assign addr[38098]= -168108346;
assign addr[38099]= -129955495;
assign addr[38100]= -91761426;
assign addr[38101]= -53538253;
assign addr[38102]= -15298099;
assign addr[38103]= 22946906;
assign addr[38104]= 61184634;
assign addr[38105]= 99402956;
assign addr[38106]= 137589750;
assign addr[38107]= 175732905;
assign addr[38108]= 213820322;
assign addr[38109]= 251839923;
assign addr[38110]= 289779648;
assign addr[38111]= 327627463;
assign addr[38112]= 365371365;
assign addr[38113]= 402999383;
assign addr[38114]= 440499581;
assign addr[38115]= 477860067;
assign addr[38116]= 515068990;
assign addr[38117]= 552114549;
assign addr[38118]= 588984994;
assign addr[38119]= 625668632;
assign addr[38120]= 662153826;
assign addr[38121]= 698429006;
assign addr[38122]= 734482665;
assign addr[38123]= 770303369;
assign addr[38124]= 805879757;
assign addr[38125]= 841200544;
assign addr[38126]= 876254528;
assign addr[38127]= 911030591;
assign addr[38128]= 945517704;
assign addr[38129]= 979704927;
assign addr[38130]= 1013581418;
assign addr[38131]= 1047136432;
assign addr[38132]= 1080359326;
assign addr[38133]= 1113239564;
assign addr[38134]= 1145766716;
assign addr[38135]= 1177930466;
assign addr[38136]= 1209720613;
assign addr[38137]= 1241127074;
assign addr[38138]= 1272139887;
assign addr[38139]= 1302749217;
assign addr[38140]= 1332945355;
assign addr[38141]= 1362718723;
assign addr[38142]= 1392059879;
assign addr[38143]= 1420959516;
assign addr[38144]= 1449408469;
assign addr[38145]= 1477397714;
assign addr[38146]= 1504918373;
assign addr[38147]= 1531961719;
assign addr[38148]= 1558519173;
assign addr[38149]= 1584582314;
assign addr[38150]= 1610142873;
assign addr[38151]= 1635192744;
assign addr[38152]= 1659723983;
assign addr[38153]= 1683728808;
assign addr[38154]= 1707199606;
assign addr[38155]= 1730128933;
assign addr[38156]= 1752509516;
assign addr[38157]= 1774334257;
assign addr[38158]= 1795596234;
assign addr[38159]= 1816288703;
assign addr[38160]= 1836405100;
assign addr[38161]= 1855939047;
assign addr[38162]= 1874884346;
assign addr[38163]= 1893234990;
assign addr[38164]= 1910985158;
assign addr[38165]= 1928129220;
assign addr[38166]= 1944661739;
assign addr[38167]= 1960577471;
assign addr[38168]= 1975871368;
assign addr[38169]= 1990538579;
assign addr[38170]= 2004574453;
assign addr[38171]= 2017974537;
assign addr[38172]= 2030734582;
assign addr[38173]= 2042850540;
assign addr[38174]= 2054318569;
assign addr[38175]= 2065135031;
assign addr[38176]= 2075296495;
assign addr[38177]= 2084799740;
assign addr[38178]= 2093641749;
assign addr[38179]= 2101819720;
assign addr[38180]= 2109331059;
assign addr[38181]= 2116173382;
assign addr[38182]= 2122344521;
assign addr[38183]= 2127842516;
assign addr[38184]= 2132665626;
assign addr[38185]= 2136812319;
assign addr[38186]= 2140281282;
assign addr[38187]= 2143071413;
assign addr[38188]= 2145181827;
assign addr[38189]= 2146611856;
assign addr[38190]= 2147361045;
assign addr[38191]= 2147429158;
assign addr[38192]= 2146816171;
assign addr[38193]= 2145522281;
assign addr[38194]= 2143547897;
assign addr[38195]= 2140893646;
assign addr[38196]= 2137560369;
assign addr[38197]= 2133549123;
assign addr[38198]= 2128861181;
assign addr[38199]= 2123498030;
assign addr[38200]= 2117461370;
assign addr[38201]= 2110753117;
assign addr[38202]= 2103375398;
assign addr[38203]= 2095330553;
assign addr[38204]= 2086621133;
assign addr[38205]= 2077249901;
assign addr[38206]= 2067219829;
assign addr[38207]= 2056534099;
assign addr[38208]= 2045196100;
assign addr[38209]= 2033209426;
assign addr[38210]= 2020577882;
assign addr[38211]= 2007305472;
assign addr[38212]= 1993396407;
assign addr[38213]= 1978855097;
assign addr[38214]= 1963686155;
assign addr[38215]= 1947894393;
assign addr[38216]= 1931484818;
assign addr[38217]= 1914462636;
assign addr[38218]= 1896833245;
assign addr[38219]= 1878602237;
assign addr[38220]= 1859775393;
assign addr[38221]= 1840358687;
assign addr[38222]= 1820358275;
assign addr[38223]= 1799780501;
assign addr[38224]= 1778631892;
assign addr[38225]= 1756919156;
assign addr[38226]= 1734649179;
assign addr[38227]= 1711829025;
assign addr[38228]= 1688465931;
assign addr[38229]= 1664567307;
assign addr[38230]= 1640140734;
assign addr[38231]= 1615193959;
assign addr[38232]= 1589734894;
assign addr[38233]= 1563771613;
assign addr[38234]= 1537312353;
assign addr[38235]= 1510365504;
assign addr[38236]= 1482939614;
assign addr[38237]= 1455043381;
assign addr[38238]= 1426685652;
assign addr[38239]= 1397875423;
assign addr[38240]= 1368621831;
assign addr[38241]= 1338934154;
assign addr[38242]= 1308821808;
assign addr[38243]= 1278294345;
assign addr[38244]= 1247361445;
assign addr[38245]= 1216032921;
assign addr[38246]= 1184318708;
assign addr[38247]= 1152228866;
assign addr[38248]= 1119773573;
assign addr[38249]= 1086963121;
assign addr[38250]= 1053807919;
assign addr[38251]= 1020318481;
assign addr[38252]= 986505429;
assign addr[38253]= 952379488;
assign addr[38254]= 917951481;
assign addr[38255]= 883232329;
assign addr[38256]= 848233042;
assign addr[38257]= 812964722;
assign addr[38258]= 777438554;
assign addr[38259]= 741665807;
assign addr[38260]= 705657826;
assign addr[38261]= 669426032;
assign addr[38262]= 632981917;
assign addr[38263]= 596337040;
assign addr[38264]= 559503022;
assign addr[38265]= 522491548;
assign addr[38266]= 485314355;
assign addr[38267]= 447983235;
assign addr[38268]= 410510029;
assign addr[38269]= 372906622;
assign addr[38270]= 335184940;
assign addr[38271]= 297356948;
assign addr[38272]= 259434643;
assign addr[38273]= 221430054;
assign addr[38274]= 183355234;
assign addr[38275]= 145222259;
assign addr[38276]= 107043224;
assign addr[38277]= 68830239;
assign addr[38278]= 30595422;
assign addr[38279]= -7649098;
assign addr[38280]= -45891193;
assign addr[38281]= -84118732;
assign addr[38282]= -122319591;
assign addr[38283]= -160481654;
assign addr[38284]= -198592817;
assign addr[38285]= -236640993;
assign addr[38286]= -274614114;
assign addr[38287]= -312500135;
assign addr[38288]= -350287041;
assign addr[38289]= -387962847;
assign addr[38290]= -425515602;
assign addr[38291]= -462933398;
assign addr[38292]= -500204365;
assign addr[38293]= -537316682;
assign addr[38294]= -574258580;
assign addr[38295]= -611018340;
assign addr[38296]= -647584304;
assign addr[38297]= -683944874;
assign addr[38298]= -720088517;
assign addr[38299]= -756003771;
assign addr[38300]= -791679244;
assign addr[38301]= -827103620;
assign addr[38302]= -862265664;
assign addr[38303]= -897154224;
assign addr[38304]= -931758235;
assign addr[38305]= -966066720;
assign addr[38306]= -1000068799;
assign addr[38307]= -1033753687;
assign addr[38308]= -1067110699;
assign addr[38309]= -1100129257;
assign addr[38310]= -1132798888;
assign addr[38311]= -1165109230;
assign addr[38312]= -1197050035;
assign addr[38313]= -1228611172;
assign addr[38314]= -1259782632;
assign addr[38315]= -1290554528;
assign addr[38316]= -1320917099;
assign addr[38317]= -1350860716;
assign addr[38318]= -1380375881;
assign addr[38319]= -1409453233;
assign addr[38320]= -1438083551;
assign addr[38321]= -1466257752;
assign addr[38322]= -1493966902;
assign addr[38323]= -1521202211;
assign addr[38324]= -1547955041;
assign addr[38325]= -1574216908;
assign addr[38326]= -1599979481;
assign addr[38327]= -1625234591;
assign addr[38328]= -1649974225;
assign addr[38329]= -1674190539;
assign addr[38330]= -1697875851;
assign addr[38331]= -1721022648;
assign addr[38332]= -1743623590;
assign addr[38333]= -1765671509;
assign addr[38334]= -1787159411;
assign addr[38335]= -1808080480;
assign addr[38336]= -1828428082;
assign addr[38337]= -1848195763;
assign addr[38338]= -1867377253;
assign addr[38339]= -1885966468;
assign addr[38340]= -1903957513;
assign addr[38341]= -1921344681;
assign addr[38342]= -1938122457;
assign addr[38343]= -1954285520;
assign addr[38344]= -1969828744;
assign addr[38345]= -1984747199;
assign addr[38346]= -1999036154;
assign addr[38347]= -2012691075;
assign addr[38348]= -2025707632;
assign addr[38349]= -2038081698;
assign addr[38350]= -2049809346;
assign addr[38351]= -2060886858;
assign addr[38352]= -2071310720;
assign addr[38353]= -2081077626;
assign addr[38354]= -2090184478;
assign addr[38355]= -2098628387;
assign addr[38356]= -2106406677;
assign addr[38357]= -2113516878;
assign addr[38358]= -2119956737;
assign addr[38359]= -2125724211;
assign addr[38360]= -2130817471;
assign addr[38361]= -2135234901;
assign addr[38362]= -2138975100;
assign addr[38363]= -2142036881;
assign addr[38364]= -2144419275;
assign addr[38365]= -2146121524;
assign addr[38366]= -2147143090;
assign addr[38367]= -2147483648;
assign addr[38368]= -2147143090;
assign addr[38369]= -2146121524;
assign addr[38370]= -2144419275;
assign addr[38371]= -2142036881;
assign addr[38372]= -2138975100;
assign addr[38373]= -2135234901;
assign addr[38374]= -2130817471;
assign addr[38375]= -2125724211;
assign addr[38376]= -2119956737;
assign addr[38377]= -2113516878;
assign addr[38378]= -2106406677;
assign addr[38379]= -2098628387;
assign addr[38380]= -2090184478;
assign addr[38381]= -2081077626;
assign addr[38382]= -2071310720;
assign addr[38383]= -2060886858;
assign addr[38384]= -2049809346;
assign addr[38385]= -2038081698;
assign addr[38386]= -2025707632;
assign addr[38387]= -2012691075;
assign addr[38388]= -1999036154;
assign addr[38389]= -1984747199;
assign addr[38390]= -1969828744;
assign addr[38391]= -1954285520;
assign addr[38392]= -1938122457;
assign addr[38393]= -1921344681;
assign addr[38394]= -1903957513;
assign addr[38395]= -1885966468;
assign addr[38396]= -1867377253;
assign addr[38397]= -1848195763;
assign addr[38398]= -1828428082;
assign addr[38399]= -1808080480;
assign addr[38400]= -1787159411;
assign addr[38401]= -1765671509;
assign addr[38402]= -1743623590;
assign addr[38403]= -1721022648;
assign addr[38404]= -1697875851;
assign addr[38405]= -1674190539;
assign addr[38406]= -1649974225;
assign addr[38407]= -1625234591;
assign addr[38408]= -1599979481;
assign addr[38409]= -1574216908;
assign addr[38410]= -1547955041;
assign addr[38411]= -1521202211;
assign addr[38412]= -1493966902;
assign addr[38413]= -1466257752;
assign addr[38414]= -1438083551;
assign addr[38415]= -1409453233;
assign addr[38416]= -1380375881;
assign addr[38417]= -1350860716;
assign addr[38418]= -1320917099;
assign addr[38419]= -1290554528;
assign addr[38420]= -1259782632;
assign addr[38421]= -1228611172;
assign addr[38422]= -1197050035;
assign addr[38423]= -1165109230;
assign addr[38424]= -1132798888;
assign addr[38425]= -1100129257;
assign addr[38426]= -1067110699;
assign addr[38427]= -1033753687;
assign addr[38428]= -1000068799;
assign addr[38429]= -966066720;
assign addr[38430]= -931758235;
assign addr[38431]= -897154224;
assign addr[38432]= -862265664;
assign addr[38433]= -827103620;
assign addr[38434]= -791679244;
assign addr[38435]= -756003771;
assign addr[38436]= -720088517;
assign addr[38437]= -683944874;
assign addr[38438]= -647584304;
assign addr[38439]= -611018340;
assign addr[38440]= -574258580;
assign addr[38441]= -537316682;
assign addr[38442]= -500204365;
assign addr[38443]= -462933398;
assign addr[38444]= -425515602;
assign addr[38445]= -387962847;
assign addr[38446]= -350287041;
assign addr[38447]= -312500135;
assign addr[38448]= -274614114;
assign addr[38449]= -236640993;
assign addr[38450]= -198592817;
assign addr[38451]= -160481654;
assign addr[38452]= -122319591;
assign addr[38453]= -84118732;
assign addr[38454]= -45891193;
assign addr[38455]= -7649098;
assign addr[38456]= 30595422;
assign addr[38457]= 68830239;
assign addr[38458]= 107043224;
assign addr[38459]= 145222259;
assign addr[38460]= 183355234;
assign addr[38461]= 221430054;
assign addr[38462]= 259434643;
assign addr[38463]= 297356948;
assign addr[38464]= 335184940;
assign addr[38465]= 372906622;
assign addr[38466]= 410510029;
assign addr[38467]= 447983235;
assign addr[38468]= 485314355;
assign addr[38469]= 522491548;
assign addr[38470]= 559503022;
assign addr[38471]= 596337040;
assign addr[38472]= 632981917;
assign addr[38473]= 669426032;
assign addr[38474]= 705657826;
assign addr[38475]= 741665807;
assign addr[38476]= 777438554;
assign addr[38477]= 812964722;
assign addr[38478]= 848233042;
assign addr[38479]= 883232329;
assign addr[38480]= 917951481;
assign addr[38481]= 952379488;
assign addr[38482]= 986505429;
assign addr[38483]= 1020318481;
assign addr[38484]= 1053807919;
assign addr[38485]= 1086963121;
assign addr[38486]= 1119773573;
assign addr[38487]= 1152228866;
assign addr[38488]= 1184318708;
assign addr[38489]= 1216032921;
assign addr[38490]= 1247361445;
assign addr[38491]= 1278294345;
assign addr[38492]= 1308821808;
assign addr[38493]= 1338934154;
assign addr[38494]= 1368621831;
assign addr[38495]= 1397875423;
assign addr[38496]= 1426685652;
assign addr[38497]= 1455043381;
assign addr[38498]= 1482939614;
assign addr[38499]= 1510365504;
assign addr[38500]= 1537312353;
assign addr[38501]= 1563771613;
assign addr[38502]= 1589734894;
assign addr[38503]= 1615193959;
assign addr[38504]= 1640140734;
assign addr[38505]= 1664567307;
assign addr[38506]= 1688465931;
assign addr[38507]= 1711829025;
assign addr[38508]= 1734649179;
assign addr[38509]= 1756919156;
assign addr[38510]= 1778631892;
assign addr[38511]= 1799780501;
assign addr[38512]= 1820358275;
assign addr[38513]= 1840358687;
assign addr[38514]= 1859775393;
assign addr[38515]= 1878602237;
assign addr[38516]= 1896833245;
assign addr[38517]= 1914462636;
assign addr[38518]= 1931484818;
assign addr[38519]= 1947894393;
assign addr[38520]= 1963686155;
assign addr[38521]= 1978855097;
assign addr[38522]= 1993396407;
assign addr[38523]= 2007305472;
assign addr[38524]= 2020577882;
assign addr[38525]= 2033209426;
assign addr[38526]= 2045196100;
assign addr[38527]= 2056534099;
assign addr[38528]= 2067219829;
assign addr[38529]= 2077249901;
assign addr[38530]= 2086621133;
assign addr[38531]= 2095330553;
assign addr[38532]= 2103375398;
assign addr[38533]= 2110753117;
assign addr[38534]= 2117461370;
assign addr[38535]= 2123498030;
assign addr[38536]= 2128861181;
assign addr[38537]= 2133549123;
assign addr[38538]= 2137560369;
assign addr[38539]= 2140893646;
assign addr[38540]= 2143547897;
assign addr[38541]= 2145522281;
assign addr[38542]= 2146816171;
assign addr[38543]= 2147429158;
assign addr[38544]= 2147361045;
assign addr[38545]= 2146611856;
assign addr[38546]= 2145181827;
assign addr[38547]= 2143071413;
assign addr[38548]= 2140281282;
assign addr[38549]= 2136812319;
assign addr[38550]= 2132665626;
assign addr[38551]= 2127842516;
assign addr[38552]= 2122344521;
assign addr[38553]= 2116173382;
assign addr[38554]= 2109331059;
assign addr[38555]= 2101819720;
assign addr[38556]= 2093641749;
assign addr[38557]= 2084799740;
assign addr[38558]= 2075296495;
assign addr[38559]= 2065135031;
assign addr[38560]= 2054318569;
assign addr[38561]= 2042850540;
assign addr[38562]= 2030734582;
assign addr[38563]= 2017974537;
assign addr[38564]= 2004574453;
assign addr[38565]= 1990538579;
assign addr[38566]= 1975871368;
assign addr[38567]= 1960577471;
assign addr[38568]= 1944661739;
assign addr[38569]= 1928129220;
assign addr[38570]= 1910985158;
assign addr[38571]= 1893234990;
assign addr[38572]= 1874884346;
assign addr[38573]= 1855939047;
assign addr[38574]= 1836405100;
assign addr[38575]= 1816288703;
assign addr[38576]= 1795596234;
assign addr[38577]= 1774334257;
assign addr[38578]= 1752509516;
assign addr[38579]= 1730128933;
assign addr[38580]= 1707199606;
assign addr[38581]= 1683728808;
assign addr[38582]= 1659723983;
assign addr[38583]= 1635192744;
assign addr[38584]= 1610142873;
assign addr[38585]= 1584582314;
assign addr[38586]= 1558519173;
assign addr[38587]= 1531961719;
assign addr[38588]= 1504918373;
assign addr[38589]= 1477397714;
assign addr[38590]= 1449408469;
assign addr[38591]= 1420959516;
assign addr[38592]= 1392059879;
assign addr[38593]= 1362718723;
assign addr[38594]= 1332945355;
assign addr[38595]= 1302749217;
assign addr[38596]= 1272139887;
assign addr[38597]= 1241127074;
assign addr[38598]= 1209720613;
assign addr[38599]= 1177930466;
assign addr[38600]= 1145766716;
assign addr[38601]= 1113239564;
assign addr[38602]= 1080359326;
assign addr[38603]= 1047136432;
assign addr[38604]= 1013581418;
assign addr[38605]= 979704927;
assign addr[38606]= 945517704;
assign addr[38607]= 911030591;
assign addr[38608]= 876254528;
assign addr[38609]= 841200544;
assign addr[38610]= 805879757;
assign addr[38611]= 770303369;
assign addr[38612]= 734482665;
assign addr[38613]= 698429006;
assign addr[38614]= 662153826;
assign addr[38615]= 625668632;
assign addr[38616]= 588984994;
assign addr[38617]= 552114549;
assign addr[38618]= 515068990;
assign addr[38619]= 477860067;
assign addr[38620]= 440499581;
assign addr[38621]= 402999383;
assign addr[38622]= 365371365;
assign addr[38623]= 327627463;
assign addr[38624]= 289779648;
assign addr[38625]= 251839923;
assign addr[38626]= 213820322;
assign addr[38627]= 175732905;
assign addr[38628]= 137589750;
assign addr[38629]= 99402956;
assign addr[38630]= 61184634;
assign addr[38631]= 22946906;
assign addr[38632]= -15298099;
assign addr[38633]= -53538253;
assign addr[38634]= -91761426;
assign addr[38635]= -129955495;
assign addr[38636]= -168108346;
assign addr[38637]= -206207878;
assign addr[38638]= -244242007;
assign addr[38639]= -282198671;
assign addr[38640]= -320065829;
assign addr[38641]= -357831473;
assign addr[38642]= -395483624;
assign addr[38643]= -433010339;
assign addr[38644]= -470399716;
assign addr[38645]= -507639898;
assign addr[38646]= -544719071;
assign addr[38647]= -581625477;
assign addr[38648]= -618347408;
assign addr[38649]= -654873219;
assign addr[38650]= -691191324;
assign addr[38651]= -727290205;
assign addr[38652]= -763158411;
assign addr[38653]= -798784567;
assign addr[38654]= -834157373;
assign addr[38655]= -869265610;
assign addr[38656]= -904098143;
assign addr[38657]= -938643924;
assign addr[38658]= -972891995;
assign addr[38659]= -1006831495;
assign addr[38660]= -1040451659;
assign addr[38661]= -1073741824;
assign addr[38662]= -1106691431;
assign addr[38663]= -1139290029;
assign addr[38664]= -1171527280;
assign addr[38665]= -1203392958;
assign addr[38666]= -1234876957;
assign addr[38667]= -1265969291;
assign addr[38668]= -1296660098;
assign addr[38669]= -1326939644;
assign addr[38670]= -1356798326;
assign addr[38671]= -1386226674;
assign addr[38672]= -1415215352;
assign addr[38673]= -1443755168;
assign addr[38674]= -1471837070;
assign addr[38675]= -1499452149;
assign addr[38676]= -1526591649;
assign addr[38677]= -1553246960;
assign addr[38678]= -1579409630;
assign addr[38679]= -1605071359;
assign addr[38680]= -1630224009;
assign addr[38681]= -1654859602;
assign addr[38682]= -1678970324;
assign addr[38683]= -1702548529;
assign addr[38684]= -1725586737;
assign addr[38685]= -1748077642;
assign addr[38686]= -1770014111;
assign addr[38687]= -1791389186;
assign addr[38688]= -1812196087;
assign addr[38689]= -1832428215;
assign addr[38690]= -1852079154;
assign addr[38691]= -1871142669;
assign addr[38692]= -1889612716;
assign addr[38693]= -1907483436;
assign addr[38694]= -1924749160;
assign addr[38695]= -1941404413;
assign addr[38696]= -1957443913;
assign addr[38697]= -1972862571;
assign addr[38698]= -1987655498;
assign addr[38699]= -2001818002;
assign addr[38700]= -2015345591;
assign addr[38701]= -2028233973;
assign addr[38702]= -2040479063;
assign addr[38703]= -2052076975;
assign addr[38704]= -2063024031;
assign addr[38705]= -2073316760;
assign addr[38706]= -2082951896;
assign addr[38707]= -2091926384;
assign addr[38708]= -2100237377;
assign addr[38709]= -2107882239;
assign addr[38710]= -2114858546;
assign addr[38711]= -2121164085;
assign addr[38712]= -2126796855;
assign addr[38713]= -2131755071;
assign addr[38714]= -2136037160;
assign addr[38715]= -2139641764;
assign addr[38716]= -2142567738;
assign addr[38717]= -2144814157;
assign addr[38718]= -2146380306;
assign addr[38719]= -2147265689;
assign addr[38720]= -2147470025;
assign addr[38721]= -2146993250;
assign addr[38722]= -2145835515;
assign addr[38723]= -2143997187;
assign addr[38724]= -2141478848;
assign addr[38725]= -2138281298;
assign addr[38726]= -2134405552;
assign addr[38727]= -2129852837;
assign addr[38728]= -2124624598;
assign addr[38729]= -2118722494;
assign addr[38730]= -2112148396;
assign addr[38731]= -2104904390;
assign addr[38732]= -2096992772;
assign addr[38733]= -2088416053;
assign addr[38734]= -2079176953;
assign addr[38735]= -2069278401;
assign addr[38736]= -2058723538;
assign addr[38737]= -2047515711;
assign addr[38738]= -2035658475;
assign addr[38739]= -2023155591;
assign addr[38740]= -2010011024;
assign addr[38741]= -1996228943;
assign addr[38742]= -1981813720;
assign addr[38743]= -1966769926;
assign addr[38744]= -1951102334;
assign addr[38745]= -1934815911;
assign addr[38746]= -1917915825;
assign addr[38747]= -1900407434;
assign addr[38748]= -1882296293;
assign addr[38749]= -1863588145;
assign addr[38750]= -1844288924;
assign addr[38751]= -1824404752;
assign addr[38752]= -1803941934;
assign addr[38753]= -1782906961;
assign addr[38754]= -1761306505;
assign addr[38755]= -1739147417;
assign addr[38756]= -1716436725;
assign addr[38757]= -1693181631;
assign addr[38758]= -1669389513;
assign addr[38759]= -1645067915;
assign addr[38760]= -1620224553;
assign addr[38761]= -1594867305;
assign addr[38762]= -1569004214;
assign addr[38763]= -1542643483;
assign addr[38764]= -1515793473;
assign addr[38765]= -1488462700;
assign addr[38766]= -1460659832;
assign addr[38767]= -1432393688;
assign addr[38768]= -1403673233;
assign addr[38769]= -1374507575;
assign addr[38770]= -1344905966;
assign addr[38771]= -1314877795;
assign addr[38772]= -1284432584;
assign addr[38773]= -1253579991;
assign addr[38774]= -1222329801;
assign addr[38775]= -1190691925;
assign addr[38776]= -1158676398;
assign addr[38777]= -1126293375;
assign addr[38778]= -1093553126;
assign addr[38779]= -1060466036;
assign addr[38780]= -1027042599;
assign addr[38781]= -993293415;
assign addr[38782]= -959229189;
assign addr[38783]= -924860725;
assign addr[38784]= -890198924;
assign addr[38785]= -855254778;
assign addr[38786]= -820039373;
assign addr[38787]= -784563876;
assign addr[38788]= -748839539;
assign addr[38789]= -712877694;
assign addr[38790]= -676689746;
assign addr[38791]= -640287172;
assign addr[38792]= -603681519;
assign addr[38793]= -566884397;
assign addr[38794]= -529907477;
assign addr[38795]= -492762486;
assign addr[38796]= -455461206;
assign addr[38797]= -418015468;
assign addr[38798]= -380437148;
assign addr[38799]= -342738165;
assign addr[38800]= -304930476;
assign addr[38801]= -267026072;
assign addr[38802]= -229036977;
assign addr[38803]= -190975237;
assign addr[38804]= -152852926;
assign addr[38805]= -114682135;
assign addr[38806]= -76474970;
assign addr[38807]= -38243550;
assign addr[38808]= 0;
assign addr[38809]= 38243550;
assign addr[38810]= 76474970;
assign addr[38811]= 114682135;
assign addr[38812]= 152852926;
assign addr[38813]= 190975237;
assign addr[38814]= 229036977;
assign addr[38815]= 267026072;
assign addr[38816]= 304930476;
assign addr[38817]= 342738165;
assign addr[38818]= 380437148;
assign addr[38819]= 418015468;
assign addr[38820]= 455461206;
assign addr[38821]= 492762486;
assign addr[38822]= 529907477;
assign addr[38823]= 566884397;
assign addr[38824]= 603681519;
assign addr[38825]= 640287172;
assign addr[38826]= 676689746;
assign addr[38827]= 712877694;
assign addr[38828]= 748839539;
assign addr[38829]= 784563876;
assign addr[38830]= 820039373;
assign addr[38831]= 855254778;
assign addr[38832]= 890198924;
assign addr[38833]= 924860725;
assign addr[38834]= 959229189;
assign addr[38835]= 993293415;
assign addr[38836]= 1027042599;
assign addr[38837]= 1060466036;
assign addr[38838]= 1093553126;
assign addr[38839]= 1126293375;
assign addr[38840]= 1158676398;
assign addr[38841]= 1190691925;
assign addr[38842]= 1222329801;
assign addr[38843]= 1253579991;
assign addr[38844]= 1284432584;
assign addr[38845]= 1314877795;
assign addr[38846]= 1344905966;
assign addr[38847]= 1374507575;
assign addr[38848]= 1403673233;
assign addr[38849]= 1432393688;
assign addr[38850]= 1460659832;
assign addr[38851]= 1488462700;
assign addr[38852]= 1515793473;
assign addr[38853]= 1542643483;
assign addr[38854]= 1569004214;
assign addr[38855]= 1594867305;
assign addr[38856]= 1620224553;
assign addr[38857]= 1645067915;
assign addr[38858]= 1669389513;
assign addr[38859]= 1693181631;
assign addr[38860]= 1716436725;
assign addr[38861]= 1739147417;
assign addr[38862]= 1761306505;
assign addr[38863]= 1782906961;
assign addr[38864]= 1803941934;
assign addr[38865]= 1824404752;
assign addr[38866]= 1844288924;
assign addr[38867]= 1863588145;
assign addr[38868]= 1882296293;
assign addr[38869]= 1900407434;
assign addr[38870]= 1917915825;
assign addr[38871]= 1934815911;
assign addr[38872]= 1951102334;
assign addr[38873]= 1966769926;
assign addr[38874]= 1981813720;
assign addr[38875]= 1996228943;
assign addr[38876]= 2010011024;
assign addr[38877]= 2023155591;
assign addr[38878]= 2035658475;
assign addr[38879]= 2047515711;
assign addr[38880]= 2058723538;
assign addr[38881]= 2069278401;
assign addr[38882]= 2079176953;
assign addr[38883]= 2088416053;
assign addr[38884]= 2096992772;
assign addr[38885]= 2104904390;
assign addr[38886]= 2112148396;
assign addr[38887]= 2118722494;
assign addr[38888]= 2124624598;
assign addr[38889]= 2129852837;
assign addr[38890]= 2134405552;
assign addr[38891]= 2138281298;
assign addr[38892]= 2141478848;
assign addr[38893]= 2143997187;
assign addr[38894]= 2145835515;
assign addr[38895]= 2146993250;
assign addr[38896]= 2147470025;
assign addr[38897]= 2147265689;
assign addr[38898]= 2146380306;
assign addr[38899]= 2144814157;
assign addr[38900]= 2142567738;
assign addr[38901]= 2139641764;
assign addr[38902]= 2136037160;
assign addr[38903]= 2131755071;
assign addr[38904]= 2126796855;
assign addr[38905]= 2121164085;
assign addr[38906]= 2114858546;
assign addr[38907]= 2107882239;
assign addr[38908]= 2100237377;
assign addr[38909]= 2091926384;
assign addr[38910]= 2082951896;
assign addr[38911]= 2073316760;
assign addr[38912]= 2063024031;
assign addr[38913]= 2052076975;
assign addr[38914]= 2040479063;
assign addr[38915]= 2028233973;
assign addr[38916]= 2015345591;
assign addr[38917]= 2001818002;
assign addr[38918]= 1987655498;
assign addr[38919]= 1972862571;
assign addr[38920]= 1957443913;
assign addr[38921]= 1941404413;
assign addr[38922]= 1924749160;
assign addr[38923]= 1907483436;
assign addr[38924]= 1889612716;
assign addr[38925]= 1871142669;
assign addr[38926]= 1852079154;
assign addr[38927]= 1832428215;
assign addr[38928]= 1812196087;
assign addr[38929]= 1791389186;
assign addr[38930]= 1770014111;
assign addr[38931]= 1748077642;
assign addr[38932]= 1725586737;
assign addr[38933]= 1702548529;
assign addr[38934]= 1678970324;
assign addr[38935]= 1654859602;
assign addr[38936]= 1630224009;
assign addr[38937]= 1605071359;
assign addr[38938]= 1579409630;
assign addr[38939]= 1553246960;
assign addr[38940]= 1526591649;
assign addr[38941]= 1499452149;
assign addr[38942]= 1471837070;
assign addr[38943]= 1443755168;
assign addr[38944]= 1415215352;
assign addr[38945]= 1386226674;
assign addr[38946]= 1356798326;
assign addr[38947]= 1326939644;
assign addr[38948]= 1296660098;
assign addr[38949]= 1265969291;
assign addr[38950]= 1234876957;
assign addr[38951]= 1203392958;
assign addr[38952]= 1171527280;
assign addr[38953]= 1139290029;
assign addr[38954]= 1106691431;
assign addr[38955]= 1073741824;
assign addr[38956]= 1040451659;
assign addr[38957]= 1006831495;
assign addr[38958]= 972891995;
assign addr[38959]= 938643924;
assign addr[38960]= 904098143;
assign addr[38961]= 869265610;
assign addr[38962]= 834157373;
assign addr[38963]= 798784567;
assign addr[38964]= 763158411;
assign addr[38965]= 727290205;
assign addr[38966]= 691191324;
assign addr[38967]= 654873219;
assign addr[38968]= 618347408;
assign addr[38969]= 581625477;
assign addr[38970]= 544719071;
assign addr[38971]= 507639898;
assign addr[38972]= 470399716;
assign addr[38973]= 433010339;
assign addr[38974]= 395483624;
assign addr[38975]= 357831473;
assign addr[38976]= 320065829;
assign addr[38977]= 282198671;
assign addr[38978]= 244242007;
assign addr[38979]= 206207878;
assign addr[38980]= 168108346;
assign addr[38981]= 129955495;
assign addr[38982]= 91761426;
assign addr[38983]= 53538253;
assign addr[38984]= 15298099;
assign addr[38985]= -22946906;
assign addr[38986]= -61184634;
assign addr[38987]= -99402956;
assign addr[38988]= -137589750;
assign addr[38989]= -175732905;
assign addr[38990]= -213820322;
assign addr[38991]= -251839923;
assign addr[38992]= -289779648;
assign addr[38993]= -327627463;
assign addr[38994]= -365371365;
assign addr[38995]= -402999383;
assign addr[38996]= -440499581;
assign addr[38997]= -477860067;
assign addr[38998]= -515068990;
assign addr[38999]= -552114549;
assign addr[39000]= -588984994;
assign addr[39001]= -625668632;
assign addr[39002]= -662153826;
assign addr[39003]= -698429006;
assign addr[39004]= -734482665;
assign addr[39005]= -770303369;
assign addr[39006]= -805879757;
assign addr[39007]= -841200544;
assign addr[39008]= -876254528;
assign addr[39009]= -911030591;
assign addr[39010]= -945517704;
assign addr[39011]= -979704927;
assign addr[39012]= -1013581418;
assign addr[39013]= -1047136432;
assign addr[39014]= -1080359326;
assign addr[39015]= -1113239564;
assign addr[39016]= -1145766716;
assign addr[39017]= -1177930466;
assign addr[39018]= -1209720613;
assign addr[39019]= -1241127074;
assign addr[39020]= -1272139887;
assign addr[39021]= -1302749217;
assign addr[39022]= -1332945355;
assign addr[39023]= -1362718723;
assign addr[39024]= -1392059879;
assign addr[39025]= -1420959516;
assign addr[39026]= -1449408469;
assign addr[39027]= -1477397714;
assign addr[39028]= -1504918373;
assign addr[39029]= -1531961719;
assign addr[39030]= -1558519173;
assign addr[39031]= -1584582314;
assign addr[39032]= -1610142873;
assign addr[39033]= -1635192744;
assign addr[39034]= -1659723983;
assign addr[39035]= -1683728808;
assign addr[39036]= -1707199606;
assign addr[39037]= -1730128933;
assign addr[39038]= -1752509516;
assign addr[39039]= -1774334257;
assign addr[39040]= -1795596234;
assign addr[39041]= -1816288703;
assign addr[39042]= -1836405100;
assign addr[39043]= -1855939047;
assign addr[39044]= -1874884346;
assign addr[39045]= -1893234990;
assign addr[39046]= -1910985158;
assign addr[39047]= -1928129220;
assign addr[39048]= -1944661739;
assign addr[39049]= -1960577471;
assign addr[39050]= -1975871368;
assign addr[39051]= -1990538579;
assign addr[39052]= -2004574453;
assign addr[39053]= -2017974537;
assign addr[39054]= -2030734582;
assign addr[39055]= -2042850540;
assign addr[39056]= -2054318569;
assign addr[39057]= -2065135031;
assign addr[39058]= -2075296495;
assign addr[39059]= -2084799740;
assign addr[39060]= -2093641749;
assign addr[39061]= -2101819720;
assign addr[39062]= -2109331059;
assign addr[39063]= -2116173382;
assign addr[39064]= -2122344521;
assign addr[39065]= -2127842516;
assign addr[39066]= -2132665626;
assign addr[39067]= -2136812319;
assign addr[39068]= -2140281282;
assign addr[39069]= -2143071413;
assign addr[39070]= -2145181827;
assign addr[39071]= -2146611856;
assign addr[39072]= -2147361045;
assign addr[39073]= -2147429158;
assign addr[39074]= -2146816171;
assign addr[39075]= -2145522281;
assign addr[39076]= -2143547897;
assign addr[39077]= -2140893646;
assign addr[39078]= -2137560369;
assign addr[39079]= -2133549123;
assign addr[39080]= -2128861181;
assign addr[39081]= -2123498030;
assign addr[39082]= -2117461370;
assign addr[39083]= -2110753117;
assign addr[39084]= -2103375398;
assign addr[39085]= -2095330553;
assign addr[39086]= -2086621133;
assign addr[39087]= -2077249901;
assign addr[39088]= -2067219829;
assign addr[39089]= -2056534099;
assign addr[39090]= -2045196100;
assign addr[39091]= -2033209426;
assign addr[39092]= -2020577882;
assign addr[39093]= -2007305472;
assign addr[39094]= -1993396407;
assign addr[39095]= -1978855097;
assign addr[39096]= -1963686155;
assign addr[39097]= -1947894393;
assign addr[39098]= -1931484818;
assign addr[39099]= -1914462636;
assign addr[39100]= -1896833245;
assign addr[39101]= -1878602237;
assign addr[39102]= -1859775393;
assign addr[39103]= -1840358687;
assign addr[39104]= -1820358275;
assign addr[39105]= -1799780501;
assign addr[39106]= -1778631892;
assign addr[39107]= -1756919156;
assign addr[39108]= -1734649179;
assign addr[39109]= -1711829025;
assign addr[39110]= -1688465931;
assign addr[39111]= -1664567307;
assign addr[39112]= -1640140734;
assign addr[39113]= -1615193959;
assign addr[39114]= -1589734894;
assign addr[39115]= -1563771613;
assign addr[39116]= -1537312353;
assign addr[39117]= -1510365504;
assign addr[39118]= -1482939614;
assign addr[39119]= -1455043381;
assign addr[39120]= -1426685652;
assign addr[39121]= -1397875423;
assign addr[39122]= -1368621831;
assign addr[39123]= -1338934154;
assign addr[39124]= -1308821808;
assign addr[39125]= -1278294345;
assign addr[39126]= -1247361445;
assign addr[39127]= -1216032921;
assign addr[39128]= -1184318708;
assign addr[39129]= -1152228866;
assign addr[39130]= -1119773573;
assign addr[39131]= -1086963121;
assign addr[39132]= -1053807919;
assign addr[39133]= -1020318481;
assign addr[39134]= -986505429;
assign addr[39135]= -952379488;
assign addr[39136]= -917951481;
assign addr[39137]= -883232329;
assign addr[39138]= -848233042;
assign addr[39139]= -812964722;
assign addr[39140]= -777438554;
assign addr[39141]= -741665807;
assign addr[39142]= -705657826;
assign addr[39143]= -669426032;
assign addr[39144]= -632981917;
assign addr[39145]= -596337040;
assign addr[39146]= -559503022;
assign addr[39147]= -522491548;
assign addr[39148]= -485314355;
assign addr[39149]= -447983235;
assign addr[39150]= -410510029;
assign addr[39151]= -372906622;
assign addr[39152]= -335184940;
assign addr[39153]= -297356948;
assign addr[39154]= -259434643;
assign addr[39155]= -221430054;
assign addr[39156]= -183355234;
assign addr[39157]= -145222259;
assign addr[39158]= -107043224;
assign addr[39159]= -68830239;
assign addr[39160]= -30595422;
assign addr[39161]= 7649098;
assign addr[39162]= 45891193;
assign addr[39163]= 84118732;
assign addr[39164]= 122319591;
assign addr[39165]= 160481654;
assign addr[39166]= 198592817;
assign addr[39167]= 236640993;
assign addr[39168]= 274614114;
assign addr[39169]= 312500135;
assign addr[39170]= 350287041;
assign addr[39171]= 387962847;
assign addr[39172]= 425515602;
assign addr[39173]= 462933398;
assign addr[39174]= 500204365;
assign addr[39175]= 537316682;
assign addr[39176]= 574258580;
assign addr[39177]= 611018340;
assign addr[39178]= 647584304;
assign addr[39179]= 683944874;
assign addr[39180]= 720088517;
assign addr[39181]= 756003771;
assign addr[39182]= 791679244;
assign addr[39183]= 827103620;
assign addr[39184]= 862265664;
assign addr[39185]= 897154224;
assign addr[39186]= 931758235;
assign addr[39187]= 966066720;
assign addr[39188]= 1000068799;
assign addr[39189]= 1033753687;
assign addr[39190]= 1067110699;
assign addr[39191]= 1100129257;
assign addr[39192]= 1132798888;
assign addr[39193]= 1165109230;
assign addr[39194]= 1197050035;
assign addr[39195]= 1228611172;
assign addr[39196]= 1259782632;
assign addr[39197]= 1290554528;
assign addr[39198]= 1320917099;
assign addr[39199]= 1350860716;
assign addr[39200]= 1380375881;
assign addr[39201]= 1409453233;
assign addr[39202]= 1438083551;
assign addr[39203]= 1466257752;
assign addr[39204]= 1493966902;
assign addr[39205]= 1521202211;
assign addr[39206]= 1547955041;
assign addr[39207]= 1574216908;
assign addr[39208]= 1599979481;
assign addr[39209]= 1625234591;
assign addr[39210]= 1649974225;
assign addr[39211]= 1674190539;
assign addr[39212]= 1697875851;
assign addr[39213]= 1721022648;
assign addr[39214]= 1743623590;
assign addr[39215]= 1765671509;
assign addr[39216]= 1787159411;
assign addr[39217]= 1808080480;
assign addr[39218]= 1828428082;
assign addr[39219]= 1848195763;
assign addr[39220]= 1867377253;
assign addr[39221]= 1885966468;
assign addr[39222]= 1903957513;
assign addr[39223]= 1921344681;
assign addr[39224]= 1938122457;
assign addr[39225]= 1954285520;
assign addr[39226]= 1969828744;
assign addr[39227]= 1984747199;
assign addr[39228]= 1999036154;
assign addr[39229]= 2012691075;
assign addr[39230]= 2025707632;
assign addr[39231]= 2038081698;
assign addr[39232]= 2049809346;
assign addr[39233]= 2060886858;
assign addr[39234]= 2071310720;
assign addr[39235]= 2081077626;
assign addr[39236]= 2090184478;
assign addr[39237]= 2098628387;
assign addr[39238]= 2106406677;
assign addr[39239]= 2113516878;
assign addr[39240]= 2119956737;
assign addr[39241]= 2125724211;
assign addr[39242]= 2130817471;
assign addr[39243]= 2135234901;
assign addr[39244]= 2138975100;
assign addr[39245]= 2142036881;
assign addr[39246]= 2144419275;
assign addr[39247]= 2146121524;
assign addr[39248]= 2147143090;
assign addr[39249]= 2147483648;
assign addr[39250]= 2147143090;
assign addr[39251]= 2146121524;
assign addr[39252]= 2144419275;
assign addr[39253]= 2142036881;
assign addr[39254]= 2138975100;
assign addr[39255]= 2135234901;
assign addr[39256]= 2130817471;
assign addr[39257]= 2125724211;
assign addr[39258]= 2119956737;
assign addr[39259]= 2113516878;
assign addr[39260]= 2106406677;
assign addr[39261]= 2098628387;
assign addr[39262]= 2090184478;
assign addr[39263]= 2081077626;
assign addr[39264]= 2071310720;
assign addr[39265]= 2060886858;
assign addr[39266]= 2049809346;
assign addr[39267]= 2038081698;
assign addr[39268]= 2025707632;
assign addr[39269]= 2012691075;
assign addr[39270]= 1999036154;
assign addr[39271]= 1984747199;
assign addr[39272]= 1969828744;
assign addr[39273]= 1954285520;
assign addr[39274]= 1938122457;
assign addr[39275]= 1921344681;
assign addr[39276]= 1903957513;
assign addr[39277]= 1885966468;
assign addr[39278]= 1867377253;
assign addr[39279]= 1848195763;
assign addr[39280]= 1828428082;
assign addr[39281]= 1808080480;
assign addr[39282]= 1787159411;
assign addr[39283]= 1765671509;
assign addr[39284]= 1743623590;
assign addr[39285]= 1721022648;
assign addr[39286]= 1697875851;
assign addr[39287]= 1674190539;
assign addr[39288]= 1649974225;
assign addr[39289]= 1625234591;
assign addr[39290]= 1599979481;
assign addr[39291]= 1574216908;
assign addr[39292]= 1547955041;
assign addr[39293]= 1521202211;
assign addr[39294]= 1493966902;
assign addr[39295]= 1466257752;
assign addr[39296]= 1438083551;
assign addr[39297]= 1409453233;
assign addr[39298]= 1380375881;
assign addr[39299]= 1350860716;
assign addr[39300]= 1320917099;
assign addr[39301]= 1290554528;
assign addr[39302]= 1259782632;
assign addr[39303]= 1228611172;
assign addr[39304]= 1197050035;
assign addr[39305]= 1165109230;
assign addr[39306]= 1132798888;
assign addr[39307]= 1100129257;
assign addr[39308]= 1067110699;
assign addr[39309]= 1033753687;
assign addr[39310]= 1000068799;
assign addr[39311]= 966066720;
assign addr[39312]= 931758235;
assign addr[39313]= 897154224;
assign addr[39314]= 862265664;
assign addr[39315]= 827103620;
assign addr[39316]= 791679244;
assign addr[39317]= 756003771;
assign addr[39318]= 720088517;
assign addr[39319]= 683944874;
assign addr[39320]= 647584304;
assign addr[39321]= 611018340;
assign addr[39322]= 574258580;
assign addr[39323]= 537316682;
assign addr[39324]= 500204365;
assign addr[39325]= 462933398;
assign addr[39326]= 425515602;
assign addr[39327]= 387962847;
assign addr[39328]= 350287041;
assign addr[39329]= 312500135;
assign addr[39330]= 274614114;
assign addr[39331]= 236640993;
assign addr[39332]= 198592817;
assign addr[39333]= 160481654;
assign addr[39334]= 122319591;
assign addr[39335]= 84118732;
assign addr[39336]= 45891193;
assign addr[39337]= 7649098;
assign addr[39338]= -30595422;
assign addr[39339]= -68830239;
assign addr[39340]= -107043224;
assign addr[39341]= -145222259;
assign addr[39342]= -183355234;
assign addr[39343]= -221430054;
assign addr[39344]= -259434643;
assign addr[39345]= -297356948;
assign addr[39346]= -335184940;
assign addr[39347]= -372906622;
assign addr[39348]= -410510029;
assign addr[39349]= -447983235;
assign addr[39350]= -485314355;
assign addr[39351]= -522491548;
assign addr[39352]= -559503022;
assign addr[39353]= -596337040;
assign addr[39354]= -632981917;
assign addr[39355]= -669426032;
assign addr[39356]= -705657826;
assign addr[39357]= -741665807;
assign addr[39358]= -777438554;
assign addr[39359]= -812964722;
assign addr[39360]= -848233042;
assign addr[39361]= -883232329;
assign addr[39362]= -917951481;
assign addr[39363]= -952379488;
assign addr[39364]= -986505429;
assign addr[39365]= -1020318481;
assign addr[39366]= -1053807919;
assign addr[39367]= -1086963121;
assign addr[39368]= -1119773573;
assign addr[39369]= -1152228866;
assign addr[39370]= -1184318708;
assign addr[39371]= -1216032921;
assign addr[39372]= -1247361445;
assign addr[39373]= -1278294345;
assign addr[39374]= -1308821808;
assign addr[39375]= -1338934154;
assign addr[39376]= -1368621831;
assign addr[39377]= -1397875423;
assign addr[39378]= -1426685652;
assign addr[39379]= -1455043381;
assign addr[39380]= -1482939614;
assign addr[39381]= -1510365504;
assign addr[39382]= -1537312353;
assign addr[39383]= -1563771613;
assign addr[39384]= -1589734894;
assign addr[39385]= -1615193959;
assign addr[39386]= -1640140734;
assign addr[39387]= -1664567307;
assign addr[39388]= -1688465931;
assign addr[39389]= -1711829025;
assign addr[39390]= -1734649179;
assign addr[39391]= -1756919156;
assign addr[39392]= -1778631892;
assign addr[39393]= -1799780501;
assign addr[39394]= -1820358275;
assign addr[39395]= -1840358687;
assign addr[39396]= -1859775393;
assign addr[39397]= -1878602237;
assign addr[39398]= -1896833245;
assign addr[39399]= -1914462636;
assign addr[39400]= -1931484818;
assign addr[39401]= -1947894393;
assign addr[39402]= -1963686155;
assign addr[39403]= -1978855097;
assign addr[39404]= -1993396407;
assign addr[39405]= -2007305472;
assign addr[39406]= -2020577882;
assign addr[39407]= -2033209426;
assign addr[39408]= -2045196100;
assign addr[39409]= -2056534099;
assign addr[39410]= -2067219829;
assign addr[39411]= -2077249901;
assign addr[39412]= -2086621133;
assign addr[39413]= -2095330553;
assign addr[39414]= -2103375398;
assign addr[39415]= -2110753117;
assign addr[39416]= -2117461370;
assign addr[39417]= -2123498030;
assign addr[39418]= -2128861181;
assign addr[39419]= -2133549123;
assign addr[39420]= -2137560369;
assign addr[39421]= -2140893646;
assign addr[39422]= -2143547897;
assign addr[39423]= -2145522281;
assign addr[39424]= -2146816171;
assign addr[39425]= -2147429158;
assign addr[39426]= -2147361045;
assign addr[39427]= -2146611856;
assign addr[39428]= -2145181827;
assign addr[39429]= -2143071413;
assign addr[39430]= -2140281282;
assign addr[39431]= -2136812319;
assign addr[39432]= -2132665626;
assign addr[39433]= -2127842516;
assign addr[39434]= -2122344521;
assign addr[39435]= -2116173382;
assign addr[39436]= -2109331059;
assign addr[39437]= -2101819720;
assign addr[39438]= -2093641749;
assign addr[39439]= -2084799740;
assign addr[39440]= -2075296495;
assign addr[39441]= -2065135031;
assign addr[39442]= -2054318569;
assign addr[39443]= -2042850540;
assign addr[39444]= -2030734582;
assign addr[39445]= -2017974537;
assign addr[39446]= -2004574453;
assign addr[39447]= -1990538579;
assign addr[39448]= -1975871368;
assign addr[39449]= -1960577471;
assign addr[39450]= -1944661739;
assign addr[39451]= -1928129220;
assign addr[39452]= -1910985158;
assign addr[39453]= -1893234990;
assign addr[39454]= -1874884346;
assign addr[39455]= -1855939047;
assign addr[39456]= -1836405100;
assign addr[39457]= -1816288703;
assign addr[39458]= -1795596234;
assign addr[39459]= -1774334257;
assign addr[39460]= -1752509516;
assign addr[39461]= -1730128933;
assign addr[39462]= -1707199606;
assign addr[39463]= -1683728808;
assign addr[39464]= -1659723983;
assign addr[39465]= -1635192744;
assign addr[39466]= -1610142873;
assign addr[39467]= -1584582314;
assign addr[39468]= -1558519173;
assign addr[39469]= -1531961719;
assign addr[39470]= -1504918373;
assign addr[39471]= -1477397714;
assign addr[39472]= -1449408469;
assign addr[39473]= -1420959516;
assign addr[39474]= -1392059879;
assign addr[39475]= -1362718723;
assign addr[39476]= -1332945355;
assign addr[39477]= -1302749217;
assign addr[39478]= -1272139887;
assign addr[39479]= -1241127074;
assign addr[39480]= -1209720613;
assign addr[39481]= -1177930466;
assign addr[39482]= -1145766716;
assign addr[39483]= -1113239564;
assign addr[39484]= -1080359326;
assign addr[39485]= -1047136432;
assign addr[39486]= -1013581418;
assign addr[39487]= -979704927;
assign addr[39488]= -945517704;
assign addr[39489]= -911030591;
assign addr[39490]= -876254528;
assign addr[39491]= -841200544;
assign addr[39492]= -805879757;
assign addr[39493]= -770303369;
assign addr[39494]= -734482665;
assign addr[39495]= -698429006;
assign addr[39496]= -662153826;
assign addr[39497]= -625668632;
assign addr[39498]= -588984994;
assign addr[39499]= -552114549;
assign addr[39500]= -515068990;
assign addr[39501]= -477860067;
assign addr[39502]= -440499581;
assign addr[39503]= -402999383;
assign addr[39504]= -365371365;
assign addr[39505]= -327627463;
assign addr[39506]= -289779648;
assign addr[39507]= -251839923;
assign addr[39508]= -213820322;
assign addr[39509]= -175732905;
assign addr[39510]= -137589750;
assign addr[39511]= -99402956;
assign addr[39512]= -61184634;
assign addr[39513]= -22946906;
assign addr[39514]= 15298099;
assign addr[39515]= 53538253;
assign addr[39516]= 91761426;
assign addr[39517]= 129955495;
assign addr[39518]= 168108346;
assign addr[39519]= 206207878;
assign addr[39520]= 244242007;
assign addr[39521]= 282198671;
assign addr[39522]= 320065829;
assign addr[39523]= 357831473;
assign addr[39524]= 395483624;
assign addr[39525]= 433010339;
assign addr[39526]= 470399716;
assign addr[39527]= 507639898;
assign addr[39528]= 544719071;
assign addr[39529]= 581625477;
assign addr[39530]= 618347408;
assign addr[39531]= 654873219;
assign addr[39532]= 691191324;
assign addr[39533]= 727290205;
assign addr[39534]= 763158411;
assign addr[39535]= 798784567;
assign addr[39536]= 834157373;
assign addr[39537]= 869265610;
assign addr[39538]= 904098143;
assign addr[39539]= 938643924;
assign addr[39540]= 972891995;
assign addr[39541]= 1006831495;
assign addr[39542]= 1040451659;
assign addr[39543]= 1073741824;
assign addr[39544]= 1106691431;
assign addr[39545]= 1139290029;
assign addr[39546]= 1171527280;
assign addr[39547]= 1203392958;
assign addr[39548]= 1234876957;
assign addr[39549]= 1265969291;
assign addr[39550]= 1296660098;
assign addr[39551]= 1326939644;
assign addr[39552]= 1356798326;
assign addr[39553]= 1386226674;
assign addr[39554]= 1415215352;
assign addr[39555]= 1443755168;
assign addr[39556]= 1471837070;
assign addr[39557]= 1499452149;
assign addr[39558]= 1526591649;
assign addr[39559]= 1553246960;
assign addr[39560]= 1579409630;
assign addr[39561]= 1605071359;
assign addr[39562]= 1630224009;
assign addr[39563]= 1654859602;
assign addr[39564]= 1678970324;
assign addr[39565]= 1702548529;
assign addr[39566]= 1725586737;
assign addr[39567]= 1748077642;
assign addr[39568]= 1770014111;
assign addr[39569]= 1791389186;
assign addr[39570]= 1812196087;
assign addr[39571]= 1832428215;
assign addr[39572]= 1852079154;
assign addr[39573]= 1871142669;
assign addr[39574]= 1889612716;
assign addr[39575]= 1907483436;
assign addr[39576]= 1924749160;
assign addr[39577]= 1941404413;
assign addr[39578]= 1957443913;
assign addr[39579]= 1972862571;
assign addr[39580]= 1987655498;
assign addr[39581]= 2001818002;
assign addr[39582]= 2015345591;
assign addr[39583]= 2028233973;
assign addr[39584]= 2040479063;
assign addr[39585]= 2052076975;
assign addr[39586]= 2063024031;
assign addr[39587]= 2073316760;
assign addr[39588]= 2082951896;
assign addr[39589]= 2091926384;
assign addr[39590]= 2100237377;
assign addr[39591]= 2107882239;
assign addr[39592]= 2114858546;
assign addr[39593]= 2121164085;
assign addr[39594]= 2126796855;
assign addr[39595]= 2131755071;
assign addr[39596]= 2136037160;
assign addr[39597]= 2139641764;
assign addr[39598]= 2142567738;
assign addr[39599]= 2144814157;
assign addr[39600]= 2146380306;
assign addr[39601]= 2147265689;
assign addr[39602]= 2147470025;
assign addr[39603]= 2146993250;
assign addr[39604]= 2145835515;
assign addr[39605]= 2143997187;
assign addr[39606]= 2141478848;
assign addr[39607]= 2138281298;
assign addr[39608]= 2134405552;
assign addr[39609]= 2129852837;
assign addr[39610]= 2124624598;
assign addr[39611]= 2118722494;
assign addr[39612]= 2112148396;
assign addr[39613]= 2104904390;
assign addr[39614]= 2096992772;
assign addr[39615]= 2088416053;
assign addr[39616]= 2079176953;
assign addr[39617]= 2069278401;
assign addr[39618]= 2058723538;
assign addr[39619]= 2047515711;
assign addr[39620]= 2035658475;
assign addr[39621]= 2023155591;
assign addr[39622]= 2010011024;
assign addr[39623]= 1996228943;
assign addr[39624]= 1981813720;
assign addr[39625]= 1966769926;
assign addr[39626]= 1951102334;
assign addr[39627]= 1934815911;
assign addr[39628]= 1917915825;
assign addr[39629]= 1900407434;
assign addr[39630]= 1882296293;
assign addr[39631]= 1863588145;
assign addr[39632]= 1844288924;
assign addr[39633]= 1824404752;
assign addr[39634]= 1803941934;
assign addr[39635]= 1782906961;
assign addr[39636]= 1761306505;
assign addr[39637]= 1739147417;
assign addr[39638]= 1716436725;
assign addr[39639]= 1693181631;
assign addr[39640]= 1669389513;
assign addr[39641]= 1645067915;
assign addr[39642]= 1620224553;
assign addr[39643]= 1594867305;
assign addr[39644]= 1569004214;
assign addr[39645]= 1542643483;
assign addr[39646]= 1515793473;
assign addr[39647]= 1488462700;
assign addr[39648]= 1460659832;
assign addr[39649]= 1432393688;
assign addr[39650]= 1403673233;
assign addr[39651]= 1374507575;
assign addr[39652]= 1344905966;
assign addr[39653]= 1314877795;
assign addr[39654]= 1284432584;
assign addr[39655]= 1253579991;
assign addr[39656]= 1222329801;
assign addr[39657]= 1190691925;
assign addr[39658]= 1158676398;
assign addr[39659]= 1126293375;
assign addr[39660]= 1093553126;
assign addr[39661]= 1060466036;
assign addr[39662]= 1027042599;
assign addr[39663]= 993293415;
assign addr[39664]= 959229189;
assign addr[39665]= 924860725;
assign addr[39666]= 890198924;
assign addr[39667]= 855254778;
assign addr[39668]= 820039373;
assign addr[39669]= 784563876;
assign addr[39670]= 748839539;
assign addr[39671]= 712877694;
assign addr[39672]= 676689746;
assign addr[39673]= 640287172;
assign addr[39674]= 603681519;
assign addr[39675]= 566884397;
assign addr[39676]= 529907477;
assign addr[39677]= 492762486;
assign addr[39678]= 455461206;
assign addr[39679]= 418015468;
assign addr[39680]= 380437148;
assign addr[39681]= 342738165;
assign addr[39682]= 304930476;
assign addr[39683]= 267026072;
assign addr[39684]= 229036977;
assign addr[39685]= 190975237;
assign addr[39686]= 152852926;
assign addr[39687]= 114682135;
assign addr[39688]= 76474970;
assign addr[39689]= 38243550;
assign addr[39690]= 0;
assign addr[39691]= -38243550;
assign addr[39692]= -76474970;
assign addr[39693]= -114682135;
assign addr[39694]= -152852926;
assign addr[39695]= -190975237;
assign addr[39696]= -229036977;
assign addr[39697]= -267026072;
assign addr[39698]= -304930476;
assign addr[39699]= -342738165;
assign addr[39700]= -380437148;
assign addr[39701]= -418015468;
assign addr[39702]= -455461206;
assign addr[39703]= -492762486;
assign addr[39704]= -529907477;
assign addr[39705]= -566884397;
assign addr[39706]= -603681519;
assign addr[39707]= -640287172;
assign addr[39708]= -676689746;
assign addr[39709]= -712877694;
assign addr[39710]= -748839539;
assign addr[39711]= -784563876;
assign addr[39712]= -820039373;
assign addr[39713]= -855254778;
assign addr[39714]= -890198924;
assign addr[39715]= -924860725;
assign addr[39716]= -959229189;
assign addr[39717]= -993293415;
assign addr[39718]= -1027042599;
assign addr[39719]= -1060466036;
assign addr[39720]= -1093553126;
assign addr[39721]= -1126293375;
assign addr[39722]= -1158676398;
assign addr[39723]= -1190691925;
assign addr[39724]= -1222329801;
assign addr[39725]= -1253579991;
assign addr[39726]= -1284432584;
assign addr[39727]= -1314877795;
assign addr[39728]= -1344905966;
assign addr[39729]= -1374507575;
assign addr[39730]= -1403673233;
assign addr[39731]= -1432393688;
assign addr[39732]= -1460659832;
assign addr[39733]= -1488462700;
assign addr[39734]= -1515793473;
assign addr[39735]= -1542643483;
assign addr[39736]= -1569004214;
assign addr[39737]= -1594867305;
assign addr[39738]= -1620224553;
assign addr[39739]= -1645067915;
assign addr[39740]= -1669389513;
assign addr[39741]= -1693181631;
assign addr[39742]= -1716436725;
assign addr[39743]= -1739147417;
assign addr[39744]= -1761306505;
assign addr[39745]= -1782906961;
assign addr[39746]= -1803941934;
assign addr[39747]= -1824404752;
assign addr[39748]= -1844288924;
assign addr[39749]= -1863588145;
assign addr[39750]= -1882296293;
assign addr[39751]= -1900407434;
assign addr[39752]= -1917915825;
assign addr[39753]= -1934815911;
assign addr[39754]= -1951102334;
assign addr[39755]= -1966769926;
assign addr[39756]= -1981813720;
assign addr[39757]= -1996228943;
assign addr[39758]= -2010011024;
assign addr[39759]= -2023155591;
assign addr[39760]= -2035658475;
assign addr[39761]= -2047515711;
assign addr[39762]= -2058723538;
assign addr[39763]= -2069278401;
assign addr[39764]= -2079176953;
assign addr[39765]= -2088416053;
assign addr[39766]= -2096992772;
assign addr[39767]= -2104904390;
assign addr[39768]= -2112148396;
assign addr[39769]= -2118722494;
assign addr[39770]= -2124624598;
assign addr[39771]= -2129852837;
assign addr[39772]= -2134405552;
assign addr[39773]= -2138281298;
assign addr[39774]= -2141478848;
assign addr[39775]= -2143997187;
assign addr[39776]= -2145835515;
assign addr[39777]= -2146993250;
assign addr[39778]= -2147470025;
assign addr[39779]= -2147265689;
assign addr[39780]= -2146380306;
assign addr[39781]= -2144814157;
assign addr[39782]= -2142567738;
assign addr[39783]= -2139641764;
assign addr[39784]= -2136037160;
assign addr[39785]= -2131755071;
assign addr[39786]= -2126796855;
assign addr[39787]= -2121164085;
assign addr[39788]= -2114858546;
assign addr[39789]= -2107882239;
assign addr[39790]= -2100237377;
assign addr[39791]= -2091926384;
assign addr[39792]= -2082951896;
assign addr[39793]= -2073316760;
assign addr[39794]= -2063024031;
assign addr[39795]= -2052076975;
assign addr[39796]= -2040479063;
assign addr[39797]= -2028233973;
assign addr[39798]= -2015345591;
assign addr[39799]= -2001818002;
assign addr[39800]= -1987655498;
assign addr[39801]= -1972862571;
assign addr[39802]= -1957443913;
assign addr[39803]= -1941404413;
assign addr[39804]= -1924749160;
assign addr[39805]= -1907483436;
assign addr[39806]= -1889612716;
assign addr[39807]= -1871142669;
assign addr[39808]= -1852079154;
assign addr[39809]= -1832428215;
assign addr[39810]= -1812196087;
assign addr[39811]= -1791389186;
assign addr[39812]= -1770014111;
assign addr[39813]= -1748077642;
assign addr[39814]= -1725586737;
assign addr[39815]= -1702548529;
assign addr[39816]= -1678970324;
assign addr[39817]= -1654859602;
assign addr[39818]= -1630224009;
assign addr[39819]= -1605071359;
assign addr[39820]= -1579409630;
assign addr[39821]= -1553246960;
assign addr[39822]= -1526591649;
assign addr[39823]= -1499452149;
assign addr[39824]= -1471837070;
assign addr[39825]= -1443755168;
assign addr[39826]= -1415215352;
assign addr[39827]= -1386226674;
assign addr[39828]= -1356798326;
assign addr[39829]= -1326939644;
assign addr[39830]= -1296660098;
assign addr[39831]= -1265969291;
assign addr[39832]= -1234876957;
assign addr[39833]= -1203392958;
assign addr[39834]= -1171527280;
assign addr[39835]= -1139290029;
assign addr[39836]= -1106691431;
assign addr[39837]= -1073741824;
assign addr[39838]= -1040451659;
assign addr[39839]= -1006831495;
assign addr[39840]= -972891995;
assign addr[39841]= -938643924;
assign addr[39842]= -904098143;
assign addr[39843]= -869265610;
assign addr[39844]= -834157373;
assign addr[39845]= -798784567;
assign addr[39846]= -763158411;
assign addr[39847]= -727290205;
assign addr[39848]= -691191324;
assign addr[39849]= -654873219;
assign addr[39850]= -618347408;
assign addr[39851]= -581625477;
assign addr[39852]= -544719071;
assign addr[39853]= -507639898;
assign addr[39854]= -470399716;
assign addr[39855]= -433010339;
assign addr[39856]= -395483624;
assign addr[39857]= -357831473;
assign addr[39858]= -320065829;
assign addr[39859]= -282198671;
assign addr[39860]= -244242007;
assign addr[39861]= -206207878;
assign addr[39862]= -168108346;
assign addr[39863]= -129955495;
assign addr[39864]= -91761426;
assign addr[39865]= -53538253;
assign addr[39866]= -15298099;
assign addr[39867]= 22946906;
assign addr[39868]= 61184634;
assign addr[39869]= 99402956;
assign addr[39870]= 137589750;
assign addr[39871]= 175732905;
assign addr[39872]= 213820322;
assign addr[39873]= 251839923;
assign addr[39874]= 289779648;
assign addr[39875]= 327627463;
assign addr[39876]= 365371365;
assign addr[39877]= 402999383;
assign addr[39878]= 440499581;
assign addr[39879]= 477860067;
assign addr[39880]= 515068990;
assign addr[39881]= 552114549;
assign addr[39882]= 588984994;
assign addr[39883]= 625668632;
assign addr[39884]= 662153826;
assign addr[39885]= 698429006;
assign addr[39886]= 734482665;
assign addr[39887]= 770303369;
assign addr[39888]= 805879757;
assign addr[39889]= 841200544;
assign addr[39890]= 876254528;
assign addr[39891]= 911030591;
assign addr[39892]= 945517704;
assign addr[39893]= 979704927;
assign addr[39894]= 1013581418;
assign addr[39895]= 1047136432;
assign addr[39896]= 1080359326;
assign addr[39897]= 1113239564;
assign addr[39898]= 1145766716;
assign addr[39899]= 1177930466;
assign addr[39900]= 1209720613;
assign addr[39901]= 1241127074;
assign addr[39902]= 1272139887;
assign addr[39903]= 1302749217;
assign addr[39904]= 1332945355;
assign addr[39905]= 1362718723;
assign addr[39906]= 1392059879;
assign addr[39907]= 1420959516;
assign addr[39908]= 1449408469;
assign addr[39909]= 1477397714;
assign addr[39910]= 1504918373;
assign addr[39911]= 1531961719;
assign addr[39912]= 1558519173;
assign addr[39913]= 1584582314;
assign addr[39914]= 1610142873;
assign addr[39915]= 1635192744;
assign addr[39916]= 1659723983;
assign addr[39917]= 1683728808;
assign addr[39918]= 1707199606;
assign addr[39919]= 1730128933;
assign addr[39920]= 1752509516;
assign addr[39921]= 1774334257;
assign addr[39922]= 1795596234;
assign addr[39923]= 1816288703;
assign addr[39924]= 1836405100;
assign addr[39925]= 1855939047;
assign addr[39926]= 1874884346;
assign addr[39927]= 1893234990;
assign addr[39928]= 1910985158;
assign addr[39929]= 1928129220;
assign addr[39930]= 1944661739;
assign addr[39931]= 1960577471;
assign addr[39932]= 1975871368;
assign addr[39933]= 1990538579;
assign addr[39934]= 2004574453;
assign addr[39935]= 2017974537;
assign addr[39936]= 2030734582;
assign addr[39937]= 2042850540;
assign addr[39938]= 2054318569;
assign addr[39939]= 2065135031;
assign addr[39940]= 2075296495;
assign addr[39941]= 2084799740;
assign addr[39942]= 2093641749;
assign addr[39943]= 2101819720;
assign addr[39944]= 2109331059;
assign addr[39945]= 2116173382;
assign addr[39946]= 2122344521;
assign addr[39947]= 2127842516;
assign addr[39948]= 2132665626;
assign addr[39949]= 2136812319;
assign addr[39950]= 2140281282;
assign addr[39951]= 2143071413;
assign addr[39952]= 2145181827;
assign addr[39953]= 2146611856;
assign addr[39954]= 2147361045;
assign addr[39955]= 2147429158;
assign addr[39956]= 2146816171;
assign addr[39957]= 2145522281;
assign addr[39958]= 2143547897;
assign addr[39959]= 2140893646;
assign addr[39960]= 2137560369;
assign addr[39961]= 2133549123;
assign addr[39962]= 2128861181;
assign addr[39963]= 2123498030;
assign addr[39964]= 2117461370;
assign addr[39965]= 2110753117;
assign addr[39966]= 2103375398;
assign addr[39967]= 2095330553;
assign addr[39968]= 2086621133;
assign addr[39969]= 2077249901;
assign addr[39970]= 2067219829;
assign addr[39971]= 2056534099;
assign addr[39972]= 2045196100;
assign addr[39973]= 2033209426;
assign addr[39974]= 2020577882;
assign addr[39975]= 2007305472;
assign addr[39976]= 1993396407;
assign addr[39977]= 1978855097;
assign addr[39978]= 1963686155;
assign addr[39979]= 1947894393;
assign addr[39980]= 1931484818;
assign addr[39981]= 1914462636;
assign addr[39982]= 1896833245;
assign addr[39983]= 1878602237;
assign addr[39984]= 1859775393;
assign addr[39985]= 1840358687;
assign addr[39986]= 1820358275;
assign addr[39987]= 1799780501;
assign addr[39988]= 1778631892;
assign addr[39989]= 1756919156;
assign addr[39990]= 1734649179;
assign addr[39991]= 1711829025;
assign addr[39992]= 1688465931;
assign addr[39993]= 1664567307;
assign addr[39994]= 1640140734;
assign addr[39995]= 1615193959;
assign addr[39996]= 1589734894;
assign addr[39997]= 1563771613;
assign addr[39998]= 1537312353;
assign addr[39999]= 1510365504;
assign addr[40000]= 1482939614;
assign addr[40001]= 1455043381;
assign addr[40002]= 1426685652;
assign addr[40003]= 1397875423;
assign addr[40004]= 1368621831;
assign addr[40005]= 1338934154;
assign addr[40006]= 1308821808;
assign addr[40007]= 1278294345;
assign addr[40008]= 1247361445;
assign addr[40009]= 1216032921;
assign addr[40010]= 1184318708;
assign addr[40011]= 1152228866;
assign addr[40012]= 1119773573;
assign addr[40013]= 1086963121;
assign addr[40014]= 1053807919;
assign addr[40015]= 1020318481;
assign addr[40016]= 986505429;
assign addr[40017]= 952379488;
assign addr[40018]= 917951481;
assign addr[40019]= 883232329;
assign addr[40020]= 848233042;
assign addr[40021]= 812964722;
assign addr[40022]= 777438554;
assign addr[40023]= 741665807;
assign addr[40024]= 705657826;
assign addr[40025]= 669426032;
assign addr[40026]= 632981917;
assign addr[40027]= 596337040;
assign addr[40028]= 559503022;
assign addr[40029]= 522491548;
assign addr[40030]= 485314355;
assign addr[40031]= 447983235;
assign addr[40032]= 410510029;
assign addr[40033]= 372906622;
assign addr[40034]= 335184940;
assign addr[40035]= 297356948;
assign addr[40036]= 259434643;
assign addr[40037]= 221430054;
assign addr[40038]= 183355234;
assign addr[40039]= 145222259;
assign addr[40040]= 107043224;
assign addr[40041]= 68830239;
assign addr[40042]= 30595422;
assign addr[40043]= -7649098;
assign addr[40044]= -45891193;
assign addr[40045]= -84118732;
assign addr[40046]= -122319591;
assign addr[40047]= -160481654;
assign addr[40048]= -198592817;
assign addr[40049]= -236640993;
assign addr[40050]= -274614114;
assign addr[40051]= -312500135;
assign addr[40052]= -350287041;
assign addr[40053]= -387962847;
assign addr[40054]= -425515602;
assign addr[40055]= -462933398;
assign addr[40056]= -500204365;
assign addr[40057]= -537316682;
assign addr[40058]= -574258580;
assign addr[40059]= -611018340;
assign addr[40060]= -647584304;
assign addr[40061]= -683944874;
assign addr[40062]= -720088517;
assign addr[40063]= -756003771;
assign addr[40064]= -791679244;
assign addr[40065]= -827103620;
assign addr[40066]= -862265664;
assign addr[40067]= -897154224;
assign addr[40068]= -931758235;
assign addr[40069]= -966066720;
assign addr[40070]= -1000068799;
assign addr[40071]= -1033753687;
assign addr[40072]= -1067110699;
assign addr[40073]= -1100129257;
assign addr[40074]= -1132798888;
assign addr[40075]= -1165109230;
assign addr[40076]= -1197050035;
assign addr[40077]= -1228611172;
assign addr[40078]= -1259782632;
assign addr[40079]= -1290554528;
assign addr[40080]= -1320917099;
assign addr[40081]= -1350860716;
assign addr[40082]= -1380375881;
assign addr[40083]= -1409453233;
assign addr[40084]= -1438083551;
assign addr[40085]= -1466257752;
assign addr[40086]= -1493966902;
assign addr[40087]= -1521202211;
assign addr[40088]= -1547955041;
assign addr[40089]= -1574216908;
assign addr[40090]= -1599979481;
assign addr[40091]= -1625234591;
assign addr[40092]= -1649974225;
assign addr[40093]= -1674190539;
assign addr[40094]= -1697875851;
assign addr[40095]= -1721022648;
assign addr[40096]= -1743623590;
assign addr[40097]= -1765671509;
assign addr[40098]= -1787159411;
assign addr[40099]= -1808080480;
assign addr[40100]= -1828428082;
assign addr[40101]= -1848195763;
assign addr[40102]= -1867377253;
assign addr[40103]= -1885966468;
assign addr[40104]= -1903957513;
assign addr[40105]= -1921344681;
assign addr[40106]= -1938122457;
assign addr[40107]= -1954285520;
assign addr[40108]= -1969828744;
assign addr[40109]= -1984747199;
assign addr[40110]= -1999036154;
assign addr[40111]= -2012691075;
assign addr[40112]= -2025707632;
assign addr[40113]= -2038081698;
assign addr[40114]= -2049809346;
assign addr[40115]= -2060886858;
assign addr[40116]= -2071310720;
assign addr[40117]= -2081077626;
assign addr[40118]= -2090184478;
assign addr[40119]= -2098628387;
assign addr[40120]= -2106406677;
assign addr[40121]= -2113516878;
assign addr[40122]= -2119956737;
assign addr[40123]= -2125724211;
assign addr[40124]= -2130817471;
assign addr[40125]= -2135234901;
assign addr[40126]= -2138975100;
assign addr[40127]= -2142036881;
assign addr[40128]= -2144419275;
assign addr[40129]= -2146121524;
assign addr[40130]= -2147143090;
assign addr[40131]= -2147483648;
assign addr[40132]= -2147143090;
assign addr[40133]= -2146121524;
assign addr[40134]= -2144419275;
assign addr[40135]= -2142036881;
assign addr[40136]= -2138975100;
assign addr[40137]= -2135234901;
assign addr[40138]= -2130817471;
assign addr[40139]= -2125724211;
assign addr[40140]= -2119956737;
assign addr[40141]= -2113516878;
assign addr[40142]= -2106406677;
assign addr[40143]= -2098628387;
assign addr[40144]= -2090184478;
assign addr[40145]= -2081077626;
assign addr[40146]= -2071310720;
assign addr[40147]= -2060886858;
assign addr[40148]= -2049809346;
assign addr[40149]= -2038081698;
assign addr[40150]= -2025707632;
assign addr[40151]= -2012691075;
assign addr[40152]= -1999036154;
assign addr[40153]= -1984747199;
assign addr[40154]= -1969828744;
assign addr[40155]= -1954285520;
assign addr[40156]= -1938122457;
assign addr[40157]= -1921344681;
assign addr[40158]= -1903957513;
assign addr[40159]= -1885966468;
assign addr[40160]= -1867377253;
assign addr[40161]= -1848195763;
assign addr[40162]= -1828428082;
assign addr[40163]= -1808080480;
assign addr[40164]= -1787159411;
assign addr[40165]= -1765671509;
assign addr[40166]= -1743623590;
assign addr[40167]= -1721022648;
assign addr[40168]= -1697875851;
assign addr[40169]= -1674190539;
assign addr[40170]= -1649974225;
assign addr[40171]= -1625234591;
assign addr[40172]= -1599979481;
assign addr[40173]= -1574216908;
assign addr[40174]= -1547955041;
assign addr[40175]= -1521202211;
assign addr[40176]= -1493966902;
assign addr[40177]= -1466257752;
assign addr[40178]= -1438083551;
assign addr[40179]= -1409453233;
assign addr[40180]= -1380375881;
assign addr[40181]= -1350860716;
assign addr[40182]= -1320917099;
assign addr[40183]= -1290554528;
assign addr[40184]= -1259782632;
assign addr[40185]= -1228611172;
assign addr[40186]= -1197050035;
assign addr[40187]= -1165109230;
assign addr[40188]= -1132798888;
assign addr[40189]= -1100129257;
assign addr[40190]= -1067110699;
assign addr[40191]= -1033753687;
assign addr[40192]= -1000068799;
assign addr[40193]= -966066720;
assign addr[40194]= -931758235;
assign addr[40195]= -897154224;
assign addr[40196]= -862265664;
assign addr[40197]= -827103620;
assign addr[40198]= -791679244;
assign addr[40199]= -756003771;
assign addr[40200]= -720088517;
assign addr[40201]= -683944874;
assign addr[40202]= -647584304;
assign addr[40203]= -611018340;
assign addr[40204]= -574258580;
assign addr[40205]= -537316682;
assign addr[40206]= -500204365;
assign addr[40207]= -462933398;
assign addr[40208]= -425515602;
assign addr[40209]= -387962847;
assign addr[40210]= -350287041;
assign addr[40211]= -312500135;
assign addr[40212]= -274614114;
assign addr[40213]= -236640993;
assign addr[40214]= -198592817;
assign addr[40215]= -160481654;
assign addr[40216]= -122319591;
assign addr[40217]= -84118732;
assign addr[40218]= -45891193;
assign addr[40219]= -7649098;
assign addr[40220]= 30595422;
assign addr[40221]= 68830239;
assign addr[40222]= 107043224;
assign addr[40223]= 145222259;
assign addr[40224]= 183355234;
assign addr[40225]= 221430054;
assign addr[40226]= 259434643;
assign addr[40227]= 297356948;
assign addr[40228]= 335184940;
assign addr[40229]= 372906622;
assign addr[40230]= 410510029;
assign addr[40231]= 447983235;
assign addr[40232]= 485314355;
assign addr[40233]= 522491548;
assign addr[40234]= 559503022;
assign addr[40235]= 596337040;
assign addr[40236]= 632981917;
assign addr[40237]= 669426032;
assign addr[40238]= 705657826;
assign addr[40239]= 741665807;
assign addr[40240]= 777438554;
assign addr[40241]= 812964722;
assign addr[40242]= 848233042;
assign addr[40243]= 883232329;
assign addr[40244]= 917951481;
assign addr[40245]= 952379488;
assign addr[40246]= 986505429;
assign addr[40247]= 1020318481;
assign addr[40248]= 1053807919;
assign addr[40249]= 1086963121;
assign addr[40250]= 1119773573;
assign addr[40251]= 1152228866;
assign addr[40252]= 1184318708;
assign addr[40253]= 1216032921;
assign addr[40254]= 1247361445;
assign addr[40255]= 1278294345;
assign addr[40256]= 1308821808;
assign addr[40257]= 1338934154;
assign addr[40258]= 1368621831;
assign addr[40259]= 1397875423;
assign addr[40260]= 1426685652;
assign addr[40261]= 1455043381;
assign addr[40262]= 1482939614;
assign addr[40263]= 1510365504;
assign addr[40264]= 1537312353;
assign addr[40265]= 1563771613;
assign addr[40266]= 1589734894;
assign addr[40267]= 1615193959;
assign addr[40268]= 1640140734;
assign addr[40269]= 1664567307;
assign addr[40270]= 1688465931;
assign addr[40271]= 1711829025;
assign addr[40272]= 1734649179;
assign addr[40273]= 1756919156;
assign addr[40274]= 1778631892;
assign addr[40275]= 1799780501;
assign addr[40276]= 1820358275;
assign addr[40277]= 1840358687;
assign addr[40278]= 1859775393;
assign addr[40279]= 1878602237;
assign addr[40280]= 1896833245;
assign addr[40281]= 1914462636;
assign addr[40282]= 1931484818;
assign addr[40283]= 1947894393;
assign addr[40284]= 1963686155;
assign addr[40285]= 1978855097;
assign addr[40286]= 1993396407;
assign addr[40287]= 2007305472;
assign addr[40288]= 2020577882;
assign addr[40289]= 2033209426;
assign addr[40290]= 2045196100;
assign addr[40291]= 2056534099;
assign addr[40292]= 2067219829;
assign addr[40293]= 2077249901;
assign addr[40294]= 2086621133;
assign addr[40295]= 2095330553;
assign addr[40296]= 2103375398;
assign addr[40297]= 2110753117;
assign addr[40298]= 2117461370;
assign addr[40299]= 2123498030;
assign addr[40300]= 2128861181;
assign addr[40301]= 2133549123;
assign addr[40302]= 2137560369;
assign addr[40303]= 2140893646;
assign addr[40304]= 2143547897;
assign addr[40305]= 2145522281;
assign addr[40306]= 2146816171;
assign addr[40307]= 2147429158;
assign addr[40308]= 2147361045;
assign addr[40309]= 2146611856;
assign addr[40310]= 2145181827;
assign addr[40311]= 2143071413;
assign addr[40312]= 2140281282;
assign addr[40313]= 2136812319;
assign addr[40314]= 2132665626;
assign addr[40315]= 2127842516;
assign addr[40316]= 2122344521;
assign addr[40317]= 2116173382;
assign addr[40318]= 2109331059;
assign addr[40319]= 2101819720;
assign addr[40320]= 2093641749;
assign addr[40321]= 2084799740;
assign addr[40322]= 2075296495;
assign addr[40323]= 2065135031;
assign addr[40324]= 2054318569;
assign addr[40325]= 2042850540;
assign addr[40326]= 2030734582;
assign addr[40327]= 2017974537;
assign addr[40328]= 2004574453;
assign addr[40329]= 1990538579;
assign addr[40330]= 1975871368;
assign addr[40331]= 1960577471;
assign addr[40332]= 1944661739;
assign addr[40333]= 1928129220;
assign addr[40334]= 1910985158;
assign addr[40335]= 1893234990;
assign addr[40336]= 1874884346;
assign addr[40337]= 1855939047;
assign addr[40338]= 1836405100;
assign addr[40339]= 1816288703;
assign addr[40340]= 1795596234;
assign addr[40341]= 1774334257;
assign addr[40342]= 1752509516;
assign addr[40343]= 1730128933;
assign addr[40344]= 1707199606;
assign addr[40345]= 1683728808;
assign addr[40346]= 1659723983;
assign addr[40347]= 1635192744;
assign addr[40348]= 1610142873;
assign addr[40349]= 1584582314;
assign addr[40350]= 1558519173;
assign addr[40351]= 1531961719;
assign addr[40352]= 1504918373;
assign addr[40353]= 1477397714;
assign addr[40354]= 1449408469;
assign addr[40355]= 1420959516;
assign addr[40356]= 1392059879;
assign addr[40357]= 1362718723;
assign addr[40358]= 1332945355;
assign addr[40359]= 1302749217;
assign addr[40360]= 1272139887;
assign addr[40361]= 1241127074;
assign addr[40362]= 1209720613;
assign addr[40363]= 1177930466;
assign addr[40364]= 1145766716;
assign addr[40365]= 1113239564;
assign addr[40366]= 1080359326;
assign addr[40367]= 1047136432;
assign addr[40368]= 1013581418;
assign addr[40369]= 979704927;
assign addr[40370]= 945517704;
assign addr[40371]= 911030591;
assign addr[40372]= 876254528;
assign addr[40373]= 841200544;
assign addr[40374]= 805879757;
assign addr[40375]= 770303369;
assign addr[40376]= 734482665;
assign addr[40377]= 698429006;
assign addr[40378]= 662153826;
assign addr[40379]= 625668632;
assign addr[40380]= 588984994;
assign addr[40381]= 552114549;
assign addr[40382]= 515068990;
assign addr[40383]= 477860067;
assign addr[40384]= 440499581;
assign addr[40385]= 402999383;
assign addr[40386]= 365371365;
assign addr[40387]= 327627463;
assign addr[40388]= 289779648;
assign addr[40389]= 251839923;
assign addr[40390]= 213820322;
assign addr[40391]= 175732905;
assign addr[40392]= 137589750;
assign addr[40393]= 99402956;
assign addr[40394]= 61184634;
assign addr[40395]= 22946906;
assign addr[40396]= -15298099;
assign addr[40397]= -53538253;
assign addr[40398]= -91761426;
assign addr[40399]= -129955495;
assign addr[40400]= -168108346;
assign addr[40401]= -206207878;
assign addr[40402]= -244242007;
assign addr[40403]= -282198671;
assign addr[40404]= -320065829;
assign addr[40405]= -357831473;
assign addr[40406]= -395483624;
assign addr[40407]= -433010339;
assign addr[40408]= -470399716;
assign addr[40409]= -507639898;
assign addr[40410]= -544719071;
assign addr[40411]= -581625477;
assign addr[40412]= -618347408;
assign addr[40413]= -654873219;
assign addr[40414]= -691191324;
assign addr[40415]= -727290205;
assign addr[40416]= -763158411;
assign addr[40417]= -798784567;
assign addr[40418]= -834157373;
assign addr[40419]= -869265610;
assign addr[40420]= -904098143;
assign addr[40421]= -938643924;
assign addr[40422]= -972891995;
assign addr[40423]= -1006831495;
assign addr[40424]= -1040451659;
assign addr[40425]= -1073741824;
assign addr[40426]= -1106691431;
assign addr[40427]= -1139290029;
assign addr[40428]= -1171527280;
assign addr[40429]= -1203392958;
assign addr[40430]= -1234876957;
assign addr[40431]= -1265969291;
assign addr[40432]= -1296660098;
assign addr[40433]= -1326939644;
assign addr[40434]= -1356798326;
assign addr[40435]= -1386226674;
assign addr[40436]= -1415215352;
assign addr[40437]= -1443755168;
assign addr[40438]= -1471837070;
assign addr[40439]= -1499452149;
assign addr[40440]= -1526591649;
assign addr[40441]= -1553246960;
assign addr[40442]= -1579409630;
assign addr[40443]= -1605071359;
assign addr[40444]= -1630224009;
assign addr[40445]= -1654859602;
assign addr[40446]= -1678970324;
assign addr[40447]= -1702548529;
assign addr[40448]= -1725586737;
assign addr[40449]= -1748077642;
assign addr[40450]= -1770014111;
assign addr[40451]= -1791389186;
assign addr[40452]= -1812196087;
assign addr[40453]= -1832428215;
assign addr[40454]= -1852079154;
assign addr[40455]= -1871142669;
assign addr[40456]= -1889612716;
assign addr[40457]= -1907483436;
assign addr[40458]= -1924749160;
assign addr[40459]= -1941404413;
assign addr[40460]= -1957443913;
assign addr[40461]= -1972862571;
assign addr[40462]= -1987655498;
assign addr[40463]= -2001818002;
assign addr[40464]= -2015345591;
assign addr[40465]= -2028233973;
assign addr[40466]= -2040479063;
assign addr[40467]= -2052076975;
assign addr[40468]= -2063024031;
assign addr[40469]= -2073316760;
assign addr[40470]= -2082951896;
assign addr[40471]= -2091926384;
assign addr[40472]= -2100237377;
assign addr[40473]= -2107882239;
assign addr[40474]= -2114858546;
assign addr[40475]= -2121164085;
assign addr[40476]= -2126796855;
assign addr[40477]= -2131755071;
assign addr[40478]= -2136037160;
assign addr[40479]= -2139641764;
assign addr[40480]= -2142567738;
assign addr[40481]= -2144814157;
assign addr[40482]= -2146380306;
assign addr[40483]= -2147265689;
assign addr[40484]= -2147470025;
assign addr[40485]= -2146993250;
assign addr[40486]= -2145835515;
assign addr[40487]= -2143997187;
assign addr[40488]= -2141478848;
assign addr[40489]= -2138281298;
assign addr[40490]= -2134405552;
assign addr[40491]= -2129852837;
assign addr[40492]= -2124624598;
assign addr[40493]= -2118722494;
assign addr[40494]= -2112148396;
assign addr[40495]= -2104904390;
assign addr[40496]= -2096992772;
assign addr[40497]= -2088416053;
assign addr[40498]= -2079176953;
assign addr[40499]= -2069278401;
assign addr[40500]= -2058723538;
assign addr[40501]= -2047515711;
assign addr[40502]= -2035658475;
assign addr[40503]= -2023155591;
assign addr[40504]= -2010011024;
assign addr[40505]= -1996228943;
assign addr[40506]= -1981813720;
assign addr[40507]= -1966769926;
assign addr[40508]= -1951102334;
assign addr[40509]= -1934815911;
assign addr[40510]= -1917915825;
assign addr[40511]= -1900407434;
assign addr[40512]= -1882296293;
assign addr[40513]= -1863588145;
assign addr[40514]= -1844288924;
assign addr[40515]= -1824404752;
assign addr[40516]= -1803941934;
assign addr[40517]= -1782906961;
assign addr[40518]= -1761306505;
assign addr[40519]= -1739147417;
assign addr[40520]= -1716436725;
assign addr[40521]= -1693181631;
assign addr[40522]= -1669389513;
assign addr[40523]= -1645067915;
assign addr[40524]= -1620224553;
assign addr[40525]= -1594867305;
assign addr[40526]= -1569004214;
assign addr[40527]= -1542643483;
assign addr[40528]= -1515793473;
assign addr[40529]= -1488462700;
assign addr[40530]= -1460659832;
assign addr[40531]= -1432393688;
assign addr[40532]= -1403673233;
assign addr[40533]= -1374507575;
assign addr[40534]= -1344905966;
assign addr[40535]= -1314877795;
assign addr[40536]= -1284432584;
assign addr[40537]= -1253579991;
assign addr[40538]= -1222329801;
assign addr[40539]= -1190691925;
assign addr[40540]= -1158676398;
assign addr[40541]= -1126293375;
assign addr[40542]= -1093553126;
assign addr[40543]= -1060466036;
assign addr[40544]= -1027042599;
assign addr[40545]= -993293415;
assign addr[40546]= -959229189;
assign addr[40547]= -924860725;
assign addr[40548]= -890198924;
assign addr[40549]= -855254778;
assign addr[40550]= -820039373;
assign addr[40551]= -784563876;
assign addr[40552]= -748839539;
assign addr[40553]= -712877694;
assign addr[40554]= -676689746;
assign addr[40555]= -640287172;
assign addr[40556]= -603681519;
assign addr[40557]= -566884397;
assign addr[40558]= -529907477;
assign addr[40559]= -492762486;
assign addr[40560]= -455461206;
assign addr[40561]= -418015468;
assign addr[40562]= -380437148;
assign addr[40563]= -342738165;
assign addr[40564]= -304930476;
assign addr[40565]= -267026072;
assign addr[40566]= -229036977;
assign addr[40567]= -190975237;
assign addr[40568]= -152852926;
assign addr[40569]= -114682135;
assign addr[40570]= -76474970;
assign addr[40571]= -38243550;
assign addr[40572]= 0;
assign addr[40573]= 38243550;
assign addr[40574]= 76474970;
assign addr[40575]= 114682135;
assign addr[40576]= 152852926;
assign addr[40577]= 190975237;
assign addr[40578]= 229036977;
assign addr[40579]= 267026072;
assign addr[40580]= 304930476;
assign addr[40581]= 342738165;
assign addr[40582]= 380437148;
assign addr[40583]= 418015468;
assign addr[40584]= 455461206;
assign addr[40585]= 492762486;
assign addr[40586]= 529907477;
assign addr[40587]= 566884397;
assign addr[40588]= 603681519;
assign addr[40589]= 640287172;
assign addr[40590]= 676689746;
assign addr[40591]= 712877694;
assign addr[40592]= 748839539;
assign addr[40593]= 784563876;
assign addr[40594]= 820039373;
assign addr[40595]= 855254778;
assign addr[40596]= 890198924;
assign addr[40597]= 924860725;
assign addr[40598]= 959229189;
assign addr[40599]= 993293415;
assign addr[40600]= 1027042599;
assign addr[40601]= 1060466036;
assign addr[40602]= 1093553126;
assign addr[40603]= 1126293375;
assign addr[40604]= 1158676398;
assign addr[40605]= 1190691925;
assign addr[40606]= 1222329801;
assign addr[40607]= 1253579991;
assign addr[40608]= 1284432584;
assign addr[40609]= 1314877795;
assign addr[40610]= 1344905966;
assign addr[40611]= 1374507575;
assign addr[40612]= 1403673233;
assign addr[40613]= 1432393688;
assign addr[40614]= 1460659832;
assign addr[40615]= 1488462700;
assign addr[40616]= 1515793473;
assign addr[40617]= 1542643483;
assign addr[40618]= 1569004214;
assign addr[40619]= 1594867305;
assign addr[40620]= 1620224553;
assign addr[40621]= 1645067915;
assign addr[40622]= 1669389513;
assign addr[40623]= 1693181631;
assign addr[40624]= 1716436725;
assign addr[40625]= 1739147417;
assign addr[40626]= 1761306505;
assign addr[40627]= 1782906961;
assign addr[40628]= 1803941934;
assign addr[40629]= 1824404752;
assign addr[40630]= 1844288924;
assign addr[40631]= 1863588145;
assign addr[40632]= 1882296293;
assign addr[40633]= 1900407434;
assign addr[40634]= 1917915825;
assign addr[40635]= 1934815911;
assign addr[40636]= 1951102334;
assign addr[40637]= 1966769926;
assign addr[40638]= 1981813720;
assign addr[40639]= 1996228943;
assign addr[40640]= 2010011024;
assign addr[40641]= 2023155591;
assign addr[40642]= 2035658475;
assign addr[40643]= 2047515711;
assign addr[40644]= 2058723538;
assign addr[40645]= 2069278401;
assign addr[40646]= 2079176953;
assign addr[40647]= 2088416053;
assign addr[40648]= 2096992772;
assign addr[40649]= 2104904390;
assign addr[40650]= 2112148396;
assign addr[40651]= 2118722494;
assign addr[40652]= 2124624598;
assign addr[40653]= 2129852837;
assign addr[40654]= 2134405552;
assign addr[40655]= 2138281298;
assign addr[40656]= 2141478848;
assign addr[40657]= 2143997187;
assign addr[40658]= 2145835515;
assign addr[40659]= 2146993250;
assign addr[40660]= 2147470025;
assign addr[40661]= 2147265689;
assign addr[40662]= 2146380306;
assign addr[40663]= 2144814157;
assign addr[40664]= 2142567738;
assign addr[40665]= 2139641764;
assign addr[40666]= 2136037160;
assign addr[40667]= 2131755071;
assign addr[40668]= 2126796855;
assign addr[40669]= 2121164085;
assign addr[40670]= 2114858546;
assign addr[40671]= 2107882239;
assign addr[40672]= 2100237377;
assign addr[40673]= 2091926384;
assign addr[40674]= 2082951896;
assign addr[40675]= 2073316760;
assign addr[40676]= 2063024031;
assign addr[40677]= 2052076975;
assign addr[40678]= 2040479063;
assign addr[40679]= 2028233973;
assign addr[40680]= 2015345591;
assign addr[40681]= 2001818002;
assign addr[40682]= 1987655498;
assign addr[40683]= 1972862571;
assign addr[40684]= 1957443913;
assign addr[40685]= 1941404413;
assign addr[40686]= 1924749160;
assign addr[40687]= 1907483436;
assign addr[40688]= 1889612716;
assign addr[40689]= 1871142669;
assign addr[40690]= 1852079154;
assign addr[40691]= 1832428215;
assign addr[40692]= 1812196087;
assign addr[40693]= 1791389186;
assign addr[40694]= 1770014111;
assign addr[40695]= 1748077642;
assign addr[40696]= 1725586737;
assign addr[40697]= 1702548529;
assign addr[40698]= 1678970324;
assign addr[40699]= 1654859602;
assign addr[40700]= 1630224009;
assign addr[40701]= 1605071359;
assign addr[40702]= 1579409630;
assign addr[40703]= 1553246960;
assign addr[40704]= 1526591649;
assign addr[40705]= 1499452149;
assign addr[40706]= 1471837070;
assign addr[40707]= 1443755168;
assign addr[40708]= 1415215352;
assign addr[40709]= 1386226674;
assign addr[40710]= 1356798326;
assign addr[40711]= 1326939644;
assign addr[40712]= 1296660098;
assign addr[40713]= 1265969291;
assign addr[40714]= 1234876957;
assign addr[40715]= 1203392958;
assign addr[40716]= 1171527280;
assign addr[40717]= 1139290029;
assign addr[40718]= 1106691431;
assign addr[40719]= 1073741824;
assign addr[40720]= 1040451659;
assign addr[40721]= 1006831495;
assign addr[40722]= 972891995;
assign addr[40723]= 938643924;
assign addr[40724]= 904098143;
assign addr[40725]= 869265610;
assign addr[40726]= 834157373;
assign addr[40727]= 798784567;
assign addr[40728]= 763158411;
assign addr[40729]= 727290205;
assign addr[40730]= 691191324;
assign addr[40731]= 654873219;
assign addr[40732]= 618347408;
assign addr[40733]= 581625477;
assign addr[40734]= 544719071;
assign addr[40735]= 507639898;
assign addr[40736]= 470399716;
assign addr[40737]= 433010339;
assign addr[40738]= 395483624;
assign addr[40739]= 357831473;
assign addr[40740]= 320065829;
assign addr[40741]= 282198671;
assign addr[40742]= 244242007;
assign addr[40743]= 206207878;
assign addr[40744]= 168108346;
assign addr[40745]= 129955495;
assign addr[40746]= 91761426;
assign addr[40747]= 53538253;
assign addr[40748]= 15298099;
assign addr[40749]= -22946906;
assign addr[40750]= -61184634;
assign addr[40751]= -99402956;
assign addr[40752]= -137589750;
assign addr[40753]= -175732905;
assign addr[40754]= -213820322;
assign addr[40755]= -251839923;
assign addr[40756]= -289779648;
assign addr[40757]= -327627463;
assign addr[40758]= -365371365;
assign addr[40759]= -402999383;
assign addr[40760]= -440499581;
assign addr[40761]= -477860067;
assign addr[40762]= -515068990;
assign addr[40763]= -552114549;
assign addr[40764]= -588984994;
assign addr[40765]= -625668632;
assign addr[40766]= -662153826;
assign addr[40767]= -698429006;
assign addr[40768]= -734482665;
assign addr[40769]= -770303369;
assign addr[40770]= -805879757;
assign addr[40771]= -841200544;
assign addr[40772]= -876254528;
assign addr[40773]= -911030591;
assign addr[40774]= -945517704;
assign addr[40775]= -979704927;
assign addr[40776]= -1013581418;
assign addr[40777]= -1047136432;
assign addr[40778]= -1080359326;
assign addr[40779]= -1113239564;
assign addr[40780]= -1145766716;
assign addr[40781]= -1177930466;
assign addr[40782]= -1209720613;
assign addr[40783]= -1241127074;
assign addr[40784]= -1272139887;
assign addr[40785]= -1302749217;
assign addr[40786]= -1332945355;
assign addr[40787]= -1362718723;
assign addr[40788]= -1392059879;
assign addr[40789]= -1420959516;
assign addr[40790]= -1449408469;
assign addr[40791]= -1477397714;
assign addr[40792]= -1504918373;
assign addr[40793]= -1531961719;
assign addr[40794]= -1558519173;
assign addr[40795]= -1584582314;
assign addr[40796]= -1610142873;
assign addr[40797]= -1635192744;
assign addr[40798]= -1659723983;
assign addr[40799]= -1683728808;
assign addr[40800]= -1707199606;
assign addr[40801]= -1730128933;
assign addr[40802]= -1752509516;
assign addr[40803]= -1774334257;
assign addr[40804]= -1795596234;
assign addr[40805]= -1816288703;
assign addr[40806]= -1836405100;
assign addr[40807]= -1855939047;
assign addr[40808]= -1874884346;
assign addr[40809]= -1893234990;
assign addr[40810]= -1910985158;
assign addr[40811]= -1928129220;
assign addr[40812]= -1944661739;
assign addr[40813]= -1960577471;
assign addr[40814]= -1975871368;
assign addr[40815]= -1990538579;
assign addr[40816]= -2004574453;
assign addr[40817]= -2017974537;
assign addr[40818]= -2030734582;
assign addr[40819]= -2042850540;
assign addr[40820]= -2054318569;
assign addr[40821]= -2065135031;
assign addr[40822]= -2075296495;
assign addr[40823]= -2084799740;
assign addr[40824]= -2093641749;
assign addr[40825]= -2101819720;
assign addr[40826]= -2109331059;
assign addr[40827]= -2116173382;
assign addr[40828]= -2122344521;
assign addr[40829]= -2127842516;
assign addr[40830]= -2132665626;
assign addr[40831]= -2136812319;
assign addr[40832]= -2140281282;
assign addr[40833]= -2143071413;
assign addr[40834]= -2145181827;
assign addr[40835]= -2146611856;
assign addr[40836]= -2147361045;
assign addr[40837]= -2147429158;
assign addr[40838]= -2146816171;
assign addr[40839]= -2145522281;
assign addr[40840]= -2143547897;
assign addr[40841]= -2140893646;
assign addr[40842]= -2137560369;
assign addr[40843]= -2133549123;
assign addr[40844]= -2128861181;
assign addr[40845]= -2123498030;
assign addr[40846]= -2117461370;
assign addr[40847]= -2110753117;
assign addr[40848]= -2103375398;
assign addr[40849]= -2095330553;
assign addr[40850]= -2086621133;
assign addr[40851]= -2077249901;
assign addr[40852]= -2067219829;
assign addr[40853]= -2056534099;
assign addr[40854]= -2045196100;
assign addr[40855]= -2033209426;
assign addr[40856]= -2020577882;
assign addr[40857]= -2007305472;
assign addr[40858]= -1993396407;
assign addr[40859]= -1978855097;
assign addr[40860]= -1963686155;
assign addr[40861]= -1947894393;
assign addr[40862]= -1931484818;
assign addr[40863]= -1914462636;
assign addr[40864]= -1896833245;
assign addr[40865]= -1878602237;
assign addr[40866]= -1859775393;
assign addr[40867]= -1840358687;
assign addr[40868]= -1820358275;
assign addr[40869]= -1799780501;
assign addr[40870]= -1778631892;
assign addr[40871]= -1756919156;
assign addr[40872]= -1734649179;
assign addr[40873]= -1711829025;
assign addr[40874]= -1688465931;
assign addr[40875]= -1664567307;
assign addr[40876]= -1640140734;
assign addr[40877]= -1615193959;
assign addr[40878]= -1589734894;
assign addr[40879]= -1563771613;
assign addr[40880]= -1537312353;
assign addr[40881]= -1510365504;
assign addr[40882]= -1482939614;
assign addr[40883]= -1455043381;
assign addr[40884]= -1426685652;
assign addr[40885]= -1397875423;
assign addr[40886]= -1368621831;
assign addr[40887]= -1338934154;
assign addr[40888]= -1308821808;
assign addr[40889]= -1278294345;
assign addr[40890]= -1247361445;
assign addr[40891]= -1216032921;
assign addr[40892]= -1184318708;
assign addr[40893]= -1152228866;
assign addr[40894]= -1119773573;
assign addr[40895]= -1086963121;
assign addr[40896]= -1053807919;
assign addr[40897]= -1020318481;
assign addr[40898]= -986505429;
assign addr[40899]= -952379488;
assign addr[40900]= -917951481;
assign addr[40901]= -883232329;
assign addr[40902]= -848233042;
assign addr[40903]= -812964722;
assign addr[40904]= -777438554;
assign addr[40905]= -741665807;
assign addr[40906]= -705657826;
assign addr[40907]= -669426032;
assign addr[40908]= -632981917;
assign addr[40909]= -596337040;
assign addr[40910]= -559503022;
assign addr[40911]= -522491548;
assign addr[40912]= -485314355;
assign addr[40913]= -447983235;
assign addr[40914]= -410510029;
assign addr[40915]= -372906622;
assign addr[40916]= -335184940;
assign addr[40917]= -297356948;
assign addr[40918]= -259434643;
assign addr[40919]= -221430054;
assign addr[40920]= -183355234;
assign addr[40921]= -145222259;
assign addr[40922]= -107043224;
assign addr[40923]= -68830239;
assign addr[40924]= -30595422;
assign addr[40925]= 7649098;
assign addr[40926]= 45891193;
assign addr[40927]= 84118732;
assign addr[40928]= 122319591;
assign addr[40929]= 160481654;
assign addr[40930]= 198592817;
assign addr[40931]= 236640993;
assign addr[40932]= 274614114;
assign addr[40933]= 312500135;
assign addr[40934]= 350287041;
assign addr[40935]= 387962847;
assign addr[40936]= 425515602;
assign addr[40937]= 462933398;
assign addr[40938]= 500204365;
assign addr[40939]= 537316682;
assign addr[40940]= 574258580;
assign addr[40941]= 611018340;
assign addr[40942]= 647584304;
assign addr[40943]= 683944874;
assign addr[40944]= 720088517;
assign addr[40945]= 756003771;
assign addr[40946]= 791679244;
assign addr[40947]= 827103620;
assign addr[40948]= 862265664;
assign addr[40949]= 897154224;
assign addr[40950]= 931758235;
assign addr[40951]= 966066720;
assign addr[40952]= 1000068799;
assign addr[40953]= 1033753687;
assign addr[40954]= 1067110699;
assign addr[40955]= 1100129257;
assign addr[40956]= 1132798888;
assign addr[40957]= 1165109230;
assign addr[40958]= 1197050035;
assign addr[40959]= 1228611172;
assign addr[40960]= 1259782632;
assign addr[40961]= 1290554528;
assign addr[40962]= 1320917099;
assign addr[40963]= 1350860716;
assign addr[40964]= 1380375881;
assign addr[40965]= 1409453233;
assign addr[40966]= 1438083551;
assign addr[40967]= 1466257752;
assign addr[40968]= 1493966902;
assign addr[40969]= 1521202211;
assign addr[40970]= 1547955041;
assign addr[40971]= 1574216908;
assign addr[40972]= 1599979481;
assign addr[40973]= 1625234591;
assign addr[40974]= 1649974225;
assign addr[40975]= 1674190539;
assign addr[40976]= 1697875851;
assign addr[40977]= 1721022648;
assign addr[40978]= 1743623590;
assign addr[40979]= 1765671509;
assign addr[40980]= 1787159411;
assign addr[40981]= 1808080480;
assign addr[40982]= 1828428082;
assign addr[40983]= 1848195763;
assign addr[40984]= 1867377253;
assign addr[40985]= 1885966468;
assign addr[40986]= 1903957513;
assign addr[40987]= 1921344681;
assign addr[40988]= 1938122457;
assign addr[40989]= 1954285520;
assign addr[40990]= 1969828744;
assign addr[40991]= 1984747199;
assign addr[40992]= 1999036154;
assign addr[40993]= 2012691075;
assign addr[40994]= 2025707632;
assign addr[40995]= 2038081698;
assign addr[40996]= 2049809346;
assign addr[40997]= 2060886858;
assign addr[40998]= 2071310720;
assign addr[40999]= 2081077626;
assign addr[41000]= 2090184478;
assign addr[41001]= 2098628387;
assign addr[41002]= 2106406677;
assign addr[41003]= 2113516878;
assign addr[41004]= 2119956737;
assign addr[41005]= 2125724211;
assign addr[41006]= 2130817471;
assign addr[41007]= 2135234901;
assign addr[41008]= 2138975100;
assign addr[41009]= 2142036881;
assign addr[41010]= 2144419275;
assign addr[41011]= 2146121524;
assign addr[41012]= 2147143090;
assign addr[41013]= 2147483648;
assign addr[41014]= 2147143090;
assign addr[41015]= 2146121524;
assign addr[41016]= 2144419275;
assign addr[41017]= 2142036881;
assign addr[41018]= 2138975100;
assign addr[41019]= 2135234901;
assign addr[41020]= 2130817471;
assign addr[41021]= 2125724211;
assign addr[41022]= 2119956737;
assign addr[41023]= 2113516878;
assign addr[41024]= 2106406677;
assign addr[41025]= 2098628387;
assign addr[41026]= 2090184478;
assign addr[41027]= 2081077626;
assign addr[41028]= 2071310720;
assign addr[41029]= 2060886858;
assign addr[41030]= 2049809346;
assign addr[41031]= 2038081698;
assign addr[41032]= 2025707632;
assign addr[41033]= 2012691075;
assign addr[41034]= 1999036154;
assign addr[41035]= 1984747199;
assign addr[41036]= 1969828744;
assign addr[41037]= 1954285520;
assign addr[41038]= 1938122457;
assign addr[41039]= 1921344681;
assign addr[41040]= 1903957513;
assign addr[41041]= 1885966468;
assign addr[41042]= 1867377253;
assign addr[41043]= 1848195763;
assign addr[41044]= 1828428082;
assign addr[41045]= 1808080480;
assign addr[41046]= 1787159411;
assign addr[41047]= 1765671509;
assign addr[41048]= 1743623590;
assign addr[41049]= 1721022648;
assign addr[41050]= 1697875851;
assign addr[41051]= 1674190539;
assign addr[41052]= 1649974225;
assign addr[41053]= 1625234591;
assign addr[41054]= 1599979481;
assign addr[41055]= 1574216908;
assign addr[41056]= 1547955041;
assign addr[41057]= 1521202211;
assign addr[41058]= 1493966902;
assign addr[41059]= 1466257752;
assign addr[41060]= 1438083551;
assign addr[41061]= 1409453233;
assign addr[41062]= 1380375881;
assign addr[41063]= 1350860716;
assign addr[41064]= 1320917099;
assign addr[41065]= 1290554528;
assign addr[41066]= 1259782632;
assign addr[41067]= 1228611172;
assign addr[41068]= 1197050035;
assign addr[41069]= 1165109230;
assign addr[41070]= 1132798888;
assign addr[41071]= 1100129257;
assign addr[41072]= 1067110699;
assign addr[41073]= 1033753687;
assign addr[41074]= 1000068799;
assign addr[41075]= 966066720;
assign addr[41076]= 931758235;
assign addr[41077]= 897154224;
assign addr[41078]= 862265664;
assign addr[41079]= 827103620;
assign addr[41080]= 791679244;
assign addr[41081]= 756003771;
assign addr[41082]= 720088517;
assign addr[41083]= 683944874;
assign addr[41084]= 647584304;
assign addr[41085]= 611018340;
assign addr[41086]= 574258580;
assign addr[41087]= 537316682;
assign addr[41088]= 500204365;
assign addr[41089]= 462933398;
assign addr[41090]= 425515602;
assign addr[41091]= 387962847;
assign addr[41092]= 350287041;
assign addr[41093]= 312500135;
assign addr[41094]= 274614114;
assign addr[41095]= 236640993;
assign addr[41096]= 198592817;
assign addr[41097]= 160481654;
assign addr[41098]= 122319591;
assign addr[41099]= 84118732;
assign addr[41100]= 45891193;
assign addr[41101]= 7649098;
assign addr[41102]= -30595422;
assign addr[41103]= -68830239;
assign addr[41104]= -107043224;
assign addr[41105]= -145222259;
assign addr[41106]= -183355234;
assign addr[41107]= -221430054;
assign addr[41108]= -259434643;
assign addr[41109]= -297356948;
assign addr[41110]= -335184940;
assign addr[41111]= -372906622;
assign addr[41112]= -410510029;
assign addr[41113]= -447983235;
assign addr[41114]= -485314355;
assign addr[41115]= -522491548;
assign addr[41116]= -559503022;
assign addr[41117]= -596337040;
assign addr[41118]= -632981917;
assign addr[41119]= -669426032;
assign addr[41120]= -705657826;
assign addr[41121]= -741665807;
assign addr[41122]= -777438554;
assign addr[41123]= -812964722;
assign addr[41124]= -848233042;
assign addr[41125]= -883232329;
assign addr[41126]= -917951481;
assign addr[41127]= -952379488;
assign addr[41128]= -986505429;
assign addr[41129]= -1020318481;
assign addr[41130]= -1053807919;
assign addr[41131]= -1086963121;
assign addr[41132]= -1119773573;
assign addr[41133]= -1152228866;
assign addr[41134]= -1184318708;
assign addr[41135]= -1216032921;
assign addr[41136]= -1247361445;
assign addr[41137]= -1278294345;
assign addr[41138]= -1308821808;
assign addr[41139]= -1338934154;
assign addr[41140]= -1368621831;
assign addr[41141]= -1397875423;
assign addr[41142]= -1426685652;
assign addr[41143]= -1455043381;
assign addr[41144]= -1482939614;
assign addr[41145]= -1510365504;
assign addr[41146]= -1537312353;
assign addr[41147]= -1563771613;
assign addr[41148]= -1589734894;
assign addr[41149]= -1615193959;
assign addr[41150]= -1640140734;
assign addr[41151]= -1664567307;
assign addr[41152]= -1688465931;
assign addr[41153]= -1711829025;
assign addr[41154]= -1734649179;
assign addr[41155]= -1756919156;
assign addr[41156]= -1778631892;
assign addr[41157]= -1799780501;
assign addr[41158]= -1820358275;
assign addr[41159]= -1840358687;
assign addr[41160]= -1859775393;
assign addr[41161]= -1878602237;
assign addr[41162]= -1896833245;
assign addr[41163]= -1914462636;
assign addr[41164]= -1931484818;
assign addr[41165]= -1947894393;
assign addr[41166]= -1963686155;
assign addr[41167]= -1978855097;
assign addr[41168]= -1993396407;
assign addr[41169]= -2007305472;
assign addr[41170]= -2020577882;
assign addr[41171]= -2033209426;
assign addr[41172]= -2045196100;
assign addr[41173]= -2056534099;
assign addr[41174]= -2067219829;
assign addr[41175]= -2077249901;
assign addr[41176]= -2086621133;
assign addr[41177]= -2095330553;
assign addr[41178]= -2103375398;
assign addr[41179]= -2110753117;
assign addr[41180]= -2117461370;
assign addr[41181]= -2123498030;
assign addr[41182]= -2128861181;
assign addr[41183]= -2133549123;
assign addr[41184]= -2137560369;
assign addr[41185]= -2140893646;
assign addr[41186]= -2143547897;
assign addr[41187]= -2145522281;
assign addr[41188]= -2146816171;
assign addr[41189]= -2147429158;
assign addr[41190]= -2147361045;
assign addr[41191]= -2146611856;
assign addr[41192]= -2145181827;
assign addr[41193]= -2143071413;
assign addr[41194]= -2140281282;
assign addr[41195]= -2136812319;
assign addr[41196]= -2132665626;
assign addr[41197]= -2127842516;
assign addr[41198]= -2122344521;
assign addr[41199]= -2116173382;
assign addr[41200]= -2109331059;
assign addr[41201]= -2101819720;
assign addr[41202]= -2093641749;
assign addr[41203]= -2084799740;
assign addr[41204]= -2075296495;
assign addr[41205]= -2065135031;
assign addr[41206]= -2054318569;
assign addr[41207]= -2042850540;
assign addr[41208]= -2030734582;
assign addr[41209]= -2017974537;
assign addr[41210]= -2004574453;
assign addr[41211]= -1990538579;
assign addr[41212]= -1975871368;
assign addr[41213]= -1960577471;
assign addr[41214]= -1944661739;
assign addr[41215]= -1928129220;
assign addr[41216]= -1910985158;
assign addr[41217]= -1893234990;
assign addr[41218]= -1874884346;
assign addr[41219]= -1855939047;
assign addr[41220]= -1836405100;
assign addr[41221]= -1816288703;
assign addr[41222]= -1795596234;
assign addr[41223]= -1774334257;
assign addr[41224]= -1752509516;
assign addr[41225]= -1730128933;
assign addr[41226]= -1707199606;
assign addr[41227]= -1683728808;
assign addr[41228]= -1659723983;
assign addr[41229]= -1635192744;
assign addr[41230]= -1610142873;
assign addr[41231]= -1584582314;
assign addr[41232]= -1558519173;
assign addr[41233]= -1531961719;
assign addr[41234]= -1504918373;
assign addr[41235]= -1477397714;
assign addr[41236]= -1449408469;
assign addr[41237]= -1420959516;
assign addr[41238]= -1392059879;
assign addr[41239]= -1362718723;
assign addr[41240]= -1332945355;
assign addr[41241]= -1302749217;
assign addr[41242]= -1272139887;
assign addr[41243]= -1241127074;
assign addr[41244]= -1209720613;
assign addr[41245]= -1177930466;
assign addr[41246]= -1145766716;
assign addr[41247]= -1113239564;
assign addr[41248]= -1080359326;
assign addr[41249]= -1047136432;
assign addr[41250]= -1013581418;
assign addr[41251]= -979704927;
assign addr[41252]= -945517704;
assign addr[41253]= -911030591;
assign addr[41254]= -876254528;
assign addr[41255]= -841200544;
assign addr[41256]= -805879757;
assign addr[41257]= -770303369;
assign addr[41258]= -734482665;
assign addr[41259]= -698429006;
assign addr[41260]= -662153826;
assign addr[41261]= -625668632;
assign addr[41262]= -588984994;
assign addr[41263]= -552114549;
assign addr[41264]= -515068990;
assign addr[41265]= -477860067;
assign addr[41266]= -440499581;
assign addr[41267]= -402999383;
assign addr[41268]= -365371365;
assign addr[41269]= -327627463;
assign addr[41270]= -289779648;
assign addr[41271]= -251839923;
assign addr[41272]= -213820322;
assign addr[41273]= -175732905;
assign addr[41274]= -137589750;
assign addr[41275]= -99402956;
assign addr[41276]= -61184634;
assign addr[41277]= -22946906;
assign addr[41278]= 15298099;
assign addr[41279]= 53538253;
assign addr[41280]= 91761426;
assign addr[41281]= 129955495;
assign addr[41282]= 168108346;
assign addr[41283]= 206207878;
assign addr[41284]= 244242007;
assign addr[41285]= 282198671;
assign addr[41286]= 320065829;
assign addr[41287]= 357831473;
assign addr[41288]= 395483624;
assign addr[41289]= 433010339;
assign addr[41290]= 470399716;
assign addr[41291]= 507639898;
assign addr[41292]= 544719071;
assign addr[41293]= 581625477;
assign addr[41294]= 618347408;
assign addr[41295]= 654873219;
assign addr[41296]= 691191324;
assign addr[41297]= 727290205;
assign addr[41298]= 763158411;
assign addr[41299]= 798784567;
assign addr[41300]= 834157373;
assign addr[41301]= 869265610;
assign addr[41302]= 904098143;
assign addr[41303]= 938643924;
assign addr[41304]= 972891995;
assign addr[41305]= 1006831495;
assign addr[41306]= 1040451659;
assign addr[41307]= 1073741824;
assign addr[41308]= 1106691431;
assign addr[41309]= 1139290029;
assign addr[41310]= 1171527280;
assign addr[41311]= 1203392958;
assign addr[41312]= 1234876957;
assign addr[41313]= 1265969291;
assign addr[41314]= 1296660098;
assign addr[41315]= 1326939644;
assign addr[41316]= 1356798326;
assign addr[41317]= 1386226674;
assign addr[41318]= 1415215352;
assign addr[41319]= 1443755168;
assign addr[41320]= 1471837070;
assign addr[41321]= 1499452149;
assign addr[41322]= 1526591649;
assign addr[41323]= 1553246960;
assign addr[41324]= 1579409630;
assign addr[41325]= 1605071359;
assign addr[41326]= 1630224009;
assign addr[41327]= 1654859602;
assign addr[41328]= 1678970324;
assign addr[41329]= 1702548529;
assign addr[41330]= 1725586737;
assign addr[41331]= 1748077642;
assign addr[41332]= 1770014111;
assign addr[41333]= 1791389186;
assign addr[41334]= 1812196087;
assign addr[41335]= 1832428215;
assign addr[41336]= 1852079154;
assign addr[41337]= 1871142669;
assign addr[41338]= 1889612716;
assign addr[41339]= 1907483436;
assign addr[41340]= 1924749160;
assign addr[41341]= 1941404413;
assign addr[41342]= 1957443913;
assign addr[41343]= 1972862571;
assign addr[41344]= 1987655498;
assign addr[41345]= 2001818002;
assign addr[41346]= 2015345591;
assign addr[41347]= 2028233973;
assign addr[41348]= 2040479063;
assign addr[41349]= 2052076975;
assign addr[41350]= 2063024031;
assign addr[41351]= 2073316760;
assign addr[41352]= 2082951896;
assign addr[41353]= 2091926384;
assign addr[41354]= 2100237377;
assign addr[41355]= 2107882239;
assign addr[41356]= 2114858546;
assign addr[41357]= 2121164085;
assign addr[41358]= 2126796855;
assign addr[41359]= 2131755071;
assign addr[41360]= 2136037160;
assign addr[41361]= 2139641764;
assign addr[41362]= 2142567738;
assign addr[41363]= 2144814157;
assign addr[41364]= 2146380306;
assign addr[41365]= 2147265689;
assign addr[41366]= 2147470025;
assign addr[41367]= 2146993250;
assign addr[41368]= 2145835515;
assign addr[41369]= 2143997187;
assign addr[41370]= 2141478848;
assign addr[41371]= 2138281298;
assign addr[41372]= 2134405552;
assign addr[41373]= 2129852837;
assign addr[41374]= 2124624598;
assign addr[41375]= 2118722494;
assign addr[41376]= 2112148396;
assign addr[41377]= 2104904390;
assign addr[41378]= 2096992772;
assign addr[41379]= 2088416053;
assign addr[41380]= 2079176953;
assign addr[41381]= 2069278401;
assign addr[41382]= 2058723538;
assign addr[41383]= 2047515711;
assign addr[41384]= 2035658475;
assign addr[41385]= 2023155591;
assign addr[41386]= 2010011024;
assign addr[41387]= 1996228943;
assign addr[41388]= 1981813720;
assign addr[41389]= 1966769926;
assign addr[41390]= 1951102334;
assign addr[41391]= 1934815911;
assign addr[41392]= 1917915825;
assign addr[41393]= 1900407434;
assign addr[41394]= 1882296293;
assign addr[41395]= 1863588145;
assign addr[41396]= 1844288924;
assign addr[41397]= 1824404752;
assign addr[41398]= 1803941934;
assign addr[41399]= 1782906961;
assign addr[41400]= 1761306505;
assign addr[41401]= 1739147417;
assign addr[41402]= 1716436725;
assign addr[41403]= 1693181631;
assign addr[41404]= 1669389513;
assign addr[41405]= 1645067915;
assign addr[41406]= 1620224553;
assign addr[41407]= 1594867305;
assign addr[41408]= 1569004214;
assign addr[41409]= 1542643483;
assign addr[41410]= 1515793473;
assign addr[41411]= 1488462700;
assign addr[41412]= 1460659832;
assign addr[41413]= 1432393688;
assign addr[41414]= 1403673233;
assign addr[41415]= 1374507575;
assign addr[41416]= 1344905966;
assign addr[41417]= 1314877795;
assign addr[41418]= 1284432584;
assign addr[41419]= 1253579991;
assign addr[41420]= 1222329801;
assign addr[41421]= 1190691925;
assign addr[41422]= 1158676398;
assign addr[41423]= 1126293375;
assign addr[41424]= 1093553126;
assign addr[41425]= 1060466036;
assign addr[41426]= 1027042599;
assign addr[41427]= 993293415;
assign addr[41428]= 959229189;
assign addr[41429]= 924860725;
assign addr[41430]= 890198924;
assign addr[41431]= 855254778;
assign addr[41432]= 820039373;
assign addr[41433]= 784563876;
assign addr[41434]= 748839539;
assign addr[41435]= 712877694;
assign addr[41436]= 676689746;
assign addr[41437]= 640287172;
assign addr[41438]= 603681519;
assign addr[41439]= 566884397;
assign addr[41440]= 529907477;
assign addr[41441]= 492762486;
assign addr[41442]= 455461206;
assign addr[41443]= 418015468;
assign addr[41444]= 380437148;
assign addr[41445]= 342738165;
assign addr[41446]= 304930476;
assign addr[41447]= 267026072;
assign addr[41448]= 229036977;
assign addr[41449]= 190975237;
assign addr[41450]= 152852926;
assign addr[41451]= 114682135;
assign addr[41452]= 76474970;
assign addr[41453]= 38243550;
assign addr[41454]= 0;
assign addr[41455]= -38243550;
assign addr[41456]= -76474970;
assign addr[41457]= -114682135;
assign addr[41458]= -152852926;
assign addr[41459]= -190975237;
assign addr[41460]= -229036977;
assign addr[41461]= -267026072;
assign addr[41462]= -304930476;
assign addr[41463]= -342738165;
assign addr[41464]= -380437148;
assign addr[41465]= -418015468;
assign addr[41466]= -455461206;
assign addr[41467]= -492762486;
assign addr[41468]= -529907477;
assign addr[41469]= -566884397;
assign addr[41470]= -603681519;
assign addr[41471]= -640287172;
assign addr[41472]= -676689746;
assign addr[41473]= -712877694;
assign addr[41474]= -748839539;
assign addr[41475]= -784563876;
assign addr[41476]= -820039373;
assign addr[41477]= -855254778;
assign addr[41478]= -890198924;
assign addr[41479]= -924860725;
assign addr[41480]= -959229189;
assign addr[41481]= -993293415;
assign addr[41482]= -1027042599;
assign addr[41483]= -1060466036;
assign addr[41484]= -1093553126;
assign addr[41485]= -1126293375;
assign addr[41486]= -1158676398;
assign addr[41487]= -1190691925;
assign addr[41488]= -1222329801;
assign addr[41489]= -1253579991;
assign addr[41490]= -1284432584;
assign addr[41491]= -1314877795;
assign addr[41492]= -1344905966;
assign addr[41493]= -1374507575;
assign addr[41494]= -1403673233;
assign addr[41495]= -1432393688;
assign addr[41496]= -1460659832;
assign addr[41497]= -1488462700;
assign addr[41498]= -1515793473;
assign addr[41499]= -1542643483;
assign addr[41500]= -1569004214;
assign addr[41501]= -1594867305;
assign addr[41502]= -1620224553;
assign addr[41503]= -1645067915;
assign addr[41504]= -1669389513;
assign addr[41505]= -1693181631;
assign addr[41506]= -1716436725;
assign addr[41507]= -1739147417;
assign addr[41508]= -1761306505;
assign addr[41509]= -1782906961;
assign addr[41510]= -1803941934;
assign addr[41511]= -1824404752;
assign addr[41512]= -1844288924;
assign addr[41513]= -1863588145;
assign addr[41514]= -1882296293;
assign addr[41515]= -1900407434;
assign addr[41516]= -1917915825;
assign addr[41517]= -1934815911;
assign addr[41518]= -1951102334;
assign addr[41519]= -1966769926;
assign addr[41520]= -1981813720;
assign addr[41521]= -1996228943;
assign addr[41522]= -2010011024;
assign addr[41523]= -2023155591;
assign addr[41524]= -2035658475;
assign addr[41525]= -2047515711;
assign addr[41526]= -2058723538;
assign addr[41527]= -2069278401;
assign addr[41528]= -2079176953;
assign addr[41529]= -2088416053;
assign addr[41530]= -2096992772;
assign addr[41531]= -2104904390;
assign addr[41532]= -2112148396;
assign addr[41533]= -2118722494;
assign addr[41534]= -2124624598;
assign addr[41535]= -2129852837;
assign addr[41536]= -2134405552;
assign addr[41537]= -2138281298;
assign addr[41538]= -2141478848;
assign addr[41539]= -2143997187;
assign addr[41540]= -2145835515;
assign addr[41541]= -2146993250;
assign addr[41542]= -2147470025;
assign addr[41543]= -2147265689;
assign addr[41544]= -2146380306;
assign addr[41545]= -2144814157;
assign addr[41546]= -2142567738;
assign addr[41547]= -2139641764;
assign addr[41548]= -2136037160;
assign addr[41549]= -2131755071;
assign addr[41550]= -2126796855;
assign addr[41551]= -2121164085;
assign addr[41552]= -2114858546;
assign addr[41553]= -2107882239;
assign addr[41554]= -2100237377;
assign addr[41555]= -2091926384;
assign addr[41556]= -2082951896;
assign addr[41557]= -2073316760;
assign addr[41558]= -2063024031;
assign addr[41559]= -2052076975;
assign addr[41560]= -2040479063;
assign addr[41561]= -2028233973;
assign addr[41562]= -2015345591;
assign addr[41563]= -2001818002;
assign addr[41564]= -1987655498;
assign addr[41565]= -1972862571;
assign addr[41566]= -1957443913;
assign addr[41567]= -1941404413;
assign addr[41568]= -1924749160;
assign addr[41569]= -1907483436;
assign addr[41570]= -1889612716;
assign addr[41571]= -1871142669;
assign addr[41572]= -1852079154;
assign addr[41573]= -1832428215;
assign addr[41574]= -1812196087;
assign addr[41575]= -1791389186;
assign addr[41576]= -1770014111;
assign addr[41577]= -1748077642;
assign addr[41578]= -1725586737;
assign addr[41579]= -1702548529;
assign addr[41580]= -1678970324;
assign addr[41581]= -1654859602;
assign addr[41582]= -1630224009;
assign addr[41583]= -1605071359;
assign addr[41584]= -1579409630;
assign addr[41585]= -1553246960;
assign addr[41586]= -1526591649;
assign addr[41587]= -1499452149;
assign addr[41588]= -1471837070;
assign addr[41589]= -1443755168;
assign addr[41590]= -1415215352;
assign addr[41591]= -1386226674;
assign addr[41592]= -1356798326;
assign addr[41593]= -1326939644;
assign addr[41594]= -1296660098;
assign addr[41595]= -1265969291;
assign addr[41596]= -1234876957;
assign addr[41597]= -1203392958;
assign addr[41598]= -1171527280;
assign addr[41599]= -1139290029;
assign addr[41600]= -1106691431;
assign addr[41601]= -1073741824;
assign addr[41602]= -1040451659;
assign addr[41603]= -1006831495;
assign addr[41604]= -972891995;
assign addr[41605]= -938643924;
assign addr[41606]= -904098143;
assign addr[41607]= -869265610;
assign addr[41608]= -834157373;
assign addr[41609]= -798784567;
assign addr[41610]= -763158411;
assign addr[41611]= -727290205;
assign addr[41612]= -691191324;
assign addr[41613]= -654873219;
assign addr[41614]= -618347408;
assign addr[41615]= -581625477;
assign addr[41616]= -544719071;
assign addr[41617]= -507639898;
assign addr[41618]= -470399716;
assign addr[41619]= -433010339;
assign addr[41620]= -395483624;
assign addr[41621]= -357831473;
assign addr[41622]= -320065829;
assign addr[41623]= -282198671;
assign addr[41624]= -244242007;
assign addr[41625]= -206207878;
assign addr[41626]= -168108346;
assign addr[41627]= -129955495;
assign addr[41628]= -91761426;
assign addr[41629]= -53538253;
assign addr[41630]= -15298099;
assign addr[41631]= 22946906;
assign addr[41632]= 61184634;
assign addr[41633]= 99402956;
assign addr[41634]= 137589750;
assign addr[41635]= 175732905;
assign addr[41636]= 213820322;
assign addr[41637]= 251839923;
assign addr[41638]= 289779648;
assign addr[41639]= 327627463;
assign addr[41640]= 365371365;
assign addr[41641]= 402999383;
assign addr[41642]= 440499581;
assign addr[41643]= 477860067;
assign addr[41644]= 515068990;
assign addr[41645]= 552114549;
assign addr[41646]= 588984994;
assign addr[41647]= 625668632;
assign addr[41648]= 662153826;
assign addr[41649]= 698429006;
assign addr[41650]= 734482665;
assign addr[41651]= 770303369;
assign addr[41652]= 805879757;
assign addr[41653]= 841200544;
assign addr[41654]= 876254528;
assign addr[41655]= 911030591;
assign addr[41656]= 945517704;
assign addr[41657]= 979704927;
assign addr[41658]= 1013581418;
assign addr[41659]= 1047136432;
assign addr[41660]= 1080359326;
assign addr[41661]= 1113239564;
assign addr[41662]= 1145766716;
assign addr[41663]= 1177930466;
assign addr[41664]= 1209720613;
assign addr[41665]= 1241127074;
assign addr[41666]= 1272139887;
assign addr[41667]= 1302749217;
assign addr[41668]= 1332945355;
assign addr[41669]= 1362718723;
assign addr[41670]= 1392059879;
assign addr[41671]= 1420959516;
assign addr[41672]= 1449408469;
assign addr[41673]= 1477397714;
assign addr[41674]= 1504918373;
assign addr[41675]= 1531961719;
assign addr[41676]= 1558519173;
assign addr[41677]= 1584582314;
assign addr[41678]= 1610142873;
assign addr[41679]= 1635192744;
assign addr[41680]= 1659723983;
assign addr[41681]= 1683728808;
assign addr[41682]= 1707199606;
assign addr[41683]= 1730128933;
assign addr[41684]= 1752509516;
assign addr[41685]= 1774334257;
assign addr[41686]= 1795596234;
assign addr[41687]= 1816288703;
assign addr[41688]= 1836405100;
assign addr[41689]= 1855939047;
assign addr[41690]= 1874884346;
assign addr[41691]= 1893234990;
assign addr[41692]= 1910985158;
assign addr[41693]= 1928129220;
assign addr[41694]= 1944661739;
assign addr[41695]= 1960577471;
assign addr[41696]= 1975871368;
assign addr[41697]= 1990538579;
assign addr[41698]= 2004574453;
assign addr[41699]= 2017974537;
assign addr[41700]= 2030734582;
assign addr[41701]= 2042850540;
assign addr[41702]= 2054318569;
assign addr[41703]= 2065135031;
assign addr[41704]= 2075296495;
assign addr[41705]= 2084799740;
assign addr[41706]= 2093641749;
assign addr[41707]= 2101819720;
assign addr[41708]= 2109331059;
assign addr[41709]= 2116173382;
assign addr[41710]= 2122344521;
assign addr[41711]= 2127842516;
assign addr[41712]= 2132665626;
assign addr[41713]= 2136812319;
assign addr[41714]= 2140281282;
assign addr[41715]= 2143071413;
assign addr[41716]= 2145181827;
assign addr[41717]= 2146611856;
assign addr[41718]= 2147361045;
assign addr[41719]= 2147429158;
assign addr[41720]= 2146816171;
assign addr[41721]= 2145522281;
assign addr[41722]= 2143547897;
assign addr[41723]= 2140893646;
assign addr[41724]= 2137560369;
assign addr[41725]= 2133549123;
assign addr[41726]= 2128861181;
assign addr[41727]= 2123498030;
assign addr[41728]= 2117461370;
assign addr[41729]= 2110753117;
assign addr[41730]= 2103375398;
assign addr[41731]= 2095330553;
assign addr[41732]= 2086621133;
assign addr[41733]= 2077249901;
assign addr[41734]= 2067219829;
assign addr[41735]= 2056534099;
assign addr[41736]= 2045196100;
assign addr[41737]= 2033209426;
assign addr[41738]= 2020577882;
assign addr[41739]= 2007305472;
assign addr[41740]= 1993396407;
assign addr[41741]= 1978855097;
assign addr[41742]= 1963686155;
assign addr[41743]= 1947894393;
assign addr[41744]= 1931484818;
assign addr[41745]= 1914462636;
assign addr[41746]= 1896833245;
assign addr[41747]= 1878602237;
assign addr[41748]= 1859775393;
assign addr[41749]= 1840358687;
assign addr[41750]= 1820358275;
assign addr[41751]= 1799780501;
assign addr[41752]= 1778631892;
assign addr[41753]= 1756919156;
assign addr[41754]= 1734649179;
assign addr[41755]= 1711829025;
assign addr[41756]= 1688465931;
assign addr[41757]= 1664567307;
assign addr[41758]= 1640140734;
assign addr[41759]= 1615193959;
assign addr[41760]= 1589734894;
assign addr[41761]= 1563771613;
assign addr[41762]= 1537312353;
assign addr[41763]= 1510365504;
assign addr[41764]= 1482939614;
assign addr[41765]= 1455043381;
assign addr[41766]= 1426685652;
assign addr[41767]= 1397875423;
assign addr[41768]= 1368621831;
assign addr[41769]= 1338934154;
assign addr[41770]= 1308821808;
assign addr[41771]= 1278294345;
assign addr[41772]= 1247361445;
assign addr[41773]= 1216032921;
assign addr[41774]= 1184318708;
assign addr[41775]= 1152228866;
assign addr[41776]= 1119773573;
assign addr[41777]= 1086963121;
assign addr[41778]= 1053807919;
assign addr[41779]= 1020318481;
assign addr[41780]= 986505429;
assign addr[41781]= 952379488;
assign addr[41782]= 917951481;
assign addr[41783]= 883232329;
assign addr[41784]= 848233042;
assign addr[41785]= 812964722;
assign addr[41786]= 777438554;
assign addr[41787]= 741665807;
assign addr[41788]= 705657826;
assign addr[41789]= 669426032;
assign addr[41790]= 632981917;
assign addr[41791]= 596337040;
assign addr[41792]= 559503022;
assign addr[41793]= 522491548;
assign addr[41794]= 485314355;
assign addr[41795]= 447983235;
assign addr[41796]= 410510029;
assign addr[41797]= 372906622;
assign addr[41798]= 335184940;
assign addr[41799]= 297356948;
assign addr[41800]= 259434643;
assign addr[41801]= 221430054;
assign addr[41802]= 183355234;
assign addr[41803]= 145222259;
assign addr[41804]= 107043224;
assign addr[41805]= 68830239;
assign addr[41806]= 30595422;
assign addr[41807]= -7649098;
assign addr[41808]= -45891193;
assign addr[41809]= -84118732;
assign addr[41810]= -122319591;
assign addr[41811]= -160481654;
assign addr[41812]= -198592817;
assign addr[41813]= -236640993;
assign addr[41814]= -274614114;
assign addr[41815]= -312500135;
assign addr[41816]= -350287041;
assign addr[41817]= -387962847;
assign addr[41818]= -425515602;
assign addr[41819]= -462933398;
assign addr[41820]= -500204365;
assign addr[41821]= -537316682;
assign addr[41822]= -574258580;
assign addr[41823]= -611018340;
assign addr[41824]= -647584304;
assign addr[41825]= -683944874;
assign addr[41826]= -720088517;
assign addr[41827]= -756003771;
assign addr[41828]= -791679244;
assign addr[41829]= -827103620;
assign addr[41830]= -862265664;
assign addr[41831]= -897154224;
assign addr[41832]= -931758235;
assign addr[41833]= -966066720;
assign addr[41834]= -1000068799;
assign addr[41835]= -1033753687;
assign addr[41836]= -1067110699;
assign addr[41837]= -1100129257;
assign addr[41838]= -1132798888;
assign addr[41839]= -1165109230;
assign addr[41840]= -1197050035;
assign addr[41841]= -1228611172;
assign addr[41842]= -1259782632;
assign addr[41843]= -1290554528;
assign addr[41844]= -1320917099;
assign addr[41845]= -1350860716;
assign addr[41846]= -1380375881;
assign addr[41847]= -1409453233;
assign addr[41848]= -1438083551;
assign addr[41849]= -1466257752;
assign addr[41850]= -1493966902;
assign addr[41851]= -1521202211;
assign addr[41852]= -1547955041;
assign addr[41853]= -1574216908;
assign addr[41854]= -1599979481;
assign addr[41855]= -1625234591;
assign addr[41856]= -1649974225;
assign addr[41857]= -1674190539;
assign addr[41858]= -1697875851;
assign addr[41859]= -1721022648;
assign addr[41860]= -1743623590;
assign addr[41861]= -1765671509;
assign addr[41862]= -1787159411;
assign addr[41863]= -1808080480;
assign addr[41864]= -1828428082;
assign addr[41865]= -1848195763;
assign addr[41866]= -1867377253;
assign addr[41867]= -1885966468;
assign addr[41868]= -1903957513;
assign addr[41869]= -1921344681;
assign addr[41870]= -1938122457;
assign addr[41871]= -1954285520;
assign addr[41872]= -1969828744;
assign addr[41873]= -1984747199;
assign addr[41874]= -1999036154;
assign addr[41875]= -2012691075;
assign addr[41876]= -2025707632;
assign addr[41877]= -2038081698;
assign addr[41878]= -2049809346;
assign addr[41879]= -2060886858;
assign addr[41880]= -2071310720;
assign addr[41881]= -2081077626;
assign addr[41882]= -2090184478;
assign addr[41883]= -2098628387;
assign addr[41884]= -2106406677;
assign addr[41885]= -2113516878;
assign addr[41886]= -2119956737;
assign addr[41887]= -2125724211;
assign addr[41888]= -2130817471;
assign addr[41889]= -2135234901;
assign addr[41890]= -2138975100;
assign addr[41891]= -2142036881;
assign addr[41892]= -2144419275;
assign addr[41893]= -2146121524;
assign addr[41894]= -2147143090;
assign addr[41895]= -2147483648;
assign addr[41896]= -2147143090;
assign addr[41897]= -2146121524;
assign addr[41898]= -2144419275;
assign addr[41899]= -2142036881;
assign addr[41900]= -2138975100;
assign addr[41901]= -2135234901;
assign addr[41902]= -2130817471;
assign addr[41903]= -2125724211;
assign addr[41904]= -2119956737;
assign addr[41905]= -2113516878;
assign addr[41906]= -2106406677;
assign addr[41907]= -2098628387;
assign addr[41908]= -2090184478;
assign addr[41909]= -2081077626;
assign addr[41910]= -2071310720;
assign addr[41911]= -2060886858;
assign addr[41912]= -2049809346;
assign addr[41913]= -2038081698;
assign addr[41914]= -2025707632;
assign addr[41915]= -2012691075;
assign addr[41916]= -1999036154;
assign addr[41917]= -1984747199;
assign addr[41918]= -1969828744;
assign addr[41919]= -1954285520;
assign addr[41920]= -1938122457;
assign addr[41921]= -1921344681;
assign addr[41922]= -1903957513;
assign addr[41923]= -1885966468;
assign addr[41924]= -1867377253;
assign addr[41925]= -1848195763;
assign addr[41926]= -1828428082;
assign addr[41927]= -1808080480;
assign addr[41928]= -1787159411;
assign addr[41929]= -1765671509;
assign addr[41930]= -1743623590;
assign addr[41931]= -1721022648;
assign addr[41932]= -1697875851;
assign addr[41933]= -1674190539;
assign addr[41934]= -1649974225;
assign addr[41935]= -1625234591;
assign addr[41936]= -1599979481;
assign addr[41937]= -1574216908;
assign addr[41938]= -1547955041;
assign addr[41939]= -1521202211;
assign addr[41940]= -1493966902;
assign addr[41941]= -1466257752;
assign addr[41942]= -1438083551;
assign addr[41943]= -1409453233;
assign addr[41944]= -1380375881;
assign addr[41945]= -1350860716;
assign addr[41946]= -1320917099;
assign addr[41947]= -1290554528;
assign addr[41948]= -1259782632;
assign addr[41949]= -1228611172;
assign addr[41950]= -1197050035;
assign addr[41951]= -1165109230;
assign addr[41952]= -1132798888;
assign addr[41953]= -1100129257;
assign addr[41954]= -1067110699;
assign addr[41955]= -1033753687;
assign addr[41956]= -1000068799;
assign addr[41957]= -966066720;
assign addr[41958]= -931758235;
assign addr[41959]= -897154224;
assign addr[41960]= -862265664;
assign addr[41961]= -827103620;
assign addr[41962]= -791679244;
assign addr[41963]= -756003771;
assign addr[41964]= -720088517;
assign addr[41965]= -683944874;
assign addr[41966]= -647584304;
assign addr[41967]= -611018340;
assign addr[41968]= -574258580;
assign addr[41969]= -537316682;
assign addr[41970]= -500204365;
assign addr[41971]= -462933398;
assign addr[41972]= -425515602;
assign addr[41973]= -387962847;
assign addr[41974]= -350287041;
assign addr[41975]= -312500135;
assign addr[41976]= -274614114;
assign addr[41977]= -236640993;
assign addr[41978]= -198592817;
assign addr[41979]= -160481654;
assign addr[41980]= -122319591;
assign addr[41981]= -84118732;
assign addr[41982]= -45891193;
assign addr[41983]= -7649098;
assign addr[41984]= 30595422;
assign addr[41985]= 68830239;
assign addr[41986]= 107043224;
assign addr[41987]= 145222259;
assign addr[41988]= 183355234;
assign addr[41989]= 221430054;
assign addr[41990]= 259434643;
assign addr[41991]= 297356948;
assign addr[41992]= 335184940;
assign addr[41993]= 372906622;
assign addr[41994]= 410510029;
assign addr[41995]= 447983235;
assign addr[41996]= 485314355;
assign addr[41997]= 522491548;
assign addr[41998]= 559503022;
assign addr[41999]= 596337040;
assign addr[42000]= 632981917;
assign addr[42001]= 669426032;
assign addr[42002]= 705657826;
assign addr[42003]= 741665807;
assign addr[42004]= 777438554;
assign addr[42005]= 812964722;
assign addr[42006]= 848233042;
assign addr[42007]= 883232329;
assign addr[42008]= 917951481;
assign addr[42009]= 952379488;
assign addr[42010]= 986505429;
assign addr[42011]= 1020318481;
assign addr[42012]= 1053807919;
assign addr[42013]= 1086963121;
assign addr[42014]= 1119773573;
assign addr[42015]= 1152228866;
assign addr[42016]= 1184318708;
assign addr[42017]= 1216032921;
assign addr[42018]= 1247361445;
assign addr[42019]= 1278294345;
assign addr[42020]= 1308821808;
assign addr[42021]= 1338934154;
assign addr[42022]= 1368621831;
assign addr[42023]= 1397875423;
assign addr[42024]= 1426685652;
assign addr[42025]= 1455043381;
assign addr[42026]= 1482939614;
assign addr[42027]= 1510365504;
assign addr[42028]= 1537312353;
assign addr[42029]= 1563771613;
assign addr[42030]= 1589734894;
assign addr[42031]= 1615193959;
assign addr[42032]= 1640140734;
assign addr[42033]= 1664567307;
assign addr[42034]= 1688465931;
assign addr[42035]= 1711829025;
assign addr[42036]= 1734649179;
assign addr[42037]= 1756919156;
assign addr[42038]= 1778631892;
assign addr[42039]= 1799780501;
assign addr[42040]= 1820358275;
assign addr[42041]= 1840358687;
assign addr[42042]= 1859775393;
assign addr[42043]= 1878602237;
assign addr[42044]= 1896833245;
assign addr[42045]= 1914462636;
assign addr[42046]= 1931484818;
assign addr[42047]= 1947894393;
assign addr[42048]= 1963686155;
assign addr[42049]= 1978855097;
assign addr[42050]= 1993396407;
assign addr[42051]= 2007305472;
assign addr[42052]= 2020577882;
assign addr[42053]= 2033209426;
assign addr[42054]= 2045196100;
assign addr[42055]= 2056534099;
assign addr[42056]= 2067219829;
assign addr[42057]= 2077249901;
assign addr[42058]= 2086621133;
assign addr[42059]= 2095330553;
assign addr[42060]= 2103375398;
assign addr[42061]= 2110753117;
assign addr[42062]= 2117461370;
assign addr[42063]= 2123498030;
assign addr[42064]= 2128861181;
assign addr[42065]= 2133549123;
assign addr[42066]= 2137560369;
assign addr[42067]= 2140893646;
assign addr[42068]= 2143547897;
assign addr[42069]= 2145522281;
assign addr[42070]= 2146816171;
assign addr[42071]= 2147429158;
assign addr[42072]= 2147361045;
assign addr[42073]= 2146611856;
assign addr[42074]= 2145181827;
assign addr[42075]= 2143071413;
assign addr[42076]= 2140281282;
assign addr[42077]= 2136812319;
assign addr[42078]= 2132665626;
assign addr[42079]= 2127842516;
assign addr[42080]= 2122344521;
assign addr[42081]= 2116173382;
assign addr[42082]= 2109331059;
assign addr[42083]= 2101819720;
assign addr[42084]= 2093641749;
assign addr[42085]= 2084799740;
assign addr[42086]= 2075296495;
assign addr[42087]= 2065135031;
assign addr[42088]= 2054318569;
assign addr[42089]= 2042850540;
assign addr[42090]= 2030734582;
assign addr[42091]= 2017974537;
assign addr[42092]= 2004574453;
assign addr[42093]= 1990538579;
assign addr[42094]= 1975871368;
assign addr[42095]= 1960577471;
assign addr[42096]= 1944661739;
assign addr[42097]= 1928129220;
assign addr[42098]= 1910985158;
assign addr[42099]= 1893234990;
assign addr[42100]= 1874884346;
assign addr[42101]= 1855939047;
assign addr[42102]= 1836405100;
assign addr[42103]= 1816288703;
assign addr[42104]= 1795596234;
assign addr[42105]= 1774334257;
assign addr[42106]= 1752509516;
assign addr[42107]= 1730128933;
assign addr[42108]= 1707199606;
assign addr[42109]= 1683728808;
assign addr[42110]= 1659723983;
assign addr[42111]= 1635192744;
assign addr[42112]= 1610142873;
assign addr[42113]= 1584582314;
assign addr[42114]= 1558519173;
assign addr[42115]= 1531961719;
assign addr[42116]= 1504918373;
assign addr[42117]= 1477397714;
assign addr[42118]= 1449408469;
assign addr[42119]= 1420959516;
assign addr[42120]= 1392059879;
assign addr[42121]= 1362718723;
assign addr[42122]= 1332945355;
assign addr[42123]= 1302749217;
assign addr[42124]= 1272139887;
assign addr[42125]= 1241127074;
assign addr[42126]= 1209720613;
assign addr[42127]= 1177930466;
assign addr[42128]= 1145766716;
assign addr[42129]= 1113239564;
assign addr[42130]= 1080359326;
assign addr[42131]= 1047136432;
assign addr[42132]= 1013581418;
assign addr[42133]= 979704927;
assign addr[42134]= 945517704;
assign addr[42135]= 911030591;
assign addr[42136]= 876254528;
assign addr[42137]= 841200544;
assign addr[42138]= 805879757;
assign addr[42139]= 770303369;
assign addr[42140]= 734482665;
assign addr[42141]= 698429006;
assign addr[42142]= 662153826;
assign addr[42143]= 625668632;
assign addr[42144]= 588984994;
assign addr[42145]= 552114549;
assign addr[42146]= 515068990;
assign addr[42147]= 477860067;
assign addr[42148]= 440499581;
assign addr[42149]= 402999383;
assign addr[42150]= 365371365;
assign addr[42151]= 327627463;
assign addr[42152]= 289779648;
assign addr[42153]= 251839923;
assign addr[42154]= 213820322;
assign addr[42155]= 175732905;
assign addr[42156]= 137589750;
assign addr[42157]= 99402956;
assign addr[42158]= 61184634;
assign addr[42159]= 22946906;
assign addr[42160]= -15298099;
assign addr[42161]= -53538253;
assign addr[42162]= -91761426;
assign addr[42163]= -129955495;
assign addr[42164]= -168108346;
assign addr[42165]= -206207878;
assign addr[42166]= -244242007;
assign addr[42167]= -282198671;
assign addr[42168]= -320065829;
assign addr[42169]= -357831473;
assign addr[42170]= -395483624;
assign addr[42171]= -433010339;
assign addr[42172]= -470399716;
assign addr[42173]= -507639898;
assign addr[42174]= -544719071;
assign addr[42175]= -581625477;
assign addr[42176]= -618347408;
assign addr[42177]= -654873219;
assign addr[42178]= -691191324;
assign addr[42179]= -727290205;
assign addr[42180]= -763158411;
assign addr[42181]= -798784567;
assign addr[42182]= -834157373;
assign addr[42183]= -869265610;
assign addr[42184]= -904098143;
assign addr[42185]= -938643924;
assign addr[42186]= -972891995;
assign addr[42187]= -1006831495;
assign addr[42188]= -1040451659;
assign addr[42189]= -1073741824;
assign addr[42190]= -1106691431;
assign addr[42191]= -1139290029;
assign addr[42192]= -1171527280;
assign addr[42193]= -1203392958;
assign addr[42194]= -1234876957;
assign addr[42195]= -1265969291;
assign addr[42196]= -1296660098;
assign addr[42197]= -1326939644;
assign addr[42198]= -1356798326;
assign addr[42199]= -1386226674;
assign addr[42200]= -1415215352;
assign addr[42201]= -1443755168;
assign addr[42202]= -1471837070;
assign addr[42203]= -1499452149;
assign addr[42204]= -1526591649;
assign addr[42205]= -1553246960;
assign addr[42206]= -1579409630;
assign addr[42207]= -1605071359;
assign addr[42208]= -1630224009;
assign addr[42209]= -1654859602;
assign addr[42210]= -1678970324;
assign addr[42211]= -1702548529;
assign addr[42212]= -1725586737;
assign addr[42213]= -1748077642;
assign addr[42214]= -1770014111;
assign addr[42215]= -1791389186;
assign addr[42216]= -1812196087;
assign addr[42217]= -1832428215;
assign addr[42218]= -1852079154;
assign addr[42219]= -1871142669;
assign addr[42220]= -1889612716;
assign addr[42221]= -1907483436;
assign addr[42222]= -1924749160;
assign addr[42223]= -1941404413;
assign addr[42224]= -1957443913;
assign addr[42225]= -1972862571;
assign addr[42226]= -1987655498;
assign addr[42227]= -2001818002;
assign addr[42228]= -2015345591;
assign addr[42229]= -2028233973;
assign addr[42230]= -2040479063;
assign addr[42231]= -2052076975;
assign addr[42232]= -2063024031;
assign addr[42233]= -2073316760;
assign addr[42234]= -2082951896;
assign addr[42235]= -2091926384;
assign addr[42236]= -2100237377;
assign addr[42237]= -2107882239;
assign addr[42238]= -2114858546;
assign addr[42239]= -2121164085;
assign addr[42240]= -2126796855;
assign addr[42241]= -2131755071;
assign addr[42242]= -2136037160;
assign addr[42243]= -2139641764;
assign addr[42244]= -2142567738;
assign addr[42245]= -2144814157;
assign addr[42246]= -2146380306;
assign addr[42247]= -2147265689;
assign addr[42248]= -2147470025;
assign addr[42249]= -2146993250;
assign addr[42250]= -2145835515;
assign addr[42251]= -2143997187;
assign addr[42252]= -2141478848;
assign addr[42253]= -2138281298;
assign addr[42254]= -2134405552;
assign addr[42255]= -2129852837;
assign addr[42256]= -2124624598;
assign addr[42257]= -2118722494;
assign addr[42258]= -2112148396;
assign addr[42259]= -2104904390;
assign addr[42260]= -2096992772;
assign addr[42261]= -2088416053;
assign addr[42262]= -2079176953;
assign addr[42263]= -2069278401;
assign addr[42264]= -2058723538;
assign addr[42265]= -2047515711;
assign addr[42266]= -2035658475;
assign addr[42267]= -2023155591;
assign addr[42268]= -2010011024;
assign addr[42269]= -1996228943;
assign addr[42270]= -1981813720;
assign addr[42271]= -1966769926;
assign addr[42272]= -1951102334;
assign addr[42273]= -1934815911;
assign addr[42274]= -1917915825;
assign addr[42275]= -1900407434;
assign addr[42276]= -1882296293;
assign addr[42277]= -1863588145;
assign addr[42278]= -1844288924;
assign addr[42279]= -1824404752;
assign addr[42280]= -1803941934;
assign addr[42281]= -1782906961;
assign addr[42282]= -1761306505;
assign addr[42283]= -1739147417;
assign addr[42284]= -1716436725;
assign addr[42285]= -1693181631;
assign addr[42286]= -1669389513;
assign addr[42287]= -1645067915;
assign addr[42288]= -1620224553;
assign addr[42289]= -1594867305;
assign addr[42290]= -1569004214;
assign addr[42291]= -1542643483;
assign addr[42292]= -1515793473;
assign addr[42293]= -1488462700;
assign addr[42294]= -1460659832;
assign addr[42295]= -1432393688;
assign addr[42296]= -1403673233;
assign addr[42297]= -1374507575;
assign addr[42298]= -1344905966;
assign addr[42299]= -1314877795;
assign addr[42300]= -1284432584;
assign addr[42301]= -1253579991;
assign addr[42302]= -1222329801;
assign addr[42303]= -1190691925;
assign addr[42304]= -1158676398;
assign addr[42305]= -1126293375;
assign addr[42306]= -1093553126;
assign addr[42307]= -1060466036;
assign addr[42308]= -1027042599;
assign addr[42309]= -993293415;
assign addr[42310]= -959229189;
assign addr[42311]= -924860725;
assign addr[42312]= -890198924;
assign addr[42313]= -855254778;
assign addr[42314]= -820039373;
assign addr[42315]= -784563876;
assign addr[42316]= -748839539;
assign addr[42317]= -712877694;
assign addr[42318]= -676689746;
assign addr[42319]= -640287172;
assign addr[42320]= -603681519;
assign addr[42321]= -566884397;
assign addr[42322]= -529907477;
assign addr[42323]= -492762486;
assign addr[42324]= -455461206;
assign addr[42325]= -418015468;
assign addr[42326]= -380437148;
assign addr[42327]= -342738165;
assign addr[42328]= -304930476;
assign addr[42329]= -267026072;
assign addr[42330]= -229036977;
assign addr[42331]= -190975237;
assign addr[42332]= -152852926;
assign addr[42333]= -114682135;
assign addr[42334]= -76474970;
assign addr[42335]= -38243550;
assign addr[42336]= 0;
assign addr[42337]= 38243550;
assign addr[42338]= 76474970;
assign addr[42339]= 114682135;
assign addr[42340]= 152852926;
assign addr[42341]= 190975237;
assign addr[42342]= 229036977;
assign addr[42343]= 267026072;
assign addr[42344]= 304930476;
assign addr[42345]= 342738165;
assign addr[42346]= 380437148;
assign addr[42347]= 418015468;
assign addr[42348]= 455461206;
assign addr[42349]= 492762486;
assign addr[42350]= 529907477;
assign addr[42351]= 566884397;
assign addr[42352]= 603681519;
assign addr[42353]= 640287172;
assign addr[42354]= 676689746;
assign addr[42355]= 712877694;
assign addr[42356]= 748839539;
assign addr[42357]= 784563876;
assign addr[42358]= 820039373;
assign addr[42359]= 855254778;
assign addr[42360]= 890198924;
assign addr[42361]= 924860725;
assign addr[42362]= 959229189;
assign addr[42363]= 993293415;
assign addr[42364]= 1027042599;
assign addr[42365]= 1060466036;
assign addr[42366]= 1093553126;
assign addr[42367]= 1126293375;
assign addr[42368]= 1158676398;
assign addr[42369]= 1190691925;
assign addr[42370]= 1222329801;
assign addr[42371]= 1253579991;
assign addr[42372]= 1284432584;
assign addr[42373]= 1314877795;
assign addr[42374]= 1344905966;
assign addr[42375]= 1374507575;
assign addr[42376]= 1403673233;
assign addr[42377]= 1432393688;
assign addr[42378]= 1460659832;
assign addr[42379]= 1488462700;
assign addr[42380]= 1515793473;
assign addr[42381]= 1542643483;
assign addr[42382]= 1569004214;
assign addr[42383]= 1594867305;
assign addr[42384]= 1620224553;
assign addr[42385]= 1645067915;
assign addr[42386]= 1669389513;
assign addr[42387]= 1693181631;
assign addr[42388]= 1716436725;
assign addr[42389]= 1739147417;
assign addr[42390]= 1761306505;
assign addr[42391]= 1782906961;
assign addr[42392]= 1803941934;
assign addr[42393]= 1824404752;
assign addr[42394]= 1844288924;
assign addr[42395]= 1863588145;
assign addr[42396]= 1882296293;
assign addr[42397]= 1900407434;
assign addr[42398]= 1917915825;
assign addr[42399]= 1934815911;
assign addr[42400]= 1951102334;
assign addr[42401]= 1966769926;
assign addr[42402]= 1981813720;
assign addr[42403]= 1996228943;
assign addr[42404]= 2010011024;
assign addr[42405]= 2023155591;
assign addr[42406]= 2035658475;
assign addr[42407]= 2047515711;
assign addr[42408]= 2058723538;
assign addr[42409]= 2069278401;
assign addr[42410]= 2079176953;
assign addr[42411]= 2088416053;
assign addr[42412]= 2096992772;
assign addr[42413]= 2104904390;
assign addr[42414]= 2112148396;
assign addr[42415]= 2118722494;
assign addr[42416]= 2124624598;
assign addr[42417]= 2129852837;
assign addr[42418]= 2134405552;
assign addr[42419]= 2138281298;
assign addr[42420]= 2141478848;
assign addr[42421]= 2143997187;
assign addr[42422]= 2145835515;
assign addr[42423]= 2146993250;
assign addr[42424]= 2147470025;
assign addr[42425]= 2147265689;
assign addr[42426]= 2146380306;
assign addr[42427]= 2144814157;
assign addr[42428]= 2142567738;
assign addr[42429]= 2139641764;
assign addr[42430]= 2136037160;
assign addr[42431]= 2131755071;
assign addr[42432]= 2126796855;
assign addr[42433]= 2121164085;
assign addr[42434]= 2114858546;
assign addr[42435]= 2107882239;
assign addr[42436]= 2100237377;
assign addr[42437]= 2091926384;
assign addr[42438]= 2082951896;
assign addr[42439]= 2073316760;
assign addr[42440]= 2063024031;
assign addr[42441]= 2052076975;
assign addr[42442]= 2040479063;
assign addr[42443]= 2028233973;
assign addr[42444]= 2015345591;
assign addr[42445]= 2001818002;
assign addr[42446]= 1987655498;
assign addr[42447]= 1972862571;
assign addr[42448]= 1957443913;
assign addr[42449]= 1941404413;
assign addr[42450]= 1924749160;
assign addr[42451]= 1907483436;
assign addr[42452]= 1889612716;
assign addr[42453]= 1871142669;
assign addr[42454]= 1852079154;
assign addr[42455]= 1832428215;
assign addr[42456]= 1812196087;
assign addr[42457]= 1791389186;
assign addr[42458]= 1770014111;
assign addr[42459]= 1748077642;
assign addr[42460]= 1725586737;
assign addr[42461]= 1702548529;
assign addr[42462]= 1678970324;
assign addr[42463]= 1654859602;
assign addr[42464]= 1630224009;
assign addr[42465]= 1605071359;
assign addr[42466]= 1579409630;
assign addr[42467]= 1553246960;
assign addr[42468]= 1526591649;
assign addr[42469]= 1499452149;
assign addr[42470]= 1471837070;
assign addr[42471]= 1443755168;
assign addr[42472]= 1415215352;
assign addr[42473]= 1386226674;
assign addr[42474]= 1356798326;
assign addr[42475]= 1326939644;
assign addr[42476]= 1296660098;
assign addr[42477]= 1265969291;
assign addr[42478]= 1234876957;
assign addr[42479]= 1203392958;
assign addr[42480]= 1171527280;
assign addr[42481]= 1139290029;
assign addr[42482]= 1106691431;
assign addr[42483]= 1073741824;
assign addr[42484]= 1040451659;
assign addr[42485]= 1006831495;
assign addr[42486]= 972891995;
assign addr[42487]= 938643924;
assign addr[42488]= 904098143;
assign addr[42489]= 869265610;
assign addr[42490]= 834157373;
assign addr[42491]= 798784567;
assign addr[42492]= 763158411;
assign addr[42493]= 727290205;
assign addr[42494]= 691191324;
assign addr[42495]= 654873219;
assign addr[42496]= 618347408;
assign addr[42497]= 581625477;
assign addr[42498]= 544719071;
assign addr[42499]= 507639898;
assign addr[42500]= 470399716;
assign addr[42501]= 433010339;
assign addr[42502]= 395483624;
assign addr[42503]= 357831473;
assign addr[42504]= 320065829;
assign addr[42505]= 282198671;
assign addr[42506]= 244242007;
assign addr[42507]= 206207878;
assign addr[42508]= 168108346;
assign addr[42509]= 129955495;
assign addr[42510]= 91761426;
assign addr[42511]= 53538253;
assign addr[42512]= 15298099;
assign addr[42513]= -22946906;
assign addr[42514]= -61184634;
assign addr[42515]= -99402956;
assign addr[42516]= -137589750;
assign addr[42517]= -175732905;
assign addr[42518]= -213820322;
assign addr[42519]= -251839923;
assign addr[42520]= -289779648;
assign addr[42521]= -327627463;
assign addr[42522]= -365371365;
assign addr[42523]= -402999383;
assign addr[42524]= -440499581;
assign addr[42525]= -477860067;
assign addr[42526]= -515068990;
assign addr[42527]= -552114549;
assign addr[42528]= -588984994;
assign addr[42529]= -625668632;
assign addr[42530]= -662153826;
assign addr[42531]= -698429006;
assign addr[42532]= -734482665;
assign addr[42533]= -770303369;
assign addr[42534]= -805879757;
assign addr[42535]= -841200544;
assign addr[42536]= -876254528;
assign addr[42537]= -911030591;
assign addr[42538]= -945517704;
assign addr[42539]= -979704927;
assign addr[42540]= -1013581418;
assign addr[42541]= -1047136432;
assign addr[42542]= -1080359326;
assign addr[42543]= -1113239564;
assign addr[42544]= -1145766716;
assign addr[42545]= -1177930466;
assign addr[42546]= -1209720613;
assign addr[42547]= -1241127074;
assign addr[42548]= -1272139887;
assign addr[42549]= -1302749217;
assign addr[42550]= -1332945355;
assign addr[42551]= -1362718723;
assign addr[42552]= -1392059879;
assign addr[42553]= -1420959516;
assign addr[42554]= -1449408469;
assign addr[42555]= -1477397714;
assign addr[42556]= -1504918373;
assign addr[42557]= -1531961719;
assign addr[42558]= -1558519173;
assign addr[42559]= -1584582314;
assign addr[42560]= -1610142873;
assign addr[42561]= -1635192744;
assign addr[42562]= -1659723983;
assign addr[42563]= -1683728808;
assign addr[42564]= -1707199606;
assign addr[42565]= -1730128933;
assign addr[42566]= -1752509516;
assign addr[42567]= -1774334257;
assign addr[42568]= -1795596234;
assign addr[42569]= -1816288703;
assign addr[42570]= -1836405100;
assign addr[42571]= -1855939047;
assign addr[42572]= -1874884346;
assign addr[42573]= -1893234990;
assign addr[42574]= -1910985158;
assign addr[42575]= -1928129220;
assign addr[42576]= -1944661739;
assign addr[42577]= -1960577471;
assign addr[42578]= -1975871368;
assign addr[42579]= -1990538579;
assign addr[42580]= -2004574453;
assign addr[42581]= -2017974537;
assign addr[42582]= -2030734582;
assign addr[42583]= -2042850540;
assign addr[42584]= -2054318569;
assign addr[42585]= -2065135031;
assign addr[42586]= -2075296495;
assign addr[42587]= -2084799740;
assign addr[42588]= -2093641749;
assign addr[42589]= -2101819720;
assign addr[42590]= -2109331059;
assign addr[42591]= -2116173382;
assign addr[42592]= -2122344521;
assign addr[42593]= -2127842516;
assign addr[42594]= -2132665626;
assign addr[42595]= -2136812319;
assign addr[42596]= -2140281282;
assign addr[42597]= -2143071413;
assign addr[42598]= -2145181827;
assign addr[42599]= -2146611856;
assign addr[42600]= -2147361045;
assign addr[42601]= -2147429158;
assign addr[42602]= -2146816171;
assign addr[42603]= -2145522281;
assign addr[42604]= -2143547897;
assign addr[42605]= -2140893646;
assign addr[42606]= -2137560369;
assign addr[42607]= -2133549123;
assign addr[42608]= -2128861181;
assign addr[42609]= -2123498030;
assign addr[42610]= -2117461370;
assign addr[42611]= -2110753117;
assign addr[42612]= -2103375398;
assign addr[42613]= -2095330553;
assign addr[42614]= -2086621133;
assign addr[42615]= -2077249901;
assign addr[42616]= -2067219829;
assign addr[42617]= -2056534099;
assign addr[42618]= -2045196100;
assign addr[42619]= -2033209426;
assign addr[42620]= -2020577882;
assign addr[42621]= -2007305472;
assign addr[42622]= -1993396407;
assign addr[42623]= -1978855097;
assign addr[42624]= -1963686155;
assign addr[42625]= -1947894393;
assign addr[42626]= -1931484818;
assign addr[42627]= -1914462636;
assign addr[42628]= -1896833245;
assign addr[42629]= -1878602237;
assign addr[42630]= -1859775393;
assign addr[42631]= -1840358687;
assign addr[42632]= -1820358275;
assign addr[42633]= -1799780501;
assign addr[42634]= -1778631892;
assign addr[42635]= -1756919156;
assign addr[42636]= -1734649179;
assign addr[42637]= -1711829025;
assign addr[42638]= -1688465931;
assign addr[42639]= -1664567307;
assign addr[42640]= -1640140734;
assign addr[42641]= -1615193959;
assign addr[42642]= -1589734894;
assign addr[42643]= -1563771613;
assign addr[42644]= -1537312353;
assign addr[42645]= -1510365504;
assign addr[42646]= -1482939614;
assign addr[42647]= -1455043381;
assign addr[42648]= -1426685652;
assign addr[42649]= -1397875423;
assign addr[42650]= -1368621831;
assign addr[42651]= -1338934154;
assign addr[42652]= -1308821808;
assign addr[42653]= -1278294345;
assign addr[42654]= -1247361445;
assign addr[42655]= -1216032921;
assign addr[42656]= -1184318708;
assign addr[42657]= -1152228866;
assign addr[42658]= -1119773573;
assign addr[42659]= -1086963121;
assign addr[42660]= -1053807919;
assign addr[42661]= -1020318481;
assign addr[42662]= -986505429;
assign addr[42663]= -952379488;
assign addr[42664]= -917951481;
assign addr[42665]= -883232329;
assign addr[42666]= -848233042;
assign addr[42667]= -812964722;
assign addr[42668]= -777438554;
assign addr[42669]= -741665807;
assign addr[42670]= -705657826;
assign addr[42671]= -669426032;
assign addr[42672]= -632981917;
assign addr[42673]= -596337040;
assign addr[42674]= -559503022;
assign addr[42675]= -522491548;
assign addr[42676]= -485314355;
assign addr[42677]= -447983235;
assign addr[42678]= -410510029;
assign addr[42679]= -372906622;
assign addr[42680]= -335184940;
assign addr[42681]= -297356948;
assign addr[42682]= -259434643;
assign addr[42683]= -221430054;
assign addr[42684]= -183355234;
assign addr[42685]= -145222259;
assign addr[42686]= -107043224;
assign addr[42687]= -68830239;
assign addr[42688]= -30595422;
assign addr[42689]= 7649098;
assign addr[42690]= 45891193;
assign addr[42691]= 84118732;
assign addr[42692]= 122319591;
assign addr[42693]= 160481654;
assign addr[42694]= 198592817;
assign addr[42695]= 236640993;
assign addr[42696]= 274614114;
assign addr[42697]= 312500135;
assign addr[42698]= 350287041;
assign addr[42699]= 387962847;
assign addr[42700]= 425515602;
assign addr[42701]= 462933398;
assign addr[42702]= 500204365;
assign addr[42703]= 537316682;
assign addr[42704]= 574258580;
assign addr[42705]= 611018340;
assign addr[42706]= 647584304;
assign addr[42707]= 683944874;
assign addr[42708]= 720088517;
assign addr[42709]= 756003771;
assign addr[42710]= 791679244;
assign addr[42711]= 827103620;
assign addr[42712]= 862265664;
assign addr[42713]= 897154224;
assign addr[42714]= 931758235;
assign addr[42715]= 966066720;
assign addr[42716]= 1000068799;
assign addr[42717]= 1033753687;
assign addr[42718]= 1067110699;
assign addr[42719]= 1100129257;
assign addr[42720]= 1132798888;
assign addr[42721]= 1165109230;
assign addr[42722]= 1197050035;
assign addr[42723]= 1228611172;
assign addr[42724]= 1259782632;
assign addr[42725]= 1290554528;
assign addr[42726]= 1320917099;
assign addr[42727]= 1350860716;
assign addr[42728]= 1380375881;
assign addr[42729]= 1409453233;
assign addr[42730]= 1438083551;
assign addr[42731]= 1466257752;
assign addr[42732]= 1493966902;
assign addr[42733]= 1521202211;
assign addr[42734]= 1547955041;
assign addr[42735]= 1574216908;
assign addr[42736]= 1599979481;
assign addr[42737]= 1625234591;
assign addr[42738]= 1649974225;
assign addr[42739]= 1674190539;
assign addr[42740]= 1697875851;
assign addr[42741]= 1721022648;
assign addr[42742]= 1743623590;
assign addr[42743]= 1765671509;
assign addr[42744]= 1787159411;
assign addr[42745]= 1808080480;
assign addr[42746]= 1828428082;
assign addr[42747]= 1848195763;
assign addr[42748]= 1867377253;
assign addr[42749]= 1885966468;
assign addr[42750]= 1903957513;
assign addr[42751]= 1921344681;
assign addr[42752]= 1938122457;
assign addr[42753]= 1954285520;
assign addr[42754]= 1969828744;
assign addr[42755]= 1984747199;
assign addr[42756]= 1999036154;
assign addr[42757]= 2012691075;
assign addr[42758]= 2025707632;
assign addr[42759]= 2038081698;
assign addr[42760]= 2049809346;
assign addr[42761]= 2060886858;
assign addr[42762]= 2071310720;
assign addr[42763]= 2081077626;
assign addr[42764]= 2090184478;
assign addr[42765]= 2098628387;
assign addr[42766]= 2106406677;
assign addr[42767]= 2113516878;
assign addr[42768]= 2119956737;
assign addr[42769]= 2125724211;
assign addr[42770]= 2130817471;
assign addr[42771]= 2135234901;
assign addr[42772]= 2138975100;
assign addr[42773]= 2142036881;
assign addr[42774]= 2144419275;
assign addr[42775]= 2146121524;
assign addr[42776]= 2147143090;
assign addr[42777]= 2147483648;
assign addr[42778]= 2147143090;
assign addr[42779]= 2146121524;
assign addr[42780]= 2144419275;
assign addr[42781]= 2142036881;
assign addr[42782]= 2138975100;
assign addr[42783]= 2135234901;
assign addr[42784]= 2130817471;
assign addr[42785]= 2125724211;
assign addr[42786]= 2119956737;
assign addr[42787]= 2113516878;
assign addr[42788]= 2106406677;
assign addr[42789]= 2098628387;
assign addr[42790]= 2090184478;
assign addr[42791]= 2081077626;
assign addr[42792]= 2071310720;
assign addr[42793]= 2060886858;
assign addr[42794]= 2049809346;
assign addr[42795]= 2038081698;
assign addr[42796]= 2025707632;
assign addr[42797]= 2012691075;
assign addr[42798]= 1999036154;
assign addr[42799]= 1984747199;
assign addr[42800]= 1969828744;
assign addr[42801]= 1954285520;
assign addr[42802]= 1938122457;
assign addr[42803]= 1921344681;
assign addr[42804]= 1903957513;
assign addr[42805]= 1885966468;
assign addr[42806]= 1867377253;
assign addr[42807]= 1848195763;
assign addr[42808]= 1828428082;
assign addr[42809]= 1808080480;
assign addr[42810]= 1787159411;
assign addr[42811]= 1765671509;
assign addr[42812]= 1743623590;
assign addr[42813]= 1721022648;
assign addr[42814]= 1697875851;
assign addr[42815]= 1674190539;
assign addr[42816]= 1649974225;
assign addr[42817]= 1625234591;
assign addr[42818]= 1599979481;
assign addr[42819]= 1574216908;
assign addr[42820]= 1547955041;
assign addr[42821]= 1521202211;
assign addr[42822]= 1493966902;
assign addr[42823]= 1466257752;
assign addr[42824]= 1438083551;
assign addr[42825]= 1409453233;
assign addr[42826]= 1380375881;
assign addr[42827]= 1350860716;
assign addr[42828]= 1320917099;
assign addr[42829]= 1290554528;
assign addr[42830]= 1259782632;
assign addr[42831]= 1228611172;
assign addr[42832]= 1197050035;
assign addr[42833]= 1165109230;
assign addr[42834]= 1132798888;
assign addr[42835]= 1100129257;
assign addr[42836]= 1067110699;
assign addr[42837]= 1033753687;
assign addr[42838]= 1000068799;
assign addr[42839]= 966066720;
assign addr[42840]= 931758235;
assign addr[42841]= 897154224;
assign addr[42842]= 862265664;
assign addr[42843]= 827103620;
assign addr[42844]= 791679244;
assign addr[42845]= 756003771;
assign addr[42846]= 720088517;
assign addr[42847]= 683944874;
assign addr[42848]= 647584304;
assign addr[42849]= 611018340;
assign addr[42850]= 574258580;
assign addr[42851]= 537316682;
assign addr[42852]= 500204365;
assign addr[42853]= 462933398;
assign addr[42854]= 425515602;
assign addr[42855]= 387962847;
assign addr[42856]= 350287041;
assign addr[42857]= 312500135;
assign addr[42858]= 274614114;
assign addr[42859]= 236640993;
assign addr[42860]= 198592817;
assign addr[42861]= 160481654;
assign addr[42862]= 122319591;
assign addr[42863]= 84118732;
assign addr[42864]= 45891193;
assign addr[42865]= 7649098;
assign addr[42866]= -30595422;
assign addr[42867]= -68830239;
assign addr[42868]= -107043224;
assign addr[42869]= -145222259;
assign addr[42870]= -183355234;
assign addr[42871]= -221430054;
assign addr[42872]= -259434643;
assign addr[42873]= -297356948;
assign addr[42874]= -335184940;
assign addr[42875]= -372906622;
assign addr[42876]= -410510029;
assign addr[42877]= -447983235;
assign addr[42878]= -485314355;
assign addr[42879]= -522491548;
assign addr[42880]= -559503022;
assign addr[42881]= -596337040;
assign addr[42882]= -632981917;
assign addr[42883]= -669426032;
assign addr[42884]= -705657826;
assign addr[42885]= -741665807;
assign addr[42886]= -777438554;
assign addr[42887]= -812964722;
assign addr[42888]= -848233042;
assign addr[42889]= -883232329;
assign addr[42890]= -917951481;
assign addr[42891]= -952379488;
assign addr[42892]= -986505429;
assign addr[42893]= -1020318481;
assign addr[42894]= -1053807919;
assign addr[42895]= -1086963121;
assign addr[42896]= -1119773573;
assign addr[42897]= -1152228866;
assign addr[42898]= -1184318708;
assign addr[42899]= -1216032921;
assign addr[42900]= -1247361445;
assign addr[42901]= -1278294345;
assign addr[42902]= -1308821808;
assign addr[42903]= -1338934154;
assign addr[42904]= -1368621831;
assign addr[42905]= -1397875423;
assign addr[42906]= -1426685652;
assign addr[42907]= -1455043381;
assign addr[42908]= -1482939614;
assign addr[42909]= -1510365504;
assign addr[42910]= -1537312353;
assign addr[42911]= -1563771613;
assign addr[42912]= -1589734894;
assign addr[42913]= -1615193959;
assign addr[42914]= -1640140734;
assign addr[42915]= -1664567307;
assign addr[42916]= -1688465931;
assign addr[42917]= -1711829025;
assign addr[42918]= -1734649179;
assign addr[42919]= -1756919156;
assign addr[42920]= -1778631892;
assign addr[42921]= -1799780501;
assign addr[42922]= -1820358275;
assign addr[42923]= -1840358687;
assign addr[42924]= -1859775393;
assign addr[42925]= -1878602237;
assign addr[42926]= -1896833245;
assign addr[42927]= -1914462636;
assign addr[42928]= -1931484818;
assign addr[42929]= -1947894393;
assign addr[42930]= -1963686155;
assign addr[42931]= -1978855097;
assign addr[42932]= -1993396407;
assign addr[42933]= -2007305472;
assign addr[42934]= -2020577882;
assign addr[42935]= -2033209426;
assign addr[42936]= -2045196100;
assign addr[42937]= -2056534099;
assign addr[42938]= -2067219829;
assign addr[42939]= -2077249901;
assign addr[42940]= -2086621133;
assign addr[42941]= -2095330553;
assign addr[42942]= -2103375398;
assign addr[42943]= -2110753117;
assign addr[42944]= -2117461370;
assign addr[42945]= -2123498030;
assign addr[42946]= -2128861181;
assign addr[42947]= -2133549123;
assign addr[42948]= -2137560369;
assign addr[42949]= -2140893646;
assign addr[42950]= -2143547897;
assign addr[42951]= -2145522281;
assign addr[42952]= -2146816171;
assign addr[42953]= -2147429158;
assign addr[42954]= -2147361045;
assign addr[42955]= -2146611856;
assign addr[42956]= -2145181827;
assign addr[42957]= -2143071413;
assign addr[42958]= -2140281282;
assign addr[42959]= -2136812319;
assign addr[42960]= -2132665626;
assign addr[42961]= -2127842516;
assign addr[42962]= -2122344521;
assign addr[42963]= -2116173382;
assign addr[42964]= -2109331059;
assign addr[42965]= -2101819720;
assign addr[42966]= -2093641749;
assign addr[42967]= -2084799740;
assign addr[42968]= -2075296495;
assign addr[42969]= -2065135031;
assign addr[42970]= -2054318569;
assign addr[42971]= -2042850540;
assign addr[42972]= -2030734582;
assign addr[42973]= -2017974537;
assign addr[42974]= -2004574453;
assign addr[42975]= -1990538579;
assign addr[42976]= -1975871368;
assign addr[42977]= -1960577471;
assign addr[42978]= -1944661739;
assign addr[42979]= -1928129220;
assign addr[42980]= -1910985158;
assign addr[42981]= -1893234990;
assign addr[42982]= -1874884346;
assign addr[42983]= -1855939047;
assign addr[42984]= -1836405100;
assign addr[42985]= -1816288703;
assign addr[42986]= -1795596234;
assign addr[42987]= -1774334257;
assign addr[42988]= -1752509516;
assign addr[42989]= -1730128933;
assign addr[42990]= -1707199606;
assign addr[42991]= -1683728808;
assign addr[42992]= -1659723983;
assign addr[42993]= -1635192744;
assign addr[42994]= -1610142873;
assign addr[42995]= -1584582314;
assign addr[42996]= -1558519173;
assign addr[42997]= -1531961719;
assign addr[42998]= -1504918373;
assign addr[42999]= -1477397714;
assign addr[43000]= -1449408469;
assign addr[43001]= -1420959516;
assign addr[43002]= -1392059879;
assign addr[43003]= -1362718723;
assign addr[43004]= -1332945355;
assign addr[43005]= -1302749217;
assign addr[43006]= -1272139887;
assign addr[43007]= -1241127074;
assign addr[43008]= -1209720613;
assign addr[43009]= -1177930466;
assign addr[43010]= -1145766716;
assign addr[43011]= -1113239564;
assign addr[43012]= -1080359326;
assign addr[43013]= -1047136432;
assign addr[43014]= -1013581418;
assign addr[43015]= -979704927;
assign addr[43016]= -945517704;
assign addr[43017]= -911030591;
assign addr[43018]= -876254528;
assign addr[43019]= -841200544;
assign addr[43020]= -805879757;
assign addr[43021]= -770303369;
assign addr[43022]= -734482665;
assign addr[43023]= -698429006;
assign addr[43024]= -662153826;
assign addr[43025]= -625668632;
assign addr[43026]= -588984994;
assign addr[43027]= -552114549;
assign addr[43028]= -515068990;
assign addr[43029]= -477860067;
assign addr[43030]= -440499581;
assign addr[43031]= -402999383;
assign addr[43032]= -365371365;
assign addr[43033]= -327627463;
assign addr[43034]= -289779648;
assign addr[43035]= -251839923;
assign addr[43036]= -213820322;
assign addr[43037]= -175732905;
assign addr[43038]= -137589750;
assign addr[43039]= -99402956;
assign addr[43040]= -61184634;
assign addr[43041]= -22946906;
assign addr[43042]= 15298099;
assign addr[43043]= 53538253;
assign addr[43044]= 91761426;
assign addr[43045]= 129955495;
assign addr[43046]= 168108346;
assign addr[43047]= 206207878;
assign addr[43048]= 244242007;
assign addr[43049]= 282198671;
assign addr[43050]= 320065829;
assign addr[43051]= 357831473;
assign addr[43052]= 395483624;
assign addr[43053]= 433010339;
assign addr[43054]= 470399716;
assign addr[43055]= 507639898;
assign addr[43056]= 544719071;
assign addr[43057]= 581625477;
assign addr[43058]= 618347408;
assign addr[43059]= 654873219;
assign addr[43060]= 691191324;
assign addr[43061]= 727290205;
assign addr[43062]= 763158411;
assign addr[43063]= 798784567;
assign addr[43064]= 834157373;
assign addr[43065]= 869265610;
assign addr[43066]= 904098143;
assign addr[43067]= 938643924;
assign addr[43068]= 972891995;
assign addr[43069]= 1006831495;
assign addr[43070]= 1040451659;
assign addr[43071]= 1073741824;
assign addr[43072]= 1106691431;
assign addr[43073]= 1139290029;
assign addr[43074]= 1171527280;
assign addr[43075]= 1203392958;
assign addr[43076]= 1234876957;
assign addr[43077]= 1265969291;
assign addr[43078]= 1296660098;
assign addr[43079]= 1326939644;
assign addr[43080]= 1356798326;
assign addr[43081]= 1386226674;
assign addr[43082]= 1415215352;
assign addr[43083]= 1443755168;
assign addr[43084]= 1471837070;
assign addr[43085]= 1499452149;
assign addr[43086]= 1526591649;
assign addr[43087]= 1553246960;
assign addr[43088]= 1579409630;
assign addr[43089]= 1605071359;
assign addr[43090]= 1630224009;
assign addr[43091]= 1654859602;
assign addr[43092]= 1678970324;
assign addr[43093]= 1702548529;
assign addr[43094]= 1725586737;
assign addr[43095]= 1748077642;
assign addr[43096]= 1770014111;
assign addr[43097]= 1791389186;
assign addr[43098]= 1812196087;
assign addr[43099]= 1832428215;
assign addr[43100]= 1852079154;
assign addr[43101]= 1871142669;
assign addr[43102]= 1889612716;
assign addr[43103]= 1907483436;
assign addr[43104]= 1924749160;
assign addr[43105]= 1941404413;
assign addr[43106]= 1957443913;
assign addr[43107]= 1972862571;
assign addr[43108]= 1987655498;
assign addr[43109]= 2001818002;
assign addr[43110]= 2015345591;
assign addr[43111]= 2028233973;
assign addr[43112]= 2040479063;
assign addr[43113]= 2052076975;
assign addr[43114]= 2063024031;
assign addr[43115]= 2073316760;
assign addr[43116]= 2082951896;
assign addr[43117]= 2091926384;
assign addr[43118]= 2100237377;
assign addr[43119]= 2107882239;
assign addr[43120]= 2114858546;
assign addr[43121]= 2121164085;
assign addr[43122]= 2126796855;
assign addr[43123]= 2131755071;
assign addr[43124]= 2136037160;
assign addr[43125]= 2139641764;
assign addr[43126]= 2142567738;
assign addr[43127]= 2144814157;
assign addr[43128]= 2146380306;
assign addr[43129]= 2147265689;
assign addr[43130]= 2147470025;
assign addr[43131]= 2146993250;
assign addr[43132]= 2145835515;
assign addr[43133]= 2143997187;
assign addr[43134]= 2141478848;
assign addr[43135]= 2138281298;
assign addr[43136]= 2134405552;
assign addr[43137]= 2129852837;
assign addr[43138]= 2124624598;
assign addr[43139]= 2118722494;
assign addr[43140]= 2112148396;
assign addr[43141]= 2104904390;
assign addr[43142]= 2096992772;
assign addr[43143]= 2088416053;
assign addr[43144]= 2079176953;
assign addr[43145]= 2069278401;
assign addr[43146]= 2058723538;
assign addr[43147]= 2047515711;
assign addr[43148]= 2035658475;
assign addr[43149]= 2023155591;
assign addr[43150]= 2010011024;
assign addr[43151]= 1996228943;
assign addr[43152]= 1981813720;
assign addr[43153]= 1966769926;
assign addr[43154]= 1951102334;
assign addr[43155]= 1934815911;
assign addr[43156]= 1917915825;
assign addr[43157]= 1900407434;
assign addr[43158]= 1882296293;
assign addr[43159]= 1863588145;
assign addr[43160]= 1844288924;
assign addr[43161]= 1824404752;
assign addr[43162]= 1803941934;
assign addr[43163]= 1782906961;
assign addr[43164]= 1761306505;
assign addr[43165]= 1739147417;
assign addr[43166]= 1716436725;
assign addr[43167]= 1693181631;
assign addr[43168]= 1669389513;
assign addr[43169]= 1645067915;
assign addr[43170]= 1620224553;
assign addr[43171]= 1594867305;
assign addr[43172]= 1569004214;
assign addr[43173]= 1542643483;
assign addr[43174]= 1515793473;
assign addr[43175]= 1488462700;
assign addr[43176]= 1460659832;
assign addr[43177]= 1432393688;
assign addr[43178]= 1403673233;
assign addr[43179]= 1374507575;
assign addr[43180]= 1344905966;
assign addr[43181]= 1314877795;
assign addr[43182]= 1284432584;
assign addr[43183]= 1253579991;
assign addr[43184]= 1222329801;
assign addr[43185]= 1190691925;
assign addr[43186]= 1158676398;
assign addr[43187]= 1126293375;
assign addr[43188]= 1093553126;
assign addr[43189]= 1060466036;
assign addr[43190]= 1027042599;
assign addr[43191]= 993293415;
assign addr[43192]= 959229189;
assign addr[43193]= 924860725;
assign addr[43194]= 890198924;
assign addr[43195]= 855254778;
assign addr[43196]= 820039373;
assign addr[43197]= 784563876;
assign addr[43198]= 748839539;
assign addr[43199]= 712877694;
assign addr[43200]= 676689746;
assign addr[43201]= 640287172;
assign addr[43202]= 603681519;
assign addr[43203]= 566884397;
assign addr[43204]= 529907477;
assign addr[43205]= 492762486;
assign addr[43206]= 455461206;
assign addr[43207]= 418015468;
assign addr[43208]= 380437148;
assign addr[43209]= 342738165;
assign addr[43210]= 304930476;
assign addr[43211]= 267026072;
assign addr[43212]= 229036977;
assign addr[43213]= 190975237;
assign addr[43214]= 152852926;
assign addr[43215]= 114682135;
assign addr[43216]= 76474970;
assign addr[43217]= 38243550;
assign addr[43218]= 0;
assign addr[43219]= -38243550;
assign addr[43220]= -76474970;
assign addr[43221]= -114682135;
assign addr[43222]= -152852926;
assign addr[43223]= -190975237;
assign addr[43224]= -229036977;
assign addr[43225]= -267026072;
assign addr[43226]= -304930476;
assign addr[43227]= -342738165;
assign addr[43228]= -380437148;
assign addr[43229]= -418015468;
assign addr[43230]= -455461206;
assign addr[43231]= -492762486;
assign addr[43232]= -529907477;
assign addr[43233]= -566884397;
assign addr[43234]= -603681519;
assign addr[43235]= -640287172;
assign addr[43236]= -676689746;
assign addr[43237]= -712877694;
assign addr[43238]= -748839539;
assign addr[43239]= -784563876;
assign addr[43240]= -820039373;
assign addr[43241]= -855254778;
assign addr[43242]= -890198924;
assign addr[43243]= -924860725;
assign addr[43244]= -959229189;
assign addr[43245]= -993293415;
assign addr[43246]= -1027042599;
assign addr[43247]= -1060466036;
assign addr[43248]= -1093553126;
assign addr[43249]= -1126293375;
assign addr[43250]= -1158676398;
assign addr[43251]= -1190691925;
assign addr[43252]= -1222329801;
assign addr[43253]= -1253579991;
assign addr[43254]= -1284432584;
assign addr[43255]= -1314877795;
assign addr[43256]= -1344905966;
assign addr[43257]= -1374507575;
assign addr[43258]= -1403673233;
assign addr[43259]= -1432393688;
assign addr[43260]= -1460659832;
assign addr[43261]= -1488462700;
assign addr[43262]= -1515793473;
assign addr[43263]= -1542643483;
assign addr[43264]= -1569004214;
assign addr[43265]= -1594867305;
assign addr[43266]= -1620224553;
assign addr[43267]= -1645067915;
assign addr[43268]= -1669389513;
assign addr[43269]= -1693181631;
assign addr[43270]= -1716436725;
assign addr[43271]= -1739147417;
assign addr[43272]= -1761306505;
assign addr[43273]= -1782906961;
assign addr[43274]= -1803941934;
assign addr[43275]= -1824404752;
assign addr[43276]= -1844288924;
assign addr[43277]= -1863588145;
assign addr[43278]= -1882296293;
assign addr[43279]= -1900407434;
assign addr[43280]= -1917915825;
assign addr[43281]= -1934815911;
assign addr[43282]= -1951102334;
assign addr[43283]= -1966769926;
assign addr[43284]= -1981813720;
assign addr[43285]= -1996228943;
assign addr[43286]= -2010011024;
assign addr[43287]= -2023155591;
assign addr[43288]= -2035658475;
assign addr[43289]= -2047515711;
assign addr[43290]= -2058723538;
assign addr[43291]= -2069278401;
assign addr[43292]= -2079176953;
assign addr[43293]= -2088416053;
assign addr[43294]= -2096992772;
assign addr[43295]= -2104904390;
assign addr[43296]= -2112148396;
assign addr[43297]= -2118722494;
assign addr[43298]= -2124624598;
assign addr[43299]= -2129852837;
assign addr[43300]= -2134405552;
assign addr[43301]= -2138281298;
assign addr[43302]= -2141478848;
assign addr[43303]= -2143997187;
assign addr[43304]= -2145835515;
assign addr[43305]= -2146993250;
assign addr[43306]= -2147470025;
assign addr[43307]= -2147265689;
assign addr[43308]= -2146380306;
assign addr[43309]= -2144814157;
assign addr[43310]= -2142567738;
assign addr[43311]= -2139641764;
assign addr[43312]= -2136037160;
assign addr[43313]= -2131755071;
assign addr[43314]= -2126796855;
assign addr[43315]= -2121164085;
assign addr[43316]= -2114858546;
assign addr[43317]= -2107882239;
assign addr[43318]= -2100237377;
assign addr[43319]= -2091926384;
assign addr[43320]= -2082951896;
assign addr[43321]= -2073316760;
assign addr[43322]= -2063024031;
assign addr[43323]= -2052076975;
assign addr[43324]= -2040479063;
assign addr[43325]= -2028233973;
assign addr[43326]= -2015345591;
assign addr[43327]= -2001818002;
assign addr[43328]= -1987655498;
assign addr[43329]= -1972862571;
assign addr[43330]= -1957443913;
assign addr[43331]= -1941404413;
assign addr[43332]= -1924749160;
assign addr[43333]= -1907483436;
assign addr[43334]= -1889612716;
assign addr[43335]= -1871142669;
assign addr[43336]= -1852079154;
assign addr[43337]= -1832428215;
assign addr[43338]= -1812196087;
assign addr[43339]= -1791389186;
assign addr[43340]= -1770014111;
assign addr[43341]= -1748077642;
assign addr[43342]= -1725586737;
assign addr[43343]= -1702548529;
assign addr[43344]= -1678970324;
assign addr[43345]= -1654859602;
assign addr[43346]= -1630224009;
assign addr[43347]= -1605071359;
assign addr[43348]= -1579409630;
assign addr[43349]= -1553246960;
assign addr[43350]= -1526591649;
assign addr[43351]= -1499452149;
assign addr[43352]= -1471837070;
assign addr[43353]= -1443755168;
assign addr[43354]= -1415215352;
assign addr[43355]= -1386226674;
assign addr[43356]= -1356798326;
assign addr[43357]= -1326939644;
assign addr[43358]= -1296660098;
assign addr[43359]= -1265969291;
assign addr[43360]= -1234876957;
assign addr[43361]= -1203392958;
assign addr[43362]= -1171527280;
assign addr[43363]= -1139290029;
assign addr[43364]= -1106691431;
assign addr[43365]= -1073741824;
assign addr[43366]= -1040451659;
assign addr[43367]= -1006831495;
assign addr[43368]= -972891995;
assign addr[43369]= -938643924;
assign addr[43370]= -904098143;
assign addr[43371]= -869265610;
assign addr[43372]= -834157373;
assign addr[43373]= -798784567;
assign addr[43374]= -763158411;
assign addr[43375]= -727290205;
assign addr[43376]= -691191324;
assign addr[43377]= -654873219;
assign addr[43378]= -618347408;
assign addr[43379]= -581625477;
assign addr[43380]= -544719071;
assign addr[43381]= -507639898;
assign addr[43382]= -470399716;
assign addr[43383]= -433010339;
assign addr[43384]= -395483624;
assign addr[43385]= -357831473;
assign addr[43386]= -320065829;
assign addr[43387]= -282198671;
assign addr[43388]= -244242007;
assign addr[43389]= -206207878;
assign addr[43390]= -168108346;
assign addr[43391]= -129955495;
assign addr[43392]= -91761426;
assign addr[43393]= -53538253;
assign addr[43394]= -15298099;
assign addr[43395]= 22946906;
assign addr[43396]= 61184634;
assign addr[43397]= 99402956;
assign addr[43398]= 137589750;
assign addr[43399]= 175732905;
assign addr[43400]= 213820322;
assign addr[43401]= 251839923;
assign addr[43402]= 289779648;
assign addr[43403]= 327627463;
assign addr[43404]= 365371365;
assign addr[43405]= 402999383;
assign addr[43406]= 440499581;
assign addr[43407]= 477860067;
assign addr[43408]= 515068990;
assign addr[43409]= 552114549;
assign addr[43410]= 588984994;
assign addr[43411]= 625668632;
assign addr[43412]= 662153826;
assign addr[43413]= 698429006;
assign addr[43414]= 734482665;
assign addr[43415]= 770303369;
assign addr[43416]= 805879757;
assign addr[43417]= 841200544;
assign addr[43418]= 876254528;
assign addr[43419]= 911030591;
assign addr[43420]= 945517704;
assign addr[43421]= 979704927;
assign addr[43422]= 1013581418;
assign addr[43423]= 1047136432;
assign addr[43424]= 1080359326;
assign addr[43425]= 1113239564;
assign addr[43426]= 1145766716;
assign addr[43427]= 1177930466;
assign addr[43428]= 1209720613;
assign addr[43429]= 1241127074;
assign addr[43430]= 1272139887;
assign addr[43431]= 1302749217;
assign addr[43432]= 1332945355;
assign addr[43433]= 1362718723;
assign addr[43434]= 1392059879;
assign addr[43435]= 1420959516;
assign addr[43436]= 1449408469;
assign addr[43437]= 1477397714;
assign addr[43438]= 1504918373;
assign addr[43439]= 1531961719;
assign addr[43440]= 1558519173;
assign addr[43441]= 1584582314;
assign addr[43442]= 1610142873;
assign addr[43443]= 1635192744;
assign addr[43444]= 1659723983;
assign addr[43445]= 1683728808;
assign addr[43446]= 1707199606;
assign addr[43447]= 1730128933;
assign addr[43448]= 1752509516;
assign addr[43449]= 1774334257;
assign addr[43450]= 1795596234;
assign addr[43451]= 1816288703;
assign addr[43452]= 1836405100;
assign addr[43453]= 1855939047;
assign addr[43454]= 1874884346;
assign addr[43455]= 1893234990;
assign addr[43456]= 1910985158;
assign addr[43457]= 1928129220;
assign addr[43458]= 1944661739;
assign addr[43459]= 1960577471;
assign addr[43460]= 1975871368;
assign addr[43461]= 1990538579;
assign addr[43462]= 2004574453;
assign addr[43463]= 2017974537;
assign addr[43464]= 2030734582;
assign addr[43465]= 2042850540;
assign addr[43466]= 2054318569;
assign addr[43467]= 2065135031;
assign addr[43468]= 2075296495;
assign addr[43469]= 2084799740;
assign addr[43470]= 2093641749;
assign addr[43471]= 2101819720;
assign addr[43472]= 2109331059;
assign addr[43473]= 2116173382;
assign addr[43474]= 2122344521;
assign addr[43475]= 2127842516;
assign addr[43476]= 2132665626;
assign addr[43477]= 2136812319;
assign addr[43478]= 2140281282;
assign addr[43479]= 2143071413;
assign addr[43480]= 2145181827;
assign addr[43481]= 2146611856;
assign addr[43482]= 2147361045;
assign addr[43483]= 2147429158;
assign addr[43484]= 2146816171;
assign addr[43485]= 2145522281;
assign addr[43486]= 2143547897;
assign addr[43487]= 2140893646;
assign addr[43488]= 2137560369;
assign addr[43489]= 2133549123;
assign addr[43490]= 2128861181;
assign addr[43491]= 2123498030;
assign addr[43492]= 2117461370;
assign addr[43493]= 2110753117;
assign addr[43494]= 2103375398;
assign addr[43495]= 2095330553;
assign addr[43496]= 2086621133;
assign addr[43497]= 2077249901;
assign addr[43498]= 2067219829;
assign addr[43499]= 2056534099;
assign addr[43500]= 2045196100;
assign addr[43501]= 2033209426;
assign addr[43502]= 2020577882;
assign addr[43503]= 2007305472;
assign addr[43504]= 1993396407;
assign addr[43505]= 1978855097;
assign addr[43506]= 1963686155;
assign addr[43507]= 1947894393;
assign addr[43508]= 1931484818;
assign addr[43509]= 1914462636;
assign addr[43510]= 1896833245;
assign addr[43511]= 1878602237;
assign addr[43512]= 1859775393;
assign addr[43513]= 1840358687;
assign addr[43514]= 1820358275;
assign addr[43515]= 1799780501;
assign addr[43516]= 1778631892;
assign addr[43517]= 1756919156;
assign addr[43518]= 1734649179;
assign addr[43519]= 1711829025;
assign addr[43520]= 1688465931;
assign addr[43521]= 1664567307;
assign addr[43522]= 1640140734;
assign addr[43523]= 1615193959;
assign addr[43524]= 1589734894;
assign addr[43525]= 1563771613;
assign addr[43526]= 1537312353;
assign addr[43527]= 1510365504;
assign addr[43528]= 1482939614;
assign addr[43529]= 1455043381;
assign addr[43530]= 1426685652;
assign addr[43531]= 1397875423;
assign addr[43532]= 1368621831;
assign addr[43533]= 1338934154;
assign addr[43534]= 1308821808;
assign addr[43535]= 1278294345;
assign addr[43536]= 1247361445;
assign addr[43537]= 1216032921;
assign addr[43538]= 1184318708;
assign addr[43539]= 1152228866;
assign addr[43540]= 1119773573;
assign addr[43541]= 1086963121;
assign addr[43542]= 1053807919;
assign addr[43543]= 1020318481;
assign addr[43544]= 986505429;
assign addr[43545]= 952379488;
assign addr[43546]= 917951481;
assign addr[43547]= 883232329;
assign addr[43548]= 848233042;
assign addr[43549]= 812964722;
assign addr[43550]= 777438554;
assign addr[43551]= 741665807;
assign addr[43552]= 705657826;
assign addr[43553]= 669426032;
assign addr[43554]= 632981917;
assign addr[43555]= 596337040;
assign addr[43556]= 559503022;
assign addr[43557]= 522491548;
assign addr[43558]= 485314355;
assign addr[43559]= 447983235;
assign addr[43560]= 410510029;
assign addr[43561]= 372906622;
assign addr[43562]= 335184940;
assign addr[43563]= 297356948;
assign addr[43564]= 259434643;
assign addr[43565]= 221430054;
assign addr[43566]= 183355234;
assign addr[43567]= 145222259;
assign addr[43568]= 107043224;
assign addr[43569]= 68830239;
assign addr[43570]= 30595422;
assign addr[43571]= -7649098;
assign addr[43572]= -45891193;
assign addr[43573]= -84118732;
assign addr[43574]= -122319591;
assign addr[43575]= -160481654;
assign addr[43576]= -198592817;
assign addr[43577]= -236640993;
assign addr[43578]= -274614114;
assign addr[43579]= -312500135;
assign addr[43580]= -350287041;
assign addr[43581]= -387962847;
assign addr[43582]= -425515602;
assign addr[43583]= -462933398;
assign addr[43584]= -500204365;
assign addr[43585]= -537316682;
assign addr[43586]= -574258580;
assign addr[43587]= -611018340;
assign addr[43588]= -647584304;
assign addr[43589]= -683944874;
assign addr[43590]= -720088517;
assign addr[43591]= -756003771;
assign addr[43592]= -791679244;
assign addr[43593]= -827103620;
assign addr[43594]= -862265664;
assign addr[43595]= -897154224;
assign addr[43596]= -931758235;
assign addr[43597]= -966066720;
assign addr[43598]= -1000068799;
assign addr[43599]= -1033753687;
assign addr[43600]= -1067110699;
assign addr[43601]= -1100129257;
assign addr[43602]= -1132798888;
assign addr[43603]= -1165109230;
assign addr[43604]= -1197050035;
assign addr[43605]= -1228611172;
assign addr[43606]= -1259782632;
assign addr[43607]= -1290554528;
assign addr[43608]= -1320917099;
assign addr[43609]= -1350860716;
assign addr[43610]= -1380375881;
assign addr[43611]= -1409453233;
assign addr[43612]= -1438083551;
assign addr[43613]= -1466257752;
assign addr[43614]= -1493966902;
assign addr[43615]= -1521202211;
assign addr[43616]= -1547955041;
assign addr[43617]= -1574216908;
assign addr[43618]= -1599979481;
assign addr[43619]= -1625234591;
assign addr[43620]= -1649974225;
assign addr[43621]= -1674190539;
assign addr[43622]= -1697875851;
assign addr[43623]= -1721022648;
assign addr[43624]= -1743623590;
assign addr[43625]= -1765671509;
assign addr[43626]= -1787159411;
assign addr[43627]= -1808080480;
assign addr[43628]= -1828428082;
assign addr[43629]= -1848195763;
assign addr[43630]= -1867377253;
assign addr[43631]= -1885966468;
assign addr[43632]= -1903957513;
assign addr[43633]= -1921344681;
assign addr[43634]= -1938122457;
assign addr[43635]= -1954285520;
assign addr[43636]= -1969828744;
assign addr[43637]= -1984747199;
assign addr[43638]= -1999036154;
assign addr[43639]= -2012691075;
assign addr[43640]= -2025707632;
assign addr[43641]= -2038081698;
assign addr[43642]= -2049809346;
assign addr[43643]= -2060886858;
assign addr[43644]= -2071310720;
assign addr[43645]= -2081077626;
assign addr[43646]= -2090184478;
assign addr[43647]= -2098628387;
assign addr[43648]= -2106406677;
assign addr[43649]= -2113516878;
assign addr[43650]= -2119956737;
assign addr[43651]= -2125724211;
assign addr[43652]= -2130817471;
assign addr[43653]= -2135234901;
assign addr[43654]= -2138975100;
assign addr[43655]= -2142036881;
assign addr[43656]= -2144419275;
assign addr[43657]= -2146121524;
assign addr[43658]= -2147143090;
assign addr[43659]= -2147483648;
assign addr[43660]= -2147143090;
assign addr[43661]= -2146121524;
assign addr[43662]= -2144419275;
assign addr[43663]= -2142036881;
assign addr[43664]= -2138975100;
assign addr[43665]= -2135234901;
assign addr[43666]= -2130817471;
assign addr[43667]= -2125724211;
assign addr[43668]= -2119956737;
assign addr[43669]= -2113516878;
assign addr[43670]= -2106406677;
assign addr[43671]= -2098628387;
assign addr[43672]= -2090184478;
assign addr[43673]= -2081077626;
assign addr[43674]= -2071310720;
assign addr[43675]= -2060886858;
assign addr[43676]= -2049809346;
assign addr[43677]= -2038081698;
assign addr[43678]= -2025707632;
assign addr[43679]= -2012691075;
assign addr[43680]= -1999036154;
assign addr[43681]= -1984747199;
assign addr[43682]= -1969828744;
assign addr[43683]= -1954285520;
assign addr[43684]= -1938122457;
assign addr[43685]= -1921344681;
assign addr[43686]= -1903957513;
assign addr[43687]= -1885966468;
assign addr[43688]= -1867377253;
assign addr[43689]= -1848195763;
assign addr[43690]= -1828428082;
assign addr[43691]= -1808080480;
assign addr[43692]= -1787159411;
assign addr[43693]= -1765671509;
assign addr[43694]= -1743623590;
assign addr[43695]= -1721022648;
assign addr[43696]= -1697875851;
assign addr[43697]= -1674190539;
assign addr[43698]= -1649974225;
assign addr[43699]= -1625234591;
assign addr[43700]= -1599979481;
assign addr[43701]= -1574216908;
assign addr[43702]= -1547955041;
assign addr[43703]= -1521202211;
assign addr[43704]= -1493966902;
assign addr[43705]= -1466257752;
assign addr[43706]= -1438083551;
assign addr[43707]= -1409453233;
assign addr[43708]= -1380375881;
assign addr[43709]= -1350860716;
assign addr[43710]= -1320917099;
assign addr[43711]= -1290554528;
assign addr[43712]= -1259782632;
assign addr[43713]= -1228611172;
assign addr[43714]= -1197050035;
assign addr[43715]= -1165109230;
assign addr[43716]= -1132798888;
assign addr[43717]= -1100129257;
assign addr[43718]= -1067110699;
assign addr[43719]= -1033753687;
assign addr[43720]= -1000068799;
assign addr[43721]= -966066720;
assign addr[43722]= -931758235;
assign addr[43723]= -897154224;
assign addr[43724]= -862265664;
assign addr[43725]= -827103620;
assign addr[43726]= -791679244;
assign addr[43727]= -756003771;
assign addr[43728]= -720088517;
assign addr[43729]= -683944874;
assign addr[43730]= -647584304;
assign addr[43731]= -611018340;
assign addr[43732]= -574258580;
assign addr[43733]= -537316682;
assign addr[43734]= -500204365;
assign addr[43735]= -462933398;
assign addr[43736]= -425515602;
assign addr[43737]= -387962847;
assign addr[43738]= -350287041;
assign addr[43739]= -312500135;
assign addr[43740]= -274614114;
assign addr[43741]= -236640993;
assign addr[43742]= -198592817;
assign addr[43743]= -160481654;
assign addr[43744]= -122319591;
assign addr[43745]= -84118732;
assign addr[43746]= -45891193;
assign addr[43747]= -7649098;
assign addr[43748]= 30595422;
assign addr[43749]= 68830239;
assign addr[43750]= 107043224;
assign addr[43751]= 145222259;
assign addr[43752]= 183355234;
assign addr[43753]= 221430054;
assign addr[43754]= 259434643;
assign addr[43755]= 297356948;
assign addr[43756]= 335184940;
assign addr[43757]= 372906622;
assign addr[43758]= 410510029;
assign addr[43759]= 447983235;
assign addr[43760]= 485314355;
assign addr[43761]= 522491548;
assign addr[43762]= 559503022;
assign addr[43763]= 596337040;
assign addr[43764]= 632981917;
assign addr[43765]= 669426032;
assign addr[43766]= 705657826;
assign addr[43767]= 741665807;
assign addr[43768]= 777438554;
assign addr[43769]= 812964722;
assign addr[43770]= 848233042;
assign addr[43771]= 883232329;
assign addr[43772]= 917951481;
assign addr[43773]= 952379488;
assign addr[43774]= 986505429;
assign addr[43775]= 1020318481;
assign addr[43776]= 1053807919;
assign addr[43777]= 1086963121;
assign addr[43778]= 1119773573;
assign addr[43779]= 1152228866;
assign addr[43780]= 1184318708;
assign addr[43781]= 1216032921;
assign addr[43782]= 1247361445;
assign addr[43783]= 1278294345;
assign addr[43784]= 1308821808;
assign addr[43785]= 1338934154;
assign addr[43786]= 1368621831;
assign addr[43787]= 1397875423;
assign addr[43788]= 1426685652;
assign addr[43789]= 1455043381;
assign addr[43790]= 1482939614;
assign addr[43791]= 1510365504;
assign addr[43792]= 1537312353;
assign addr[43793]= 1563771613;
assign addr[43794]= 1589734894;
assign addr[43795]= 1615193959;
assign addr[43796]= 1640140734;
assign addr[43797]= 1664567307;
assign addr[43798]= 1688465931;
assign addr[43799]= 1711829025;
assign addr[43800]= 1734649179;
assign addr[43801]= 1756919156;
assign addr[43802]= 1778631892;
assign addr[43803]= 1799780501;
assign addr[43804]= 1820358275;
assign addr[43805]= 1840358687;
assign addr[43806]= 1859775393;
assign addr[43807]= 1878602237;
assign addr[43808]= 1896833245;
assign addr[43809]= 1914462636;
assign addr[43810]= 1931484818;
assign addr[43811]= 1947894393;
assign addr[43812]= 1963686155;
assign addr[43813]= 1978855097;
assign addr[43814]= 1993396407;
assign addr[43815]= 2007305472;
assign addr[43816]= 2020577882;
assign addr[43817]= 2033209426;
assign addr[43818]= 2045196100;
assign addr[43819]= 2056534099;
assign addr[43820]= 2067219829;
assign addr[43821]= 2077249901;
assign addr[43822]= 2086621133;
assign addr[43823]= 2095330553;
assign addr[43824]= 2103375398;
assign addr[43825]= 2110753117;
assign addr[43826]= 2117461370;
assign addr[43827]= 2123498030;
assign addr[43828]= 2128861181;
assign addr[43829]= 2133549123;
assign addr[43830]= 2137560369;
assign addr[43831]= 2140893646;
assign addr[43832]= 2143547897;
assign addr[43833]= 2145522281;
assign addr[43834]= 2146816171;
assign addr[43835]= 2147429158;
assign addr[43836]= 2147361045;
assign addr[43837]= 2146611856;
assign addr[43838]= 2145181827;
assign addr[43839]= 2143071413;
assign addr[43840]= 2140281282;
assign addr[43841]= 2136812319;
assign addr[43842]= 2132665626;
assign addr[43843]= 2127842516;
assign addr[43844]= 2122344521;
assign addr[43845]= 2116173382;
assign addr[43846]= 2109331059;
assign addr[43847]= 2101819720;
assign addr[43848]= 2093641749;
assign addr[43849]= 2084799740;
assign addr[43850]= 2075296495;
assign addr[43851]= 2065135031;
assign addr[43852]= 2054318569;
assign addr[43853]= 2042850540;
assign addr[43854]= 2030734582;
assign addr[43855]= 2017974537;
assign addr[43856]= 2004574453;
assign addr[43857]= 1990538579;
assign addr[43858]= 1975871368;
assign addr[43859]= 1960577471;
assign addr[43860]= 1944661739;
assign addr[43861]= 1928129220;
assign addr[43862]= 1910985158;
assign addr[43863]= 1893234990;
assign addr[43864]= 1874884346;
assign addr[43865]= 1855939047;
assign addr[43866]= 1836405100;
assign addr[43867]= 1816288703;
assign addr[43868]= 1795596234;
assign addr[43869]= 1774334257;
assign addr[43870]= 1752509516;
assign addr[43871]= 1730128933;
assign addr[43872]= 1707199606;
assign addr[43873]= 1683728808;
assign addr[43874]= 1659723983;
assign addr[43875]= 1635192744;
assign addr[43876]= 1610142873;
assign addr[43877]= 1584582314;
assign addr[43878]= 1558519173;
assign addr[43879]= 1531961719;
assign addr[43880]= 1504918373;
assign addr[43881]= 1477397714;
assign addr[43882]= 1449408469;
assign addr[43883]= 1420959516;
assign addr[43884]= 1392059879;
assign addr[43885]= 1362718723;
assign addr[43886]= 1332945355;
assign addr[43887]= 1302749217;
assign addr[43888]= 1272139887;
assign addr[43889]= 1241127074;
assign addr[43890]= 1209720613;
assign addr[43891]= 1177930466;
assign addr[43892]= 1145766716;
assign addr[43893]= 1113239564;
assign addr[43894]= 1080359326;
assign addr[43895]= 1047136432;
assign addr[43896]= 1013581418;
assign addr[43897]= 979704927;
assign addr[43898]= 945517704;
assign addr[43899]= 911030591;
assign addr[43900]= 876254528;
assign addr[43901]= 841200544;
assign addr[43902]= 805879757;
assign addr[43903]= 770303369;
assign addr[43904]= 734482665;
assign addr[43905]= 698429006;
assign addr[43906]= 662153826;
assign addr[43907]= 625668632;
assign addr[43908]= 588984994;
assign addr[43909]= 552114549;
assign addr[43910]= 515068990;
assign addr[43911]= 477860067;
assign addr[43912]= 440499581;
assign addr[43913]= 402999383;
assign addr[43914]= 365371365;
assign addr[43915]= 327627463;
assign addr[43916]= 289779648;
assign addr[43917]= 251839923;
assign addr[43918]= 213820322;
assign addr[43919]= 175732905;
assign addr[43920]= 137589750;
assign addr[43921]= 99402956;
assign addr[43922]= 61184634;
assign addr[43923]= 22946906;
assign addr[43924]= -15298099;
assign addr[43925]= -53538253;
assign addr[43926]= -91761426;
assign addr[43927]= -129955495;
assign addr[43928]= -168108346;
assign addr[43929]= -206207878;
assign addr[43930]= -244242007;
assign addr[43931]= -282198671;
assign addr[43932]= -320065829;
assign addr[43933]= -357831473;
assign addr[43934]= -395483624;
assign addr[43935]= -433010339;
assign addr[43936]= -470399716;
assign addr[43937]= -507639898;
assign addr[43938]= -544719071;
assign addr[43939]= -581625477;
assign addr[43940]= -618347408;
assign addr[43941]= -654873219;
assign addr[43942]= -691191324;
assign addr[43943]= -727290205;
assign addr[43944]= -763158411;
assign addr[43945]= -798784567;
assign addr[43946]= -834157373;
assign addr[43947]= -869265610;
assign addr[43948]= -904098143;
assign addr[43949]= -938643924;
assign addr[43950]= -972891995;
assign addr[43951]= -1006831495;
assign addr[43952]= -1040451659;
assign addr[43953]= -1073741824;
assign addr[43954]= -1106691431;
assign addr[43955]= -1139290029;
assign addr[43956]= -1171527280;
assign addr[43957]= -1203392958;
assign addr[43958]= -1234876957;
assign addr[43959]= -1265969291;
assign addr[43960]= -1296660098;
assign addr[43961]= -1326939644;
assign addr[43962]= -1356798326;
assign addr[43963]= -1386226674;
assign addr[43964]= -1415215352;
assign addr[43965]= -1443755168;
assign addr[43966]= -1471837070;
assign addr[43967]= -1499452149;
assign addr[43968]= -1526591649;
assign addr[43969]= -1553246960;
assign addr[43970]= -1579409630;
assign addr[43971]= -1605071359;
assign addr[43972]= -1630224009;
assign addr[43973]= -1654859602;
assign addr[43974]= -1678970324;
assign addr[43975]= -1702548529;
assign addr[43976]= -1725586737;
assign addr[43977]= -1748077642;
assign addr[43978]= -1770014111;
assign addr[43979]= -1791389186;
assign addr[43980]= -1812196087;
assign addr[43981]= -1832428215;
assign addr[43982]= -1852079154;
assign addr[43983]= -1871142669;
assign addr[43984]= -1889612716;
assign addr[43985]= -1907483436;
assign addr[43986]= -1924749160;
assign addr[43987]= -1941404413;
assign addr[43988]= -1957443913;
assign addr[43989]= -1972862571;
assign addr[43990]= -1987655498;
assign addr[43991]= -2001818002;
assign addr[43992]= -2015345591;
assign addr[43993]= -2028233973;
assign addr[43994]= -2040479063;
assign addr[43995]= -2052076975;
assign addr[43996]= -2063024031;
assign addr[43997]= -2073316760;
assign addr[43998]= -2082951896;
assign addr[43999]= -2091926384;
assign addr[44000]= -2100237377;
assign addr[44001]= -2107882239;
assign addr[44002]= -2114858546;
assign addr[44003]= -2121164085;
assign addr[44004]= -2126796855;
assign addr[44005]= -2131755071;
assign addr[44006]= -2136037160;
assign addr[44007]= -2139641764;
assign addr[44008]= -2142567738;
assign addr[44009]= -2144814157;
assign addr[44010]= -2146380306;
assign addr[44011]= -2147265689;
assign addr[44012]= -2147470025;
assign addr[44013]= -2146993250;
assign addr[44014]= -2145835515;
assign addr[44015]= -2143997187;
assign addr[44016]= -2141478848;
assign addr[44017]= -2138281298;
assign addr[44018]= -2134405552;
assign addr[44019]= -2129852837;
assign addr[44020]= -2124624598;
assign addr[44021]= -2118722494;
assign addr[44022]= -2112148396;
assign addr[44023]= -2104904390;
assign addr[44024]= -2096992772;
assign addr[44025]= -2088416053;
assign addr[44026]= -2079176953;
assign addr[44027]= -2069278401;
assign addr[44028]= -2058723538;
assign addr[44029]= -2047515711;
assign addr[44030]= -2035658475;
assign addr[44031]= -2023155591;
assign addr[44032]= -2010011024;
assign addr[44033]= -1996228943;
assign addr[44034]= -1981813720;
assign addr[44035]= -1966769926;
assign addr[44036]= -1951102334;
assign addr[44037]= -1934815911;
assign addr[44038]= -1917915825;
assign addr[44039]= -1900407434;
assign addr[44040]= -1882296293;
assign addr[44041]= -1863588145;
assign addr[44042]= -1844288924;
assign addr[44043]= -1824404752;
assign addr[44044]= -1803941934;
assign addr[44045]= -1782906961;
assign addr[44046]= -1761306505;
assign addr[44047]= -1739147417;
assign addr[44048]= -1716436725;
assign addr[44049]= -1693181631;
assign addr[44050]= -1669389513;
assign addr[44051]= -1645067915;
assign addr[44052]= -1620224553;
assign addr[44053]= -1594867305;
assign addr[44054]= -1569004214;
assign addr[44055]= -1542643483;
assign addr[44056]= -1515793473;
assign addr[44057]= -1488462700;
assign addr[44058]= -1460659832;
assign addr[44059]= -1432393688;
assign addr[44060]= -1403673233;
assign addr[44061]= -1374507575;
assign addr[44062]= -1344905966;
assign addr[44063]= -1314877795;
assign addr[44064]= -1284432584;
assign addr[44065]= -1253579991;
assign addr[44066]= -1222329801;
assign addr[44067]= -1190691925;
assign addr[44068]= -1158676398;
assign addr[44069]= -1126293375;
assign addr[44070]= -1093553126;
assign addr[44071]= -1060466036;
assign addr[44072]= -1027042599;
assign addr[44073]= -993293415;
assign addr[44074]= -959229189;
assign addr[44075]= -924860725;
assign addr[44076]= -890198924;
assign addr[44077]= -855254778;
assign addr[44078]= -820039373;
assign addr[44079]= -784563876;
assign addr[44080]= -748839539;
assign addr[44081]= -712877694;
assign addr[44082]= -676689746;
assign addr[44083]= -640287172;
assign addr[44084]= -603681519;
assign addr[44085]= -566884397;
assign addr[44086]= -529907477;
assign addr[44087]= -492762486;
assign addr[44088]= -455461206;
assign addr[44089]= -418015468;
assign addr[44090]= -380437148;
assign addr[44091]= -342738165;
assign addr[44092]= -304930476;
assign addr[44093]= -267026072;
assign addr[44094]= -229036977;
assign addr[44095]= -190975237;
assign addr[44096]= -152852926;
assign addr[44097]= -114682135;
assign addr[44098]= -76474970;
assign addr[44099]= -38243550;
assign addr[44100]= 0;
assign addr[44101]= 38243550;
assign addr[44102]= 76474970;
assign addr[44103]= 114682135;
assign addr[44104]= 152852926;
assign addr[44105]= 190975237;
assign addr[44106]= 229036977;
assign addr[44107]= 267026072;
assign addr[44108]= 304930476;
assign addr[44109]= 342738165;
assign addr[44110]= 380437148;
assign addr[44111]= 418015468;
assign addr[44112]= 455461206;
assign addr[44113]= 492762486;
assign addr[44114]= 529907477;
assign addr[44115]= 566884397;
assign addr[44116]= 603681519;
assign addr[44117]= 640287172;
assign addr[44118]= 676689746;
assign addr[44119]= 712877694;
assign addr[44120]= 748839539;
assign addr[44121]= 784563876;
assign addr[44122]= 820039373;
assign addr[44123]= 855254778;
assign addr[44124]= 890198924;
assign addr[44125]= 924860725;
assign addr[44126]= 959229189;
assign addr[44127]= 993293415;
assign addr[44128]= 1027042599;
assign addr[44129]= 1060466036;
assign addr[44130]= 1093553126;
assign addr[44131]= 1126293375;
assign addr[44132]= 1158676398;
assign addr[44133]= 1190691925;
assign addr[44134]= 1222329801;
assign addr[44135]= 1253579991;
assign addr[44136]= 1284432584;
assign addr[44137]= 1314877795;
assign addr[44138]= 1344905966;
assign addr[44139]= 1374507575;
assign addr[44140]= 1403673233;
assign addr[44141]= 1432393688;
assign addr[44142]= 1460659832;
assign addr[44143]= 1488462700;
assign addr[44144]= 1515793473;
assign addr[44145]= 1542643483;
assign addr[44146]= 1569004214;
assign addr[44147]= 1594867305;
assign addr[44148]= 1620224553;
assign addr[44149]= 1645067915;
assign addr[44150]= 1669389513;
assign addr[44151]= 1693181631;
assign addr[44152]= 1716436725;
assign addr[44153]= 1739147417;
assign addr[44154]= 1761306505;
assign addr[44155]= 1782906961;
assign addr[44156]= 1803941934;
assign addr[44157]= 1824404752;
assign addr[44158]= 1844288924;
assign addr[44159]= 1863588145;
assign addr[44160]= 1882296293;
assign addr[44161]= 1900407434;
assign addr[44162]= 1917915825;
assign addr[44163]= 1934815911;
assign addr[44164]= 1951102334;
assign addr[44165]= 1966769926;
assign addr[44166]= 1981813720;
assign addr[44167]= 1996228943;
assign addr[44168]= 2010011024;
assign addr[44169]= 2023155591;
assign addr[44170]= 2035658475;
assign addr[44171]= 2047515711;
assign addr[44172]= 2058723538;
assign addr[44173]= 2069278401;
assign addr[44174]= 2079176953;
assign addr[44175]= 2088416053;
assign addr[44176]= 2096992772;
assign addr[44177]= 2104904390;
assign addr[44178]= 2112148396;
assign addr[44179]= 2118722494;
assign addr[44180]= 2124624598;
assign addr[44181]= 2129852837;
assign addr[44182]= 2134405552;
assign addr[44183]= 2138281298;
assign addr[44184]= 2141478848;
assign addr[44185]= 2143997187;
assign addr[44186]= 2145835515;
assign addr[44187]= 2146993250;
assign addr[44188]= 2147470025;
assign addr[44189]= 2147265689;
assign addr[44190]= 2146380306;
assign addr[44191]= 2144814157;
assign addr[44192]= 2142567738;
assign addr[44193]= 2139641764;
assign addr[44194]= 2136037160;
assign addr[44195]= 2131755071;
assign addr[44196]= 2126796855;
assign addr[44197]= 2121164085;
assign addr[44198]= 2114858546;
assign addr[44199]= 2107882239;
assign addr[44200]= 2100237377;
assign addr[44201]= 2091926384;
assign addr[44202]= 2082951896;
assign addr[44203]= 2073316760;
assign addr[44204]= 2063024031;
assign addr[44205]= 2052076975;
assign addr[44206]= 2040479063;
assign addr[44207]= 2028233973;
assign addr[44208]= 2015345591;
assign addr[44209]= 2001818002;
assign addr[44210]= 1987655498;
assign addr[44211]= 1972862571;
assign addr[44212]= 1957443913;
assign addr[44213]= 1941404413;
assign addr[44214]= 1924749160;
assign addr[44215]= 1907483436;
assign addr[44216]= 1889612716;
assign addr[44217]= 1871142669;
assign addr[44218]= 1852079154;
assign addr[44219]= 1832428215;
assign addr[44220]= 1812196087;
assign addr[44221]= 1791389186;
assign addr[44222]= 1770014111;
assign addr[44223]= 1748077642;
assign addr[44224]= 1725586737;
assign addr[44225]= 1702548529;
assign addr[44226]= 1678970324;
assign addr[44227]= 1654859602;
assign addr[44228]= 1630224009;
assign addr[44229]= 1605071359;
assign addr[44230]= 1579409630;
assign addr[44231]= 1553246960;
assign addr[44232]= 1526591649;
assign addr[44233]= 1499452149;
assign addr[44234]= 1471837070;
assign addr[44235]= 1443755168;
assign addr[44236]= 1415215352;
assign addr[44237]= 1386226674;
assign addr[44238]= 1356798326;
assign addr[44239]= 1326939644;
assign addr[44240]= 1296660098;
assign addr[44241]= 1265969291;
assign addr[44242]= 1234876957;
assign addr[44243]= 1203392958;
assign addr[44244]= 1171527280;
assign addr[44245]= 1139290029;
assign addr[44246]= 1106691431;
assign addr[44247]= 1073741824;
assign addr[44248]= 1040451659;
assign addr[44249]= 1006831495;
assign addr[44250]= 972891995;
assign addr[44251]= 938643924;
assign addr[44252]= 904098143;
assign addr[44253]= 869265610;
assign addr[44254]= 834157373;
assign addr[44255]= 798784567;
assign addr[44256]= 763158411;
assign addr[44257]= 727290205;
assign addr[44258]= 691191324;
assign addr[44259]= 654873219;
assign addr[44260]= 618347408;
assign addr[44261]= 581625477;
assign addr[44262]= 544719071;
assign addr[44263]= 507639898;
assign addr[44264]= 470399716;
assign addr[44265]= 433010339;
assign addr[44266]= 395483624;
assign addr[44267]= 357831473;
assign addr[44268]= 320065829;
assign addr[44269]= 282198671;
assign addr[44270]= 244242007;
assign addr[44271]= 206207878;
assign addr[44272]= 168108346;
assign addr[44273]= 129955495;
assign addr[44274]= 91761426;
assign addr[44275]= 53538253;
assign addr[44276]= 15298099;
assign addr[44277]= -22946906;
assign addr[44278]= -61184634;
assign addr[44279]= -99402956;
assign addr[44280]= -137589750;
assign addr[44281]= -175732905;
assign addr[44282]= -213820322;
assign addr[44283]= -251839923;
assign addr[44284]= -289779648;
assign addr[44285]= -327627463;
assign addr[44286]= -365371365;
assign addr[44287]= -402999383;
assign addr[44288]= -440499581;
assign addr[44289]= -477860067;
assign addr[44290]= -515068990;
assign addr[44291]= -552114549;
assign addr[44292]= -588984994;
assign addr[44293]= -625668632;
assign addr[44294]= -662153826;
assign addr[44295]= -698429006;
assign addr[44296]= -734482665;
assign addr[44297]= -770303369;
assign addr[44298]= -805879757;
assign addr[44299]= -841200544;
assign addr[44300]= -876254528;
assign addr[44301]= -911030591;
assign addr[44302]= -945517704;
assign addr[44303]= -979704927;
assign addr[44304]= -1013581418;
assign addr[44305]= -1047136432;
assign addr[44306]= -1080359326;
assign addr[44307]= -1113239564;
assign addr[44308]= -1145766716;
assign addr[44309]= -1177930466;
assign addr[44310]= -1209720613;
assign addr[44311]= -1241127074;
assign addr[44312]= -1272139887;
assign addr[44313]= -1302749217;
assign addr[44314]= -1332945355;
assign addr[44315]= -1362718723;
assign addr[44316]= -1392059879;
assign addr[44317]= -1420959516;
assign addr[44318]= -1449408469;
assign addr[44319]= -1477397714;
assign addr[44320]= -1504918373;
assign addr[44321]= -1531961719;
assign addr[44322]= -1558519173;
assign addr[44323]= -1584582314;
assign addr[44324]= -1610142873;
assign addr[44325]= -1635192744;
assign addr[44326]= -1659723983;
assign addr[44327]= -1683728808;
assign addr[44328]= -1707199606;
assign addr[44329]= -1730128933;
assign addr[44330]= -1752509516;
assign addr[44331]= -1774334257;
assign addr[44332]= -1795596234;
assign addr[44333]= -1816288703;
assign addr[44334]= -1836405100;
assign addr[44335]= -1855939047;
assign addr[44336]= -1874884346;
assign addr[44337]= -1893234990;
assign addr[44338]= -1910985158;
assign addr[44339]= -1928129220;
assign addr[44340]= -1944661739;
assign addr[44341]= -1960577471;
assign addr[44342]= -1975871368;
assign addr[44343]= -1990538579;
assign addr[44344]= -2004574453;
assign addr[44345]= -2017974537;
assign addr[44346]= -2030734582;
assign addr[44347]= -2042850540;
assign addr[44348]= -2054318569;
assign addr[44349]= -2065135031;
assign addr[44350]= -2075296495;
assign addr[44351]= -2084799740;
assign addr[44352]= -2093641749;
assign addr[44353]= -2101819720;
assign addr[44354]= -2109331059;
assign addr[44355]= -2116173382;
assign addr[44356]= -2122344521;
assign addr[44357]= -2127842516;
assign addr[44358]= -2132665626;
assign addr[44359]= -2136812319;
assign addr[44360]= -2140281282;
assign addr[44361]= -2143071413;
assign addr[44362]= -2145181827;
assign addr[44363]= -2146611856;
assign addr[44364]= -2147361045;
assign addr[44365]= -2147429158;
assign addr[44366]= -2146816171;
assign addr[44367]= -2145522281;
assign addr[44368]= -2143547897;
assign addr[44369]= -2140893646;
assign addr[44370]= -2137560369;
assign addr[44371]= -2133549123;
assign addr[44372]= -2128861181;
assign addr[44373]= -2123498030;
assign addr[44374]= -2117461370;
assign addr[44375]= -2110753117;
assign addr[44376]= -2103375398;
assign addr[44377]= -2095330553;
assign addr[44378]= -2086621133;
assign addr[44379]= -2077249901;
assign addr[44380]= -2067219829;
assign addr[44381]= -2056534099;
assign addr[44382]= -2045196100;
assign addr[44383]= -2033209426;
assign addr[44384]= -2020577882;
assign addr[44385]= -2007305472;
assign addr[44386]= -1993396407;
assign addr[44387]= -1978855097;
assign addr[44388]= -1963686155;
assign addr[44389]= -1947894393;
assign addr[44390]= -1931484818;
assign addr[44391]= -1914462636;
assign addr[44392]= -1896833245;
assign addr[44393]= -1878602237;
assign addr[44394]= -1859775393;
assign addr[44395]= -1840358687;
assign addr[44396]= -1820358275;
assign addr[44397]= -1799780501;
assign addr[44398]= -1778631892;
assign addr[44399]= -1756919156;
assign addr[44400]= -1734649179;
assign addr[44401]= -1711829025;
assign addr[44402]= -1688465931;
assign addr[44403]= -1664567307;
assign addr[44404]= -1640140734;
assign addr[44405]= -1615193959;
assign addr[44406]= -1589734894;
assign addr[44407]= -1563771613;
assign addr[44408]= -1537312353;
assign addr[44409]= -1510365504;
assign addr[44410]= -1482939614;
assign addr[44411]= -1455043381;
assign addr[44412]= -1426685652;
assign addr[44413]= -1397875423;
assign addr[44414]= -1368621831;
assign addr[44415]= -1338934154;
assign addr[44416]= -1308821808;
assign addr[44417]= -1278294345;
assign addr[44418]= -1247361445;
assign addr[44419]= -1216032921;
assign addr[44420]= -1184318708;
assign addr[44421]= -1152228866;
assign addr[44422]= -1119773573;
assign addr[44423]= -1086963121;
assign addr[44424]= -1053807919;
assign addr[44425]= -1020318481;
assign addr[44426]= -986505429;
assign addr[44427]= -952379488;
assign addr[44428]= -917951481;
assign addr[44429]= -883232329;
assign addr[44430]= -848233042;
assign addr[44431]= -812964722;
assign addr[44432]= -777438554;
assign addr[44433]= -741665807;
assign addr[44434]= -705657826;
assign addr[44435]= -669426032;
assign addr[44436]= -632981917;
assign addr[44437]= -596337040;
assign addr[44438]= -559503022;
assign addr[44439]= -522491548;
assign addr[44440]= -485314355;
assign addr[44441]= -447983235;
assign addr[44442]= -410510029;
assign addr[44443]= -372906622;
assign addr[44444]= -335184940;
assign addr[44445]= -297356948;
assign addr[44446]= -259434643;
assign addr[44447]= -221430054;
assign addr[44448]= -183355234;
assign addr[44449]= -145222259;
assign addr[44450]= -107043224;
assign addr[44451]= -68830239;
assign addr[44452]= -30595422;
assign addr[44453]= 7649098;
assign addr[44454]= 45891193;
assign addr[44455]= 84118732;
assign addr[44456]= 122319591;
assign addr[44457]= 160481654;
assign addr[44458]= 198592817;
assign addr[44459]= 236640993;
assign addr[44460]= 274614114;
assign addr[44461]= 312500135;
assign addr[44462]= 350287041;
assign addr[44463]= 387962847;
assign addr[44464]= 425515602;
assign addr[44465]= 462933398;
assign addr[44466]= 500204365;
assign addr[44467]= 537316682;
assign addr[44468]= 574258580;
assign addr[44469]= 611018340;
assign addr[44470]= 647584304;
assign addr[44471]= 683944874;
assign addr[44472]= 720088517;
assign addr[44473]= 756003771;
assign addr[44474]= 791679244;
assign addr[44475]= 827103620;
assign addr[44476]= 862265664;
assign addr[44477]= 897154224;
assign addr[44478]= 931758235;
assign addr[44479]= 966066720;
assign addr[44480]= 1000068799;
assign addr[44481]= 1033753687;
assign addr[44482]= 1067110699;
assign addr[44483]= 1100129257;
assign addr[44484]= 1132798888;
assign addr[44485]= 1165109230;
assign addr[44486]= 1197050035;
assign addr[44487]= 1228611172;
assign addr[44488]= 1259782632;
assign addr[44489]= 1290554528;
assign addr[44490]= 1320917099;
assign addr[44491]= 1350860716;
assign addr[44492]= 1380375881;
assign addr[44493]= 1409453233;
assign addr[44494]= 1438083551;
assign addr[44495]= 1466257752;
assign addr[44496]= 1493966902;
assign addr[44497]= 1521202211;
assign addr[44498]= 1547955041;
assign addr[44499]= 1574216908;
assign addr[44500]= 1599979481;
assign addr[44501]= 1625234591;
assign addr[44502]= 1649974225;
assign addr[44503]= 1674190539;
assign addr[44504]= 1697875851;
assign addr[44505]= 1721022648;
assign addr[44506]= 1743623590;
assign addr[44507]= 1765671509;
assign addr[44508]= 1787159411;
assign addr[44509]= 1808080480;
assign addr[44510]= 1828428082;
assign addr[44511]= 1848195763;
assign addr[44512]= 1867377253;
assign addr[44513]= 1885966468;
assign addr[44514]= 1903957513;
assign addr[44515]= 1921344681;
assign addr[44516]= 1938122457;
assign addr[44517]= 1954285520;
assign addr[44518]= 1969828744;
assign addr[44519]= 1984747199;
assign addr[44520]= 1999036154;
assign addr[44521]= 2012691075;
assign addr[44522]= 2025707632;
assign addr[44523]= 2038081698;
assign addr[44524]= 2049809346;
assign addr[44525]= 2060886858;
assign addr[44526]= 2071310720;
assign addr[44527]= 2081077626;
assign addr[44528]= 2090184478;
assign addr[44529]= 2098628387;
assign addr[44530]= 2106406677;
assign addr[44531]= 2113516878;
assign addr[44532]= 2119956737;
assign addr[44533]= 2125724211;
assign addr[44534]= 2130817471;
assign addr[44535]= 2135234901;
assign addr[44536]= 2138975100;
assign addr[44537]= 2142036881;
assign addr[44538]= 2144419275;
assign addr[44539]= 2146121524;
assign addr[44540]= 2147143090;
assign addr[44541]= 2147483648;
assign addr[44542]= 2147143090;
assign addr[44543]= 2146121524;
assign addr[44544]= 2144419275;
assign addr[44545]= 2142036881;
assign addr[44546]= 2138975100;
assign addr[44547]= 2135234901;
assign addr[44548]= 2130817471;
assign addr[44549]= 2125724211;
assign addr[44550]= 2119956737;
assign addr[44551]= 2113516878;
assign addr[44552]= 2106406677;
assign addr[44553]= 2098628387;
assign addr[44554]= 2090184478;
assign addr[44555]= 2081077626;
assign addr[44556]= 2071310720;
assign addr[44557]= 2060886858;
assign addr[44558]= 2049809346;
assign addr[44559]= 2038081698;
assign addr[44560]= 2025707632;
assign addr[44561]= 2012691075;
assign addr[44562]= 1999036154;
assign addr[44563]= 1984747199;
assign addr[44564]= 1969828744;
assign addr[44565]= 1954285520;
assign addr[44566]= 1938122457;
assign addr[44567]= 1921344681;
assign addr[44568]= 1903957513;
assign addr[44569]= 1885966468;
assign addr[44570]= 1867377253;
assign addr[44571]= 1848195763;
assign addr[44572]= 1828428082;
assign addr[44573]= 1808080480;
assign addr[44574]= 1787159411;
assign addr[44575]= 1765671509;
assign addr[44576]= 1743623590;
assign addr[44577]= 1721022648;
assign addr[44578]= 1697875851;
assign addr[44579]= 1674190539;
assign addr[44580]= 1649974225;
assign addr[44581]= 1625234591;
assign addr[44582]= 1599979481;
assign addr[44583]= 1574216908;
assign addr[44584]= 1547955041;
assign addr[44585]= 1521202211;
assign addr[44586]= 1493966902;
assign addr[44587]= 1466257752;
assign addr[44588]= 1438083551;
assign addr[44589]= 1409453233;
assign addr[44590]= 1380375881;
assign addr[44591]= 1350860716;
assign addr[44592]= 1320917099;
assign addr[44593]= 1290554528;
assign addr[44594]= 1259782632;
assign addr[44595]= 1228611172;
assign addr[44596]= 1197050035;
assign addr[44597]= 1165109230;
assign addr[44598]= 1132798888;
assign addr[44599]= 1100129257;
assign addr[44600]= 1067110699;
assign addr[44601]= 1033753687;
assign addr[44602]= 1000068799;
assign addr[44603]= 966066720;
assign addr[44604]= 931758235;
assign addr[44605]= 897154224;
assign addr[44606]= 862265664;
assign addr[44607]= 827103620;
assign addr[44608]= 791679244;
assign addr[44609]= 756003771;
assign addr[44610]= 720088517;
assign addr[44611]= 683944874;
assign addr[44612]= 647584304;
assign addr[44613]= 611018340;
assign addr[44614]= 574258580;
assign addr[44615]= 537316682;
assign addr[44616]= 500204365;
assign addr[44617]= 462933398;
assign addr[44618]= 425515602;
assign addr[44619]= 387962847;
assign addr[44620]= 350287041;
assign addr[44621]= 312500135;
assign addr[44622]= 274614114;
assign addr[44623]= 236640993;
assign addr[44624]= 198592817;
assign addr[44625]= 160481654;
assign addr[44626]= 122319591;
assign addr[44627]= 84118732;
assign addr[44628]= 45891193;
assign addr[44629]= 7649098;
assign addr[44630]= -30595422;
assign addr[44631]= -68830239;
assign addr[44632]= -107043224;
assign addr[44633]= -145222259;
assign addr[44634]= -183355234;
assign addr[44635]= -221430054;
assign addr[44636]= -259434643;
assign addr[44637]= -297356948;
assign addr[44638]= -335184940;
assign addr[44639]= -372906622;
assign addr[44640]= -410510029;
assign addr[44641]= -447983235;
assign addr[44642]= -485314355;
assign addr[44643]= -522491548;
assign addr[44644]= -559503022;
assign addr[44645]= -596337040;
assign addr[44646]= -632981917;
assign addr[44647]= -669426032;
assign addr[44648]= -705657826;
assign addr[44649]= -741665807;
assign addr[44650]= -777438554;
assign addr[44651]= -812964722;
assign addr[44652]= -848233042;
assign addr[44653]= -883232329;
assign addr[44654]= -917951481;
assign addr[44655]= -952379488;
assign addr[44656]= -986505429;
assign addr[44657]= -1020318481;
assign addr[44658]= -1053807919;
assign addr[44659]= -1086963121;
assign addr[44660]= -1119773573;
assign addr[44661]= -1152228866;
assign addr[44662]= -1184318708;
assign addr[44663]= -1216032921;
assign addr[44664]= -1247361445;
assign addr[44665]= -1278294345;
assign addr[44666]= -1308821808;
assign addr[44667]= -1338934154;
assign addr[44668]= -1368621831;
assign addr[44669]= -1397875423;
assign addr[44670]= -1426685652;
assign addr[44671]= -1455043381;
assign addr[44672]= -1482939614;
assign addr[44673]= -1510365504;
assign addr[44674]= -1537312353;
assign addr[44675]= -1563771613;
assign addr[44676]= -1589734894;
assign addr[44677]= -1615193959;
assign addr[44678]= -1640140734;
assign addr[44679]= -1664567307;
assign addr[44680]= -1688465931;
assign addr[44681]= -1711829025;
assign addr[44682]= -1734649179;
assign addr[44683]= -1756919156;
assign addr[44684]= -1778631892;
assign addr[44685]= -1799780501;
assign addr[44686]= -1820358275;
assign addr[44687]= -1840358687;
assign addr[44688]= -1859775393;
assign addr[44689]= -1878602237;
assign addr[44690]= -1896833245;
assign addr[44691]= -1914462636;
assign addr[44692]= -1931484818;
assign addr[44693]= -1947894393;
assign addr[44694]= -1963686155;
assign addr[44695]= -1978855097;
assign addr[44696]= -1993396407;
assign addr[44697]= -2007305472;
assign addr[44698]= -2020577882;
assign addr[44699]= -2033209426;
assign addr[44700]= -2045196100;
assign addr[44701]= -2056534099;
assign addr[44702]= -2067219829;
assign addr[44703]= -2077249901;
assign addr[44704]= -2086621133;
assign addr[44705]= -2095330553;
assign addr[44706]= -2103375398;
assign addr[44707]= -2110753117;
assign addr[44708]= -2117461370;
assign addr[44709]= -2123498030;
assign addr[44710]= -2128861181;
assign addr[44711]= -2133549123;
assign addr[44712]= -2137560369;
assign addr[44713]= -2140893646;
assign addr[44714]= -2143547897;
assign addr[44715]= -2145522281;
assign addr[44716]= -2146816171;
assign addr[44717]= -2147429158;
assign addr[44718]= -2147361045;
assign addr[44719]= -2146611856;
assign addr[44720]= -2145181827;
assign addr[44721]= -2143071413;
assign addr[44722]= -2140281282;
assign addr[44723]= -2136812319;
assign addr[44724]= -2132665626;
assign addr[44725]= -2127842516;
assign addr[44726]= -2122344521;
assign addr[44727]= -2116173382;
assign addr[44728]= -2109331059;
assign addr[44729]= -2101819720;
assign addr[44730]= -2093641749;
assign addr[44731]= -2084799740;
assign addr[44732]= -2075296495;
assign addr[44733]= -2065135031;
assign addr[44734]= -2054318569;
assign addr[44735]= -2042850540;
assign addr[44736]= -2030734582;
assign addr[44737]= -2017974537;
assign addr[44738]= -2004574453;
assign addr[44739]= -1990538579;
assign addr[44740]= -1975871368;
assign addr[44741]= -1960577471;
assign addr[44742]= -1944661739;
assign addr[44743]= -1928129220;
assign addr[44744]= -1910985158;
assign addr[44745]= -1893234990;
assign addr[44746]= -1874884346;
assign addr[44747]= -1855939047;
assign addr[44748]= -1836405100;
assign addr[44749]= -1816288703;
assign addr[44750]= -1795596234;
assign addr[44751]= -1774334257;
assign addr[44752]= -1752509516;
assign addr[44753]= -1730128933;
assign addr[44754]= -1707199606;
assign addr[44755]= -1683728808;
assign addr[44756]= -1659723983;
assign addr[44757]= -1635192744;
assign addr[44758]= -1610142873;
assign addr[44759]= -1584582314;
assign addr[44760]= -1558519173;
assign addr[44761]= -1531961719;
assign addr[44762]= -1504918373;
assign addr[44763]= -1477397714;
assign addr[44764]= -1449408469;
assign addr[44765]= -1420959516;
assign addr[44766]= -1392059879;
assign addr[44767]= -1362718723;
assign addr[44768]= -1332945355;
assign addr[44769]= -1302749217;
assign addr[44770]= -1272139887;
assign addr[44771]= -1241127074;
assign addr[44772]= -1209720613;
assign addr[44773]= -1177930466;
assign addr[44774]= -1145766716;
assign addr[44775]= -1113239564;
assign addr[44776]= -1080359326;
assign addr[44777]= -1047136432;
assign addr[44778]= -1013581418;
assign addr[44779]= -979704927;
assign addr[44780]= -945517704;
assign addr[44781]= -911030591;
assign addr[44782]= -876254528;
assign addr[44783]= -841200544;
assign addr[44784]= -805879757;
assign addr[44785]= -770303369;
assign addr[44786]= -734482665;
assign addr[44787]= -698429006;
assign addr[44788]= -662153826;
assign addr[44789]= -625668632;
assign addr[44790]= -588984994;
assign addr[44791]= -552114549;
assign addr[44792]= -515068990;
assign addr[44793]= -477860067;
assign addr[44794]= -440499581;
assign addr[44795]= -402999383;
assign addr[44796]= -365371365;
assign addr[44797]= -327627463;
assign addr[44798]= -289779648;
assign addr[44799]= -251839923;
assign addr[44800]= -213820322;
assign addr[44801]= -175732905;
assign addr[44802]= -137589750;
assign addr[44803]= -99402956;
assign addr[44804]= -61184634;
assign addr[44805]= -22946906;
assign addr[44806]= 15298099;
assign addr[44807]= 53538253;
assign addr[44808]= 91761426;
assign addr[44809]= 129955495;
assign addr[44810]= 168108346;
assign addr[44811]= 206207878;
assign addr[44812]= 244242007;
assign addr[44813]= 282198671;
assign addr[44814]= 320065829;
assign addr[44815]= 357831473;
assign addr[44816]= 395483624;
assign addr[44817]= 433010339;
assign addr[44818]= 470399716;
assign addr[44819]= 507639898;
assign addr[44820]= 544719071;
assign addr[44821]= 581625477;
assign addr[44822]= 618347408;
assign addr[44823]= 654873219;
assign addr[44824]= 691191324;
assign addr[44825]= 727290205;
assign addr[44826]= 763158411;
assign addr[44827]= 798784567;
assign addr[44828]= 834157373;
assign addr[44829]= 869265610;
assign addr[44830]= 904098143;
assign addr[44831]= 938643924;
assign addr[44832]= 972891995;
assign addr[44833]= 1006831495;
assign addr[44834]= 1040451659;
assign addr[44835]= 1073741824;
assign addr[44836]= 1106691431;
assign addr[44837]= 1139290029;
assign addr[44838]= 1171527280;
assign addr[44839]= 1203392958;
assign addr[44840]= 1234876957;
assign addr[44841]= 1265969291;
assign addr[44842]= 1296660098;
assign addr[44843]= 1326939644;
assign addr[44844]= 1356798326;
assign addr[44845]= 1386226674;
assign addr[44846]= 1415215352;
assign addr[44847]= 1443755168;
assign addr[44848]= 1471837070;
assign addr[44849]= 1499452149;
assign addr[44850]= 1526591649;
assign addr[44851]= 1553246960;
assign addr[44852]= 1579409630;
assign addr[44853]= 1605071359;
assign addr[44854]= 1630224009;
assign addr[44855]= 1654859602;
assign addr[44856]= 1678970324;
assign addr[44857]= 1702548529;
assign addr[44858]= 1725586737;
assign addr[44859]= 1748077642;
assign addr[44860]= 1770014111;
assign addr[44861]= 1791389186;
assign addr[44862]= 1812196087;
assign addr[44863]= 1832428215;
assign addr[44864]= 1852079154;
assign addr[44865]= 1871142669;
assign addr[44866]= 1889612716;
assign addr[44867]= 1907483436;
assign addr[44868]= 1924749160;
assign addr[44869]= 1941404413;
assign addr[44870]= 1957443913;
assign addr[44871]= 1972862571;
assign addr[44872]= 1987655498;
assign addr[44873]= 2001818002;
assign addr[44874]= 2015345591;
assign addr[44875]= 2028233973;
assign addr[44876]= 2040479063;
assign addr[44877]= 2052076975;
assign addr[44878]= 2063024031;
assign addr[44879]= 2073316760;
assign addr[44880]= 2082951896;
assign addr[44881]= 2091926384;
assign addr[44882]= 2100237377;
assign addr[44883]= 2107882239;
assign addr[44884]= 2114858546;
assign addr[44885]= 2121164085;
assign addr[44886]= 2126796855;
assign addr[44887]= 2131755071;
assign addr[44888]= 2136037160;
assign addr[44889]= 2139641764;
assign addr[44890]= 2142567738;
assign addr[44891]= 2144814157;
assign addr[44892]= 2146380306;
assign addr[44893]= 2147265689;
assign addr[44894]= 2147470025;
assign addr[44895]= 2146993250;
assign addr[44896]= 2145835515;
assign addr[44897]= 2143997187;
assign addr[44898]= 2141478848;
assign addr[44899]= 2138281298;
assign addr[44900]= 2134405552;
assign addr[44901]= 2129852837;
assign addr[44902]= 2124624598;
assign addr[44903]= 2118722494;
assign addr[44904]= 2112148396;
assign addr[44905]= 2104904390;
assign addr[44906]= 2096992772;
assign addr[44907]= 2088416053;
assign addr[44908]= 2079176953;
assign addr[44909]= 2069278401;
assign addr[44910]= 2058723538;
assign addr[44911]= 2047515711;
assign addr[44912]= 2035658475;
assign addr[44913]= 2023155591;
assign addr[44914]= 2010011024;
assign addr[44915]= 1996228943;
assign addr[44916]= 1981813720;
assign addr[44917]= 1966769926;
assign addr[44918]= 1951102334;
assign addr[44919]= 1934815911;
assign addr[44920]= 1917915825;
assign addr[44921]= 1900407434;
assign addr[44922]= 1882296293;
assign addr[44923]= 1863588145;
assign addr[44924]= 1844288924;
assign addr[44925]= 1824404752;
assign addr[44926]= 1803941934;
assign addr[44927]= 1782906961;
assign addr[44928]= 1761306505;
assign addr[44929]= 1739147417;
assign addr[44930]= 1716436725;
assign addr[44931]= 1693181631;
assign addr[44932]= 1669389513;
assign addr[44933]= 1645067915;
assign addr[44934]= 1620224553;
assign addr[44935]= 1594867305;
assign addr[44936]= 1569004214;
assign addr[44937]= 1542643483;
assign addr[44938]= 1515793473;
assign addr[44939]= 1488462700;
assign addr[44940]= 1460659832;
assign addr[44941]= 1432393688;
assign addr[44942]= 1403673233;
assign addr[44943]= 1374507575;
assign addr[44944]= 1344905966;
assign addr[44945]= 1314877795;
assign addr[44946]= 1284432584;
assign addr[44947]= 1253579991;
assign addr[44948]= 1222329801;
assign addr[44949]= 1190691925;
assign addr[44950]= 1158676398;
assign addr[44951]= 1126293375;
assign addr[44952]= 1093553126;
assign addr[44953]= 1060466036;
assign addr[44954]= 1027042599;
assign addr[44955]= 993293415;
assign addr[44956]= 959229189;
assign addr[44957]= 924860725;
assign addr[44958]= 890198924;
assign addr[44959]= 855254778;
assign addr[44960]= 820039373;
assign addr[44961]= 784563876;
assign addr[44962]= 748839539;
assign addr[44963]= 712877694;
assign addr[44964]= 676689746;
assign addr[44965]= 640287172;
assign addr[44966]= 603681519;
assign addr[44967]= 566884397;
assign addr[44968]= 529907477;
assign addr[44969]= 492762486;
assign addr[44970]= 455461206;
assign addr[44971]= 418015468;
assign addr[44972]= 380437148;
assign addr[44973]= 342738165;
assign addr[44974]= 304930476;
assign addr[44975]= 267026072;
assign addr[44976]= 229036977;
assign addr[44977]= 190975237;
assign addr[44978]= 152852926;
assign addr[44979]= 114682135;
assign addr[44980]= 76474970;
assign addr[44981]= 38243550;
assign addr[44982]= 0;
assign addr[44983]= -38243550;
assign addr[44984]= -76474970;
assign addr[44985]= -114682135;
assign addr[44986]= -152852926;
assign addr[44987]= -190975237;
assign addr[44988]= -229036977;
assign addr[44989]= -267026072;
assign addr[44990]= -304930476;
assign addr[44991]= -342738165;
assign addr[44992]= -380437148;
assign addr[44993]= -418015468;
assign addr[44994]= -455461206;
assign addr[44995]= -492762486;
assign addr[44996]= -529907477;
assign addr[44997]= -566884397;
assign addr[44998]= -603681519;
assign addr[44999]= -640287172;
assign addr[45000]= -676689746;
assign addr[45001]= -712877694;
assign addr[45002]= -748839539;
assign addr[45003]= -784563876;
assign addr[45004]= -820039373;
assign addr[45005]= -855254778;
assign addr[45006]= -890198924;
assign addr[45007]= -924860725;
assign addr[45008]= -959229189;
assign addr[45009]= -993293415;
assign addr[45010]= -1027042599;
assign addr[45011]= -1060466036;
assign addr[45012]= -1093553126;
assign addr[45013]= -1126293375;
assign addr[45014]= -1158676398;
assign addr[45015]= -1190691925;
assign addr[45016]= -1222329801;
assign addr[45017]= -1253579991;
assign addr[45018]= -1284432584;
assign addr[45019]= -1314877795;
assign addr[45020]= -1344905966;
assign addr[45021]= -1374507575;
assign addr[45022]= -1403673233;
assign addr[45023]= -1432393688;
assign addr[45024]= -1460659832;
assign addr[45025]= -1488462700;
assign addr[45026]= -1515793473;
assign addr[45027]= -1542643483;
assign addr[45028]= -1569004214;
assign addr[45029]= -1594867305;
assign addr[45030]= -1620224553;
assign addr[45031]= -1645067915;
assign addr[45032]= -1669389513;
assign addr[45033]= -1693181631;
assign addr[45034]= -1716436725;
assign addr[45035]= -1739147417;
assign addr[45036]= -1761306505;
assign addr[45037]= -1782906961;
assign addr[45038]= -1803941934;
assign addr[45039]= -1824404752;
assign addr[45040]= -1844288924;
assign addr[45041]= -1863588145;
assign addr[45042]= -1882296293;
assign addr[45043]= -1900407434;
assign addr[45044]= -1917915825;
assign addr[45045]= -1934815911;
assign addr[45046]= -1951102334;
assign addr[45047]= -1966769926;
assign addr[45048]= -1981813720;
assign addr[45049]= -1996228943;
assign addr[45050]= -2010011024;
assign addr[45051]= -2023155591;
assign addr[45052]= -2035658475;
assign addr[45053]= -2047515711;
assign addr[45054]= -2058723538;
assign addr[45055]= -2069278401;
assign addr[45056]= -2079176953;
assign addr[45057]= -2088416053;
assign addr[45058]= -2096992772;
assign addr[45059]= -2104904390;
assign addr[45060]= -2112148396;
assign addr[45061]= -2118722494;
assign addr[45062]= -2124624598;
assign addr[45063]= -2129852837;
assign addr[45064]= -2134405552;
assign addr[45065]= -2138281298;
assign addr[45066]= -2141478848;
assign addr[45067]= -2143997187;
assign addr[45068]= -2145835515;
assign addr[45069]= -2146993250;
assign addr[45070]= -2147470025;
assign addr[45071]= -2147265689;
assign addr[45072]= -2146380306;
assign addr[45073]= -2144814157;
assign addr[45074]= -2142567738;
assign addr[45075]= -2139641764;
assign addr[45076]= -2136037160;
assign addr[45077]= -2131755071;
assign addr[45078]= -2126796855;
assign addr[45079]= -2121164085;
assign addr[45080]= -2114858546;
assign addr[45081]= -2107882239;
assign addr[45082]= -2100237377;
assign addr[45083]= -2091926384;
assign addr[45084]= -2082951896;
assign addr[45085]= -2073316760;
assign addr[45086]= -2063024031;
assign addr[45087]= -2052076975;
assign addr[45088]= -2040479063;
assign addr[45089]= -2028233973;
assign addr[45090]= -2015345591;
assign addr[45091]= -2001818002;
assign addr[45092]= -1987655498;
assign addr[45093]= -1972862571;
assign addr[45094]= -1957443913;
assign addr[45095]= -1941404413;
assign addr[45096]= -1924749160;
assign addr[45097]= -1907483436;
assign addr[45098]= -1889612716;
assign addr[45099]= -1871142669;
assign addr[45100]= -1852079154;
assign addr[45101]= -1832428215;
assign addr[45102]= -1812196087;
assign addr[45103]= -1791389186;
assign addr[45104]= -1770014111;
assign addr[45105]= -1748077642;
assign addr[45106]= -1725586737;
assign addr[45107]= -1702548529;
assign addr[45108]= -1678970324;
assign addr[45109]= -1654859602;
assign addr[45110]= -1630224009;
assign addr[45111]= -1605071359;
assign addr[45112]= -1579409630;
assign addr[45113]= -1553246960;
assign addr[45114]= -1526591649;
assign addr[45115]= -1499452149;
assign addr[45116]= -1471837070;
assign addr[45117]= -1443755168;
assign addr[45118]= -1415215352;
assign addr[45119]= -1386226674;
assign addr[45120]= -1356798326;
assign addr[45121]= -1326939644;
assign addr[45122]= -1296660098;
assign addr[45123]= -1265969291;
assign addr[45124]= -1234876957;
assign addr[45125]= -1203392958;
assign addr[45126]= -1171527280;
assign addr[45127]= -1139290029;
assign addr[45128]= -1106691431;
assign addr[45129]= -1073741824;
assign addr[45130]= -1040451659;
assign addr[45131]= -1006831495;
assign addr[45132]= -972891995;
assign addr[45133]= -938643924;
assign addr[45134]= -904098143;
assign addr[45135]= -869265610;
assign addr[45136]= -834157373;
assign addr[45137]= -798784567;
assign addr[45138]= -763158411;
assign addr[45139]= -727290205;
assign addr[45140]= -691191324;
assign addr[45141]= -654873219;
assign addr[45142]= -618347408;
assign addr[45143]= -581625477;
assign addr[45144]= -544719071;
assign addr[45145]= -507639898;
assign addr[45146]= -470399716;
assign addr[45147]= -433010339;
assign addr[45148]= -395483624;
assign addr[45149]= -357831473;
assign addr[45150]= -320065829;
assign addr[45151]= -282198671;
assign addr[45152]= -244242007;
assign addr[45153]= -206207878;
assign addr[45154]= -168108346;
assign addr[45155]= -129955495;
assign addr[45156]= -91761426;
assign addr[45157]= -53538253;
assign addr[45158]= -15298099;
assign addr[45159]= 22946906;
assign addr[45160]= 61184634;
assign addr[45161]= 99402956;
assign addr[45162]= 137589750;
assign addr[45163]= 175732905;
assign addr[45164]= 213820322;
assign addr[45165]= 251839923;
assign addr[45166]= 289779648;
assign addr[45167]= 327627463;
assign addr[45168]= 365371365;
assign addr[45169]= 402999383;
assign addr[45170]= 440499581;
assign addr[45171]= 477860067;
assign addr[45172]= 515068990;
assign addr[45173]= 552114549;
assign addr[45174]= 588984994;
assign addr[45175]= 625668632;
assign addr[45176]= 662153826;
assign addr[45177]= 698429006;
assign addr[45178]= 734482665;
assign addr[45179]= 770303369;
assign addr[45180]= 805879757;
assign addr[45181]= 841200544;
assign addr[45182]= 876254528;
assign addr[45183]= 911030591;
assign addr[45184]= 945517704;
assign addr[45185]= 979704927;
assign addr[45186]= 1013581418;
assign addr[45187]= 1047136432;
assign addr[45188]= 1080359326;
assign addr[45189]= 1113239564;
assign addr[45190]= 1145766716;
assign addr[45191]= 1177930466;
assign addr[45192]= 1209720613;
assign addr[45193]= 1241127074;
assign addr[45194]= 1272139887;
assign addr[45195]= 1302749217;
assign addr[45196]= 1332945355;
assign addr[45197]= 1362718723;
assign addr[45198]= 1392059879;
assign addr[45199]= 1420959516;
assign addr[45200]= 1449408469;
assign addr[45201]= 1477397714;
assign addr[45202]= 1504918373;
assign addr[45203]= 1531961719;
assign addr[45204]= 1558519173;
assign addr[45205]= 1584582314;
assign addr[45206]= 1610142873;
assign addr[45207]= 1635192744;
assign addr[45208]= 1659723983;
assign addr[45209]= 1683728808;
assign addr[45210]= 1707199606;
assign addr[45211]= 1730128933;
assign addr[45212]= 1752509516;
assign addr[45213]= 1774334257;
assign addr[45214]= 1795596234;
assign addr[45215]= 1816288703;
assign addr[45216]= 1836405100;
assign addr[45217]= 1855939047;
assign addr[45218]= 1874884346;
assign addr[45219]= 1893234990;
assign addr[45220]= 1910985158;
assign addr[45221]= 1928129220;
assign addr[45222]= 1944661739;
assign addr[45223]= 1960577471;
assign addr[45224]= 1975871368;
assign addr[45225]= 1990538579;
assign addr[45226]= 2004574453;
assign addr[45227]= 2017974537;
assign addr[45228]= 2030734582;
assign addr[45229]= 2042850540;
assign addr[45230]= 2054318569;
assign addr[45231]= 2065135031;
assign addr[45232]= 2075296495;
assign addr[45233]= 2084799740;
assign addr[45234]= 2093641749;
assign addr[45235]= 2101819720;
assign addr[45236]= 2109331059;
assign addr[45237]= 2116173382;
assign addr[45238]= 2122344521;
assign addr[45239]= 2127842516;
assign addr[45240]= 2132665626;
assign addr[45241]= 2136812319;
assign addr[45242]= 2140281282;
assign addr[45243]= 2143071413;
assign addr[45244]= 2145181827;
assign addr[45245]= 2146611856;
assign addr[45246]= 2147361045;
assign addr[45247]= 2147429158;
assign addr[45248]= 2146816171;
assign addr[45249]= 2145522281;
assign addr[45250]= 2143547897;
assign addr[45251]= 2140893646;
assign addr[45252]= 2137560369;
assign addr[45253]= 2133549123;
assign addr[45254]= 2128861181;
assign addr[45255]= 2123498030;
assign addr[45256]= 2117461370;
assign addr[45257]= 2110753117;
assign addr[45258]= 2103375398;
assign addr[45259]= 2095330553;
assign addr[45260]= 2086621133;
assign addr[45261]= 2077249901;
assign addr[45262]= 2067219829;
assign addr[45263]= 2056534099;
assign addr[45264]= 2045196100;
assign addr[45265]= 2033209426;
assign addr[45266]= 2020577882;
assign addr[45267]= 2007305472;
assign addr[45268]= 1993396407;
assign addr[45269]= 1978855097;
assign addr[45270]= 1963686155;
assign addr[45271]= 1947894393;
assign addr[45272]= 1931484818;
assign addr[45273]= 1914462636;
assign addr[45274]= 1896833245;
assign addr[45275]= 1878602237;
assign addr[45276]= 1859775393;
assign addr[45277]= 1840358687;
assign addr[45278]= 1820358275;
assign addr[45279]= 1799780501;
assign addr[45280]= 1778631892;
assign addr[45281]= 1756919156;
assign addr[45282]= 1734649179;
assign addr[45283]= 1711829025;
assign addr[45284]= 1688465931;
assign addr[45285]= 1664567307;
assign addr[45286]= 1640140734;
assign addr[45287]= 1615193959;
assign addr[45288]= 1589734894;
assign addr[45289]= 1563771613;
assign addr[45290]= 1537312353;
assign addr[45291]= 1510365504;
assign addr[45292]= 1482939614;
assign addr[45293]= 1455043381;
assign addr[45294]= 1426685652;
assign addr[45295]= 1397875423;
assign addr[45296]= 1368621831;
assign addr[45297]= 1338934154;
assign addr[45298]= 1308821808;
assign addr[45299]= 1278294345;
assign addr[45300]= 1247361445;
assign addr[45301]= 1216032921;
assign addr[45302]= 1184318708;
assign addr[45303]= 1152228866;
assign addr[45304]= 1119773573;
assign addr[45305]= 1086963121;
assign addr[45306]= 1053807919;
assign addr[45307]= 1020318481;
assign addr[45308]= 986505429;
assign addr[45309]= 952379488;
assign addr[45310]= 917951481;
assign addr[45311]= 883232329;
assign addr[45312]= 848233042;
assign addr[45313]= 812964722;
assign addr[45314]= 777438554;
assign addr[45315]= 741665807;
assign addr[45316]= 705657826;
assign addr[45317]= 669426032;
assign addr[45318]= 632981917;
assign addr[45319]= 596337040;
assign addr[45320]= 559503022;
assign addr[45321]= 522491548;
assign addr[45322]= 485314355;
assign addr[45323]= 447983235;
assign addr[45324]= 410510029;
assign addr[45325]= 372906622;
assign addr[45326]= 335184940;
assign addr[45327]= 297356948;
assign addr[45328]= 259434643;
assign addr[45329]= 221430054;
assign addr[45330]= 183355234;
assign addr[45331]= 145222259;
assign addr[45332]= 107043224;
assign addr[45333]= 68830239;
assign addr[45334]= 30595422;
assign addr[45335]= -7649098;
assign addr[45336]= -45891193;
assign addr[45337]= -84118732;
assign addr[45338]= -122319591;
assign addr[45339]= -160481654;
assign addr[45340]= -198592817;
assign addr[45341]= -236640993;
assign addr[45342]= -274614114;
assign addr[45343]= -312500135;
assign addr[45344]= -350287041;
assign addr[45345]= -387962847;
assign addr[45346]= -425515602;
assign addr[45347]= -462933398;
assign addr[45348]= -500204365;
assign addr[45349]= -537316682;
assign addr[45350]= -574258580;
assign addr[45351]= -611018340;
assign addr[45352]= -647584304;
assign addr[45353]= -683944874;
assign addr[45354]= -720088517;
assign addr[45355]= -756003771;
assign addr[45356]= -791679244;
assign addr[45357]= -827103620;
assign addr[45358]= -862265664;
assign addr[45359]= -897154224;
assign addr[45360]= -931758235;
assign addr[45361]= -966066720;
assign addr[45362]= -1000068799;
assign addr[45363]= -1033753687;
assign addr[45364]= -1067110699;
assign addr[45365]= -1100129257;
assign addr[45366]= -1132798888;
assign addr[45367]= -1165109230;
assign addr[45368]= -1197050035;
assign addr[45369]= -1228611172;
assign addr[45370]= -1259782632;
assign addr[45371]= -1290554528;
assign addr[45372]= -1320917099;
assign addr[45373]= -1350860716;
assign addr[45374]= -1380375881;
assign addr[45375]= -1409453233;
assign addr[45376]= -1438083551;
assign addr[45377]= -1466257752;
assign addr[45378]= -1493966902;
assign addr[45379]= -1521202211;
assign addr[45380]= -1547955041;
assign addr[45381]= -1574216908;
assign addr[45382]= -1599979481;
assign addr[45383]= -1625234591;
assign addr[45384]= -1649974225;
assign addr[45385]= -1674190539;
assign addr[45386]= -1697875851;
assign addr[45387]= -1721022648;
assign addr[45388]= -1743623590;
assign addr[45389]= -1765671509;
assign addr[45390]= -1787159411;
assign addr[45391]= -1808080480;
assign addr[45392]= -1828428082;
assign addr[45393]= -1848195763;
assign addr[45394]= -1867377253;
assign addr[45395]= -1885966468;
assign addr[45396]= -1903957513;
assign addr[45397]= -1921344681;
assign addr[45398]= -1938122457;
assign addr[45399]= -1954285520;
assign addr[45400]= -1969828744;
assign addr[45401]= -1984747199;
assign addr[45402]= -1999036154;
assign addr[45403]= -2012691075;
assign addr[45404]= -2025707632;
assign addr[45405]= -2038081698;
assign addr[45406]= -2049809346;
assign addr[45407]= -2060886858;
assign addr[45408]= -2071310720;
assign addr[45409]= -2081077626;
assign addr[45410]= -2090184478;
assign addr[45411]= -2098628387;
assign addr[45412]= -2106406677;
assign addr[45413]= -2113516878;
assign addr[45414]= -2119956737;
assign addr[45415]= -2125724211;
assign addr[45416]= -2130817471;
assign addr[45417]= -2135234901;
assign addr[45418]= -2138975100;
assign addr[45419]= -2142036881;
assign addr[45420]= -2144419275;
assign addr[45421]= -2146121524;
assign addr[45422]= -2147143090;
assign addr[45423]= -2147483648;
assign addr[45424]= -2147143090;
assign addr[45425]= -2146121524;
assign addr[45426]= -2144419275;
assign addr[45427]= -2142036881;
assign addr[45428]= -2138975100;
assign addr[45429]= -2135234901;
assign addr[45430]= -2130817471;
assign addr[45431]= -2125724211;
assign addr[45432]= -2119956737;
assign addr[45433]= -2113516878;
assign addr[45434]= -2106406677;
assign addr[45435]= -2098628387;
assign addr[45436]= -2090184478;
assign addr[45437]= -2081077626;
assign addr[45438]= -2071310720;
assign addr[45439]= -2060886858;
assign addr[45440]= -2049809346;
assign addr[45441]= -2038081698;
assign addr[45442]= -2025707632;
assign addr[45443]= -2012691075;
assign addr[45444]= -1999036154;
assign addr[45445]= -1984747199;
assign addr[45446]= -1969828744;
assign addr[45447]= -1954285520;
assign addr[45448]= -1938122457;
assign addr[45449]= -1921344681;
assign addr[45450]= -1903957513;
assign addr[45451]= -1885966468;
assign addr[45452]= -1867377253;
assign addr[45453]= -1848195763;
assign addr[45454]= -1828428082;
assign addr[45455]= -1808080480;
assign addr[45456]= -1787159411;
assign addr[45457]= -1765671509;
assign addr[45458]= -1743623590;
assign addr[45459]= -1721022648;
assign addr[45460]= -1697875851;
assign addr[45461]= -1674190539;
assign addr[45462]= -1649974225;
assign addr[45463]= -1625234591;
assign addr[45464]= -1599979481;
assign addr[45465]= -1574216908;
assign addr[45466]= -1547955041;
assign addr[45467]= -1521202211;
assign addr[45468]= -1493966902;
assign addr[45469]= -1466257752;
assign addr[45470]= -1438083551;
assign addr[45471]= -1409453233;
assign addr[45472]= -1380375881;
assign addr[45473]= -1350860716;
assign addr[45474]= -1320917099;
assign addr[45475]= -1290554528;
assign addr[45476]= -1259782632;
assign addr[45477]= -1228611172;
assign addr[45478]= -1197050035;
assign addr[45479]= -1165109230;
assign addr[45480]= -1132798888;
assign addr[45481]= -1100129257;
assign addr[45482]= -1067110699;
assign addr[45483]= -1033753687;
assign addr[45484]= -1000068799;
assign addr[45485]= -966066720;
assign addr[45486]= -931758235;
assign addr[45487]= -897154224;
assign addr[45488]= -862265664;
assign addr[45489]= -827103620;
assign addr[45490]= -791679244;
assign addr[45491]= -756003771;
assign addr[45492]= -720088517;
assign addr[45493]= -683944874;
assign addr[45494]= -647584304;
assign addr[45495]= -611018340;
assign addr[45496]= -574258580;
assign addr[45497]= -537316682;
assign addr[45498]= -500204365;
assign addr[45499]= -462933398;
assign addr[45500]= -425515602;
assign addr[45501]= -387962847;
assign addr[45502]= -350287041;
assign addr[45503]= -312500135;
assign addr[45504]= -274614114;
assign addr[45505]= -236640993;
assign addr[45506]= -198592817;
assign addr[45507]= -160481654;
assign addr[45508]= -122319591;
assign addr[45509]= -84118732;
assign addr[45510]= -45891193;
assign addr[45511]= -7649098;
assign addr[45512]= 30595422;
assign addr[45513]= 68830239;
assign addr[45514]= 107043224;
assign addr[45515]= 145222259;
assign addr[45516]= 183355234;
assign addr[45517]= 221430054;
assign addr[45518]= 259434643;
assign addr[45519]= 297356948;
assign addr[45520]= 335184940;
assign addr[45521]= 372906622;
assign addr[45522]= 410510029;
assign addr[45523]= 447983235;
assign addr[45524]= 485314355;
assign addr[45525]= 522491548;
assign addr[45526]= 559503022;
assign addr[45527]= 596337040;
assign addr[45528]= 632981917;
assign addr[45529]= 669426032;
assign addr[45530]= 705657826;
assign addr[45531]= 741665807;
assign addr[45532]= 777438554;
assign addr[45533]= 812964722;
assign addr[45534]= 848233042;
assign addr[45535]= 883232329;
assign addr[45536]= 917951481;
assign addr[45537]= 952379488;
assign addr[45538]= 986505429;
assign addr[45539]= 1020318481;
assign addr[45540]= 1053807919;
assign addr[45541]= 1086963121;
assign addr[45542]= 1119773573;
assign addr[45543]= 1152228866;
assign addr[45544]= 1184318708;
assign addr[45545]= 1216032921;
assign addr[45546]= 1247361445;
assign addr[45547]= 1278294345;
assign addr[45548]= 1308821808;
assign addr[45549]= 1338934154;
assign addr[45550]= 1368621831;
assign addr[45551]= 1397875423;
assign addr[45552]= 1426685652;
assign addr[45553]= 1455043381;
assign addr[45554]= 1482939614;
assign addr[45555]= 1510365504;
assign addr[45556]= 1537312353;
assign addr[45557]= 1563771613;
assign addr[45558]= 1589734894;
assign addr[45559]= 1615193959;
assign addr[45560]= 1640140734;
assign addr[45561]= 1664567307;
assign addr[45562]= 1688465931;
assign addr[45563]= 1711829025;
assign addr[45564]= 1734649179;
assign addr[45565]= 1756919156;
assign addr[45566]= 1778631892;
assign addr[45567]= 1799780501;
assign addr[45568]= 1820358275;
assign addr[45569]= 1840358687;
assign addr[45570]= 1859775393;
assign addr[45571]= 1878602237;
assign addr[45572]= 1896833245;
assign addr[45573]= 1914462636;
assign addr[45574]= 1931484818;
assign addr[45575]= 1947894393;
assign addr[45576]= 1963686155;
assign addr[45577]= 1978855097;
assign addr[45578]= 1993396407;
assign addr[45579]= 2007305472;
assign addr[45580]= 2020577882;
assign addr[45581]= 2033209426;
assign addr[45582]= 2045196100;
assign addr[45583]= 2056534099;
assign addr[45584]= 2067219829;
assign addr[45585]= 2077249901;
assign addr[45586]= 2086621133;
assign addr[45587]= 2095330553;
assign addr[45588]= 2103375398;
assign addr[45589]= 2110753117;
assign addr[45590]= 2117461370;
assign addr[45591]= 2123498030;
assign addr[45592]= 2128861181;
assign addr[45593]= 2133549123;
assign addr[45594]= 2137560369;
assign addr[45595]= 2140893646;
assign addr[45596]= 2143547897;
assign addr[45597]= 2145522281;
assign addr[45598]= 2146816171;
assign addr[45599]= 2147429158;
assign addr[45600]= 2147361045;
assign addr[45601]= 2146611856;
assign addr[45602]= 2145181827;
assign addr[45603]= 2143071413;
assign addr[45604]= 2140281282;
assign addr[45605]= 2136812319;
assign addr[45606]= 2132665626;
assign addr[45607]= 2127842516;
assign addr[45608]= 2122344521;
assign addr[45609]= 2116173382;
assign addr[45610]= 2109331059;
assign addr[45611]= 2101819720;
assign addr[45612]= 2093641749;
assign addr[45613]= 2084799740;
assign addr[45614]= 2075296495;
assign addr[45615]= 2065135031;
assign addr[45616]= 2054318569;
assign addr[45617]= 2042850540;
assign addr[45618]= 2030734582;
assign addr[45619]= 2017974537;
assign addr[45620]= 2004574453;
assign addr[45621]= 1990538579;
assign addr[45622]= 1975871368;
assign addr[45623]= 1960577471;
assign addr[45624]= 1944661739;
assign addr[45625]= 1928129220;
assign addr[45626]= 1910985158;
assign addr[45627]= 1893234990;
assign addr[45628]= 1874884346;
assign addr[45629]= 1855939047;
assign addr[45630]= 1836405100;
assign addr[45631]= 1816288703;
assign addr[45632]= 1795596234;
assign addr[45633]= 1774334257;
assign addr[45634]= 1752509516;
assign addr[45635]= 1730128933;
assign addr[45636]= 1707199606;
assign addr[45637]= 1683728808;
assign addr[45638]= 1659723983;
assign addr[45639]= 1635192744;
assign addr[45640]= 1610142873;
assign addr[45641]= 1584582314;
assign addr[45642]= 1558519173;
assign addr[45643]= 1531961719;
assign addr[45644]= 1504918373;
assign addr[45645]= 1477397714;
assign addr[45646]= 1449408469;
assign addr[45647]= 1420959516;
assign addr[45648]= 1392059879;
assign addr[45649]= 1362718723;
assign addr[45650]= 1332945355;
assign addr[45651]= 1302749217;
assign addr[45652]= 1272139887;
assign addr[45653]= 1241127074;
assign addr[45654]= 1209720613;
assign addr[45655]= 1177930466;
assign addr[45656]= 1145766716;
assign addr[45657]= 1113239564;
assign addr[45658]= 1080359326;
assign addr[45659]= 1047136432;
assign addr[45660]= 1013581418;
assign addr[45661]= 979704927;
assign addr[45662]= 945517704;
assign addr[45663]= 911030591;
assign addr[45664]= 876254528;
assign addr[45665]= 841200544;
assign addr[45666]= 805879757;
assign addr[45667]= 770303369;
assign addr[45668]= 734482665;
assign addr[45669]= 698429006;
assign addr[45670]= 662153826;
assign addr[45671]= 625668632;
assign addr[45672]= 588984994;
assign addr[45673]= 552114549;
assign addr[45674]= 515068990;
assign addr[45675]= 477860067;
assign addr[45676]= 440499581;
assign addr[45677]= 402999383;
assign addr[45678]= 365371365;
assign addr[45679]= 327627463;
assign addr[45680]= 289779648;
assign addr[45681]= 251839923;
assign addr[45682]= 213820322;
assign addr[45683]= 175732905;
assign addr[45684]= 137589750;
assign addr[45685]= 99402956;
assign addr[45686]= 61184634;
assign addr[45687]= 22946906;
assign addr[45688]= -15298099;
assign addr[45689]= -53538253;
assign addr[45690]= -91761426;
assign addr[45691]= -129955495;
assign addr[45692]= -168108346;
assign addr[45693]= -206207878;
assign addr[45694]= -244242007;
assign addr[45695]= -282198671;
assign addr[45696]= -320065829;
assign addr[45697]= -357831473;
assign addr[45698]= -395483624;
assign addr[45699]= -433010339;
assign addr[45700]= -470399716;
assign addr[45701]= -507639898;
assign addr[45702]= -544719071;
assign addr[45703]= -581625477;
assign addr[45704]= -618347408;
assign addr[45705]= -654873219;
assign addr[45706]= -691191324;
assign addr[45707]= -727290205;
assign addr[45708]= -763158411;
assign addr[45709]= -798784567;
assign addr[45710]= -834157373;
assign addr[45711]= -869265610;
assign addr[45712]= -904098143;
assign addr[45713]= -938643924;
assign addr[45714]= -972891995;
assign addr[45715]= -1006831495;
assign addr[45716]= -1040451659;
assign addr[45717]= -1073741824;
assign addr[45718]= -1106691431;
assign addr[45719]= -1139290029;
assign addr[45720]= -1171527280;
assign addr[45721]= -1203392958;
assign addr[45722]= -1234876957;
assign addr[45723]= -1265969291;
assign addr[45724]= -1296660098;
assign addr[45725]= -1326939644;
assign addr[45726]= -1356798326;
assign addr[45727]= -1386226674;
assign addr[45728]= -1415215352;
assign addr[45729]= -1443755168;
assign addr[45730]= -1471837070;
assign addr[45731]= -1499452149;
assign addr[45732]= -1526591649;
assign addr[45733]= -1553246960;
assign addr[45734]= -1579409630;
assign addr[45735]= -1605071359;
assign addr[45736]= -1630224009;
assign addr[45737]= -1654859602;
assign addr[45738]= -1678970324;
assign addr[45739]= -1702548529;
assign addr[45740]= -1725586737;
assign addr[45741]= -1748077642;
assign addr[45742]= -1770014111;
assign addr[45743]= -1791389186;
assign addr[45744]= -1812196087;
assign addr[45745]= -1832428215;
assign addr[45746]= -1852079154;
assign addr[45747]= -1871142669;
assign addr[45748]= -1889612716;
assign addr[45749]= -1907483436;
assign addr[45750]= -1924749160;
assign addr[45751]= -1941404413;
assign addr[45752]= -1957443913;
assign addr[45753]= -1972862571;
assign addr[45754]= -1987655498;
assign addr[45755]= -2001818002;
assign addr[45756]= -2015345591;
assign addr[45757]= -2028233973;
assign addr[45758]= -2040479063;
assign addr[45759]= -2052076975;
assign addr[45760]= -2063024031;
assign addr[45761]= -2073316760;
assign addr[45762]= -2082951896;
assign addr[45763]= -2091926384;
assign addr[45764]= -2100237377;
assign addr[45765]= -2107882239;
assign addr[45766]= -2114858546;
assign addr[45767]= -2121164085;
assign addr[45768]= -2126796855;
assign addr[45769]= -2131755071;
assign addr[45770]= -2136037160;
assign addr[45771]= -2139641764;
assign addr[45772]= -2142567738;
assign addr[45773]= -2144814157;
assign addr[45774]= -2146380306;
assign addr[45775]= -2147265689;
assign addr[45776]= -2147470025;
assign addr[45777]= -2146993250;
assign addr[45778]= -2145835515;
assign addr[45779]= -2143997187;
assign addr[45780]= -2141478848;
assign addr[45781]= -2138281298;
assign addr[45782]= -2134405552;
assign addr[45783]= -2129852837;
assign addr[45784]= -2124624598;
assign addr[45785]= -2118722494;
assign addr[45786]= -2112148396;
assign addr[45787]= -2104904390;
assign addr[45788]= -2096992772;
assign addr[45789]= -2088416053;
assign addr[45790]= -2079176953;
assign addr[45791]= -2069278401;
assign addr[45792]= -2058723538;
assign addr[45793]= -2047515711;
assign addr[45794]= -2035658475;
assign addr[45795]= -2023155591;
assign addr[45796]= -2010011024;
assign addr[45797]= -1996228943;
assign addr[45798]= -1981813720;
assign addr[45799]= -1966769926;
assign addr[45800]= -1951102334;
assign addr[45801]= -1934815911;
assign addr[45802]= -1917915825;
assign addr[45803]= -1900407434;
assign addr[45804]= -1882296293;
assign addr[45805]= -1863588145;
assign addr[45806]= -1844288924;
assign addr[45807]= -1824404752;
assign addr[45808]= -1803941934;
assign addr[45809]= -1782906961;
assign addr[45810]= -1761306505;
assign addr[45811]= -1739147417;
assign addr[45812]= -1716436725;
assign addr[45813]= -1693181631;
assign addr[45814]= -1669389513;
assign addr[45815]= -1645067915;
assign addr[45816]= -1620224553;
assign addr[45817]= -1594867305;
assign addr[45818]= -1569004214;
assign addr[45819]= -1542643483;
assign addr[45820]= -1515793473;
assign addr[45821]= -1488462700;
assign addr[45822]= -1460659832;
assign addr[45823]= -1432393688;
assign addr[45824]= -1403673233;
assign addr[45825]= -1374507575;
assign addr[45826]= -1344905966;
assign addr[45827]= -1314877795;
assign addr[45828]= -1284432584;
assign addr[45829]= -1253579991;
assign addr[45830]= -1222329801;
assign addr[45831]= -1190691925;
assign addr[45832]= -1158676398;
assign addr[45833]= -1126293375;
assign addr[45834]= -1093553126;
assign addr[45835]= -1060466036;
assign addr[45836]= -1027042599;
assign addr[45837]= -993293415;
assign addr[45838]= -959229189;
assign addr[45839]= -924860725;
assign addr[45840]= -890198924;
assign addr[45841]= -855254778;
assign addr[45842]= -820039373;
assign addr[45843]= -784563876;
assign addr[45844]= -748839539;
assign addr[45845]= -712877694;
assign addr[45846]= -676689746;
assign addr[45847]= -640287172;
assign addr[45848]= -603681519;
assign addr[45849]= -566884397;
assign addr[45850]= -529907477;
assign addr[45851]= -492762486;
assign addr[45852]= -455461206;
assign addr[45853]= -418015468;
assign addr[45854]= -380437148;
assign addr[45855]= -342738165;
assign addr[45856]= -304930476;
assign addr[45857]= -267026072;
assign addr[45858]= -229036977;
assign addr[45859]= -190975237;
assign addr[45860]= -152852926;
assign addr[45861]= -114682135;
assign addr[45862]= -76474970;
assign addr[45863]= -38243550;
assign addr[45864]= 0;
assign addr[45865]= 38243550;
assign addr[45866]= 76474970;
assign addr[45867]= 114682135;
assign addr[45868]= 152852926;
assign addr[45869]= 190975237;
assign addr[45870]= 229036977;
assign addr[45871]= 267026072;
assign addr[45872]= 304930476;
assign addr[45873]= 342738165;
assign addr[45874]= 380437148;
assign addr[45875]= 418015468;
assign addr[45876]= 455461206;
assign addr[45877]= 492762486;
assign addr[45878]= 529907477;
assign addr[45879]= 566884397;
assign addr[45880]= 603681519;
assign addr[45881]= 640287172;
assign addr[45882]= 676689746;
assign addr[45883]= 712877694;
assign addr[45884]= 748839539;
assign addr[45885]= 784563876;
assign addr[45886]= 820039373;
assign addr[45887]= 855254778;
assign addr[45888]= 890198924;
assign addr[45889]= 924860725;
assign addr[45890]= 959229189;
assign addr[45891]= 993293415;
assign addr[45892]= 1027042599;
assign addr[45893]= 1060466036;
assign addr[45894]= 1093553126;
assign addr[45895]= 1126293375;
assign addr[45896]= 1158676398;
assign addr[45897]= 1190691925;
assign addr[45898]= 1222329801;
assign addr[45899]= 1253579991;
assign addr[45900]= 1284432584;
assign addr[45901]= 1314877795;
assign addr[45902]= 1344905966;
assign addr[45903]= 1374507575;
assign addr[45904]= 1403673233;
assign addr[45905]= 1432393688;
assign addr[45906]= 1460659832;
assign addr[45907]= 1488462700;
assign addr[45908]= 1515793473;
assign addr[45909]= 1542643483;
assign addr[45910]= 1569004214;
assign addr[45911]= 1594867305;
assign addr[45912]= 1620224553;
assign addr[45913]= 1645067915;
assign addr[45914]= 1669389513;
assign addr[45915]= 1693181631;
assign addr[45916]= 1716436725;
assign addr[45917]= 1739147417;
assign addr[45918]= 1761306505;
assign addr[45919]= 1782906961;
assign addr[45920]= 1803941934;
assign addr[45921]= 1824404752;
assign addr[45922]= 1844288924;
assign addr[45923]= 1863588145;
assign addr[45924]= 1882296293;
assign addr[45925]= 1900407434;
assign addr[45926]= 1917915825;
assign addr[45927]= 1934815911;
assign addr[45928]= 1951102334;
assign addr[45929]= 1966769926;
assign addr[45930]= 1981813720;
assign addr[45931]= 1996228943;
assign addr[45932]= 2010011024;
assign addr[45933]= 2023155591;
assign addr[45934]= 2035658475;
assign addr[45935]= 2047515711;
assign addr[45936]= 2058723538;
assign addr[45937]= 2069278401;
assign addr[45938]= 2079176953;
assign addr[45939]= 2088416053;
assign addr[45940]= 2096992772;
assign addr[45941]= 2104904390;
assign addr[45942]= 2112148396;
assign addr[45943]= 2118722494;
assign addr[45944]= 2124624598;
assign addr[45945]= 2129852837;
assign addr[45946]= 2134405552;
assign addr[45947]= 2138281298;
assign addr[45948]= 2141478848;
assign addr[45949]= 2143997187;
assign addr[45950]= 2145835515;
assign addr[45951]= 2146993250;
assign addr[45952]= 2147470025;
assign addr[45953]= 2147265689;
assign addr[45954]= 2146380306;
assign addr[45955]= 2144814157;
assign addr[45956]= 2142567738;
assign addr[45957]= 2139641764;
assign addr[45958]= 2136037160;
assign addr[45959]= 2131755071;
assign addr[45960]= 2126796855;
assign addr[45961]= 2121164085;
assign addr[45962]= 2114858546;
assign addr[45963]= 2107882239;
assign addr[45964]= 2100237377;
assign addr[45965]= 2091926384;
assign addr[45966]= 2082951896;
assign addr[45967]= 2073316760;
assign addr[45968]= 2063024031;
assign addr[45969]= 2052076975;
assign addr[45970]= 2040479063;
assign addr[45971]= 2028233973;
assign addr[45972]= 2015345591;
assign addr[45973]= 2001818002;
assign addr[45974]= 1987655498;
assign addr[45975]= 1972862571;
assign addr[45976]= 1957443913;
assign addr[45977]= 1941404413;
assign addr[45978]= 1924749160;
assign addr[45979]= 1907483436;
assign addr[45980]= 1889612716;
assign addr[45981]= 1871142669;
assign addr[45982]= 1852079154;
assign addr[45983]= 1832428215;
assign addr[45984]= 1812196087;
assign addr[45985]= 1791389186;
assign addr[45986]= 1770014111;
assign addr[45987]= 1748077642;
assign addr[45988]= 1725586737;
assign addr[45989]= 1702548529;
assign addr[45990]= 1678970324;
assign addr[45991]= 1654859602;
assign addr[45992]= 1630224009;
assign addr[45993]= 1605071359;
assign addr[45994]= 1579409630;
assign addr[45995]= 1553246960;
assign addr[45996]= 1526591649;
assign addr[45997]= 1499452149;
assign addr[45998]= 1471837070;
assign addr[45999]= 1443755168;
assign addr[46000]= 1415215352;
assign addr[46001]= 1386226674;
assign addr[46002]= 1356798326;
assign addr[46003]= 1326939644;
assign addr[46004]= 1296660098;
assign addr[46005]= 1265969291;
assign addr[46006]= 1234876957;
assign addr[46007]= 1203392958;
assign addr[46008]= 1171527280;
assign addr[46009]= 1139290029;
assign addr[46010]= 1106691431;
assign addr[46011]= 1073741824;
assign addr[46012]= 1040451659;
assign addr[46013]= 1006831495;
assign addr[46014]= 972891995;
assign addr[46015]= 938643924;
assign addr[46016]= 904098143;
assign addr[46017]= 869265610;
assign addr[46018]= 834157373;
assign addr[46019]= 798784567;
assign addr[46020]= 763158411;
assign addr[46021]= 727290205;
assign addr[46022]= 691191324;
assign addr[46023]= 654873219;
assign addr[46024]= 618347408;
assign addr[46025]= 581625477;
assign addr[46026]= 544719071;
assign addr[46027]= 507639898;
assign addr[46028]= 470399716;
assign addr[46029]= 433010339;
assign addr[46030]= 395483624;
assign addr[46031]= 357831473;
assign addr[46032]= 320065829;
assign addr[46033]= 282198671;
assign addr[46034]= 244242007;
assign addr[46035]= 206207878;
assign addr[46036]= 168108346;
assign addr[46037]= 129955495;
assign addr[46038]= 91761426;
assign addr[46039]= 53538253;
assign addr[46040]= 15298099;
assign addr[46041]= -22946906;
assign addr[46042]= -61184634;
assign addr[46043]= -99402956;
assign addr[46044]= -137589750;
assign addr[46045]= -175732905;
assign addr[46046]= -213820322;
assign addr[46047]= -251839923;
assign addr[46048]= -289779648;
assign addr[46049]= -327627463;
assign addr[46050]= -365371365;
assign addr[46051]= -402999383;
assign addr[46052]= -440499581;
assign addr[46053]= -477860067;
assign addr[46054]= -515068990;
assign addr[46055]= -552114549;
assign addr[46056]= -588984994;
assign addr[46057]= -625668632;
assign addr[46058]= -662153826;
assign addr[46059]= -698429006;
assign addr[46060]= -734482665;
assign addr[46061]= -770303369;
assign addr[46062]= -805879757;
assign addr[46063]= -841200544;
assign addr[46064]= -876254528;
assign addr[46065]= -911030591;
assign addr[46066]= -945517704;
assign addr[46067]= -979704927;
assign addr[46068]= -1013581418;
assign addr[46069]= -1047136432;
assign addr[46070]= -1080359326;
assign addr[46071]= -1113239564;
assign addr[46072]= -1145766716;
assign addr[46073]= -1177930466;
assign addr[46074]= -1209720613;
assign addr[46075]= -1241127074;
assign addr[46076]= -1272139887;
assign addr[46077]= -1302749217;
assign addr[46078]= -1332945355;
assign addr[46079]= -1362718723;
assign addr[46080]= -1392059879;
assign addr[46081]= -1420959516;
assign addr[46082]= -1449408469;
assign addr[46083]= -1477397714;
assign addr[46084]= -1504918373;
assign addr[46085]= -1531961719;
assign addr[46086]= -1558519173;
assign addr[46087]= -1584582314;
assign addr[46088]= -1610142873;
assign addr[46089]= -1635192744;
assign addr[46090]= -1659723983;
assign addr[46091]= -1683728808;
assign addr[46092]= -1707199606;
assign addr[46093]= -1730128933;
assign addr[46094]= -1752509516;
assign addr[46095]= -1774334257;
assign addr[46096]= -1795596234;
assign addr[46097]= -1816288703;
assign addr[46098]= -1836405100;
assign addr[46099]= -1855939047;
assign addr[46100]= -1874884346;
assign addr[46101]= -1893234990;
assign addr[46102]= -1910985158;
assign addr[46103]= -1928129220;
assign addr[46104]= -1944661739;
assign addr[46105]= -1960577471;
assign addr[46106]= -1975871368;
assign addr[46107]= -1990538579;
assign addr[46108]= -2004574453;
assign addr[46109]= -2017974537;
assign addr[46110]= -2030734582;
assign addr[46111]= -2042850540;
assign addr[46112]= -2054318569;
assign addr[46113]= -2065135031;
assign addr[46114]= -2075296495;
assign addr[46115]= -2084799740;
assign addr[46116]= -2093641749;
assign addr[46117]= -2101819720;
assign addr[46118]= -2109331059;
assign addr[46119]= -2116173382;
assign addr[46120]= -2122344521;
assign addr[46121]= -2127842516;
assign addr[46122]= -2132665626;
assign addr[46123]= -2136812319;
assign addr[46124]= -2140281282;
assign addr[46125]= -2143071413;
assign addr[46126]= -2145181827;
assign addr[46127]= -2146611856;
assign addr[46128]= -2147361045;
assign addr[46129]= -2147429158;
assign addr[46130]= -2146816171;
assign addr[46131]= -2145522281;
assign addr[46132]= -2143547897;
assign addr[46133]= -2140893646;
assign addr[46134]= -2137560369;
assign addr[46135]= -2133549123;
assign addr[46136]= -2128861181;
assign addr[46137]= -2123498030;
assign addr[46138]= -2117461370;
assign addr[46139]= -2110753117;
assign addr[46140]= -2103375398;
assign addr[46141]= -2095330553;
assign addr[46142]= -2086621133;
assign addr[46143]= -2077249901;
assign addr[46144]= -2067219829;
assign addr[46145]= -2056534099;
assign addr[46146]= -2045196100;
assign addr[46147]= -2033209426;
assign addr[46148]= -2020577882;
assign addr[46149]= -2007305472;
assign addr[46150]= -1993396407;
assign addr[46151]= -1978855097;
assign addr[46152]= -1963686155;
assign addr[46153]= -1947894393;
assign addr[46154]= -1931484818;
assign addr[46155]= -1914462636;
assign addr[46156]= -1896833245;
assign addr[46157]= -1878602237;
assign addr[46158]= -1859775393;
assign addr[46159]= -1840358687;
assign addr[46160]= -1820358275;
assign addr[46161]= -1799780501;
assign addr[46162]= -1778631892;
assign addr[46163]= -1756919156;
assign addr[46164]= -1734649179;
assign addr[46165]= -1711829025;
assign addr[46166]= -1688465931;
assign addr[46167]= -1664567307;
assign addr[46168]= -1640140734;
assign addr[46169]= -1615193959;
assign addr[46170]= -1589734894;
assign addr[46171]= -1563771613;
assign addr[46172]= -1537312353;
assign addr[46173]= -1510365504;
assign addr[46174]= -1482939614;
assign addr[46175]= -1455043381;
assign addr[46176]= -1426685652;
assign addr[46177]= -1397875423;
assign addr[46178]= -1368621831;
assign addr[46179]= -1338934154;
assign addr[46180]= -1308821808;
assign addr[46181]= -1278294345;
assign addr[46182]= -1247361445;
assign addr[46183]= -1216032921;
assign addr[46184]= -1184318708;
assign addr[46185]= -1152228866;
assign addr[46186]= -1119773573;
assign addr[46187]= -1086963121;
assign addr[46188]= -1053807919;
assign addr[46189]= -1020318481;
assign addr[46190]= -986505429;
assign addr[46191]= -952379488;
assign addr[46192]= -917951481;
assign addr[46193]= -883232329;
assign addr[46194]= -848233042;
assign addr[46195]= -812964722;
assign addr[46196]= -777438554;
assign addr[46197]= -741665807;
assign addr[46198]= -705657826;
assign addr[46199]= -669426032;
assign addr[46200]= -632981917;
assign addr[46201]= -596337040;
assign addr[46202]= -559503022;
assign addr[46203]= -522491548;
assign addr[46204]= -485314355;
assign addr[46205]= -447983235;
assign addr[46206]= -410510029;
assign addr[46207]= -372906622;
assign addr[46208]= -335184940;
assign addr[46209]= -297356948;
assign addr[46210]= -259434643;
assign addr[46211]= -221430054;
assign addr[46212]= -183355234;
assign addr[46213]= -145222259;
assign addr[46214]= -107043224;
assign addr[46215]= -68830239;
assign addr[46216]= -30595422;
assign addr[46217]= 7649098;
assign addr[46218]= 45891193;
assign addr[46219]= 84118732;
assign addr[46220]= 122319591;
assign addr[46221]= 160481654;
assign addr[46222]= 198592817;
assign addr[46223]= 236640993;
assign addr[46224]= 274614114;
assign addr[46225]= 312500135;
assign addr[46226]= 350287041;
assign addr[46227]= 387962847;
assign addr[46228]= 425515602;
assign addr[46229]= 462933398;
assign addr[46230]= 500204365;
assign addr[46231]= 537316682;
assign addr[46232]= 574258580;
assign addr[46233]= 611018340;
assign addr[46234]= 647584304;
assign addr[46235]= 683944874;
assign addr[46236]= 720088517;
assign addr[46237]= 756003771;
assign addr[46238]= 791679244;
assign addr[46239]= 827103620;
assign addr[46240]= 862265664;
assign addr[46241]= 897154224;
assign addr[46242]= 931758235;
assign addr[46243]= 966066720;
assign addr[46244]= 1000068799;
assign addr[46245]= 1033753687;
assign addr[46246]= 1067110699;
assign addr[46247]= 1100129257;
assign addr[46248]= 1132798888;
assign addr[46249]= 1165109230;
assign addr[46250]= 1197050035;
assign addr[46251]= 1228611172;
assign addr[46252]= 1259782632;
assign addr[46253]= 1290554528;
assign addr[46254]= 1320917099;
assign addr[46255]= 1350860716;
assign addr[46256]= 1380375881;
assign addr[46257]= 1409453233;
assign addr[46258]= 1438083551;
assign addr[46259]= 1466257752;
assign addr[46260]= 1493966902;
assign addr[46261]= 1521202211;
assign addr[46262]= 1547955041;
assign addr[46263]= 1574216908;
assign addr[46264]= 1599979481;
assign addr[46265]= 1625234591;
assign addr[46266]= 1649974225;
assign addr[46267]= 1674190539;
assign addr[46268]= 1697875851;
assign addr[46269]= 1721022648;
assign addr[46270]= 1743623590;
assign addr[46271]= 1765671509;
assign addr[46272]= 1787159411;
assign addr[46273]= 1808080480;
assign addr[46274]= 1828428082;
assign addr[46275]= 1848195763;
assign addr[46276]= 1867377253;
assign addr[46277]= 1885966468;
assign addr[46278]= 1903957513;
assign addr[46279]= 1921344681;
assign addr[46280]= 1938122457;
assign addr[46281]= 1954285520;
assign addr[46282]= 1969828744;
assign addr[46283]= 1984747199;
assign addr[46284]= 1999036154;
assign addr[46285]= 2012691075;
assign addr[46286]= 2025707632;
assign addr[46287]= 2038081698;
assign addr[46288]= 2049809346;
assign addr[46289]= 2060886858;
assign addr[46290]= 2071310720;
assign addr[46291]= 2081077626;
assign addr[46292]= 2090184478;
assign addr[46293]= 2098628387;
assign addr[46294]= 2106406677;
assign addr[46295]= 2113516878;
assign addr[46296]= 2119956737;
assign addr[46297]= 2125724211;
assign addr[46298]= 2130817471;
assign addr[46299]= 2135234901;
assign addr[46300]= 2138975100;
assign addr[46301]= 2142036881;
assign addr[46302]= 2144419275;
assign addr[46303]= 2146121524;
assign addr[46304]= 2147143090;
assign addr[46305]= 2147483648;
assign addr[46306]= 2147143090;
assign addr[46307]= 2146121524;
assign addr[46308]= 2144419275;
assign addr[46309]= 2142036881;
assign addr[46310]= 2138975100;
assign addr[46311]= 2135234901;
assign addr[46312]= 2130817471;
assign addr[46313]= 2125724211;
assign addr[46314]= 2119956737;
assign addr[46315]= 2113516878;
assign addr[46316]= 2106406677;
assign addr[46317]= 2098628387;
assign addr[46318]= 2090184478;
assign addr[46319]= 2081077626;
assign addr[46320]= 2071310720;
assign addr[46321]= 2060886858;
assign addr[46322]= 2049809346;
assign addr[46323]= 2038081698;
assign addr[46324]= 2025707632;
assign addr[46325]= 2012691075;
assign addr[46326]= 1999036154;
assign addr[46327]= 1984747199;
assign addr[46328]= 1969828744;
assign addr[46329]= 1954285520;
assign addr[46330]= 1938122457;
assign addr[46331]= 1921344681;
assign addr[46332]= 1903957513;
assign addr[46333]= 1885966468;
assign addr[46334]= 1867377253;
assign addr[46335]= 1848195763;
assign addr[46336]= 1828428082;
assign addr[46337]= 1808080480;
assign addr[46338]= 1787159411;
assign addr[46339]= 1765671509;
assign addr[46340]= 1743623590;
assign addr[46341]= 1721022648;
assign addr[46342]= 1697875851;
assign addr[46343]= 1674190539;
assign addr[46344]= 1649974225;
assign addr[46345]= 1625234591;
assign addr[46346]= 1599979481;
assign addr[46347]= 1574216908;
assign addr[46348]= 1547955041;
assign addr[46349]= 1521202211;
assign addr[46350]= 1493966902;
assign addr[46351]= 1466257752;
assign addr[46352]= 1438083551;
assign addr[46353]= 1409453233;
assign addr[46354]= 1380375881;
assign addr[46355]= 1350860716;
assign addr[46356]= 1320917099;
assign addr[46357]= 1290554528;
assign addr[46358]= 1259782632;
assign addr[46359]= 1228611172;
assign addr[46360]= 1197050035;
assign addr[46361]= 1165109230;
assign addr[46362]= 1132798888;
assign addr[46363]= 1100129257;
assign addr[46364]= 1067110699;
assign addr[46365]= 1033753687;
assign addr[46366]= 1000068799;
assign addr[46367]= 966066720;
assign addr[46368]= 931758235;
assign addr[46369]= 897154224;
assign addr[46370]= 862265664;
assign addr[46371]= 827103620;
assign addr[46372]= 791679244;
assign addr[46373]= 756003771;
assign addr[46374]= 720088517;
assign addr[46375]= 683944874;
assign addr[46376]= 647584304;
assign addr[46377]= 611018340;
assign addr[46378]= 574258580;
assign addr[46379]= 537316682;
assign addr[46380]= 500204365;
assign addr[46381]= 462933398;
assign addr[46382]= 425515602;
assign addr[46383]= 387962847;
assign addr[46384]= 350287041;
assign addr[46385]= 312500135;
assign addr[46386]= 274614114;
assign addr[46387]= 236640993;
assign addr[46388]= 198592817;
assign addr[46389]= 160481654;
assign addr[46390]= 122319591;
assign addr[46391]= 84118732;
assign addr[46392]= 45891193;
assign addr[46393]= 7649098;
assign addr[46394]= -30595422;
assign addr[46395]= -68830239;
assign addr[46396]= -107043224;
assign addr[46397]= -145222259;
assign addr[46398]= -183355234;
assign addr[46399]= -221430054;
assign addr[46400]= -259434643;
assign addr[46401]= -297356948;
assign addr[46402]= -335184940;
assign addr[46403]= -372906622;
assign addr[46404]= -410510029;
assign addr[46405]= -447983235;
assign addr[46406]= -485314355;
assign addr[46407]= -522491548;
assign addr[46408]= -559503022;
assign addr[46409]= -596337040;
assign addr[46410]= -632981917;
assign addr[46411]= -669426032;
assign addr[46412]= -705657826;
assign addr[46413]= -741665807;
assign addr[46414]= -777438554;
assign addr[46415]= -812964722;
assign addr[46416]= -848233042;
assign addr[46417]= -883232329;
assign addr[46418]= -917951481;
assign addr[46419]= -952379488;
assign addr[46420]= -986505429;
assign addr[46421]= -1020318481;
assign addr[46422]= -1053807919;
assign addr[46423]= -1086963121;
assign addr[46424]= -1119773573;
assign addr[46425]= -1152228866;
assign addr[46426]= -1184318708;
assign addr[46427]= -1216032921;
assign addr[46428]= -1247361445;
assign addr[46429]= -1278294345;
assign addr[46430]= -1308821808;
assign addr[46431]= -1338934154;
assign addr[46432]= -1368621831;
assign addr[46433]= -1397875423;
assign addr[46434]= -1426685652;
assign addr[46435]= -1455043381;
assign addr[46436]= -1482939614;
assign addr[46437]= -1510365504;
assign addr[46438]= -1537312353;
assign addr[46439]= -1563771613;
assign addr[46440]= -1589734894;
assign addr[46441]= -1615193959;
assign addr[46442]= -1640140734;
assign addr[46443]= -1664567307;
assign addr[46444]= -1688465931;
assign addr[46445]= -1711829025;
assign addr[46446]= -1734649179;
assign addr[46447]= -1756919156;
assign addr[46448]= -1778631892;
assign addr[46449]= -1799780501;
assign addr[46450]= -1820358275;
assign addr[46451]= -1840358687;
assign addr[46452]= -1859775393;
assign addr[46453]= -1878602237;
assign addr[46454]= -1896833245;
assign addr[46455]= -1914462636;
assign addr[46456]= -1931484818;
assign addr[46457]= -1947894393;
assign addr[46458]= -1963686155;
assign addr[46459]= -1978855097;
assign addr[46460]= -1993396407;
assign addr[46461]= -2007305472;
assign addr[46462]= -2020577882;
assign addr[46463]= -2033209426;
assign addr[46464]= -2045196100;
assign addr[46465]= -2056534099;
assign addr[46466]= -2067219829;
assign addr[46467]= -2077249901;
assign addr[46468]= -2086621133;
assign addr[46469]= -2095330553;
assign addr[46470]= -2103375398;
assign addr[46471]= -2110753117;
assign addr[46472]= -2117461370;
assign addr[46473]= -2123498030;
assign addr[46474]= -2128861181;
assign addr[46475]= -2133549123;
assign addr[46476]= -2137560369;
assign addr[46477]= -2140893646;
assign addr[46478]= -2143547897;
assign addr[46479]= -2145522281;
assign addr[46480]= -2146816171;
assign addr[46481]= -2147429158;
assign addr[46482]= -2147361045;
assign addr[46483]= -2146611856;
assign addr[46484]= -2145181827;
assign addr[46485]= -2143071413;
assign addr[46486]= -2140281282;
assign addr[46487]= -2136812319;
assign addr[46488]= -2132665626;
assign addr[46489]= -2127842516;
assign addr[46490]= -2122344521;
assign addr[46491]= -2116173382;
assign addr[46492]= -2109331059;
assign addr[46493]= -2101819720;
assign addr[46494]= -2093641749;
assign addr[46495]= -2084799740;
assign addr[46496]= -2075296495;
assign addr[46497]= -2065135031;
assign addr[46498]= -2054318569;
assign addr[46499]= -2042850540;
assign addr[46500]= -2030734582;
assign addr[46501]= -2017974537;
assign addr[46502]= -2004574453;
assign addr[46503]= -1990538579;
assign addr[46504]= -1975871368;
assign addr[46505]= -1960577471;
assign addr[46506]= -1944661739;
assign addr[46507]= -1928129220;
assign addr[46508]= -1910985158;
assign addr[46509]= -1893234990;
assign addr[46510]= -1874884346;
assign addr[46511]= -1855939047;
assign addr[46512]= -1836405100;
assign addr[46513]= -1816288703;
assign addr[46514]= -1795596234;
assign addr[46515]= -1774334257;
assign addr[46516]= -1752509516;
assign addr[46517]= -1730128933;
assign addr[46518]= -1707199606;
assign addr[46519]= -1683728808;
assign addr[46520]= -1659723983;
assign addr[46521]= -1635192744;
assign addr[46522]= -1610142873;
assign addr[46523]= -1584582314;
assign addr[46524]= -1558519173;
assign addr[46525]= -1531961719;
assign addr[46526]= -1504918373;
assign addr[46527]= -1477397714;
assign addr[46528]= -1449408469;
assign addr[46529]= -1420959516;
assign addr[46530]= -1392059879;
assign addr[46531]= -1362718723;
assign addr[46532]= -1332945355;
assign addr[46533]= -1302749217;
assign addr[46534]= -1272139887;
assign addr[46535]= -1241127074;
assign addr[46536]= -1209720613;
assign addr[46537]= -1177930466;
assign addr[46538]= -1145766716;
assign addr[46539]= -1113239564;
assign addr[46540]= -1080359326;
assign addr[46541]= -1047136432;
assign addr[46542]= -1013581418;
assign addr[46543]= -979704927;
assign addr[46544]= -945517704;
assign addr[46545]= -911030591;
assign addr[46546]= -876254528;
assign addr[46547]= -841200544;
assign addr[46548]= -805879757;
assign addr[46549]= -770303369;
assign addr[46550]= -734482665;
assign addr[46551]= -698429006;
assign addr[46552]= -662153826;
assign addr[46553]= -625668632;
assign addr[46554]= -588984994;
assign addr[46555]= -552114549;
assign addr[46556]= -515068990;
assign addr[46557]= -477860067;
assign addr[46558]= -440499581;
assign addr[46559]= -402999383;
assign addr[46560]= -365371365;
assign addr[46561]= -327627463;
assign addr[46562]= -289779648;
assign addr[46563]= -251839923;
assign addr[46564]= -213820322;
assign addr[46565]= -175732905;
assign addr[46566]= -137589750;
assign addr[46567]= -99402956;
assign addr[46568]= -61184634;
assign addr[46569]= -22946906;
assign addr[46570]= 15298099;
assign addr[46571]= 53538253;
assign addr[46572]= 91761426;
assign addr[46573]= 129955495;
assign addr[46574]= 168108346;
assign addr[46575]= 206207878;
assign addr[46576]= 244242007;
assign addr[46577]= 282198671;
assign addr[46578]= 320065829;
assign addr[46579]= 357831473;
assign addr[46580]= 395483624;
assign addr[46581]= 433010339;
assign addr[46582]= 470399716;
assign addr[46583]= 507639898;
assign addr[46584]= 544719071;
assign addr[46585]= 581625477;
assign addr[46586]= 618347408;
assign addr[46587]= 654873219;
assign addr[46588]= 691191324;
assign addr[46589]= 727290205;
assign addr[46590]= 763158411;
assign addr[46591]= 798784567;
assign addr[46592]= 834157373;
assign addr[46593]= 869265610;
assign addr[46594]= 904098143;
assign addr[46595]= 938643924;
assign addr[46596]= 972891995;
assign addr[46597]= 1006831495;
assign addr[46598]= 1040451659;
assign addr[46599]= 1073741824;
assign addr[46600]= 1106691431;
assign addr[46601]= 1139290029;
assign addr[46602]= 1171527280;
assign addr[46603]= 1203392958;
assign addr[46604]= 1234876957;
assign addr[46605]= 1265969291;
assign addr[46606]= 1296660098;
assign addr[46607]= 1326939644;
assign addr[46608]= 1356798326;
assign addr[46609]= 1386226674;
assign addr[46610]= 1415215352;
assign addr[46611]= 1443755168;
assign addr[46612]= 1471837070;
assign addr[46613]= 1499452149;
assign addr[46614]= 1526591649;
assign addr[46615]= 1553246960;
assign addr[46616]= 1579409630;
assign addr[46617]= 1605071359;
assign addr[46618]= 1630224009;
assign addr[46619]= 1654859602;
assign addr[46620]= 1678970324;
assign addr[46621]= 1702548529;
assign addr[46622]= 1725586737;
assign addr[46623]= 1748077642;
assign addr[46624]= 1770014111;
assign addr[46625]= 1791389186;
assign addr[46626]= 1812196087;
assign addr[46627]= 1832428215;
assign addr[46628]= 1852079154;
assign addr[46629]= 1871142669;
assign addr[46630]= 1889612716;
assign addr[46631]= 1907483436;
assign addr[46632]= 1924749160;
assign addr[46633]= 1941404413;
assign addr[46634]= 1957443913;
assign addr[46635]= 1972862571;
assign addr[46636]= 1987655498;
assign addr[46637]= 2001818002;
assign addr[46638]= 2015345591;
assign addr[46639]= 2028233973;
assign addr[46640]= 2040479063;
assign addr[46641]= 2052076975;
assign addr[46642]= 2063024031;
assign addr[46643]= 2073316760;
assign addr[46644]= 2082951896;
assign addr[46645]= 2091926384;
assign addr[46646]= 2100237377;
assign addr[46647]= 2107882239;
assign addr[46648]= 2114858546;
assign addr[46649]= 2121164085;
assign addr[46650]= 2126796855;
assign addr[46651]= 2131755071;
assign addr[46652]= 2136037160;
assign addr[46653]= 2139641764;
assign addr[46654]= 2142567738;
assign addr[46655]= 2144814157;
assign addr[46656]= 2146380306;
assign addr[46657]= 2147265689;
assign addr[46658]= 2147470025;
assign addr[46659]= 2146993250;
assign addr[46660]= 2145835515;
assign addr[46661]= 2143997187;
assign addr[46662]= 2141478848;
assign addr[46663]= 2138281298;
assign addr[46664]= 2134405552;
assign addr[46665]= 2129852837;
assign addr[46666]= 2124624598;
assign addr[46667]= 2118722494;
assign addr[46668]= 2112148396;
assign addr[46669]= 2104904390;
assign addr[46670]= 2096992772;
assign addr[46671]= 2088416053;
assign addr[46672]= 2079176953;
assign addr[46673]= 2069278401;
assign addr[46674]= 2058723538;
assign addr[46675]= 2047515711;
assign addr[46676]= 2035658475;
assign addr[46677]= 2023155591;
assign addr[46678]= 2010011024;
assign addr[46679]= 1996228943;
assign addr[46680]= 1981813720;
assign addr[46681]= 1966769926;
assign addr[46682]= 1951102334;
assign addr[46683]= 1934815911;
assign addr[46684]= 1917915825;
assign addr[46685]= 1900407434;
assign addr[46686]= 1882296293;
assign addr[46687]= 1863588145;
assign addr[46688]= 1844288924;
assign addr[46689]= 1824404752;
assign addr[46690]= 1803941934;
assign addr[46691]= 1782906961;
assign addr[46692]= 1761306505;
assign addr[46693]= 1739147417;
assign addr[46694]= 1716436725;
assign addr[46695]= 1693181631;
assign addr[46696]= 1669389513;
assign addr[46697]= 1645067915;
assign addr[46698]= 1620224553;
assign addr[46699]= 1594867305;
assign addr[46700]= 1569004214;
assign addr[46701]= 1542643483;
assign addr[46702]= 1515793473;
assign addr[46703]= 1488462700;
assign addr[46704]= 1460659832;
assign addr[46705]= 1432393688;
assign addr[46706]= 1403673233;
assign addr[46707]= 1374507575;
assign addr[46708]= 1344905966;
assign addr[46709]= 1314877795;
assign addr[46710]= 1284432584;
assign addr[46711]= 1253579991;
assign addr[46712]= 1222329801;
assign addr[46713]= 1190691925;
assign addr[46714]= 1158676398;
assign addr[46715]= 1126293375;
assign addr[46716]= 1093553126;
assign addr[46717]= 1060466036;
assign addr[46718]= 1027042599;
assign addr[46719]= 993293415;
assign addr[46720]= 959229189;
assign addr[46721]= 924860725;
assign addr[46722]= 890198924;
assign addr[46723]= 855254778;
assign addr[46724]= 820039373;
assign addr[46725]= 784563876;
assign addr[46726]= 748839539;
assign addr[46727]= 712877694;
assign addr[46728]= 676689746;
assign addr[46729]= 640287172;
assign addr[46730]= 603681519;
assign addr[46731]= 566884397;
assign addr[46732]= 529907477;
assign addr[46733]= 492762486;
assign addr[46734]= 455461206;
assign addr[46735]= 418015468;
assign addr[46736]= 380437148;
assign addr[46737]= 342738165;
assign addr[46738]= 304930476;
assign addr[46739]= 267026072;
assign addr[46740]= 229036977;
assign addr[46741]= 190975237;
assign addr[46742]= 152852926;
assign addr[46743]= 114682135;
assign addr[46744]= 76474970;
assign addr[46745]= 38243550;
assign addr[46746]= 0;
assign addr[46747]= -38243550;
assign addr[46748]= -76474970;
assign addr[46749]= -114682135;
assign addr[46750]= -152852926;
assign addr[46751]= -190975237;
assign addr[46752]= -229036977;
assign addr[46753]= -267026072;
assign addr[46754]= -304930476;
assign addr[46755]= -342738165;
assign addr[46756]= -380437148;
assign addr[46757]= -418015468;
assign addr[46758]= -455461206;
assign addr[46759]= -492762486;
assign addr[46760]= -529907477;
assign addr[46761]= -566884397;
assign addr[46762]= -603681519;
assign addr[46763]= -640287172;
assign addr[46764]= -676689746;
assign addr[46765]= -712877694;
assign addr[46766]= -748839539;
assign addr[46767]= -784563876;
assign addr[46768]= -820039373;
assign addr[46769]= -855254778;
assign addr[46770]= -890198924;
assign addr[46771]= -924860725;
assign addr[46772]= -959229189;
assign addr[46773]= -993293415;
assign addr[46774]= -1027042599;
assign addr[46775]= -1060466036;
assign addr[46776]= -1093553126;
assign addr[46777]= -1126293375;
assign addr[46778]= -1158676398;
assign addr[46779]= -1190691925;
assign addr[46780]= -1222329801;
assign addr[46781]= -1253579991;
assign addr[46782]= -1284432584;
assign addr[46783]= -1314877795;
assign addr[46784]= -1344905966;
assign addr[46785]= -1374507575;
assign addr[46786]= -1403673233;
assign addr[46787]= -1432393688;
assign addr[46788]= -1460659832;
assign addr[46789]= -1488462700;
assign addr[46790]= -1515793473;
assign addr[46791]= -1542643483;
assign addr[46792]= -1569004214;
assign addr[46793]= -1594867305;
assign addr[46794]= -1620224553;
assign addr[46795]= -1645067915;
assign addr[46796]= -1669389513;
assign addr[46797]= -1693181631;
assign addr[46798]= -1716436725;
assign addr[46799]= -1739147417;
assign addr[46800]= -1761306505;
assign addr[46801]= -1782906961;
assign addr[46802]= -1803941934;
assign addr[46803]= -1824404752;
assign addr[46804]= -1844288924;
assign addr[46805]= -1863588145;
assign addr[46806]= -1882296293;
assign addr[46807]= -1900407434;
assign addr[46808]= -1917915825;
assign addr[46809]= -1934815911;
assign addr[46810]= -1951102334;
assign addr[46811]= -1966769926;
assign addr[46812]= -1981813720;
assign addr[46813]= -1996228943;
assign addr[46814]= -2010011024;
assign addr[46815]= -2023155591;
assign addr[46816]= -2035658475;
assign addr[46817]= -2047515711;
assign addr[46818]= -2058723538;
assign addr[46819]= -2069278401;
assign addr[46820]= -2079176953;
assign addr[46821]= -2088416053;
assign addr[46822]= -2096992772;
assign addr[46823]= -2104904390;
assign addr[46824]= -2112148396;
assign addr[46825]= -2118722494;
assign addr[46826]= -2124624598;
assign addr[46827]= -2129852837;
assign addr[46828]= -2134405552;
assign addr[46829]= -2138281298;
assign addr[46830]= -2141478848;
assign addr[46831]= -2143997187;
assign addr[46832]= -2145835515;
assign addr[46833]= -2146993250;
assign addr[46834]= -2147470025;
assign addr[46835]= -2147265689;
assign addr[46836]= -2146380306;
assign addr[46837]= -2144814157;
assign addr[46838]= -2142567738;
assign addr[46839]= -2139641764;
assign addr[46840]= -2136037160;
assign addr[46841]= -2131755071;
assign addr[46842]= -2126796855;
assign addr[46843]= -2121164085;
assign addr[46844]= -2114858546;
assign addr[46845]= -2107882239;
assign addr[46846]= -2100237377;
assign addr[46847]= -2091926384;
assign addr[46848]= -2082951896;
assign addr[46849]= -2073316760;
assign addr[46850]= -2063024031;
assign addr[46851]= -2052076975;
assign addr[46852]= -2040479063;
assign addr[46853]= -2028233973;
assign addr[46854]= -2015345591;
assign addr[46855]= -2001818002;
assign addr[46856]= -1987655498;
assign addr[46857]= -1972862571;
assign addr[46858]= -1957443913;
assign addr[46859]= -1941404413;
assign addr[46860]= -1924749160;
assign addr[46861]= -1907483436;
assign addr[46862]= -1889612716;
assign addr[46863]= -1871142669;
assign addr[46864]= -1852079154;
assign addr[46865]= -1832428215;
assign addr[46866]= -1812196087;
assign addr[46867]= -1791389186;
assign addr[46868]= -1770014111;
assign addr[46869]= -1748077642;
assign addr[46870]= -1725586737;
assign addr[46871]= -1702548529;
assign addr[46872]= -1678970324;
assign addr[46873]= -1654859602;
assign addr[46874]= -1630224009;
assign addr[46875]= -1605071359;
assign addr[46876]= -1579409630;
assign addr[46877]= -1553246960;
assign addr[46878]= -1526591649;
assign addr[46879]= -1499452149;
assign addr[46880]= -1471837070;
assign addr[46881]= -1443755168;
assign addr[46882]= -1415215352;
assign addr[46883]= -1386226674;
assign addr[46884]= -1356798326;
assign addr[46885]= -1326939644;
assign addr[46886]= -1296660098;
assign addr[46887]= -1265969291;
assign addr[46888]= -1234876957;
assign addr[46889]= -1203392958;
assign addr[46890]= -1171527280;
assign addr[46891]= -1139290029;
assign addr[46892]= -1106691431;
assign addr[46893]= -1073741824;
assign addr[46894]= -1040451659;
assign addr[46895]= -1006831495;
assign addr[46896]= -972891995;
assign addr[46897]= -938643924;
assign addr[46898]= -904098143;
assign addr[46899]= -869265610;
assign addr[46900]= -834157373;
assign addr[46901]= -798784567;
assign addr[46902]= -763158411;
assign addr[46903]= -727290205;
assign addr[46904]= -691191324;
assign addr[46905]= -654873219;
assign addr[46906]= -618347408;
assign addr[46907]= -581625477;
assign addr[46908]= -544719071;
assign addr[46909]= -507639898;
assign addr[46910]= -470399716;
assign addr[46911]= -433010339;
assign addr[46912]= -395483624;
assign addr[46913]= -357831473;
assign addr[46914]= -320065829;
assign addr[46915]= -282198671;
assign addr[46916]= -244242007;
assign addr[46917]= -206207878;
assign addr[46918]= -168108346;
assign addr[46919]= -129955495;
assign addr[46920]= -91761426;
assign addr[46921]= -53538253;
assign addr[46922]= -15298099;
assign addr[46923]= 22946906;
assign addr[46924]= 61184634;
assign addr[46925]= 99402956;
assign addr[46926]= 137589750;
assign addr[46927]= 175732905;
assign addr[46928]= 213820322;
assign addr[46929]= 251839923;
assign addr[46930]= 289779648;
assign addr[46931]= 327627463;
assign addr[46932]= 365371365;
assign addr[46933]= 402999383;
assign addr[46934]= 440499581;
assign addr[46935]= 477860067;
assign addr[46936]= 515068990;
assign addr[46937]= 552114549;
assign addr[46938]= 588984994;
assign addr[46939]= 625668632;
assign addr[46940]= 662153826;
assign addr[46941]= 698429006;
assign addr[46942]= 734482665;
assign addr[46943]= 770303369;
assign addr[46944]= 805879757;
assign addr[46945]= 841200544;
assign addr[46946]= 876254528;
assign addr[46947]= 911030591;
assign addr[46948]= 945517704;
assign addr[46949]= 979704927;
assign addr[46950]= 1013581418;
assign addr[46951]= 1047136432;
assign addr[46952]= 1080359326;
assign addr[46953]= 1113239564;
assign addr[46954]= 1145766716;
assign addr[46955]= 1177930466;
assign addr[46956]= 1209720613;
assign addr[46957]= 1241127074;
assign addr[46958]= 1272139887;
assign addr[46959]= 1302749217;
assign addr[46960]= 1332945355;
assign addr[46961]= 1362718723;
assign addr[46962]= 1392059879;
assign addr[46963]= 1420959516;
assign addr[46964]= 1449408469;
assign addr[46965]= 1477397714;
assign addr[46966]= 1504918373;
assign addr[46967]= 1531961719;
assign addr[46968]= 1558519173;
assign addr[46969]= 1584582314;
assign addr[46970]= 1610142873;
assign addr[46971]= 1635192744;
assign addr[46972]= 1659723983;
assign addr[46973]= 1683728808;
assign addr[46974]= 1707199606;
assign addr[46975]= 1730128933;
assign addr[46976]= 1752509516;
assign addr[46977]= 1774334257;
assign addr[46978]= 1795596234;
assign addr[46979]= 1816288703;
assign addr[46980]= 1836405100;
assign addr[46981]= 1855939047;
assign addr[46982]= 1874884346;
assign addr[46983]= 1893234990;
assign addr[46984]= 1910985158;
assign addr[46985]= 1928129220;
assign addr[46986]= 1944661739;
assign addr[46987]= 1960577471;
assign addr[46988]= 1975871368;
assign addr[46989]= 1990538579;
assign addr[46990]= 2004574453;
assign addr[46991]= 2017974537;
assign addr[46992]= 2030734582;
assign addr[46993]= 2042850540;
assign addr[46994]= 2054318569;
assign addr[46995]= 2065135031;
assign addr[46996]= 2075296495;
assign addr[46997]= 2084799740;
assign addr[46998]= 2093641749;
assign addr[46999]= 2101819720;
assign addr[47000]= 2109331059;
assign addr[47001]= 2116173382;
assign addr[47002]= 2122344521;
assign addr[47003]= 2127842516;
assign addr[47004]= 2132665626;
assign addr[47005]= 2136812319;
assign addr[47006]= 2140281282;
assign addr[47007]= 2143071413;
assign addr[47008]= 2145181827;
assign addr[47009]= 2146611856;
assign addr[47010]= 2147361045;
assign addr[47011]= 2147429158;
assign addr[47012]= 2146816171;
assign addr[47013]= 2145522281;
assign addr[47014]= 2143547897;
assign addr[47015]= 2140893646;
assign addr[47016]= 2137560369;
assign addr[47017]= 2133549123;
assign addr[47018]= 2128861181;
assign addr[47019]= 2123498030;
assign addr[47020]= 2117461370;
assign addr[47021]= 2110753117;
assign addr[47022]= 2103375398;
assign addr[47023]= 2095330553;
assign addr[47024]= 2086621133;
assign addr[47025]= 2077249901;
assign addr[47026]= 2067219829;
assign addr[47027]= 2056534099;
assign addr[47028]= 2045196100;
assign addr[47029]= 2033209426;
assign addr[47030]= 2020577882;
assign addr[47031]= 2007305472;
assign addr[47032]= 1993396407;
assign addr[47033]= 1978855097;
assign addr[47034]= 1963686155;
assign addr[47035]= 1947894393;
assign addr[47036]= 1931484818;
assign addr[47037]= 1914462636;
assign addr[47038]= 1896833245;
assign addr[47039]= 1878602237;
assign addr[47040]= 1859775393;
assign addr[47041]= 1840358687;
assign addr[47042]= 1820358275;
assign addr[47043]= 1799780501;
assign addr[47044]= 1778631892;
assign addr[47045]= 1756919156;
assign addr[47046]= 1734649179;
assign addr[47047]= 1711829025;
assign addr[47048]= 1688465931;
assign addr[47049]= 1664567307;
assign addr[47050]= 1640140734;
assign addr[47051]= 1615193959;
assign addr[47052]= 1589734894;
assign addr[47053]= 1563771613;
assign addr[47054]= 1537312353;
assign addr[47055]= 1510365504;
assign addr[47056]= 1482939614;
assign addr[47057]= 1455043381;
assign addr[47058]= 1426685652;
assign addr[47059]= 1397875423;
assign addr[47060]= 1368621831;
assign addr[47061]= 1338934154;
assign addr[47062]= 1308821808;
assign addr[47063]= 1278294345;
assign addr[47064]= 1247361445;
assign addr[47065]= 1216032921;
assign addr[47066]= 1184318708;
assign addr[47067]= 1152228866;
assign addr[47068]= 1119773573;
assign addr[47069]= 1086963121;
assign addr[47070]= 1053807919;
assign addr[47071]= 1020318481;
assign addr[47072]= 986505429;
assign addr[47073]= 952379488;
assign addr[47074]= 917951481;
assign addr[47075]= 883232329;
assign addr[47076]= 848233042;
assign addr[47077]= 812964722;
assign addr[47078]= 777438554;
assign addr[47079]= 741665807;
assign addr[47080]= 705657826;
assign addr[47081]= 669426032;
assign addr[47082]= 632981917;
assign addr[47083]= 596337040;
assign addr[47084]= 559503022;
assign addr[47085]= 522491548;
assign addr[47086]= 485314355;
assign addr[47087]= 447983235;
assign addr[47088]= 410510029;
assign addr[47089]= 372906622;
assign addr[47090]= 335184940;
assign addr[47091]= 297356948;
assign addr[47092]= 259434643;
assign addr[47093]= 221430054;
assign addr[47094]= 183355234;
assign addr[47095]= 145222259;
assign addr[47096]= 107043224;
assign addr[47097]= 68830239;
assign addr[47098]= 30595422;
assign addr[47099]= -7649098;
assign addr[47100]= -45891193;
assign addr[47101]= -84118732;
assign addr[47102]= -122319591;
assign addr[47103]= -160481654;
assign addr[47104]= -198592817;
assign addr[47105]= -236640993;
assign addr[47106]= -274614114;
assign addr[47107]= -312500135;
assign addr[47108]= -350287041;
assign addr[47109]= -387962847;
assign addr[47110]= -425515602;
assign addr[47111]= -462933398;
assign addr[47112]= -500204365;
assign addr[47113]= -537316682;
assign addr[47114]= -574258580;
assign addr[47115]= -611018340;
assign addr[47116]= -647584304;
assign addr[47117]= -683944874;
assign addr[47118]= -720088517;
assign addr[47119]= -756003771;
assign addr[47120]= -791679244;
assign addr[47121]= -827103620;
assign addr[47122]= -862265664;
assign addr[47123]= -897154224;
assign addr[47124]= -931758235;
assign addr[47125]= -966066720;
assign addr[47126]= -1000068799;
assign addr[47127]= -1033753687;
assign addr[47128]= -1067110699;
assign addr[47129]= -1100129257;
assign addr[47130]= -1132798888;
assign addr[47131]= -1165109230;
assign addr[47132]= -1197050035;
assign addr[47133]= -1228611172;
assign addr[47134]= -1259782632;
assign addr[47135]= -1290554528;
assign addr[47136]= -1320917099;
assign addr[47137]= -1350860716;
assign addr[47138]= -1380375881;
assign addr[47139]= -1409453233;
assign addr[47140]= -1438083551;
assign addr[47141]= -1466257752;
assign addr[47142]= -1493966902;
assign addr[47143]= -1521202211;
assign addr[47144]= -1547955041;
assign addr[47145]= -1574216908;
assign addr[47146]= -1599979481;
assign addr[47147]= -1625234591;
assign addr[47148]= -1649974225;
assign addr[47149]= -1674190539;
assign addr[47150]= -1697875851;
assign addr[47151]= -1721022648;
assign addr[47152]= -1743623590;
assign addr[47153]= -1765671509;
assign addr[47154]= -1787159411;
assign addr[47155]= -1808080480;
assign addr[47156]= -1828428082;
assign addr[47157]= -1848195763;
assign addr[47158]= -1867377253;
assign addr[47159]= -1885966468;
assign addr[47160]= -1903957513;
assign addr[47161]= -1921344681;
assign addr[47162]= -1938122457;
assign addr[47163]= -1954285520;
assign addr[47164]= -1969828744;
assign addr[47165]= -1984747199;
assign addr[47166]= -1999036154;
assign addr[47167]= -2012691075;
assign addr[47168]= -2025707632;
assign addr[47169]= -2038081698;
assign addr[47170]= -2049809346;
assign addr[47171]= -2060886858;
assign addr[47172]= -2071310720;
assign addr[47173]= -2081077626;
assign addr[47174]= -2090184478;
assign addr[47175]= -2098628387;
assign addr[47176]= -2106406677;
assign addr[47177]= -2113516878;
assign addr[47178]= -2119956737;
assign addr[47179]= -2125724211;
assign addr[47180]= -2130817471;
assign addr[47181]= -2135234901;
assign addr[47182]= -2138975100;
assign addr[47183]= -2142036881;
assign addr[47184]= -2144419275;
assign addr[47185]= -2146121524;
assign addr[47186]= -2147143090;
assign addr[47187]= -2147483648;
assign addr[47188]= -2147143090;
assign addr[47189]= -2146121524;
assign addr[47190]= -2144419275;
assign addr[47191]= -2142036881;
assign addr[47192]= -2138975100;
assign addr[47193]= -2135234901;
assign addr[47194]= -2130817471;
assign addr[47195]= -2125724211;
assign addr[47196]= -2119956737;
assign addr[47197]= -2113516878;
assign addr[47198]= -2106406677;
assign addr[47199]= -2098628387;
assign addr[47200]= -2090184478;
assign addr[47201]= -2081077626;
assign addr[47202]= -2071310720;
assign addr[47203]= -2060886858;
assign addr[47204]= -2049809346;
assign addr[47205]= -2038081698;
assign addr[47206]= -2025707632;
assign addr[47207]= -2012691075;
assign addr[47208]= -1999036154;
assign addr[47209]= -1984747199;
assign addr[47210]= -1969828744;
assign addr[47211]= -1954285520;
assign addr[47212]= -1938122457;
assign addr[47213]= -1921344681;
assign addr[47214]= -1903957513;
assign addr[47215]= -1885966468;
assign addr[47216]= -1867377253;
assign addr[47217]= -1848195763;
assign addr[47218]= -1828428082;
assign addr[47219]= -1808080480;
assign addr[47220]= -1787159411;
assign addr[47221]= -1765671509;
assign addr[47222]= -1743623590;
assign addr[47223]= -1721022648;
assign addr[47224]= -1697875851;
assign addr[47225]= -1674190539;
assign addr[47226]= -1649974225;
assign addr[47227]= -1625234591;
assign addr[47228]= -1599979481;
assign addr[47229]= -1574216908;
assign addr[47230]= -1547955041;
assign addr[47231]= -1521202211;
assign addr[47232]= -1493966902;
assign addr[47233]= -1466257752;
assign addr[47234]= -1438083551;
assign addr[47235]= -1409453233;
assign addr[47236]= -1380375881;
assign addr[47237]= -1350860716;
assign addr[47238]= -1320917099;
assign addr[47239]= -1290554528;
assign addr[47240]= -1259782632;
assign addr[47241]= -1228611172;
assign addr[47242]= -1197050035;
assign addr[47243]= -1165109230;
assign addr[47244]= -1132798888;
assign addr[47245]= -1100129257;
assign addr[47246]= -1067110699;
assign addr[47247]= -1033753687;
assign addr[47248]= -1000068799;
assign addr[47249]= -966066720;
assign addr[47250]= -931758235;
assign addr[47251]= -897154224;
assign addr[47252]= -862265664;
assign addr[47253]= -827103620;
assign addr[47254]= -791679244;
assign addr[47255]= -756003771;
assign addr[47256]= -720088517;
assign addr[47257]= -683944874;
assign addr[47258]= -647584304;
assign addr[47259]= -611018340;
assign addr[47260]= -574258580;
assign addr[47261]= -537316682;
assign addr[47262]= -500204365;
assign addr[47263]= -462933398;
assign addr[47264]= -425515602;
assign addr[47265]= -387962847;
assign addr[47266]= -350287041;
assign addr[47267]= -312500135;
assign addr[47268]= -274614114;
assign addr[47269]= -236640993;
assign addr[47270]= -198592817;
assign addr[47271]= -160481654;
assign addr[47272]= -122319591;
assign addr[47273]= -84118732;
assign addr[47274]= -45891193;
assign addr[47275]= -7649098;
assign addr[47276]= 30595422;
assign addr[47277]= 68830239;
assign addr[47278]= 107043224;
assign addr[47279]= 145222259;
assign addr[47280]= 183355234;
assign addr[47281]= 221430054;
assign addr[47282]= 259434643;
assign addr[47283]= 297356948;
assign addr[47284]= 335184940;
assign addr[47285]= 372906622;
assign addr[47286]= 410510029;
assign addr[47287]= 447983235;
assign addr[47288]= 485314355;
assign addr[47289]= 522491548;
assign addr[47290]= 559503022;
assign addr[47291]= 596337040;
assign addr[47292]= 632981917;
assign addr[47293]= 669426032;
assign addr[47294]= 705657826;
assign addr[47295]= 741665807;
assign addr[47296]= 777438554;
assign addr[47297]= 812964722;
assign addr[47298]= 848233042;
assign addr[47299]= 883232329;
assign addr[47300]= 917951481;
assign addr[47301]= 952379488;
assign addr[47302]= 986505429;
assign addr[47303]= 1020318481;
assign addr[47304]= 1053807919;
assign addr[47305]= 1086963121;
assign addr[47306]= 1119773573;
assign addr[47307]= 1152228866;
assign addr[47308]= 1184318708;
assign addr[47309]= 1216032921;
assign addr[47310]= 1247361445;
assign addr[47311]= 1278294345;
assign addr[47312]= 1308821808;
assign addr[47313]= 1338934154;
assign addr[47314]= 1368621831;
assign addr[47315]= 1397875423;
assign addr[47316]= 1426685652;
assign addr[47317]= 1455043381;
assign addr[47318]= 1482939614;
assign addr[47319]= 1510365504;
assign addr[47320]= 1537312353;
assign addr[47321]= 1563771613;
assign addr[47322]= 1589734894;
assign addr[47323]= 1615193959;
assign addr[47324]= 1640140734;
assign addr[47325]= 1664567307;
assign addr[47326]= 1688465931;
assign addr[47327]= 1711829025;
assign addr[47328]= 1734649179;
assign addr[47329]= 1756919156;
assign addr[47330]= 1778631892;
assign addr[47331]= 1799780501;
assign addr[47332]= 1820358275;
assign addr[47333]= 1840358687;
assign addr[47334]= 1859775393;
assign addr[47335]= 1878602237;
assign addr[47336]= 1896833245;
assign addr[47337]= 1914462636;
assign addr[47338]= 1931484818;
assign addr[47339]= 1947894393;
assign addr[47340]= 1963686155;
assign addr[47341]= 1978855097;
assign addr[47342]= 1993396407;
assign addr[47343]= 2007305472;
assign addr[47344]= 2020577882;
assign addr[47345]= 2033209426;
assign addr[47346]= 2045196100;
assign addr[47347]= 2056534099;
assign addr[47348]= 2067219829;
assign addr[47349]= 2077249901;
assign addr[47350]= 2086621133;
assign addr[47351]= 2095330553;
assign addr[47352]= 2103375398;
assign addr[47353]= 2110753117;
assign addr[47354]= 2117461370;
assign addr[47355]= 2123498030;
assign addr[47356]= 2128861181;
assign addr[47357]= 2133549123;
assign addr[47358]= 2137560369;
assign addr[47359]= 2140893646;
assign addr[47360]= 2143547897;
assign addr[47361]= 2145522281;
assign addr[47362]= 2146816171;
assign addr[47363]= 2147429158;
assign addr[47364]= 2147361045;
assign addr[47365]= 2146611856;
assign addr[47366]= 2145181827;
assign addr[47367]= 2143071413;
assign addr[47368]= 2140281282;
assign addr[47369]= 2136812319;
assign addr[47370]= 2132665626;
assign addr[47371]= 2127842516;
assign addr[47372]= 2122344521;
assign addr[47373]= 2116173382;
assign addr[47374]= 2109331059;
assign addr[47375]= 2101819720;
assign addr[47376]= 2093641749;
assign addr[47377]= 2084799740;
assign addr[47378]= 2075296495;
assign addr[47379]= 2065135031;
assign addr[47380]= 2054318569;
assign addr[47381]= 2042850540;
assign addr[47382]= 2030734582;
assign addr[47383]= 2017974537;
assign addr[47384]= 2004574453;
assign addr[47385]= 1990538579;
assign addr[47386]= 1975871368;
assign addr[47387]= 1960577471;
assign addr[47388]= 1944661739;
assign addr[47389]= 1928129220;
assign addr[47390]= 1910985158;
assign addr[47391]= 1893234990;
assign addr[47392]= 1874884346;
assign addr[47393]= 1855939047;
assign addr[47394]= 1836405100;
assign addr[47395]= 1816288703;
assign addr[47396]= 1795596234;
assign addr[47397]= 1774334257;
assign addr[47398]= 1752509516;
assign addr[47399]= 1730128933;
assign addr[47400]= 1707199606;
assign addr[47401]= 1683728808;
assign addr[47402]= 1659723983;
assign addr[47403]= 1635192744;
assign addr[47404]= 1610142873;
assign addr[47405]= 1584582314;
assign addr[47406]= 1558519173;
assign addr[47407]= 1531961719;
assign addr[47408]= 1504918373;
assign addr[47409]= 1477397714;
assign addr[47410]= 1449408469;
assign addr[47411]= 1420959516;
assign addr[47412]= 1392059879;
assign addr[47413]= 1362718723;
assign addr[47414]= 1332945355;
assign addr[47415]= 1302749217;
assign addr[47416]= 1272139887;
assign addr[47417]= 1241127074;
assign addr[47418]= 1209720613;
assign addr[47419]= 1177930466;
assign addr[47420]= 1145766716;
assign addr[47421]= 1113239564;
assign addr[47422]= 1080359326;
assign addr[47423]= 1047136432;
assign addr[47424]= 1013581418;
assign addr[47425]= 979704927;
assign addr[47426]= 945517704;
assign addr[47427]= 911030591;
assign addr[47428]= 876254528;
assign addr[47429]= 841200544;
assign addr[47430]= 805879757;
assign addr[47431]= 770303369;
assign addr[47432]= 734482665;
assign addr[47433]= 698429006;
assign addr[47434]= 662153826;
assign addr[47435]= 625668632;
assign addr[47436]= 588984994;
assign addr[47437]= 552114549;
assign addr[47438]= 515068990;
assign addr[47439]= 477860067;
assign addr[47440]= 440499581;
assign addr[47441]= 402999383;
assign addr[47442]= 365371365;
assign addr[47443]= 327627463;
assign addr[47444]= 289779648;
assign addr[47445]= 251839923;
assign addr[47446]= 213820322;
assign addr[47447]= 175732905;
assign addr[47448]= 137589750;
assign addr[47449]= 99402956;
assign addr[47450]= 61184634;
assign addr[47451]= 22946906;
assign addr[47452]= -15298099;
assign addr[47453]= -53538253;
assign addr[47454]= -91761426;
assign addr[47455]= -129955495;
assign addr[47456]= -168108346;
assign addr[47457]= -206207878;
assign addr[47458]= -244242007;
assign addr[47459]= -282198671;
assign addr[47460]= -320065829;
assign addr[47461]= -357831473;
assign addr[47462]= -395483624;
assign addr[47463]= -433010339;
assign addr[47464]= -470399716;
assign addr[47465]= -507639898;
assign addr[47466]= -544719071;
assign addr[47467]= -581625477;
assign addr[47468]= -618347408;
assign addr[47469]= -654873219;
assign addr[47470]= -691191324;
assign addr[47471]= -727290205;
assign addr[47472]= -763158411;
assign addr[47473]= -798784567;
assign addr[47474]= -834157373;
assign addr[47475]= -869265610;
assign addr[47476]= -904098143;
assign addr[47477]= -938643924;
assign addr[47478]= -972891995;
assign addr[47479]= -1006831495;
assign addr[47480]= -1040451659;
assign addr[47481]= -1073741824;
assign addr[47482]= -1106691431;
assign addr[47483]= -1139290029;
assign addr[47484]= -1171527280;
assign addr[47485]= -1203392958;
assign addr[47486]= -1234876957;
assign addr[47487]= -1265969291;
assign addr[47488]= -1296660098;
assign addr[47489]= -1326939644;
assign addr[47490]= -1356798326;
assign addr[47491]= -1386226674;
assign addr[47492]= -1415215352;
assign addr[47493]= -1443755168;
assign addr[47494]= -1471837070;
assign addr[47495]= -1499452149;
assign addr[47496]= -1526591649;
assign addr[47497]= -1553246960;
assign addr[47498]= -1579409630;
assign addr[47499]= -1605071359;
assign addr[47500]= -1630224009;
assign addr[47501]= -1654859602;
assign addr[47502]= -1678970324;
assign addr[47503]= -1702548529;
assign addr[47504]= -1725586737;
assign addr[47505]= -1748077642;
assign addr[47506]= -1770014111;
assign addr[47507]= -1791389186;
assign addr[47508]= -1812196087;
assign addr[47509]= -1832428215;
assign addr[47510]= -1852079154;
assign addr[47511]= -1871142669;
assign addr[47512]= -1889612716;
assign addr[47513]= -1907483436;
assign addr[47514]= -1924749160;
assign addr[47515]= -1941404413;
assign addr[47516]= -1957443913;
assign addr[47517]= -1972862571;
assign addr[47518]= -1987655498;
assign addr[47519]= -2001818002;
assign addr[47520]= -2015345591;
assign addr[47521]= -2028233973;
assign addr[47522]= -2040479063;
assign addr[47523]= -2052076975;
assign addr[47524]= -2063024031;
assign addr[47525]= -2073316760;
assign addr[47526]= -2082951896;
assign addr[47527]= -2091926384;
assign addr[47528]= -2100237377;
assign addr[47529]= -2107882239;
assign addr[47530]= -2114858546;
assign addr[47531]= -2121164085;
assign addr[47532]= -2126796855;
assign addr[47533]= -2131755071;
assign addr[47534]= -2136037160;
assign addr[47535]= -2139641764;
assign addr[47536]= -2142567738;
assign addr[47537]= -2144814157;
assign addr[47538]= -2146380306;
assign addr[47539]= -2147265689;
assign addr[47540]= -2147470025;
assign addr[47541]= -2146993250;
assign addr[47542]= -2145835515;
assign addr[47543]= -2143997187;
assign addr[47544]= -2141478848;
assign addr[47545]= -2138281298;
assign addr[47546]= -2134405552;
assign addr[47547]= -2129852837;
assign addr[47548]= -2124624598;
assign addr[47549]= -2118722494;
assign addr[47550]= -2112148396;
assign addr[47551]= -2104904390;
assign addr[47552]= -2096992772;
assign addr[47553]= -2088416053;
assign addr[47554]= -2079176953;
assign addr[47555]= -2069278401;
assign addr[47556]= -2058723538;
assign addr[47557]= -2047515711;
assign addr[47558]= -2035658475;
assign addr[47559]= -2023155591;
assign addr[47560]= -2010011024;
assign addr[47561]= -1996228943;
assign addr[47562]= -1981813720;
assign addr[47563]= -1966769926;
assign addr[47564]= -1951102334;
assign addr[47565]= -1934815911;
assign addr[47566]= -1917915825;
assign addr[47567]= -1900407434;
assign addr[47568]= -1882296293;
assign addr[47569]= -1863588145;
assign addr[47570]= -1844288924;
assign addr[47571]= -1824404752;
assign addr[47572]= -1803941934;
assign addr[47573]= -1782906961;
assign addr[47574]= -1761306505;
assign addr[47575]= -1739147417;
assign addr[47576]= -1716436725;
assign addr[47577]= -1693181631;
assign addr[47578]= -1669389513;
assign addr[47579]= -1645067915;
assign addr[47580]= -1620224553;
assign addr[47581]= -1594867305;
assign addr[47582]= -1569004214;
assign addr[47583]= -1542643483;
assign addr[47584]= -1515793473;
assign addr[47585]= -1488462700;
assign addr[47586]= -1460659832;
assign addr[47587]= -1432393688;
assign addr[47588]= -1403673233;
assign addr[47589]= -1374507575;
assign addr[47590]= -1344905966;
assign addr[47591]= -1314877795;
assign addr[47592]= -1284432584;
assign addr[47593]= -1253579991;
assign addr[47594]= -1222329801;
assign addr[47595]= -1190691925;
assign addr[47596]= -1158676398;
assign addr[47597]= -1126293375;
assign addr[47598]= -1093553126;
assign addr[47599]= -1060466036;
assign addr[47600]= -1027042599;
assign addr[47601]= -993293415;
assign addr[47602]= -959229189;
assign addr[47603]= -924860725;
assign addr[47604]= -890198924;
assign addr[47605]= -855254778;
assign addr[47606]= -820039373;
assign addr[47607]= -784563876;
assign addr[47608]= -748839539;
assign addr[47609]= -712877694;
assign addr[47610]= -676689746;
assign addr[47611]= -640287172;
assign addr[47612]= -603681519;
assign addr[47613]= -566884397;
assign addr[47614]= -529907477;
assign addr[47615]= -492762486;
assign addr[47616]= -455461206;
assign addr[47617]= -418015468;
assign addr[47618]= -380437148;
assign addr[47619]= -342738165;
assign addr[47620]= -304930476;
assign addr[47621]= -267026072;
assign addr[47622]= -229036977;
assign addr[47623]= -190975237;
assign addr[47624]= -152852926;
assign addr[47625]= -114682135;
assign addr[47626]= -76474970;
assign addr[47627]= -38243550;
assign addr[47628]= 0;
assign addr[47629]= 38243550;
assign addr[47630]= 76474970;
assign addr[47631]= 114682135;
assign addr[47632]= 152852926;
assign addr[47633]= 190975237;
assign addr[47634]= 229036977;
assign addr[47635]= 267026072;
assign addr[47636]= 304930476;
assign addr[47637]= 342738165;
assign addr[47638]= 380437148;
assign addr[47639]= 418015468;
assign addr[47640]= 455461206;
assign addr[47641]= 492762486;
assign addr[47642]= 529907477;
assign addr[47643]= 566884397;
assign addr[47644]= 603681519;
assign addr[47645]= 640287172;
assign addr[47646]= 676689746;
assign addr[47647]= 712877694;
assign addr[47648]= 748839539;
assign addr[47649]= 784563876;
assign addr[47650]= 820039373;
assign addr[47651]= 855254778;
assign addr[47652]= 890198924;
assign addr[47653]= 924860725;
assign addr[47654]= 959229189;
assign addr[47655]= 993293415;
assign addr[47656]= 1027042599;
assign addr[47657]= 1060466036;
assign addr[47658]= 1093553126;
assign addr[47659]= 1126293375;
assign addr[47660]= 1158676398;
assign addr[47661]= 1190691925;
assign addr[47662]= 1222329801;
assign addr[47663]= 1253579991;
assign addr[47664]= 1284432584;
assign addr[47665]= 1314877795;
assign addr[47666]= 1344905966;
assign addr[47667]= 1374507575;
assign addr[47668]= 1403673233;
assign addr[47669]= 1432393688;
assign addr[47670]= 1460659832;
assign addr[47671]= 1488462700;
assign addr[47672]= 1515793473;
assign addr[47673]= 1542643483;
assign addr[47674]= 1569004214;
assign addr[47675]= 1594867305;
assign addr[47676]= 1620224553;
assign addr[47677]= 1645067915;
assign addr[47678]= 1669389513;
assign addr[47679]= 1693181631;
assign addr[47680]= 1716436725;
assign addr[47681]= 1739147417;
assign addr[47682]= 1761306505;
assign addr[47683]= 1782906961;
assign addr[47684]= 1803941934;
assign addr[47685]= 1824404752;
assign addr[47686]= 1844288924;
assign addr[47687]= 1863588145;
assign addr[47688]= 1882296293;
assign addr[47689]= 1900407434;
assign addr[47690]= 1917915825;
assign addr[47691]= 1934815911;
assign addr[47692]= 1951102334;
assign addr[47693]= 1966769926;
assign addr[47694]= 1981813720;
assign addr[47695]= 1996228943;
assign addr[47696]= 2010011024;
assign addr[47697]= 2023155591;
assign addr[47698]= 2035658475;
assign addr[47699]= 2047515711;
assign addr[47700]= 2058723538;
assign addr[47701]= 2069278401;
assign addr[47702]= 2079176953;
assign addr[47703]= 2088416053;
assign addr[47704]= 2096992772;
assign addr[47705]= 2104904390;
assign addr[47706]= 2112148396;
assign addr[47707]= 2118722494;
assign addr[47708]= 2124624598;
assign addr[47709]= 2129852837;
assign addr[47710]= 2134405552;
assign addr[47711]= 2138281298;
assign addr[47712]= 2141478848;
assign addr[47713]= 2143997187;
assign addr[47714]= 2145835515;
assign addr[47715]= 2146993250;
assign addr[47716]= 2147470025;
assign addr[47717]= 2147265689;
assign addr[47718]= 2146380306;
assign addr[47719]= 2144814157;
assign addr[47720]= 2142567738;
assign addr[47721]= 2139641764;
assign addr[47722]= 2136037160;
assign addr[47723]= 2131755071;
assign addr[47724]= 2126796855;
assign addr[47725]= 2121164085;
assign addr[47726]= 2114858546;
assign addr[47727]= 2107882239;
assign addr[47728]= 2100237377;
assign addr[47729]= 2091926384;
assign addr[47730]= 2082951896;
assign addr[47731]= 2073316760;
assign addr[47732]= 2063024031;
assign addr[47733]= 2052076975;
assign addr[47734]= 2040479063;
assign addr[47735]= 2028233973;
assign addr[47736]= 2015345591;
assign addr[47737]= 2001818002;
assign addr[47738]= 1987655498;
assign addr[47739]= 1972862571;
assign addr[47740]= 1957443913;
assign addr[47741]= 1941404413;
assign addr[47742]= 1924749160;
assign addr[47743]= 1907483436;
assign addr[47744]= 1889612716;
assign addr[47745]= 1871142669;
assign addr[47746]= 1852079154;
assign addr[47747]= 1832428215;
assign addr[47748]= 1812196087;
assign addr[47749]= 1791389186;
assign addr[47750]= 1770014111;
assign addr[47751]= 1748077642;
assign addr[47752]= 1725586737;
assign addr[47753]= 1702548529;
assign addr[47754]= 1678970324;
assign addr[47755]= 1654859602;
assign addr[47756]= 1630224009;
assign addr[47757]= 1605071359;
assign addr[47758]= 1579409630;
assign addr[47759]= 1553246960;
assign addr[47760]= 1526591649;
assign addr[47761]= 1499452149;
assign addr[47762]= 1471837070;
assign addr[47763]= 1443755168;
assign addr[47764]= 1415215352;
assign addr[47765]= 1386226674;
assign addr[47766]= 1356798326;
assign addr[47767]= 1326939644;
assign addr[47768]= 1296660098;
assign addr[47769]= 1265969291;
assign addr[47770]= 1234876957;
assign addr[47771]= 1203392958;
assign addr[47772]= 1171527280;
assign addr[47773]= 1139290029;
assign addr[47774]= 1106691431;
assign addr[47775]= 1073741824;
assign addr[47776]= 1040451659;
assign addr[47777]= 1006831495;
assign addr[47778]= 972891995;
assign addr[47779]= 938643924;
assign addr[47780]= 904098143;
assign addr[47781]= 869265610;
assign addr[47782]= 834157373;
assign addr[47783]= 798784567;
assign addr[47784]= 763158411;
assign addr[47785]= 727290205;
assign addr[47786]= 691191324;
assign addr[47787]= 654873219;
assign addr[47788]= 618347408;
assign addr[47789]= 581625477;
assign addr[47790]= 544719071;
assign addr[47791]= 507639898;
assign addr[47792]= 470399716;
assign addr[47793]= 433010339;
assign addr[47794]= 395483624;
assign addr[47795]= 357831473;
assign addr[47796]= 320065829;
assign addr[47797]= 282198671;
assign addr[47798]= 244242007;
assign addr[47799]= 206207878;
assign addr[47800]= 168108346;
assign addr[47801]= 129955495;
assign addr[47802]= 91761426;
assign addr[47803]= 53538253;
assign addr[47804]= 15298099;
assign addr[47805]= -22946906;
assign addr[47806]= -61184634;
assign addr[47807]= -99402956;
assign addr[47808]= -137589750;
assign addr[47809]= -175732905;
assign addr[47810]= -213820322;
assign addr[47811]= -251839923;
assign addr[47812]= -289779648;
assign addr[47813]= -327627463;
assign addr[47814]= -365371365;
assign addr[47815]= -402999383;
assign addr[47816]= -440499581;
assign addr[47817]= -477860067;
assign addr[47818]= -515068990;
assign addr[47819]= -552114549;
assign addr[47820]= -588984994;
assign addr[47821]= -625668632;
assign addr[47822]= -662153826;
assign addr[47823]= -698429006;
assign addr[47824]= -734482665;
assign addr[47825]= -770303369;
assign addr[47826]= -805879757;
assign addr[47827]= -841200544;
assign addr[47828]= -876254528;
assign addr[47829]= -911030591;
assign addr[47830]= -945517704;
assign addr[47831]= -979704927;
assign addr[47832]= -1013581418;
assign addr[47833]= -1047136432;
assign addr[47834]= -1080359326;
assign addr[47835]= -1113239564;
assign addr[47836]= -1145766716;
assign addr[47837]= -1177930466;
assign addr[47838]= -1209720613;
assign addr[47839]= -1241127074;
assign addr[47840]= -1272139887;
assign addr[47841]= -1302749217;
assign addr[47842]= -1332945355;
assign addr[47843]= -1362718723;
assign addr[47844]= -1392059879;
assign addr[47845]= -1420959516;
assign addr[47846]= -1449408469;
assign addr[47847]= -1477397714;
assign addr[47848]= -1504918373;
assign addr[47849]= -1531961719;
assign addr[47850]= -1558519173;
assign addr[47851]= -1584582314;
assign addr[47852]= -1610142873;
assign addr[47853]= -1635192744;
assign addr[47854]= -1659723983;
assign addr[47855]= -1683728808;
assign addr[47856]= -1707199606;
assign addr[47857]= -1730128933;
assign addr[47858]= -1752509516;
assign addr[47859]= -1774334257;
assign addr[47860]= -1795596234;
assign addr[47861]= -1816288703;
assign addr[47862]= -1836405100;
assign addr[47863]= -1855939047;
assign addr[47864]= -1874884346;
assign addr[47865]= -1893234990;
assign addr[47866]= -1910985158;
assign addr[47867]= -1928129220;
assign addr[47868]= -1944661739;
assign addr[47869]= -1960577471;
assign addr[47870]= -1975871368;
assign addr[47871]= -1990538579;
assign addr[47872]= -2004574453;
assign addr[47873]= -2017974537;
assign addr[47874]= -2030734582;
assign addr[47875]= -2042850540;
assign addr[47876]= -2054318569;
assign addr[47877]= -2065135031;
assign addr[47878]= -2075296495;
assign addr[47879]= -2084799740;
assign addr[47880]= -2093641749;
assign addr[47881]= -2101819720;
assign addr[47882]= -2109331059;
assign addr[47883]= -2116173382;
assign addr[47884]= -2122344521;
assign addr[47885]= -2127842516;
assign addr[47886]= -2132665626;
assign addr[47887]= -2136812319;
assign addr[47888]= -2140281282;
assign addr[47889]= -2143071413;
assign addr[47890]= -2145181827;
assign addr[47891]= -2146611856;
assign addr[47892]= -2147361045;
assign addr[47893]= -2147429158;
assign addr[47894]= -2146816171;
assign addr[47895]= -2145522281;
assign addr[47896]= -2143547897;
assign addr[47897]= -2140893646;
assign addr[47898]= -2137560369;
assign addr[47899]= -2133549123;
assign addr[47900]= -2128861181;
assign addr[47901]= -2123498030;
assign addr[47902]= -2117461370;
assign addr[47903]= -2110753117;
assign addr[47904]= -2103375398;
assign addr[47905]= -2095330553;
assign addr[47906]= -2086621133;
assign addr[47907]= -2077249901;
assign addr[47908]= -2067219829;
assign addr[47909]= -2056534099;
assign addr[47910]= -2045196100;
assign addr[47911]= -2033209426;
assign addr[47912]= -2020577882;
assign addr[47913]= -2007305472;
assign addr[47914]= -1993396407;
assign addr[47915]= -1978855097;
assign addr[47916]= -1963686155;
assign addr[47917]= -1947894393;
assign addr[47918]= -1931484818;
assign addr[47919]= -1914462636;
assign addr[47920]= -1896833245;
assign addr[47921]= -1878602237;
assign addr[47922]= -1859775393;
assign addr[47923]= -1840358687;
assign addr[47924]= -1820358275;
assign addr[47925]= -1799780501;
assign addr[47926]= -1778631892;
assign addr[47927]= -1756919156;
assign addr[47928]= -1734649179;
assign addr[47929]= -1711829025;
assign addr[47930]= -1688465931;
assign addr[47931]= -1664567307;
assign addr[47932]= -1640140734;
assign addr[47933]= -1615193959;
assign addr[47934]= -1589734894;
assign addr[47935]= -1563771613;
assign addr[47936]= -1537312353;
assign addr[47937]= -1510365504;
assign addr[47938]= -1482939614;
assign addr[47939]= -1455043381;
assign addr[47940]= -1426685652;
assign addr[47941]= -1397875423;
assign addr[47942]= -1368621831;
assign addr[47943]= -1338934154;
assign addr[47944]= -1308821808;
assign addr[47945]= -1278294345;
assign addr[47946]= -1247361445;
assign addr[47947]= -1216032921;
assign addr[47948]= -1184318708;
assign addr[47949]= -1152228866;
assign addr[47950]= -1119773573;
assign addr[47951]= -1086963121;
assign addr[47952]= -1053807919;
assign addr[47953]= -1020318481;
assign addr[47954]= -986505429;
assign addr[47955]= -952379488;
assign addr[47956]= -917951481;
assign addr[47957]= -883232329;
assign addr[47958]= -848233042;
assign addr[47959]= -812964722;
assign addr[47960]= -777438554;
assign addr[47961]= -741665807;
assign addr[47962]= -705657826;
assign addr[47963]= -669426032;
assign addr[47964]= -632981917;
assign addr[47965]= -596337040;
assign addr[47966]= -559503022;
assign addr[47967]= -522491548;
assign addr[47968]= -485314355;
assign addr[47969]= -447983235;
assign addr[47970]= -410510029;
assign addr[47971]= -372906622;
assign addr[47972]= -335184940;
assign addr[47973]= -297356948;
assign addr[47974]= -259434643;
assign addr[47975]= -221430054;
assign addr[47976]= -183355234;
assign addr[47977]= -145222259;
assign addr[47978]= -107043224;
assign addr[47979]= -68830239;
assign addr[47980]= -30595422;
assign addr[47981]= 7649098;
assign addr[47982]= 45891193;
assign addr[47983]= 84118732;
assign addr[47984]= 122319591;
assign addr[47985]= 160481654;
assign addr[47986]= 198592817;
assign addr[47987]= 236640993;
assign addr[47988]= 274614114;
assign addr[47989]= 312500135;
assign addr[47990]= 350287041;
assign addr[47991]= 387962847;
assign addr[47992]= 425515602;
assign addr[47993]= 462933398;
assign addr[47994]= 500204365;
assign addr[47995]= 537316682;
assign addr[47996]= 574258580;
assign addr[47997]= 611018340;
assign addr[47998]= 647584304;
assign addr[47999]= 683944874;
assign addr[48000]= 720088517;
assign addr[48001]= 756003771;
assign addr[48002]= 791679244;
assign addr[48003]= 827103620;
assign addr[48004]= 862265664;
assign addr[48005]= 897154224;
assign addr[48006]= 931758235;
assign addr[48007]= 966066720;
assign addr[48008]= 1000068799;
assign addr[48009]= 1033753687;
assign addr[48010]= 1067110699;
assign addr[48011]= 1100129257;
assign addr[48012]= 1132798888;
assign addr[48013]= 1165109230;
assign addr[48014]= 1197050035;
assign addr[48015]= 1228611172;
assign addr[48016]= 1259782632;
assign addr[48017]= 1290554528;
assign addr[48018]= 1320917099;
assign addr[48019]= 1350860716;
assign addr[48020]= 1380375881;
assign addr[48021]= 1409453233;
assign addr[48022]= 1438083551;
assign addr[48023]= 1466257752;
assign addr[48024]= 1493966902;
assign addr[48025]= 1521202211;
assign addr[48026]= 1547955041;
assign addr[48027]= 1574216908;
assign addr[48028]= 1599979481;
assign addr[48029]= 1625234591;
assign addr[48030]= 1649974225;
assign addr[48031]= 1674190539;
assign addr[48032]= 1697875851;
assign addr[48033]= 1721022648;
assign addr[48034]= 1743623590;
assign addr[48035]= 1765671509;
assign addr[48036]= 1787159411;
assign addr[48037]= 1808080480;
assign addr[48038]= 1828428082;
assign addr[48039]= 1848195763;
assign addr[48040]= 1867377253;
assign addr[48041]= 1885966468;
assign addr[48042]= 1903957513;
assign addr[48043]= 1921344681;
assign addr[48044]= 1938122457;
assign addr[48045]= 1954285520;
assign addr[48046]= 1969828744;
assign addr[48047]= 1984747199;
assign addr[48048]= 1999036154;
assign addr[48049]= 2012691075;
assign addr[48050]= 2025707632;
assign addr[48051]= 2038081698;
assign addr[48052]= 2049809346;
assign addr[48053]= 2060886858;
assign addr[48054]= 2071310720;
assign addr[48055]= 2081077626;
assign addr[48056]= 2090184478;
assign addr[48057]= 2098628387;
assign addr[48058]= 2106406677;
assign addr[48059]= 2113516878;
assign addr[48060]= 2119956737;
assign addr[48061]= 2125724211;
assign addr[48062]= 2130817471;
assign addr[48063]= 2135234901;
assign addr[48064]= 2138975100;
assign addr[48065]= 2142036881;
assign addr[48066]= 2144419275;
assign addr[48067]= 2146121524;
assign addr[48068]= 2147143090;
assign addr[48069]= 2147483648;
assign addr[48070]= 2147143090;
assign addr[48071]= 2146121524;
assign addr[48072]= 2144419275;
assign addr[48073]= 2142036881;
assign addr[48074]= 2138975100;
assign addr[48075]= 2135234901;
assign addr[48076]= 2130817471;
assign addr[48077]= 2125724211;
assign addr[48078]= 2119956737;
assign addr[48079]= 2113516878;
assign addr[48080]= 2106406677;
assign addr[48081]= 2098628387;
assign addr[48082]= 2090184478;
assign addr[48083]= 2081077626;
assign addr[48084]= 2071310720;
assign addr[48085]= 2060886858;
assign addr[48086]= 2049809346;
assign addr[48087]= 2038081698;
assign addr[48088]= 2025707632;
assign addr[48089]= 2012691075;
assign addr[48090]= 1999036154;
assign addr[48091]= 1984747199;
assign addr[48092]= 1969828744;
assign addr[48093]= 1954285520;
assign addr[48094]= 1938122457;
assign addr[48095]= 1921344681;
assign addr[48096]= 1903957513;
assign addr[48097]= 1885966468;
assign addr[48098]= 1867377253;
assign addr[48099]= 1848195763;
assign addr[48100]= 1828428082;
assign addr[48101]= 1808080480;
assign addr[48102]= 1787159411;
assign addr[48103]= 1765671509;
assign addr[48104]= 1743623590;
assign addr[48105]= 1721022648;
assign addr[48106]= 1697875851;
assign addr[48107]= 1674190539;
assign addr[48108]= 1649974225;
assign addr[48109]= 1625234591;
assign addr[48110]= 1599979481;
assign addr[48111]= 1574216908;
assign addr[48112]= 1547955041;
assign addr[48113]= 1521202211;
assign addr[48114]= 1493966902;
assign addr[48115]= 1466257752;
assign addr[48116]= 1438083551;
assign addr[48117]= 1409453233;
assign addr[48118]= 1380375881;
assign addr[48119]= 1350860716;
assign addr[48120]= 1320917099;
assign addr[48121]= 1290554528;
assign addr[48122]= 1259782632;
assign addr[48123]= 1228611172;
assign addr[48124]= 1197050035;
assign addr[48125]= 1165109230;
assign addr[48126]= 1132798888;
assign addr[48127]= 1100129257;
assign addr[48128]= 1067110699;
assign addr[48129]= 1033753687;
assign addr[48130]= 1000068799;
assign addr[48131]= 966066720;
assign addr[48132]= 931758235;
assign addr[48133]= 897154224;
assign addr[48134]= 862265664;
assign addr[48135]= 827103620;
assign addr[48136]= 791679244;
assign addr[48137]= 756003771;
assign addr[48138]= 720088517;
assign addr[48139]= 683944874;
assign addr[48140]= 647584304;
assign addr[48141]= 611018340;
assign addr[48142]= 574258580;
assign addr[48143]= 537316682;
assign addr[48144]= 500204365;
assign addr[48145]= 462933398;
assign addr[48146]= 425515602;
assign addr[48147]= 387962847;
assign addr[48148]= 350287041;
assign addr[48149]= 312500135;
assign addr[48150]= 274614114;
assign addr[48151]= 236640993;
assign addr[48152]= 198592817;
assign addr[48153]= 160481654;
assign addr[48154]= 122319591;
assign addr[48155]= 84118732;
assign addr[48156]= 45891193;
assign addr[48157]= 7649098;
assign addr[48158]= -30595422;
assign addr[48159]= -68830239;
assign addr[48160]= -107043224;
assign addr[48161]= -145222259;
assign addr[48162]= -183355234;
assign addr[48163]= -221430054;
assign addr[48164]= -259434643;
assign addr[48165]= -297356948;
assign addr[48166]= -335184940;
assign addr[48167]= -372906622;
assign addr[48168]= -410510029;
assign addr[48169]= -447983235;
assign addr[48170]= -485314355;
assign addr[48171]= -522491548;
assign addr[48172]= -559503022;
assign addr[48173]= -596337040;
assign addr[48174]= -632981917;
assign addr[48175]= -669426032;
assign addr[48176]= -705657826;
assign addr[48177]= -741665807;
assign addr[48178]= -777438554;
assign addr[48179]= -812964722;
assign addr[48180]= -848233042;
assign addr[48181]= -883232329;
assign addr[48182]= -917951481;
assign addr[48183]= -952379488;
assign addr[48184]= -986505429;
assign addr[48185]= -1020318481;
assign addr[48186]= -1053807919;
assign addr[48187]= -1086963121;
assign addr[48188]= -1119773573;
assign addr[48189]= -1152228866;
assign addr[48190]= -1184318708;
assign addr[48191]= -1216032921;
assign addr[48192]= -1247361445;
assign addr[48193]= -1278294345;
assign addr[48194]= -1308821808;
assign addr[48195]= -1338934154;
assign addr[48196]= -1368621831;
assign addr[48197]= -1397875423;
assign addr[48198]= -1426685652;
assign addr[48199]= -1455043381;
assign addr[48200]= -1482939614;
assign addr[48201]= -1510365504;
assign addr[48202]= -1537312353;
assign addr[48203]= -1563771613;
assign addr[48204]= -1589734894;
assign addr[48205]= -1615193959;
assign addr[48206]= -1640140734;
assign addr[48207]= -1664567307;
assign addr[48208]= -1688465931;
assign addr[48209]= -1711829025;
assign addr[48210]= -1734649179;
assign addr[48211]= -1756919156;
assign addr[48212]= -1778631892;
assign addr[48213]= -1799780501;
assign addr[48214]= -1820358275;
assign addr[48215]= -1840358687;
assign addr[48216]= -1859775393;
assign addr[48217]= -1878602237;
assign addr[48218]= -1896833245;
assign addr[48219]= -1914462636;
assign addr[48220]= -1931484818;
assign addr[48221]= -1947894393;
assign addr[48222]= -1963686155;
assign addr[48223]= -1978855097;
assign addr[48224]= -1993396407;
assign addr[48225]= -2007305472;
assign addr[48226]= -2020577882;
assign addr[48227]= -2033209426;
assign addr[48228]= -2045196100;
assign addr[48229]= -2056534099;
assign addr[48230]= -2067219829;
assign addr[48231]= -2077249901;
assign addr[48232]= -2086621133;
assign addr[48233]= -2095330553;
assign addr[48234]= -2103375398;
assign addr[48235]= -2110753117;
assign addr[48236]= -2117461370;
assign addr[48237]= -2123498030;
assign addr[48238]= -2128861181;
assign addr[48239]= -2133549123;
assign addr[48240]= -2137560369;
assign addr[48241]= -2140893646;
assign addr[48242]= -2143547897;
assign addr[48243]= -2145522281;
assign addr[48244]= -2146816171;
assign addr[48245]= -2147429158;
assign addr[48246]= -2147361045;
assign addr[48247]= -2146611856;
assign addr[48248]= -2145181827;
assign addr[48249]= -2143071413;
assign addr[48250]= -2140281282;
assign addr[48251]= -2136812319;
assign addr[48252]= -2132665626;
assign addr[48253]= -2127842516;
assign addr[48254]= -2122344521;
assign addr[48255]= -2116173382;
assign addr[48256]= -2109331059;
assign addr[48257]= -2101819720;
assign addr[48258]= -2093641749;
assign addr[48259]= -2084799740;
assign addr[48260]= -2075296495;
assign addr[48261]= -2065135031;
assign addr[48262]= -2054318569;
assign addr[48263]= -2042850540;
assign addr[48264]= -2030734582;
assign addr[48265]= -2017974537;
assign addr[48266]= -2004574453;
assign addr[48267]= -1990538579;
assign addr[48268]= -1975871368;
assign addr[48269]= -1960577471;
assign addr[48270]= -1944661739;
assign addr[48271]= -1928129220;
assign addr[48272]= -1910985158;
assign addr[48273]= -1893234990;
assign addr[48274]= -1874884346;
assign addr[48275]= -1855939047;
assign addr[48276]= -1836405100;
assign addr[48277]= -1816288703;
assign addr[48278]= -1795596234;
assign addr[48279]= -1774334257;
assign addr[48280]= -1752509516;
assign addr[48281]= -1730128933;
assign addr[48282]= -1707199606;
assign addr[48283]= -1683728808;
assign addr[48284]= -1659723983;
assign addr[48285]= -1635192744;
assign addr[48286]= -1610142873;
assign addr[48287]= -1584582314;
assign addr[48288]= -1558519173;
assign addr[48289]= -1531961719;
assign addr[48290]= -1504918373;
assign addr[48291]= -1477397714;
assign addr[48292]= -1449408469;
assign addr[48293]= -1420959516;
assign addr[48294]= -1392059879;
assign addr[48295]= -1362718723;
assign addr[48296]= -1332945355;
assign addr[48297]= -1302749217;
assign addr[48298]= -1272139887;
assign addr[48299]= -1241127074;
assign addr[48300]= -1209720613;
assign addr[48301]= -1177930466;
assign addr[48302]= -1145766716;
assign addr[48303]= -1113239564;
assign addr[48304]= -1080359326;
assign addr[48305]= -1047136432;
assign addr[48306]= -1013581418;
assign addr[48307]= -979704927;
assign addr[48308]= -945517704;
assign addr[48309]= -911030591;
assign addr[48310]= -876254528;
assign addr[48311]= -841200544;
assign addr[48312]= -805879757;
assign addr[48313]= -770303369;
assign addr[48314]= -734482665;
assign addr[48315]= -698429006;
assign addr[48316]= -662153826;
assign addr[48317]= -625668632;
assign addr[48318]= -588984994;
assign addr[48319]= -552114549;
assign addr[48320]= -515068990;
assign addr[48321]= -477860067;
assign addr[48322]= -440499581;
assign addr[48323]= -402999383;
assign addr[48324]= -365371365;
assign addr[48325]= -327627463;
assign addr[48326]= -289779648;
assign addr[48327]= -251839923;
assign addr[48328]= -213820322;
assign addr[48329]= -175732905;
assign addr[48330]= -137589750;
assign addr[48331]= -99402956;
assign addr[48332]= -61184634;
assign addr[48333]= -22946906;
assign addr[48334]= 15298099;
assign addr[48335]= 53538253;
assign addr[48336]= 91761426;
assign addr[48337]= 129955495;
assign addr[48338]= 168108346;
assign addr[48339]= 206207878;
assign addr[48340]= 244242007;
assign addr[48341]= 282198671;
assign addr[48342]= 320065829;
assign addr[48343]= 357831473;
assign addr[48344]= 395483624;
assign addr[48345]= 433010339;
assign addr[48346]= 470399716;
assign addr[48347]= 507639898;
assign addr[48348]= 544719071;
assign addr[48349]= 581625477;
assign addr[48350]= 618347408;
assign addr[48351]= 654873219;
assign addr[48352]= 691191324;
assign addr[48353]= 727290205;
assign addr[48354]= 763158411;
assign addr[48355]= 798784567;
assign addr[48356]= 834157373;
assign addr[48357]= 869265610;
assign addr[48358]= 904098143;
assign addr[48359]= 938643924;
assign addr[48360]= 972891995;
assign addr[48361]= 1006831495;
assign addr[48362]= 1040451659;
assign addr[48363]= 1073741824;
assign addr[48364]= 1106691431;
assign addr[48365]= 1139290029;
assign addr[48366]= 1171527280;
assign addr[48367]= 1203392958;
assign addr[48368]= 1234876957;
assign addr[48369]= 1265969291;
assign addr[48370]= 1296660098;
assign addr[48371]= 1326939644;
assign addr[48372]= 1356798326;
assign addr[48373]= 1386226674;
assign addr[48374]= 1415215352;
assign addr[48375]= 1443755168;
assign addr[48376]= 1471837070;
assign addr[48377]= 1499452149;
assign addr[48378]= 1526591649;
assign addr[48379]= 1553246960;
assign addr[48380]= 1579409630;
assign addr[48381]= 1605071359;
assign addr[48382]= 1630224009;
assign addr[48383]= 1654859602;
assign addr[48384]= 1678970324;
assign addr[48385]= 1702548529;
assign addr[48386]= 1725586737;
assign addr[48387]= 1748077642;
assign addr[48388]= 1770014111;
assign addr[48389]= 1791389186;
assign addr[48390]= 1812196087;
assign addr[48391]= 1832428215;
assign addr[48392]= 1852079154;
assign addr[48393]= 1871142669;
assign addr[48394]= 1889612716;
assign addr[48395]= 1907483436;
assign addr[48396]= 1924749160;
assign addr[48397]= 1941404413;
assign addr[48398]= 1957443913;
assign addr[48399]= 1972862571;
assign addr[48400]= 1987655498;
assign addr[48401]= 2001818002;
assign addr[48402]= 2015345591;
assign addr[48403]= 2028233973;
assign addr[48404]= 2040479063;
assign addr[48405]= 2052076975;
assign addr[48406]= 2063024031;
assign addr[48407]= 2073316760;
assign addr[48408]= 2082951896;
assign addr[48409]= 2091926384;
assign addr[48410]= 2100237377;
assign addr[48411]= 2107882239;
assign addr[48412]= 2114858546;
assign addr[48413]= 2121164085;
assign addr[48414]= 2126796855;
assign addr[48415]= 2131755071;
assign addr[48416]= 2136037160;
assign addr[48417]= 2139641764;
assign addr[48418]= 2142567738;
assign addr[48419]= 2144814157;
assign addr[48420]= 2146380306;
assign addr[48421]= 2147265689;
assign addr[48422]= 2147470025;
assign addr[48423]= 2146993250;
assign addr[48424]= 2145835515;
assign addr[48425]= 2143997187;
assign addr[48426]= 2141478848;
assign addr[48427]= 2138281298;
assign addr[48428]= 2134405552;
assign addr[48429]= 2129852837;
assign addr[48430]= 2124624598;
assign addr[48431]= 2118722494;
assign addr[48432]= 2112148396;
assign addr[48433]= 2104904390;
assign addr[48434]= 2096992772;
assign addr[48435]= 2088416053;
assign addr[48436]= 2079176953;
assign addr[48437]= 2069278401;
assign addr[48438]= 2058723538;
assign addr[48439]= 2047515711;
assign addr[48440]= 2035658475;
assign addr[48441]= 2023155591;
assign addr[48442]= 2010011024;
assign addr[48443]= 1996228943;
assign addr[48444]= 1981813720;
assign addr[48445]= 1966769926;
assign addr[48446]= 1951102334;
assign addr[48447]= 1934815911;
assign addr[48448]= 1917915825;
assign addr[48449]= 1900407434;
assign addr[48450]= 1882296293;
assign addr[48451]= 1863588145;
assign addr[48452]= 1844288924;
assign addr[48453]= 1824404752;
assign addr[48454]= 1803941934;
assign addr[48455]= 1782906961;
assign addr[48456]= 1761306505;
assign addr[48457]= 1739147417;
assign addr[48458]= 1716436725;
assign addr[48459]= 1693181631;
assign addr[48460]= 1669389513;
assign addr[48461]= 1645067915;
assign addr[48462]= 1620224553;
assign addr[48463]= 1594867305;
assign addr[48464]= 1569004214;
assign addr[48465]= 1542643483;
assign addr[48466]= 1515793473;
assign addr[48467]= 1488462700;
assign addr[48468]= 1460659832;
assign addr[48469]= 1432393688;
assign addr[48470]= 1403673233;
assign addr[48471]= 1374507575;
assign addr[48472]= 1344905966;
assign addr[48473]= 1314877795;
assign addr[48474]= 1284432584;
assign addr[48475]= 1253579991;
assign addr[48476]= 1222329801;
assign addr[48477]= 1190691925;
assign addr[48478]= 1158676398;
assign addr[48479]= 1126293375;
assign addr[48480]= 1093553126;
assign addr[48481]= 1060466036;
assign addr[48482]= 1027042599;
assign addr[48483]= 993293415;
assign addr[48484]= 959229189;
assign addr[48485]= 924860725;
assign addr[48486]= 890198924;
assign addr[48487]= 855254778;
assign addr[48488]= 820039373;
assign addr[48489]= 784563876;
assign addr[48490]= 748839539;
assign addr[48491]= 712877694;
assign addr[48492]= 676689746;
assign addr[48493]= 640287172;
assign addr[48494]= 603681519;
assign addr[48495]= 566884397;
assign addr[48496]= 529907477;
assign addr[48497]= 492762486;
assign addr[48498]= 455461206;
assign addr[48499]= 418015468;
assign addr[48500]= 380437148;
assign addr[48501]= 342738165;
assign addr[48502]= 304930476;
assign addr[48503]= 267026072;
assign addr[48504]= 229036977;
assign addr[48505]= 190975237;
assign addr[48506]= 152852926;
assign addr[48507]= 114682135;
assign addr[48508]= 76474970;
assign addr[48509]= 38243550;
assign addr[48510]= 0;
assign addr[48511]= -38243550;
assign addr[48512]= -76474970;
assign addr[48513]= -114682135;
assign addr[48514]= -152852926;
assign addr[48515]= -190975237;
assign addr[48516]= -229036977;
assign addr[48517]= -267026072;
assign addr[48518]= -304930476;
assign addr[48519]= -342738165;
assign addr[48520]= -380437148;
assign addr[48521]= -418015468;
assign addr[48522]= -455461206;
assign addr[48523]= -492762486;
assign addr[48524]= -529907477;
assign addr[48525]= -566884397;
assign addr[48526]= -603681519;
assign addr[48527]= -640287172;
assign addr[48528]= -676689746;
assign addr[48529]= -712877694;
assign addr[48530]= -748839539;
assign addr[48531]= -784563876;
assign addr[48532]= -820039373;
assign addr[48533]= -855254778;
assign addr[48534]= -890198924;
assign addr[48535]= -924860725;
assign addr[48536]= -959229189;
assign addr[48537]= -993293415;
assign addr[48538]= -1027042599;
assign addr[48539]= -1060466036;
assign addr[48540]= -1093553126;
assign addr[48541]= -1126293375;
assign addr[48542]= -1158676398;
assign addr[48543]= -1190691925;
assign addr[48544]= -1222329801;
assign addr[48545]= -1253579991;
assign addr[48546]= -1284432584;
assign addr[48547]= -1314877795;
assign addr[48548]= -1344905966;
assign addr[48549]= -1374507575;
assign addr[48550]= -1403673233;
assign addr[48551]= -1432393688;
assign addr[48552]= -1460659832;
assign addr[48553]= -1488462700;
assign addr[48554]= -1515793473;
assign addr[48555]= -1542643483;
assign addr[48556]= -1569004214;
assign addr[48557]= -1594867305;
assign addr[48558]= -1620224553;
assign addr[48559]= -1645067915;
assign addr[48560]= -1669389513;
assign addr[48561]= -1693181631;
assign addr[48562]= -1716436725;
assign addr[48563]= -1739147417;
assign addr[48564]= -1761306505;
assign addr[48565]= -1782906961;
assign addr[48566]= -1803941934;
assign addr[48567]= -1824404752;
assign addr[48568]= -1844288924;
assign addr[48569]= -1863588145;
assign addr[48570]= -1882296293;
assign addr[48571]= -1900407434;
assign addr[48572]= -1917915825;
assign addr[48573]= -1934815911;
assign addr[48574]= -1951102334;
assign addr[48575]= -1966769926;
assign addr[48576]= -1981813720;
assign addr[48577]= -1996228943;
assign addr[48578]= -2010011024;
assign addr[48579]= -2023155591;
assign addr[48580]= -2035658475;
assign addr[48581]= -2047515711;
assign addr[48582]= -2058723538;
assign addr[48583]= -2069278401;
assign addr[48584]= -2079176953;
assign addr[48585]= -2088416053;
assign addr[48586]= -2096992772;
assign addr[48587]= -2104904390;
assign addr[48588]= -2112148396;
assign addr[48589]= -2118722494;
assign addr[48590]= -2124624598;
assign addr[48591]= -2129852837;
assign addr[48592]= -2134405552;
assign addr[48593]= -2138281298;
assign addr[48594]= -2141478848;
assign addr[48595]= -2143997187;
assign addr[48596]= -2145835515;
assign addr[48597]= -2146993250;
assign addr[48598]= -2147470025;
assign addr[48599]= -2147265689;
assign addr[48600]= -2146380306;
assign addr[48601]= -2144814157;
assign addr[48602]= -2142567738;
assign addr[48603]= -2139641764;
assign addr[48604]= -2136037160;
assign addr[48605]= -2131755071;
assign addr[48606]= -2126796855;
assign addr[48607]= -2121164085;
assign addr[48608]= -2114858546;
assign addr[48609]= -2107882239;
assign addr[48610]= -2100237377;
assign addr[48611]= -2091926384;
assign addr[48612]= -2082951896;
assign addr[48613]= -2073316760;
assign addr[48614]= -2063024031;
assign addr[48615]= -2052076975;
assign addr[48616]= -2040479063;
assign addr[48617]= -2028233973;
assign addr[48618]= -2015345591;
assign addr[48619]= -2001818002;
assign addr[48620]= -1987655498;
assign addr[48621]= -1972862571;
assign addr[48622]= -1957443913;
assign addr[48623]= -1941404413;
assign addr[48624]= -1924749160;
assign addr[48625]= -1907483436;
assign addr[48626]= -1889612716;
assign addr[48627]= -1871142669;
assign addr[48628]= -1852079154;
assign addr[48629]= -1832428215;
assign addr[48630]= -1812196087;
assign addr[48631]= -1791389186;
assign addr[48632]= -1770014111;
assign addr[48633]= -1748077642;
assign addr[48634]= -1725586737;
assign addr[48635]= -1702548529;
assign addr[48636]= -1678970324;
assign addr[48637]= -1654859602;
assign addr[48638]= -1630224009;
assign addr[48639]= -1605071359;
assign addr[48640]= -1579409630;
assign addr[48641]= -1553246960;
assign addr[48642]= -1526591649;
assign addr[48643]= -1499452149;
assign addr[48644]= -1471837070;
assign addr[48645]= -1443755168;
assign addr[48646]= -1415215352;
assign addr[48647]= -1386226674;
assign addr[48648]= -1356798326;
assign addr[48649]= -1326939644;
assign addr[48650]= -1296660098;
assign addr[48651]= -1265969291;
assign addr[48652]= -1234876957;
assign addr[48653]= -1203392958;
assign addr[48654]= -1171527280;
assign addr[48655]= -1139290029;
assign addr[48656]= -1106691431;
assign addr[48657]= -1073741824;
assign addr[48658]= -1040451659;
assign addr[48659]= -1006831495;
assign addr[48660]= -972891995;
assign addr[48661]= -938643924;
assign addr[48662]= -904098143;
assign addr[48663]= -869265610;
assign addr[48664]= -834157373;
assign addr[48665]= -798784567;
assign addr[48666]= -763158411;
assign addr[48667]= -727290205;
assign addr[48668]= -691191324;
assign addr[48669]= -654873219;
assign addr[48670]= -618347408;
assign addr[48671]= -581625477;
assign addr[48672]= -544719071;
assign addr[48673]= -507639898;
assign addr[48674]= -470399716;
assign addr[48675]= -433010339;
assign addr[48676]= -395483624;
assign addr[48677]= -357831473;
assign addr[48678]= -320065829;
assign addr[48679]= -282198671;
assign addr[48680]= -244242007;
assign addr[48681]= -206207878;
assign addr[48682]= -168108346;
assign addr[48683]= -129955495;
assign addr[48684]= -91761426;
assign addr[48685]= -53538253;
assign addr[48686]= -15298099;
assign addr[48687]= 22946906;
assign addr[48688]= 61184634;
assign addr[48689]= 99402956;
assign addr[48690]= 137589750;
assign addr[48691]= 175732905;
assign addr[48692]= 213820322;
assign addr[48693]= 251839923;
assign addr[48694]= 289779648;
assign addr[48695]= 327627463;
assign addr[48696]= 365371365;
assign addr[48697]= 402999383;
assign addr[48698]= 440499581;
assign addr[48699]= 477860067;
assign addr[48700]= 515068990;
assign addr[48701]= 552114549;
assign addr[48702]= 588984994;
assign addr[48703]= 625668632;
assign addr[48704]= 662153826;
assign addr[48705]= 698429006;
assign addr[48706]= 734482665;
assign addr[48707]= 770303369;
assign addr[48708]= 805879757;
assign addr[48709]= 841200544;
assign addr[48710]= 876254528;
assign addr[48711]= 911030591;
assign addr[48712]= 945517704;
assign addr[48713]= 979704927;
assign addr[48714]= 1013581418;
assign addr[48715]= 1047136432;
assign addr[48716]= 1080359326;
assign addr[48717]= 1113239564;
assign addr[48718]= 1145766716;
assign addr[48719]= 1177930466;
assign addr[48720]= 1209720613;
assign addr[48721]= 1241127074;
assign addr[48722]= 1272139887;
assign addr[48723]= 1302749217;
assign addr[48724]= 1332945355;
assign addr[48725]= 1362718723;
assign addr[48726]= 1392059879;
assign addr[48727]= 1420959516;
assign addr[48728]= 1449408469;
assign addr[48729]= 1477397714;
assign addr[48730]= 1504918373;
assign addr[48731]= 1531961719;
assign addr[48732]= 1558519173;
assign addr[48733]= 1584582314;
assign addr[48734]= 1610142873;
assign addr[48735]= 1635192744;
assign addr[48736]= 1659723983;
assign addr[48737]= 1683728808;
assign addr[48738]= 1707199606;
assign addr[48739]= 1730128933;
assign addr[48740]= 1752509516;
assign addr[48741]= 1774334257;
assign addr[48742]= 1795596234;
assign addr[48743]= 1816288703;
assign addr[48744]= 1836405100;
assign addr[48745]= 1855939047;
assign addr[48746]= 1874884346;
assign addr[48747]= 1893234990;
assign addr[48748]= 1910985158;
assign addr[48749]= 1928129220;
assign addr[48750]= 1944661739;
assign addr[48751]= 1960577471;
assign addr[48752]= 1975871368;
assign addr[48753]= 1990538579;
assign addr[48754]= 2004574453;
assign addr[48755]= 2017974537;
assign addr[48756]= 2030734582;
assign addr[48757]= 2042850540;
assign addr[48758]= 2054318569;
assign addr[48759]= 2065135031;
assign addr[48760]= 2075296495;
assign addr[48761]= 2084799740;
assign addr[48762]= 2093641749;
assign addr[48763]= 2101819720;
assign addr[48764]= 2109331059;
assign addr[48765]= 2116173382;
assign addr[48766]= 2122344521;
assign addr[48767]= 2127842516;
assign addr[48768]= 2132665626;
assign addr[48769]= 2136812319;
assign addr[48770]= 2140281282;
assign addr[48771]= 2143071413;
assign addr[48772]= 2145181827;
assign addr[48773]= 2146611856;
assign addr[48774]= 2147361045;
assign addr[48775]= 2147429158;
assign addr[48776]= 2146816171;
assign addr[48777]= 2145522281;
assign addr[48778]= 2143547897;
assign addr[48779]= 2140893646;
assign addr[48780]= 2137560369;
assign addr[48781]= 2133549123;
assign addr[48782]= 2128861181;
assign addr[48783]= 2123498030;
assign addr[48784]= 2117461370;
assign addr[48785]= 2110753117;
assign addr[48786]= 2103375398;
assign addr[48787]= 2095330553;
assign addr[48788]= 2086621133;
assign addr[48789]= 2077249901;
assign addr[48790]= 2067219829;
assign addr[48791]= 2056534099;
assign addr[48792]= 2045196100;
assign addr[48793]= 2033209426;
assign addr[48794]= 2020577882;
assign addr[48795]= 2007305472;
assign addr[48796]= 1993396407;
assign addr[48797]= 1978855097;
assign addr[48798]= 1963686155;
assign addr[48799]= 1947894393;
assign addr[48800]= 1931484818;
assign addr[48801]= 1914462636;
assign addr[48802]= 1896833245;
assign addr[48803]= 1878602237;
assign addr[48804]= 1859775393;
assign addr[48805]= 1840358687;
assign addr[48806]= 1820358275;
assign addr[48807]= 1799780501;
assign addr[48808]= 1778631892;
assign addr[48809]= 1756919156;
assign addr[48810]= 1734649179;
assign addr[48811]= 1711829025;
assign addr[48812]= 1688465931;
assign addr[48813]= 1664567307;
assign addr[48814]= 1640140734;
assign addr[48815]= 1615193959;
assign addr[48816]= 1589734894;
assign addr[48817]= 1563771613;
assign addr[48818]= 1537312353;
assign addr[48819]= 1510365504;
assign addr[48820]= 1482939614;
assign addr[48821]= 1455043381;
assign addr[48822]= 1426685652;
assign addr[48823]= 1397875423;
assign addr[48824]= 1368621831;
assign addr[48825]= 1338934154;
assign addr[48826]= 1308821808;
assign addr[48827]= 1278294345;
assign addr[48828]= 1247361445;
assign addr[48829]= 1216032921;
assign addr[48830]= 1184318708;
assign addr[48831]= 1152228866;
assign addr[48832]= 1119773573;
assign addr[48833]= 1086963121;
assign addr[48834]= 1053807919;
assign addr[48835]= 1020318481;
assign addr[48836]= 986505429;
assign addr[48837]= 952379488;
assign addr[48838]= 917951481;
assign addr[48839]= 883232329;
assign addr[48840]= 848233042;
assign addr[48841]= 812964722;
assign addr[48842]= 777438554;
assign addr[48843]= 741665807;
assign addr[48844]= 705657826;
assign addr[48845]= 669426032;
assign addr[48846]= 632981917;
assign addr[48847]= 596337040;
assign addr[48848]= 559503022;
assign addr[48849]= 522491548;
assign addr[48850]= 485314355;
assign addr[48851]= 447983235;
assign addr[48852]= 410510029;
assign addr[48853]= 372906622;
assign addr[48854]= 335184940;
assign addr[48855]= 297356948;
assign addr[48856]= 259434643;
assign addr[48857]= 221430054;
assign addr[48858]= 183355234;
assign addr[48859]= 145222259;
assign addr[48860]= 107043224;
assign addr[48861]= 68830239;
assign addr[48862]= 30595422;
assign addr[48863]= -7649098;
assign addr[48864]= -45891193;
assign addr[48865]= -84118732;
assign addr[48866]= -122319591;
assign addr[48867]= -160481654;
assign addr[48868]= -198592817;
assign addr[48869]= -236640993;
assign addr[48870]= -274614114;
assign addr[48871]= -312500135;
assign addr[48872]= -350287041;
assign addr[48873]= -387962847;
assign addr[48874]= -425515602;
assign addr[48875]= -462933398;
assign addr[48876]= -500204365;
assign addr[48877]= -537316682;
assign addr[48878]= -574258580;
assign addr[48879]= -611018340;
assign addr[48880]= -647584304;
assign addr[48881]= -683944874;
assign addr[48882]= -720088517;
assign addr[48883]= -756003771;
assign addr[48884]= -791679244;
assign addr[48885]= -827103620;
assign addr[48886]= -862265664;
assign addr[48887]= -897154224;
assign addr[48888]= -931758235;
assign addr[48889]= -966066720;
assign addr[48890]= -1000068799;
assign addr[48891]= -1033753687;
assign addr[48892]= -1067110699;
assign addr[48893]= -1100129257;
assign addr[48894]= -1132798888;
assign addr[48895]= -1165109230;
assign addr[48896]= -1197050035;
assign addr[48897]= -1228611172;
assign addr[48898]= -1259782632;
assign addr[48899]= -1290554528;
assign addr[48900]= -1320917099;
assign addr[48901]= -1350860716;
assign addr[48902]= -1380375881;
assign addr[48903]= -1409453233;
assign addr[48904]= -1438083551;
assign addr[48905]= -1466257752;
assign addr[48906]= -1493966902;
assign addr[48907]= -1521202211;
assign addr[48908]= -1547955041;
assign addr[48909]= -1574216908;
assign addr[48910]= -1599979481;
assign addr[48911]= -1625234591;
assign addr[48912]= -1649974225;
assign addr[48913]= -1674190539;
assign addr[48914]= -1697875851;
assign addr[48915]= -1721022648;
assign addr[48916]= -1743623590;
assign addr[48917]= -1765671509;
assign addr[48918]= -1787159411;
assign addr[48919]= -1808080480;
assign addr[48920]= -1828428082;
assign addr[48921]= -1848195763;
assign addr[48922]= -1867377253;
assign addr[48923]= -1885966468;
assign addr[48924]= -1903957513;
assign addr[48925]= -1921344681;
assign addr[48926]= -1938122457;
assign addr[48927]= -1954285520;
assign addr[48928]= -1969828744;
assign addr[48929]= -1984747199;
assign addr[48930]= -1999036154;
assign addr[48931]= -2012691075;
assign addr[48932]= -2025707632;
assign addr[48933]= -2038081698;
assign addr[48934]= -2049809346;
assign addr[48935]= -2060886858;
assign addr[48936]= -2071310720;
assign addr[48937]= -2081077626;
assign addr[48938]= -2090184478;
assign addr[48939]= -2098628387;
assign addr[48940]= -2106406677;
assign addr[48941]= -2113516878;
assign addr[48942]= -2119956737;
assign addr[48943]= -2125724211;
assign addr[48944]= -2130817471;
assign addr[48945]= -2135234901;
assign addr[48946]= -2138975100;
assign addr[48947]= -2142036881;
assign addr[48948]= -2144419275;
assign addr[48949]= -2146121524;
assign addr[48950]= -2147143090;
assign addr[48951]= -2147483648;
assign addr[48952]= -2147143090;
assign addr[48953]= -2146121524;
assign addr[48954]= -2144419275;
assign addr[48955]= -2142036881;
assign addr[48956]= -2138975100;
assign addr[48957]= -2135234901;
assign addr[48958]= -2130817471;
assign addr[48959]= -2125724211;
assign addr[48960]= -2119956737;
assign addr[48961]= -2113516878;
assign addr[48962]= -2106406677;
assign addr[48963]= -2098628387;
assign addr[48964]= -2090184478;
assign addr[48965]= -2081077626;
assign addr[48966]= -2071310720;
assign addr[48967]= -2060886858;
assign addr[48968]= -2049809346;
assign addr[48969]= -2038081698;
assign addr[48970]= -2025707632;
assign addr[48971]= -2012691075;
assign addr[48972]= -1999036154;
assign addr[48973]= -1984747199;
assign addr[48974]= -1969828744;
assign addr[48975]= -1954285520;
assign addr[48976]= -1938122457;
assign addr[48977]= -1921344681;
assign addr[48978]= -1903957513;
assign addr[48979]= -1885966468;
assign addr[48980]= -1867377253;
assign addr[48981]= -1848195763;
assign addr[48982]= -1828428082;
assign addr[48983]= -1808080480;
assign addr[48984]= -1787159411;
assign addr[48985]= -1765671509;
assign addr[48986]= -1743623590;
assign addr[48987]= -1721022648;
assign addr[48988]= -1697875851;
assign addr[48989]= -1674190539;
assign addr[48990]= -1649974225;
assign addr[48991]= -1625234591;
assign addr[48992]= -1599979481;
assign addr[48993]= -1574216908;
assign addr[48994]= -1547955041;
assign addr[48995]= -1521202211;
assign addr[48996]= -1493966902;
assign addr[48997]= -1466257752;
assign addr[48998]= -1438083551;
assign addr[48999]= -1409453233;
assign addr[49000]= -1380375881;
assign addr[49001]= -1350860716;
assign addr[49002]= -1320917099;
assign addr[49003]= -1290554528;
assign addr[49004]= -1259782632;
assign addr[49005]= -1228611172;
assign addr[49006]= -1197050035;
assign addr[49007]= -1165109230;
assign addr[49008]= -1132798888;
assign addr[49009]= -1100129257;
assign addr[49010]= -1067110699;
assign addr[49011]= -1033753687;
assign addr[49012]= -1000068799;
assign addr[49013]= -966066720;
assign addr[49014]= -931758235;
assign addr[49015]= -897154224;
assign addr[49016]= -862265664;
assign addr[49017]= -827103620;
assign addr[49018]= -791679244;
assign addr[49019]= -756003771;
assign addr[49020]= -720088517;
assign addr[49021]= -683944874;
assign addr[49022]= -647584304;
assign addr[49023]= -611018340;
assign addr[49024]= -574258580;
assign addr[49025]= -537316682;
assign addr[49026]= -500204365;
assign addr[49027]= -462933398;
assign addr[49028]= -425515602;
assign addr[49029]= -387962847;
assign addr[49030]= -350287041;
assign addr[49031]= -312500135;
assign addr[49032]= -274614114;
assign addr[49033]= -236640993;
assign addr[49034]= -198592817;
assign addr[49035]= -160481654;
assign addr[49036]= -122319591;
assign addr[49037]= -84118732;
assign addr[49038]= -45891193;
assign addr[49039]= -7649098;
assign addr[49040]= 30595422;
assign addr[49041]= 68830239;
assign addr[49042]= 107043224;
assign addr[49043]= 145222259;
assign addr[49044]= 183355234;
assign addr[49045]= 221430054;
assign addr[49046]= 259434643;
assign addr[49047]= 297356948;
assign addr[49048]= 335184940;
assign addr[49049]= 372906622;
assign addr[49050]= 410510029;
assign addr[49051]= 447983235;
assign addr[49052]= 485314355;
assign addr[49053]= 522491548;
assign addr[49054]= 559503022;
assign addr[49055]= 596337040;
assign addr[49056]= 632981917;
assign addr[49057]= 669426032;
assign addr[49058]= 705657826;
assign addr[49059]= 741665807;
assign addr[49060]= 777438554;
assign addr[49061]= 812964722;
assign addr[49062]= 848233042;
assign addr[49063]= 883232329;
assign addr[49064]= 917951481;
assign addr[49065]= 952379488;
assign addr[49066]= 986505429;
assign addr[49067]= 1020318481;
assign addr[49068]= 1053807919;
assign addr[49069]= 1086963121;
assign addr[49070]= 1119773573;
assign addr[49071]= 1152228866;
assign addr[49072]= 1184318708;
assign addr[49073]= 1216032921;
assign addr[49074]= 1247361445;
assign addr[49075]= 1278294345;
assign addr[49076]= 1308821808;
assign addr[49077]= 1338934154;
assign addr[49078]= 1368621831;
assign addr[49079]= 1397875423;
assign addr[49080]= 1426685652;
assign addr[49081]= 1455043381;
assign addr[49082]= 1482939614;
assign addr[49083]= 1510365504;
assign addr[49084]= 1537312353;
assign addr[49085]= 1563771613;
assign addr[49086]= 1589734894;
assign addr[49087]= 1615193959;
assign addr[49088]= 1640140734;
assign addr[49089]= 1664567307;
assign addr[49090]= 1688465931;
assign addr[49091]= 1711829025;
assign addr[49092]= 1734649179;
assign addr[49093]= 1756919156;
assign addr[49094]= 1778631892;
assign addr[49095]= 1799780501;
assign addr[49096]= 1820358275;
assign addr[49097]= 1840358687;
assign addr[49098]= 1859775393;
assign addr[49099]= 1878602237;
assign addr[49100]= 1896833245;
assign addr[49101]= 1914462636;
assign addr[49102]= 1931484818;
assign addr[49103]= 1947894393;
assign addr[49104]= 1963686155;
assign addr[49105]= 1978855097;
assign addr[49106]= 1993396407;
assign addr[49107]= 2007305472;
assign addr[49108]= 2020577882;
assign addr[49109]= 2033209426;
assign addr[49110]= 2045196100;
assign addr[49111]= 2056534099;
assign addr[49112]= 2067219829;
assign addr[49113]= 2077249901;
assign addr[49114]= 2086621133;
assign addr[49115]= 2095330553;
assign addr[49116]= 2103375398;
assign addr[49117]= 2110753117;
assign addr[49118]= 2117461370;
assign addr[49119]= 2123498030;
assign addr[49120]= 2128861181;
assign addr[49121]= 2133549123;
assign addr[49122]= 2137560369;
assign addr[49123]= 2140893646;
assign addr[49124]= 2143547897;
assign addr[49125]= 2145522281;
assign addr[49126]= 2146816171;
assign addr[49127]= 2147429158;
assign addr[49128]= 2147361045;
assign addr[49129]= 2146611856;
assign addr[49130]= 2145181827;
assign addr[49131]= 2143071413;
assign addr[49132]= 2140281282;
assign addr[49133]= 2136812319;
assign addr[49134]= 2132665626;
assign addr[49135]= 2127842516;
assign addr[49136]= 2122344521;
assign addr[49137]= 2116173382;
assign addr[49138]= 2109331059;
assign addr[49139]= 2101819720;
assign addr[49140]= 2093641749;
assign addr[49141]= 2084799740;
assign addr[49142]= 2075296495;
assign addr[49143]= 2065135031;
assign addr[49144]= 2054318569;
assign addr[49145]= 2042850540;
assign addr[49146]= 2030734582;
assign addr[49147]= 2017974537;
assign addr[49148]= 2004574453;
assign addr[49149]= 1990538579;
assign addr[49150]= 1975871368;
assign addr[49151]= 1960577471;
assign addr[49152]= 1944661739;
assign addr[49153]= 1928129220;
assign addr[49154]= 1910985158;
assign addr[49155]= 1893234990;
assign addr[49156]= 1874884346;
assign addr[49157]= 1855939047;
assign addr[49158]= 1836405100;
assign addr[49159]= 1816288703;
assign addr[49160]= 1795596234;
assign addr[49161]= 1774334257;
assign addr[49162]= 1752509516;
assign addr[49163]= 1730128933;
assign addr[49164]= 1707199606;
assign addr[49165]= 1683728808;
assign addr[49166]= 1659723983;
assign addr[49167]= 1635192744;
assign addr[49168]= 1610142873;
assign addr[49169]= 1584582314;
assign addr[49170]= 1558519173;
assign addr[49171]= 1531961719;
assign addr[49172]= 1504918373;
assign addr[49173]= 1477397714;
assign addr[49174]= 1449408469;
assign addr[49175]= 1420959516;
assign addr[49176]= 1392059879;
assign addr[49177]= 1362718723;
assign addr[49178]= 1332945355;
assign addr[49179]= 1302749217;
assign addr[49180]= 1272139887;
assign addr[49181]= 1241127074;
assign addr[49182]= 1209720613;
assign addr[49183]= 1177930466;
assign addr[49184]= 1145766716;
assign addr[49185]= 1113239564;
assign addr[49186]= 1080359326;
assign addr[49187]= 1047136432;
assign addr[49188]= 1013581418;
assign addr[49189]= 979704927;
assign addr[49190]= 945517704;
assign addr[49191]= 911030591;
assign addr[49192]= 876254528;
assign addr[49193]= 841200544;
assign addr[49194]= 805879757;
assign addr[49195]= 770303369;
assign addr[49196]= 734482665;
assign addr[49197]= 698429006;
assign addr[49198]= 662153826;
assign addr[49199]= 625668632;
assign addr[49200]= 588984994;
assign addr[49201]= 552114549;
assign addr[49202]= 515068990;
assign addr[49203]= 477860067;
assign addr[49204]= 440499581;
assign addr[49205]= 402999383;
assign addr[49206]= 365371365;
assign addr[49207]= 327627463;
assign addr[49208]= 289779648;
assign addr[49209]= 251839923;
assign addr[49210]= 213820322;
assign addr[49211]= 175732905;
assign addr[49212]= 137589750;
assign addr[49213]= 99402956;
assign addr[49214]= 61184634;
assign addr[49215]= 22946906;
assign addr[49216]= -15298099;
assign addr[49217]= -53538253;
assign addr[49218]= -91761426;
assign addr[49219]= -129955495;
assign addr[49220]= -168108346;
assign addr[49221]= -206207878;
assign addr[49222]= -244242007;
assign addr[49223]= -282198671;
assign addr[49224]= -320065829;
assign addr[49225]= -357831473;
assign addr[49226]= -395483624;
assign addr[49227]= -433010339;
assign addr[49228]= -470399716;
assign addr[49229]= -507639898;
assign addr[49230]= -544719071;
assign addr[49231]= -581625477;
assign addr[49232]= -618347408;
assign addr[49233]= -654873219;
assign addr[49234]= -691191324;
assign addr[49235]= -727290205;
assign addr[49236]= -763158411;
assign addr[49237]= -798784567;
assign addr[49238]= -834157373;
assign addr[49239]= -869265610;
assign addr[49240]= -904098143;
assign addr[49241]= -938643924;
assign addr[49242]= -972891995;
assign addr[49243]= -1006831495;
assign addr[49244]= -1040451659;
assign addr[49245]= -1073741824;
assign addr[49246]= -1106691431;
assign addr[49247]= -1139290029;
assign addr[49248]= -1171527280;
assign addr[49249]= -1203392958;
assign addr[49250]= -1234876957;
assign addr[49251]= -1265969291;
assign addr[49252]= -1296660098;
assign addr[49253]= -1326939644;
assign addr[49254]= -1356798326;
assign addr[49255]= -1386226674;
assign addr[49256]= -1415215352;
assign addr[49257]= -1443755168;
assign addr[49258]= -1471837070;
assign addr[49259]= -1499452149;
assign addr[49260]= -1526591649;
assign addr[49261]= -1553246960;
assign addr[49262]= -1579409630;
assign addr[49263]= -1605071359;
assign addr[49264]= -1630224009;
assign addr[49265]= -1654859602;
assign addr[49266]= -1678970324;
assign addr[49267]= -1702548529;
assign addr[49268]= -1725586737;
assign addr[49269]= -1748077642;
assign addr[49270]= -1770014111;
assign addr[49271]= -1791389186;
assign addr[49272]= -1812196087;
assign addr[49273]= -1832428215;
assign addr[49274]= -1852079154;
assign addr[49275]= -1871142669;
assign addr[49276]= -1889612716;
assign addr[49277]= -1907483436;
assign addr[49278]= -1924749160;
assign addr[49279]= -1941404413;
assign addr[49280]= -1957443913;
assign addr[49281]= -1972862571;
assign addr[49282]= -1987655498;
assign addr[49283]= -2001818002;
assign addr[49284]= -2015345591;
assign addr[49285]= -2028233973;
assign addr[49286]= -2040479063;
assign addr[49287]= -2052076975;
assign addr[49288]= -2063024031;
assign addr[49289]= -2073316760;
assign addr[49290]= -2082951896;
assign addr[49291]= -2091926384;
assign addr[49292]= -2100237377;
assign addr[49293]= -2107882239;
assign addr[49294]= -2114858546;
assign addr[49295]= -2121164085;
assign addr[49296]= -2126796855;
assign addr[49297]= -2131755071;
assign addr[49298]= -2136037160;
assign addr[49299]= -2139641764;
assign addr[49300]= -2142567738;
assign addr[49301]= -2144814157;
assign addr[49302]= -2146380306;
assign addr[49303]= -2147265689;
assign addr[49304]= -2147470025;
assign addr[49305]= -2146993250;
assign addr[49306]= -2145835515;
assign addr[49307]= -2143997187;
assign addr[49308]= -2141478848;
assign addr[49309]= -2138281298;
assign addr[49310]= -2134405552;
assign addr[49311]= -2129852837;
assign addr[49312]= -2124624598;
assign addr[49313]= -2118722494;
assign addr[49314]= -2112148396;
assign addr[49315]= -2104904390;
assign addr[49316]= -2096992772;
assign addr[49317]= -2088416053;
assign addr[49318]= -2079176953;
assign addr[49319]= -2069278401;
assign addr[49320]= -2058723538;
assign addr[49321]= -2047515711;
assign addr[49322]= -2035658475;
assign addr[49323]= -2023155591;
assign addr[49324]= -2010011024;
assign addr[49325]= -1996228943;
assign addr[49326]= -1981813720;
assign addr[49327]= -1966769926;
assign addr[49328]= -1951102334;
assign addr[49329]= -1934815911;
assign addr[49330]= -1917915825;
assign addr[49331]= -1900407434;
assign addr[49332]= -1882296293;
assign addr[49333]= -1863588145;
assign addr[49334]= -1844288924;
assign addr[49335]= -1824404752;
assign addr[49336]= -1803941934;
assign addr[49337]= -1782906961;
assign addr[49338]= -1761306505;
assign addr[49339]= -1739147417;
assign addr[49340]= -1716436725;
assign addr[49341]= -1693181631;
assign addr[49342]= -1669389513;
assign addr[49343]= -1645067915;
assign addr[49344]= -1620224553;
assign addr[49345]= -1594867305;
assign addr[49346]= -1569004214;
assign addr[49347]= -1542643483;
assign addr[49348]= -1515793473;
assign addr[49349]= -1488462700;
assign addr[49350]= -1460659832;
assign addr[49351]= -1432393688;
assign addr[49352]= -1403673233;
assign addr[49353]= -1374507575;
assign addr[49354]= -1344905966;
assign addr[49355]= -1314877795;
assign addr[49356]= -1284432584;
assign addr[49357]= -1253579991;
assign addr[49358]= -1222329801;
assign addr[49359]= -1190691925;
assign addr[49360]= -1158676398;
assign addr[49361]= -1126293375;
assign addr[49362]= -1093553126;
assign addr[49363]= -1060466036;
assign addr[49364]= -1027042599;
assign addr[49365]= -993293415;
assign addr[49366]= -959229189;
assign addr[49367]= -924860725;
assign addr[49368]= -890198924;
assign addr[49369]= -855254778;
assign addr[49370]= -820039373;
assign addr[49371]= -784563876;
assign addr[49372]= -748839539;
assign addr[49373]= -712877694;
assign addr[49374]= -676689746;
assign addr[49375]= -640287172;
assign addr[49376]= -603681519;
assign addr[49377]= -566884397;
assign addr[49378]= -529907477;
assign addr[49379]= -492762486;
assign addr[49380]= -455461206;
assign addr[49381]= -418015468;
assign addr[49382]= -380437148;
assign addr[49383]= -342738165;
assign addr[49384]= -304930476;
assign addr[49385]= -267026072;
assign addr[49386]= -229036977;
assign addr[49387]= -190975237;
assign addr[49388]= -152852926;
assign addr[49389]= -114682135;
assign addr[49390]= -76474970;
assign addr[49391]= -38243550;
assign addr[49392]= 0;
assign addr[49393]= 38243550;
assign addr[49394]= 76474970;
assign addr[49395]= 114682135;
assign addr[49396]= 152852926;
assign addr[49397]= 190975237;
assign addr[49398]= 229036977;
assign addr[49399]= 267026072;
assign addr[49400]= 304930476;
assign addr[49401]= 342738165;
assign addr[49402]= 380437148;
assign addr[49403]= 418015468;
assign addr[49404]= 455461206;
assign addr[49405]= 492762486;
assign addr[49406]= 529907477;
assign addr[49407]= 566884397;
assign addr[49408]= 603681519;
assign addr[49409]= 640287172;
assign addr[49410]= 676689746;
assign addr[49411]= 712877694;
assign addr[49412]= 748839539;
assign addr[49413]= 784563876;
assign addr[49414]= 820039373;
assign addr[49415]= 855254778;
assign addr[49416]= 890198924;
assign addr[49417]= 924860725;
assign addr[49418]= 959229189;
assign addr[49419]= 993293415;
assign addr[49420]= 1027042599;
assign addr[49421]= 1060466036;
assign addr[49422]= 1093553126;
assign addr[49423]= 1126293375;
assign addr[49424]= 1158676398;
assign addr[49425]= 1190691925;
assign addr[49426]= 1222329801;
assign addr[49427]= 1253579991;
assign addr[49428]= 1284432584;
assign addr[49429]= 1314877795;
assign addr[49430]= 1344905966;
assign addr[49431]= 1374507575;
assign addr[49432]= 1403673233;
assign addr[49433]= 1432393688;
assign addr[49434]= 1460659832;
assign addr[49435]= 1488462700;
assign addr[49436]= 1515793473;
assign addr[49437]= 1542643483;
assign addr[49438]= 1569004214;
assign addr[49439]= 1594867305;
assign addr[49440]= 1620224553;
assign addr[49441]= 1645067915;
assign addr[49442]= 1669389513;
assign addr[49443]= 1693181631;
assign addr[49444]= 1716436725;
assign addr[49445]= 1739147417;
assign addr[49446]= 1761306505;
assign addr[49447]= 1782906961;
assign addr[49448]= 1803941934;
assign addr[49449]= 1824404752;
assign addr[49450]= 1844288924;
assign addr[49451]= 1863588145;
assign addr[49452]= 1882296293;
assign addr[49453]= 1900407434;
assign addr[49454]= 1917915825;
assign addr[49455]= 1934815911;
assign addr[49456]= 1951102334;
assign addr[49457]= 1966769926;
assign addr[49458]= 1981813720;
assign addr[49459]= 1996228943;
assign addr[49460]= 2010011024;
assign addr[49461]= 2023155591;
assign addr[49462]= 2035658475;
assign addr[49463]= 2047515711;
assign addr[49464]= 2058723538;
assign addr[49465]= 2069278401;
assign addr[49466]= 2079176953;
assign addr[49467]= 2088416053;
assign addr[49468]= 2096992772;
assign addr[49469]= 2104904390;
assign addr[49470]= 2112148396;
assign addr[49471]= 2118722494;
assign addr[49472]= 2124624598;
assign addr[49473]= 2129852837;
assign addr[49474]= 2134405552;
assign addr[49475]= 2138281298;
assign addr[49476]= 2141478848;
assign addr[49477]= 2143997187;
assign addr[49478]= 2145835515;
assign addr[49479]= 2146993250;
assign addr[49480]= 2147470025;
assign addr[49481]= 2147265689;
assign addr[49482]= 2146380306;
assign addr[49483]= 2144814157;
assign addr[49484]= 2142567738;
assign addr[49485]= 2139641764;
assign addr[49486]= 2136037160;
assign addr[49487]= 2131755071;
assign addr[49488]= 2126796855;
assign addr[49489]= 2121164085;
assign addr[49490]= 2114858546;
assign addr[49491]= 2107882239;
assign addr[49492]= 2100237377;
assign addr[49493]= 2091926384;
assign addr[49494]= 2082951896;
assign addr[49495]= 2073316760;
assign addr[49496]= 2063024031;
assign addr[49497]= 2052076975;
assign addr[49498]= 2040479063;
assign addr[49499]= 2028233973;
assign addr[49500]= 2015345591;
assign addr[49501]= 2001818002;
assign addr[49502]= 1987655498;
assign addr[49503]= 1972862571;
assign addr[49504]= 1957443913;
assign addr[49505]= 1941404413;
assign addr[49506]= 1924749160;
assign addr[49507]= 1907483436;
assign addr[49508]= 1889612716;
assign addr[49509]= 1871142669;
assign addr[49510]= 1852079154;
assign addr[49511]= 1832428215;
assign addr[49512]= 1812196087;
assign addr[49513]= 1791389186;
assign addr[49514]= 1770014111;
assign addr[49515]= 1748077642;
assign addr[49516]= 1725586737;
assign addr[49517]= 1702548529;
assign addr[49518]= 1678970324;
assign addr[49519]= 1654859602;
assign addr[49520]= 1630224009;
assign addr[49521]= 1605071359;
assign addr[49522]= 1579409630;
assign addr[49523]= 1553246960;
assign addr[49524]= 1526591649;
assign addr[49525]= 1499452149;
assign addr[49526]= 1471837070;
assign addr[49527]= 1443755168;
assign addr[49528]= 1415215352;
assign addr[49529]= 1386226674;
assign addr[49530]= 1356798326;
assign addr[49531]= 1326939644;
assign addr[49532]= 1296660098;
assign addr[49533]= 1265969291;
assign addr[49534]= 1234876957;
assign addr[49535]= 1203392958;
assign addr[49536]= 1171527280;
assign addr[49537]= 1139290029;
assign addr[49538]= 1106691431;
assign addr[49539]= 1073741824;
assign addr[49540]= 1040451659;
assign addr[49541]= 1006831495;
assign addr[49542]= 972891995;
assign addr[49543]= 938643924;
assign addr[49544]= 904098143;
assign addr[49545]= 869265610;
assign addr[49546]= 834157373;
assign addr[49547]= 798784567;
assign addr[49548]= 763158411;
assign addr[49549]= 727290205;
assign addr[49550]= 691191324;
assign addr[49551]= 654873219;
assign addr[49552]= 618347408;
assign addr[49553]= 581625477;
assign addr[49554]= 544719071;
assign addr[49555]= 507639898;
assign addr[49556]= 470399716;
assign addr[49557]= 433010339;
assign addr[49558]= 395483624;
assign addr[49559]= 357831473;
assign addr[49560]= 320065829;
assign addr[49561]= 282198671;
assign addr[49562]= 244242007;
assign addr[49563]= 206207878;
assign addr[49564]= 168108346;
assign addr[49565]= 129955495;
assign addr[49566]= 91761426;
assign addr[49567]= 53538253;
assign addr[49568]= 15298099;
assign addr[49569]= -22946906;
assign addr[49570]= -61184634;
assign addr[49571]= -99402956;
assign addr[49572]= -137589750;
assign addr[49573]= -175732905;
assign addr[49574]= -213820322;
assign addr[49575]= -251839923;
assign addr[49576]= -289779648;
assign addr[49577]= -327627463;
assign addr[49578]= -365371365;
assign addr[49579]= -402999383;
assign addr[49580]= -440499581;
assign addr[49581]= -477860067;
assign addr[49582]= -515068990;
assign addr[49583]= -552114549;
assign addr[49584]= -588984994;
assign addr[49585]= -625668632;
assign addr[49586]= -662153826;
assign addr[49587]= -698429006;
assign addr[49588]= -734482665;
assign addr[49589]= -770303369;
assign addr[49590]= -805879757;
assign addr[49591]= -841200544;
assign addr[49592]= -876254528;
assign addr[49593]= -911030591;
assign addr[49594]= -945517704;
assign addr[49595]= -979704927;
assign addr[49596]= -1013581418;
assign addr[49597]= -1047136432;
assign addr[49598]= -1080359326;
assign addr[49599]= -1113239564;
assign addr[49600]= -1145766716;
assign addr[49601]= -1177930466;
assign addr[49602]= -1209720613;
assign addr[49603]= -1241127074;
assign addr[49604]= -1272139887;
assign addr[49605]= -1302749217;
assign addr[49606]= -1332945355;
assign addr[49607]= -1362718723;
assign addr[49608]= -1392059879;
assign addr[49609]= -1420959516;
assign addr[49610]= -1449408469;
assign addr[49611]= -1477397714;
assign addr[49612]= -1504918373;
assign addr[49613]= -1531961719;
assign addr[49614]= -1558519173;
assign addr[49615]= -1584582314;
assign addr[49616]= -1610142873;
assign addr[49617]= -1635192744;
assign addr[49618]= -1659723983;
assign addr[49619]= -1683728808;
assign addr[49620]= -1707199606;
assign addr[49621]= -1730128933;
assign addr[49622]= -1752509516;
assign addr[49623]= -1774334257;
assign addr[49624]= -1795596234;
assign addr[49625]= -1816288703;
assign addr[49626]= -1836405100;
assign addr[49627]= -1855939047;
assign addr[49628]= -1874884346;
assign addr[49629]= -1893234990;
assign addr[49630]= -1910985158;
assign addr[49631]= -1928129220;
assign addr[49632]= -1944661739;
assign addr[49633]= -1960577471;
assign addr[49634]= -1975871368;
assign addr[49635]= -1990538579;
assign addr[49636]= -2004574453;
assign addr[49637]= -2017974537;
assign addr[49638]= -2030734582;
assign addr[49639]= -2042850540;
assign addr[49640]= -2054318569;
assign addr[49641]= -2065135031;
assign addr[49642]= -2075296495;
assign addr[49643]= -2084799740;
assign addr[49644]= -2093641749;
assign addr[49645]= -2101819720;
assign addr[49646]= -2109331059;
assign addr[49647]= -2116173382;
assign addr[49648]= -2122344521;
assign addr[49649]= -2127842516;
assign addr[49650]= -2132665626;
assign addr[49651]= -2136812319;
assign addr[49652]= -2140281282;
assign addr[49653]= -2143071413;
assign addr[49654]= -2145181827;
assign addr[49655]= -2146611856;
assign addr[49656]= -2147361045;
assign addr[49657]= -2147429158;
assign addr[49658]= -2146816171;
assign addr[49659]= -2145522281;
assign addr[49660]= -2143547897;
assign addr[49661]= -2140893646;
assign addr[49662]= -2137560369;
assign addr[49663]= -2133549123;
assign addr[49664]= -2128861181;
assign addr[49665]= -2123498030;
assign addr[49666]= -2117461370;
assign addr[49667]= -2110753117;
assign addr[49668]= -2103375398;
assign addr[49669]= -2095330553;
assign addr[49670]= -2086621133;
assign addr[49671]= -2077249901;
assign addr[49672]= -2067219829;
assign addr[49673]= -2056534099;
assign addr[49674]= -2045196100;
assign addr[49675]= -2033209426;
assign addr[49676]= -2020577882;
assign addr[49677]= -2007305472;
assign addr[49678]= -1993396407;
assign addr[49679]= -1978855097;
assign addr[49680]= -1963686155;
assign addr[49681]= -1947894393;
assign addr[49682]= -1931484818;
assign addr[49683]= -1914462636;
assign addr[49684]= -1896833245;
assign addr[49685]= -1878602237;
assign addr[49686]= -1859775393;
assign addr[49687]= -1840358687;
assign addr[49688]= -1820358275;
assign addr[49689]= -1799780501;
assign addr[49690]= -1778631892;
assign addr[49691]= -1756919156;
assign addr[49692]= -1734649179;
assign addr[49693]= -1711829025;
assign addr[49694]= -1688465931;
assign addr[49695]= -1664567307;
assign addr[49696]= -1640140734;
assign addr[49697]= -1615193959;
assign addr[49698]= -1589734894;
assign addr[49699]= -1563771613;
assign addr[49700]= -1537312353;
assign addr[49701]= -1510365504;
assign addr[49702]= -1482939614;
assign addr[49703]= -1455043381;
assign addr[49704]= -1426685652;
assign addr[49705]= -1397875423;
assign addr[49706]= -1368621831;
assign addr[49707]= -1338934154;
assign addr[49708]= -1308821808;
assign addr[49709]= -1278294345;
assign addr[49710]= -1247361445;
assign addr[49711]= -1216032921;
assign addr[49712]= -1184318708;
assign addr[49713]= -1152228866;
assign addr[49714]= -1119773573;
assign addr[49715]= -1086963121;
assign addr[49716]= -1053807919;
assign addr[49717]= -1020318481;
assign addr[49718]= -986505429;
assign addr[49719]= -952379488;
assign addr[49720]= -917951481;
assign addr[49721]= -883232329;
assign addr[49722]= -848233042;
assign addr[49723]= -812964722;
assign addr[49724]= -777438554;
assign addr[49725]= -741665807;
assign addr[49726]= -705657826;
assign addr[49727]= -669426032;
assign addr[49728]= -632981917;
assign addr[49729]= -596337040;
assign addr[49730]= -559503022;
assign addr[49731]= -522491548;
assign addr[49732]= -485314355;
assign addr[49733]= -447983235;
assign addr[49734]= -410510029;
assign addr[49735]= -372906622;
assign addr[49736]= -335184940;
assign addr[49737]= -297356948;
assign addr[49738]= -259434643;
assign addr[49739]= -221430054;
assign addr[49740]= -183355234;
assign addr[49741]= -145222259;
assign addr[49742]= -107043224;
assign addr[49743]= -68830239;
assign addr[49744]= -30595422;
assign addr[49745]= 7649098;
assign addr[49746]= 45891193;
assign addr[49747]= 84118732;
assign addr[49748]= 122319591;
assign addr[49749]= 160481654;
assign addr[49750]= 198592817;
assign addr[49751]= 236640993;
assign addr[49752]= 274614114;
assign addr[49753]= 312500135;
assign addr[49754]= 350287041;
assign addr[49755]= 387962847;
assign addr[49756]= 425515602;
assign addr[49757]= 462933398;
assign addr[49758]= 500204365;
assign addr[49759]= 537316682;
assign addr[49760]= 574258580;
assign addr[49761]= 611018340;
assign addr[49762]= 647584304;
assign addr[49763]= 683944874;
assign addr[49764]= 720088517;
assign addr[49765]= 756003771;
assign addr[49766]= 791679244;
assign addr[49767]= 827103620;
assign addr[49768]= 862265664;
assign addr[49769]= 897154224;
assign addr[49770]= 931758235;
assign addr[49771]= 966066720;
assign addr[49772]= 1000068799;
assign addr[49773]= 1033753687;
assign addr[49774]= 1067110699;
assign addr[49775]= 1100129257;
assign addr[49776]= 1132798888;
assign addr[49777]= 1165109230;
assign addr[49778]= 1197050035;
assign addr[49779]= 1228611172;
assign addr[49780]= 1259782632;
assign addr[49781]= 1290554528;
assign addr[49782]= 1320917099;
assign addr[49783]= 1350860716;
assign addr[49784]= 1380375881;
assign addr[49785]= 1409453233;
assign addr[49786]= 1438083551;
assign addr[49787]= 1466257752;
assign addr[49788]= 1493966902;
assign addr[49789]= 1521202211;
assign addr[49790]= 1547955041;
assign addr[49791]= 1574216908;
assign addr[49792]= 1599979481;
assign addr[49793]= 1625234591;
assign addr[49794]= 1649974225;
assign addr[49795]= 1674190539;
assign addr[49796]= 1697875851;
assign addr[49797]= 1721022648;
assign addr[49798]= 1743623590;
assign addr[49799]= 1765671509;
assign addr[49800]= 1787159411;
assign addr[49801]= 1808080480;
assign addr[49802]= 1828428082;
assign addr[49803]= 1848195763;
assign addr[49804]= 1867377253;
assign addr[49805]= 1885966468;
assign addr[49806]= 1903957513;
assign addr[49807]= 1921344681;
assign addr[49808]= 1938122457;
assign addr[49809]= 1954285520;
assign addr[49810]= 1969828744;
assign addr[49811]= 1984747199;
assign addr[49812]= 1999036154;
assign addr[49813]= 2012691075;
assign addr[49814]= 2025707632;
assign addr[49815]= 2038081698;
assign addr[49816]= 2049809346;
assign addr[49817]= 2060886858;
assign addr[49818]= 2071310720;
assign addr[49819]= 2081077626;
assign addr[49820]= 2090184478;
assign addr[49821]= 2098628387;
assign addr[49822]= 2106406677;
assign addr[49823]= 2113516878;
assign addr[49824]= 2119956737;
assign addr[49825]= 2125724211;
assign addr[49826]= 2130817471;
assign addr[49827]= 2135234901;
assign addr[49828]= 2138975100;
assign addr[49829]= 2142036881;
assign addr[49830]= 2144419275;
assign addr[49831]= 2146121524;
assign addr[49832]= 2147143090;
assign addr[49833]= 2147483648;
assign addr[49834]= 2147143090;
assign addr[49835]= 2146121524;
assign addr[49836]= 2144419275;
assign addr[49837]= 2142036881;
assign addr[49838]= 2138975100;
assign addr[49839]= 2135234901;
assign addr[49840]= 2130817471;
assign addr[49841]= 2125724211;
assign addr[49842]= 2119956737;
assign addr[49843]= 2113516878;
assign addr[49844]= 2106406677;
assign addr[49845]= 2098628387;
assign addr[49846]= 2090184478;
assign addr[49847]= 2081077626;
assign addr[49848]= 2071310720;
assign addr[49849]= 2060886858;
assign addr[49850]= 2049809346;
assign addr[49851]= 2038081698;
assign addr[49852]= 2025707632;
assign addr[49853]= 2012691075;
assign addr[49854]= 1999036154;
assign addr[49855]= 1984747199;
assign addr[49856]= 1969828744;
assign addr[49857]= 1954285520;
assign addr[49858]= 1938122457;
assign addr[49859]= 1921344681;
assign addr[49860]= 1903957513;
assign addr[49861]= 1885966468;
assign addr[49862]= 1867377253;
assign addr[49863]= 1848195763;
assign addr[49864]= 1828428082;
assign addr[49865]= 1808080480;
assign addr[49866]= 1787159411;
assign addr[49867]= 1765671509;
assign addr[49868]= 1743623590;
assign addr[49869]= 1721022648;
assign addr[49870]= 1697875851;
assign addr[49871]= 1674190539;
assign addr[49872]= 1649974225;
assign addr[49873]= 1625234591;
assign addr[49874]= 1599979481;
assign addr[49875]= 1574216908;
assign addr[49876]= 1547955041;
assign addr[49877]= 1521202211;
assign addr[49878]= 1493966902;
assign addr[49879]= 1466257752;
assign addr[49880]= 1438083551;
assign addr[49881]= 1409453233;
assign addr[49882]= 1380375881;
assign addr[49883]= 1350860716;
assign addr[49884]= 1320917099;
assign addr[49885]= 1290554528;
assign addr[49886]= 1259782632;
assign addr[49887]= 1228611172;
assign addr[49888]= 1197050035;
assign addr[49889]= 1165109230;
assign addr[49890]= 1132798888;
assign addr[49891]= 1100129257;
assign addr[49892]= 1067110699;
assign addr[49893]= 1033753687;
assign addr[49894]= 1000068799;
assign addr[49895]= 966066720;
assign addr[49896]= 931758235;
assign addr[49897]= 897154224;
assign addr[49898]= 862265664;
assign addr[49899]= 827103620;
assign addr[49900]= 791679244;
assign addr[49901]= 756003771;
assign addr[49902]= 720088517;
assign addr[49903]= 683944874;
assign addr[49904]= 647584304;
assign addr[49905]= 611018340;
assign addr[49906]= 574258580;
assign addr[49907]= 537316682;
assign addr[49908]= 500204365;
assign addr[49909]= 462933398;
assign addr[49910]= 425515602;
assign addr[49911]= 387962847;
assign addr[49912]= 350287041;
assign addr[49913]= 312500135;
assign addr[49914]= 274614114;
assign addr[49915]= 236640993;
assign addr[49916]= 198592817;
assign addr[49917]= 160481654;
assign addr[49918]= 122319591;
assign addr[49919]= 84118732;
assign addr[49920]= 45891193;
assign addr[49921]= 7649098;
assign addr[49922]= -30595422;
assign addr[49923]= -68830239;
assign addr[49924]= -107043224;
assign addr[49925]= -145222259;
assign addr[49926]= -183355234;
assign addr[49927]= -221430054;
assign addr[49928]= -259434643;
assign addr[49929]= -297356948;
assign addr[49930]= -335184940;
assign addr[49931]= -372906622;
assign addr[49932]= -410510029;
assign addr[49933]= -447983235;
assign addr[49934]= -485314355;
assign addr[49935]= -522491548;
assign addr[49936]= -559503022;
assign addr[49937]= -596337040;
assign addr[49938]= -632981917;
assign addr[49939]= -669426032;
assign addr[49940]= -705657826;
assign addr[49941]= -741665807;
assign addr[49942]= -777438554;
assign addr[49943]= -812964722;
assign addr[49944]= -848233042;
assign addr[49945]= -883232329;
assign addr[49946]= -917951481;
assign addr[49947]= -952379488;
assign addr[49948]= -986505429;
assign addr[49949]= -1020318481;
assign addr[49950]= -1053807919;
assign addr[49951]= -1086963121;
assign addr[49952]= -1119773573;
assign addr[49953]= -1152228866;
assign addr[49954]= -1184318708;
assign addr[49955]= -1216032921;
assign addr[49956]= -1247361445;
assign addr[49957]= -1278294345;
assign addr[49958]= -1308821808;
assign addr[49959]= -1338934154;
assign addr[49960]= -1368621831;
assign addr[49961]= -1397875423;
assign addr[49962]= -1426685652;
assign addr[49963]= -1455043381;
assign addr[49964]= -1482939614;
assign addr[49965]= -1510365504;
assign addr[49966]= -1537312353;
assign addr[49967]= -1563771613;
assign addr[49968]= -1589734894;
assign addr[49969]= -1615193959;
assign addr[49970]= -1640140734;
assign addr[49971]= -1664567307;
assign addr[49972]= -1688465931;
assign addr[49973]= -1711829025;
assign addr[49974]= -1734649179;
assign addr[49975]= -1756919156;
assign addr[49976]= -1778631892;
assign addr[49977]= -1799780501;
assign addr[49978]= -1820358275;
assign addr[49979]= -1840358687;
assign addr[49980]= -1859775393;
assign addr[49981]= -1878602237;
assign addr[49982]= -1896833245;
assign addr[49983]= -1914462636;
assign addr[49984]= -1931484818;
assign addr[49985]= -1947894393;
assign addr[49986]= -1963686155;
assign addr[49987]= -1978855097;
assign addr[49988]= -1993396407;
assign addr[49989]= -2007305472;
assign addr[49990]= -2020577882;
assign addr[49991]= -2033209426;
assign addr[49992]= -2045196100;
assign addr[49993]= -2056534099;
assign addr[49994]= -2067219829;
assign addr[49995]= -2077249901;
assign addr[49996]= -2086621133;
assign addr[49997]= -2095330553;
assign addr[49998]= -2103375398;
assign addr[49999]= -2110753117;
assign addr[50000]= -2117461370;
assign addr[50001]= -2123498030;
assign addr[50002]= -2128861181;
assign addr[50003]= -2133549123;
assign addr[50004]= -2137560369;
assign addr[50005]= -2140893646;
assign addr[50006]= -2143547897;
assign addr[50007]= -2145522281;
assign addr[50008]= -2146816171;
assign addr[50009]= -2147429158;
assign addr[50010]= -2147361045;
assign addr[50011]= -2146611856;
assign addr[50012]= -2145181827;
assign addr[50013]= -2143071413;
assign addr[50014]= -2140281282;
assign addr[50015]= -2136812319;
assign addr[50016]= -2132665626;
assign addr[50017]= -2127842516;
assign addr[50018]= -2122344521;
assign addr[50019]= -2116173382;
assign addr[50020]= -2109331059;
assign addr[50021]= -2101819720;
assign addr[50022]= -2093641749;
assign addr[50023]= -2084799740;
assign addr[50024]= -2075296495;
assign addr[50025]= -2065135031;
assign addr[50026]= -2054318569;
assign addr[50027]= -2042850540;
assign addr[50028]= -2030734582;
assign addr[50029]= -2017974537;
assign addr[50030]= -2004574453;
assign addr[50031]= -1990538579;
assign addr[50032]= -1975871368;
assign addr[50033]= -1960577471;
assign addr[50034]= -1944661739;
assign addr[50035]= -1928129220;
assign addr[50036]= -1910985158;
assign addr[50037]= -1893234990;
assign addr[50038]= -1874884346;
assign addr[50039]= -1855939047;
assign addr[50040]= -1836405100;
assign addr[50041]= -1816288703;
assign addr[50042]= -1795596234;
assign addr[50043]= -1774334257;
assign addr[50044]= -1752509516;
assign addr[50045]= -1730128933;
assign addr[50046]= -1707199606;
assign addr[50047]= -1683728808;
assign addr[50048]= -1659723983;
assign addr[50049]= -1635192744;
assign addr[50050]= -1610142873;
assign addr[50051]= -1584582314;
assign addr[50052]= -1558519173;
assign addr[50053]= -1531961719;
assign addr[50054]= -1504918373;
assign addr[50055]= -1477397714;
assign addr[50056]= -1449408469;
assign addr[50057]= -1420959516;
assign addr[50058]= -1392059879;
assign addr[50059]= -1362718723;
assign addr[50060]= -1332945355;
assign addr[50061]= -1302749217;
assign addr[50062]= -1272139887;
assign addr[50063]= -1241127074;
assign addr[50064]= -1209720613;
assign addr[50065]= -1177930466;
assign addr[50066]= -1145766716;
assign addr[50067]= -1113239564;
assign addr[50068]= -1080359326;
assign addr[50069]= -1047136432;
assign addr[50070]= -1013581418;
assign addr[50071]= -979704927;
assign addr[50072]= -945517704;
assign addr[50073]= -911030591;
assign addr[50074]= -876254528;
assign addr[50075]= -841200544;
assign addr[50076]= -805879757;
assign addr[50077]= -770303369;
assign addr[50078]= -734482665;
assign addr[50079]= -698429006;
assign addr[50080]= -662153826;
assign addr[50081]= -625668632;
assign addr[50082]= -588984994;
assign addr[50083]= -552114549;
assign addr[50084]= -515068990;
assign addr[50085]= -477860067;
assign addr[50086]= -440499581;
assign addr[50087]= -402999383;
assign addr[50088]= -365371365;
assign addr[50089]= -327627463;
assign addr[50090]= -289779648;
assign addr[50091]= -251839923;
assign addr[50092]= -213820322;
assign addr[50093]= -175732905;
assign addr[50094]= -137589750;
assign addr[50095]= -99402956;
assign addr[50096]= -61184634;
assign addr[50097]= -22946906;
assign addr[50098]= 15298099;
assign addr[50099]= 53538253;
assign addr[50100]= 91761426;
assign addr[50101]= 129955495;
assign addr[50102]= 168108346;
assign addr[50103]= 206207878;
assign addr[50104]= 244242007;
assign addr[50105]= 282198671;
assign addr[50106]= 320065829;
assign addr[50107]= 357831473;
assign addr[50108]= 395483624;
assign addr[50109]= 433010339;
assign addr[50110]= 470399716;
assign addr[50111]= 507639898;
assign addr[50112]= 544719071;
assign addr[50113]= 581625477;
assign addr[50114]= 618347408;
assign addr[50115]= 654873219;
assign addr[50116]= 691191324;
assign addr[50117]= 727290205;
assign addr[50118]= 763158411;
assign addr[50119]= 798784567;
assign addr[50120]= 834157373;
assign addr[50121]= 869265610;
assign addr[50122]= 904098143;
assign addr[50123]= 938643924;
assign addr[50124]= 972891995;
assign addr[50125]= 1006831495;
assign addr[50126]= 1040451659;
assign addr[50127]= 1073741824;
assign addr[50128]= 1106691431;
assign addr[50129]= 1139290029;
assign addr[50130]= 1171527280;
assign addr[50131]= 1203392958;
assign addr[50132]= 1234876957;
assign addr[50133]= 1265969291;
assign addr[50134]= 1296660098;
assign addr[50135]= 1326939644;
assign addr[50136]= 1356798326;
assign addr[50137]= 1386226674;
assign addr[50138]= 1415215352;
assign addr[50139]= 1443755168;
assign addr[50140]= 1471837070;
assign addr[50141]= 1499452149;
assign addr[50142]= 1526591649;
assign addr[50143]= 1553246960;
assign addr[50144]= 1579409630;
assign addr[50145]= 1605071359;
assign addr[50146]= 1630224009;
assign addr[50147]= 1654859602;
assign addr[50148]= 1678970324;
assign addr[50149]= 1702548529;
assign addr[50150]= 1725586737;
assign addr[50151]= 1748077642;
assign addr[50152]= 1770014111;
assign addr[50153]= 1791389186;
assign addr[50154]= 1812196087;
assign addr[50155]= 1832428215;
assign addr[50156]= 1852079154;
assign addr[50157]= 1871142669;
assign addr[50158]= 1889612716;
assign addr[50159]= 1907483436;
assign addr[50160]= 1924749160;
assign addr[50161]= 1941404413;
assign addr[50162]= 1957443913;
assign addr[50163]= 1972862571;
assign addr[50164]= 1987655498;
assign addr[50165]= 2001818002;
assign addr[50166]= 2015345591;
assign addr[50167]= 2028233973;
assign addr[50168]= 2040479063;
assign addr[50169]= 2052076975;
assign addr[50170]= 2063024031;
assign addr[50171]= 2073316760;
assign addr[50172]= 2082951896;
assign addr[50173]= 2091926384;
assign addr[50174]= 2100237377;
assign addr[50175]= 2107882239;
assign addr[50176]= 2114858546;
assign addr[50177]= 2121164085;
assign addr[50178]= 2126796855;
assign addr[50179]= 2131755071;
assign addr[50180]= 2136037160;
assign addr[50181]= 2139641764;
assign addr[50182]= 2142567738;
assign addr[50183]= 2144814157;
assign addr[50184]= 2146380306;
assign addr[50185]= 2147265689;
assign addr[50186]= 2147470025;
assign addr[50187]= 2146993250;
assign addr[50188]= 2145835515;
assign addr[50189]= 2143997187;
assign addr[50190]= 2141478848;
assign addr[50191]= 2138281298;
assign addr[50192]= 2134405552;
assign addr[50193]= 2129852837;
assign addr[50194]= 2124624598;
assign addr[50195]= 2118722494;
assign addr[50196]= 2112148396;
assign addr[50197]= 2104904390;
assign addr[50198]= 2096992772;
assign addr[50199]= 2088416053;
assign addr[50200]= 2079176953;
assign addr[50201]= 2069278401;
assign addr[50202]= 2058723538;
assign addr[50203]= 2047515711;
assign addr[50204]= 2035658475;
assign addr[50205]= 2023155591;
assign addr[50206]= 2010011024;
assign addr[50207]= 1996228943;
assign addr[50208]= 1981813720;
assign addr[50209]= 1966769926;
assign addr[50210]= 1951102334;
assign addr[50211]= 1934815911;
assign addr[50212]= 1917915825;
assign addr[50213]= 1900407434;
assign addr[50214]= 1882296293;
assign addr[50215]= 1863588145;
assign addr[50216]= 1844288924;
assign addr[50217]= 1824404752;
assign addr[50218]= 1803941934;
assign addr[50219]= 1782906961;
assign addr[50220]= 1761306505;
assign addr[50221]= 1739147417;
assign addr[50222]= 1716436725;
assign addr[50223]= 1693181631;
assign addr[50224]= 1669389513;
assign addr[50225]= 1645067915;
assign addr[50226]= 1620224553;
assign addr[50227]= 1594867305;
assign addr[50228]= 1569004214;
assign addr[50229]= 1542643483;
assign addr[50230]= 1515793473;
assign addr[50231]= 1488462700;
assign addr[50232]= 1460659832;
assign addr[50233]= 1432393688;
assign addr[50234]= 1403673233;
assign addr[50235]= 1374507575;
assign addr[50236]= 1344905966;
assign addr[50237]= 1314877795;
assign addr[50238]= 1284432584;
assign addr[50239]= 1253579991;
assign addr[50240]= 1222329801;
assign addr[50241]= 1190691925;
assign addr[50242]= 1158676398;
assign addr[50243]= 1126293375;
assign addr[50244]= 1093553126;
assign addr[50245]= 1060466036;
assign addr[50246]= 1027042599;
assign addr[50247]= 993293415;
assign addr[50248]= 959229189;
assign addr[50249]= 924860725;
assign addr[50250]= 890198924;
assign addr[50251]= 855254778;
assign addr[50252]= 820039373;
assign addr[50253]= 784563876;
assign addr[50254]= 748839539;
assign addr[50255]= 712877694;
assign addr[50256]= 676689746;
assign addr[50257]= 640287172;
assign addr[50258]= 603681519;
assign addr[50259]= 566884397;
assign addr[50260]= 529907477;
assign addr[50261]= 492762486;
assign addr[50262]= 455461206;
assign addr[50263]= 418015468;
assign addr[50264]= 380437148;
assign addr[50265]= 342738165;
assign addr[50266]= 304930476;
assign addr[50267]= 267026072;
assign addr[50268]= 229036977;
assign addr[50269]= 190975237;
assign addr[50270]= 152852926;
assign addr[50271]= 114682135;
assign addr[50272]= 76474970;
assign addr[50273]= 38243550;
assign addr[50274]= 0;
assign addr[50275]= -38243550;
assign addr[50276]= -76474970;
assign addr[50277]= -114682135;
assign addr[50278]= -152852926;
assign addr[50279]= -190975237;
assign addr[50280]= -229036977;
assign addr[50281]= -267026072;
assign addr[50282]= -304930476;
assign addr[50283]= -342738165;
assign addr[50284]= -380437148;
assign addr[50285]= -418015468;
assign addr[50286]= -455461206;
assign addr[50287]= -492762486;
assign addr[50288]= -529907477;
assign addr[50289]= -566884397;
assign addr[50290]= -603681519;
assign addr[50291]= -640287172;
assign addr[50292]= -676689746;
assign addr[50293]= -712877694;
assign addr[50294]= -748839539;
assign addr[50295]= -784563876;
assign addr[50296]= -820039373;
assign addr[50297]= -855254778;
assign addr[50298]= -890198924;
assign addr[50299]= -924860725;
assign addr[50300]= -959229189;
assign addr[50301]= -993293415;
assign addr[50302]= -1027042599;
assign addr[50303]= -1060466036;
assign addr[50304]= -1093553126;
assign addr[50305]= -1126293375;
assign addr[50306]= -1158676398;
assign addr[50307]= -1190691925;
assign addr[50308]= -1222329801;
assign addr[50309]= -1253579991;
assign addr[50310]= -1284432584;
assign addr[50311]= -1314877795;
assign addr[50312]= -1344905966;
assign addr[50313]= -1374507575;
assign addr[50314]= -1403673233;
assign addr[50315]= -1432393688;
assign addr[50316]= -1460659832;
assign addr[50317]= -1488462700;
assign addr[50318]= -1515793473;
assign addr[50319]= -1542643483;
assign addr[50320]= -1569004214;
assign addr[50321]= -1594867305;
assign addr[50322]= -1620224553;
assign addr[50323]= -1645067915;
assign addr[50324]= -1669389513;
assign addr[50325]= -1693181631;
assign addr[50326]= -1716436725;
assign addr[50327]= -1739147417;
assign addr[50328]= -1761306505;
assign addr[50329]= -1782906961;
assign addr[50330]= -1803941934;
assign addr[50331]= -1824404752;
assign addr[50332]= -1844288924;
assign addr[50333]= -1863588145;
assign addr[50334]= -1882296293;
assign addr[50335]= -1900407434;
assign addr[50336]= -1917915825;
assign addr[50337]= -1934815911;
assign addr[50338]= -1951102334;
assign addr[50339]= -1966769926;
assign addr[50340]= -1981813720;
assign addr[50341]= -1996228943;
assign addr[50342]= -2010011024;
assign addr[50343]= -2023155591;
assign addr[50344]= -2035658475;
assign addr[50345]= -2047515711;
assign addr[50346]= -2058723538;
assign addr[50347]= -2069278401;
assign addr[50348]= -2079176953;
assign addr[50349]= -2088416053;
assign addr[50350]= -2096992772;
assign addr[50351]= -2104904390;
assign addr[50352]= -2112148396;
assign addr[50353]= -2118722494;
assign addr[50354]= -2124624598;
assign addr[50355]= -2129852837;
assign addr[50356]= -2134405552;
assign addr[50357]= -2138281298;
assign addr[50358]= -2141478848;
assign addr[50359]= -2143997187;
assign addr[50360]= -2145835515;
assign addr[50361]= -2146993250;
assign addr[50362]= -2147470025;
assign addr[50363]= -2147265689;
assign addr[50364]= -2146380306;
assign addr[50365]= -2144814157;
assign addr[50366]= -2142567738;
assign addr[50367]= -2139641764;
assign addr[50368]= -2136037160;
assign addr[50369]= -2131755071;
assign addr[50370]= -2126796855;
assign addr[50371]= -2121164085;
assign addr[50372]= -2114858546;
assign addr[50373]= -2107882239;
assign addr[50374]= -2100237377;
assign addr[50375]= -2091926384;
assign addr[50376]= -2082951896;
assign addr[50377]= -2073316760;
assign addr[50378]= -2063024031;
assign addr[50379]= -2052076975;
assign addr[50380]= -2040479063;
assign addr[50381]= -2028233973;
assign addr[50382]= -2015345591;
assign addr[50383]= -2001818002;
assign addr[50384]= -1987655498;
assign addr[50385]= -1972862571;
assign addr[50386]= -1957443913;
assign addr[50387]= -1941404413;
assign addr[50388]= -1924749160;
assign addr[50389]= -1907483436;
assign addr[50390]= -1889612716;
assign addr[50391]= -1871142669;
assign addr[50392]= -1852079154;
assign addr[50393]= -1832428215;
assign addr[50394]= -1812196087;
assign addr[50395]= -1791389186;
assign addr[50396]= -1770014111;
assign addr[50397]= -1748077642;
assign addr[50398]= -1725586737;
assign addr[50399]= -1702548529;
assign addr[50400]= -1678970324;
assign addr[50401]= -1654859602;
assign addr[50402]= -1630224009;
assign addr[50403]= -1605071359;
assign addr[50404]= -1579409630;
assign addr[50405]= -1553246960;
assign addr[50406]= -1526591649;
assign addr[50407]= -1499452149;
assign addr[50408]= -1471837070;
assign addr[50409]= -1443755168;
assign addr[50410]= -1415215352;
assign addr[50411]= -1386226674;
assign addr[50412]= -1356798326;
assign addr[50413]= -1326939644;
assign addr[50414]= -1296660098;
assign addr[50415]= -1265969291;
assign addr[50416]= -1234876957;
assign addr[50417]= -1203392958;
assign addr[50418]= -1171527280;
assign addr[50419]= -1139290029;
assign addr[50420]= -1106691431;
assign addr[50421]= -1073741824;
assign addr[50422]= -1040451659;
assign addr[50423]= -1006831495;
assign addr[50424]= -972891995;
assign addr[50425]= -938643924;
assign addr[50426]= -904098143;
assign addr[50427]= -869265610;
assign addr[50428]= -834157373;
assign addr[50429]= -798784567;
assign addr[50430]= -763158411;
assign addr[50431]= -727290205;
assign addr[50432]= -691191324;
assign addr[50433]= -654873219;
assign addr[50434]= -618347408;
assign addr[50435]= -581625477;
assign addr[50436]= -544719071;
assign addr[50437]= -507639898;
assign addr[50438]= -470399716;
assign addr[50439]= -433010339;
assign addr[50440]= -395483624;
assign addr[50441]= -357831473;
assign addr[50442]= -320065829;
assign addr[50443]= -282198671;
assign addr[50444]= -244242007;
assign addr[50445]= -206207878;
assign addr[50446]= -168108346;
assign addr[50447]= -129955495;
assign addr[50448]= -91761426;
assign addr[50449]= -53538253;
assign addr[50450]= -15298099;
assign addr[50451]= 22946906;
assign addr[50452]= 61184634;
assign addr[50453]= 99402956;
assign addr[50454]= 137589750;
assign addr[50455]= 175732905;
assign addr[50456]= 213820322;
assign addr[50457]= 251839923;
assign addr[50458]= 289779648;
assign addr[50459]= 327627463;
assign addr[50460]= 365371365;
assign addr[50461]= 402999383;
assign addr[50462]= 440499581;
assign addr[50463]= 477860067;
assign addr[50464]= 515068990;
assign addr[50465]= 552114549;
assign addr[50466]= 588984994;
assign addr[50467]= 625668632;
assign addr[50468]= 662153826;
assign addr[50469]= 698429006;
assign addr[50470]= 734482665;
assign addr[50471]= 770303369;
assign addr[50472]= 805879757;
assign addr[50473]= 841200544;
assign addr[50474]= 876254528;
assign addr[50475]= 911030591;
assign addr[50476]= 945517704;
assign addr[50477]= 979704927;
assign addr[50478]= 1013581418;
assign addr[50479]= 1047136432;
assign addr[50480]= 1080359326;
assign addr[50481]= 1113239564;
assign addr[50482]= 1145766716;
assign addr[50483]= 1177930466;
assign addr[50484]= 1209720613;
assign addr[50485]= 1241127074;
assign addr[50486]= 1272139887;
assign addr[50487]= 1302749217;
assign addr[50488]= 1332945355;
assign addr[50489]= 1362718723;
assign addr[50490]= 1392059879;
assign addr[50491]= 1420959516;
assign addr[50492]= 1449408469;
assign addr[50493]= 1477397714;
assign addr[50494]= 1504918373;
assign addr[50495]= 1531961719;
assign addr[50496]= 1558519173;
assign addr[50497]= 1584582314;
assign addr[50498]= 1610142873;
assign addr[50499]= 1635192744;
assign addr[50500]= 1659723983;
assign addr[50501]= 1683728808;
assign addr[50502]= 1707199606;
assign addr[50503]= 1730128933;
assign addr[50504]= 1752509516;
assign addr[50505]= 1774334257;
assign addr[50506]= 1795596234;
assign addr[50507]= 1816288703;
assign addr[50508]= 1836405100;
assign addr[50509]= 1855939047;
assign addr[50510]= 1874884346;
assign addr[50511]= 1893234990;
assign addr[50512]= 1910985158;
assign addr[50513]= 1928129220;
assign addr[50514]= 1944661739;
assign addr[50515]= 1960577471;
assign addr[50516]= 1975871368;
assign addr[50517]= 1990538579;
assign addr[50518]= 2004574453;
assign addr[50519]= 2017974537;
assign addr[50520]= 2030734582;
assign addr[50521]= 2042850540;
assign addr[50522]= 2054318569;
assign addr[50523]= 2065135031;
assign addr[50524]= 2075296495;
assign addr[50525]= 2084799740;
assign addr[50526]= 2093641749;
assign addr[50527]= 2101819720;
assign addr[50528]= 2109331059;
assign addr[50529]= 2116173382;
assign addr[50530]= 2122344521;
assign addr[50531]= 2127842516;
assign addr[50532]= 2132665626;
assign addr[50533]= 2136812319;
assign addr[50534]= 2140281282;
assign addr[50535]= 2143071413;
assign addr[50536]= 2145181827;
assign addr[50537]= 2146611856;
assign addr[50538]= 2147361045;
assign addr[50539]= 2147429158;
assign addr[50540]= 2146816171;
assign addr[50541]= 2145522281;
assign addr[50542]= 2143547897;
assign addr[50543]= 2140893646;
assign addr[50544]= 2137560369;
assign addr[50545]= 2133549123;
assign addr[50546]= 2128861181;
assign addr[50547]= 2123498030;
assign addr[50548]= 2117461370;
assign addr[50549]= 2110753117;
assign addr[50550]= 2103375398;
assign addr[50551]= 2095330553;
assign addr[50552]= 2086621133;
assign addr[50553]= 2077249901;
assign addr[50554]= 2067219829;
assign addr[50555]= 2056534099;
assign addr[50556]= 2045196100;
assign addr[50557]= 2033209426;
assign addr[50558]= 2020577882;
assign addr[50559]= 2007305472;
assign addr[50560]= 1993396407;
assign addr[50561]= 1978855097;
assign addr[50562]= 1963686155;
assign addr[50563]= 1947894393;
assign addr[50564]= 1931484818;
assign addr[50565]= 1914462636;
assign addr[50566]= 1896833245;
assign addr[50567]= 1878602237;
assign addr[50568]= 1859775393;
assign addr[50569]= 1840358687;
assign addr[50570]= 1820358275;
assign addr[50571]= 1799780501;
assign addr[50572]= 1778631892;
assign addr[50573]= 1756919156;
assign addr[50574]= 1734649179;
assign addr[50575]= 1711829025;
assign addr[50576]= 1688465931;
assign addr[50577]= 1664567307;
assign addr[50578]= 1640140734;
assign addr[50579]= 1615193959;
assign addr[50580]= 1589734894;
assign addr[50581]= 1563771613;
assign addr[50582]= 1537312353;
assign addr[50583]= 1510365504;
assign addr[50584]= 1482939614;
assign addr[50585]= 1455043381;
assign addr[50586]= 1426685652;
assign addr[50587]= 1397875423;
assign addr[50588]= 1368621831;
assign addr[50589]= 1338934154;
assign addr[50590]= 1308821808;
assign addr[50591]= 1278294345;
assign addr[50592]= 1247361445;
assign addr[50593]= 1216032921;
assign addr[50594]= 1184318708;
assign addr[50595]= 1152228866;
assign addr[50596]= 1119773573;
assign addr[50597]= 1086963121;
assign addr[50598]= 1053807919;
assign addr[50599]= 1020318481;
assign addr[50600]= 986505429;
assign addr[50601]= 952379488;
assign addr[50602]= 917951481;
assign addr[50603]= 883232329;
assign addr[50604]= 848233042;
assign addr[50605]= 812964722;
assign addr[50606]= 777438554;
assign addr[50607]= 741665807;
assign addr[50608]= 705657826;
assign addr[50609]= 669426032;
assign addr[50610]= 632981917;
assign addr[50611]= 596337040;
assign addr[50612]= 559503022;
assign addr[50613]= 522491548;
assign addr[50614]= 485314355;
assign addr[50615]= 447983235;
assign addr[50616]= 410510029;
assign addr[50617]= 372906622;
assign addr[50618]= 335184940;
assign addr[50619]= 297356948;
assign addr[50620]= 259434643;
assign addr[50621]= 221430054;
assign addr[50622]= 183355234;
assign addr[50623]= 145222259;
assign addr[50624]= 107043224;
assign addr[50625]= 68830239;
assign addr[50626]= 30595422;
assign addr[50627]= -7649098;
assign addr[50628]= -45891193;
assign addr[50629]= -84118732;
assign addr[50630]= -122319591;
assign addr[50631]= -160481654;
assign addr[50632]= -198592817;
assign addr[50633]= -236640993;
assign addr[50634]= -274614114;
assign addr[50635]= -312500135;
assign addr[50636]= -350287041;
assign addr[50637]= -387962847;
assign addr[50638]= -425515602;
assign addr[50639]= -462933398;
assign addr[50640]= -500204365;
assign addr[50641]= -537316682;
assign addr[50642]= -574258580;
assign addr[50643]= -611018340;
assign addr[50644]= -647584304;
assign addr[50645]= -683944874;
assign addr[50646]= -720088517;
assign addr[50647]= -756003771;
assign addr[50648]= -791679244;
assign addr[50649]= -827103620;
assign addr[50650]= -862265664;
assign addr[50651]= -897154224;
assign addr[50652]= -931758235;
assign addr[50653]= -966066720;
assign addr[50654]= -1000068799;
assign addr[50655]= -1033753687;
assign addr[50656]= -1067110699;
assign addr[50657]= -1100129257;
assign addr[50658]= -1132798888;
assign addr[50659]= -1165109230;
assign addr[50660]= -1197050035;
assign addr[50661]= -1228611172;
assign addr[50662]= -1259782632;
assign addr[50663]= -1290554528;
assign addr[50664]= -1320917099;
assign addr[50665]= -1350860716;
assign addr[50666]= -1380375881;
assign addr[50667]= -1409453233;
assign addr[50668]= -1438083551;
assign addr[50669]= -1466257752;
assign addr[50670]= -1493966902;
assign addr[50671]= -1521202211;
assign addr[50672]= -1547955041;
assign addr[50673]= -1574216908;
assign addr[50674]= -1599979481;
assign addr[50675]= -1625234591;
assign addr[50676]= -1649974225;
assign addr[50677]= -1674190539;
assign addr[50678]= -1697875851;
assign addr[50679]= -1721022648;
assign addr[50680]= -1743623590;
assign addr[50681]= -1765671509;
assign addr[50682]= -1787159411;
assign addr[50683]= -1808080480;
assign addr[50684]= -1828428082;
assign addr[50685]= -1848195763;
assign addr[50686]= -1867377253;
assign addr[50687]= -1885966468;
assign addr[50688]= -1903957513;
assign addr[50689]= -1921344681;
assign addr[50690]= -1938122457;
assign addr[50691]= -1954285520;
assign addr[50692]= -1969828744;
assign addr[50693]= -1984747199;
assign addr[50694]= -1999036154;
assign addr[50695]= -2012691075;
assign addr[50696]= -2025707632;
assign addr[50697]= -2038081698;
assign addr[50698]= -2049809346;
assign addr[50699]= -2060886858;
assign addr[50700]= -2071310720;
assign addr[50701]= -2081077626;
assign addr[50702]= -2090184478;
assign addr[50703]= -2098628387;
assign addr[50704]= -2106406677;
assign addr[50705]= -2113516878;
assign addr[50706]= -2119956737;
assign addr[50707]= -2125724211;
assign addr[50708]= -2130817471;
assign addr[50709]= -2135234901;
assign addr[50710]= -2138975100;
assign addr[50711]= -2142036881;
assign addr[50712]= -2144419275;
assign addr[50713]= -2146121524;
assign addr[50714]= -2147143090;
assign addr[50715]= -2147483648;
assign addr[50716]= -2147143090;
assign addr[50717]= -2146121524;
assign addr[50718]= -2144419275;
assign addr[50719]= -2142036881;
assign addr[50720]= -2138975100;
assign addr[50721]= -2135234901;
assign addr[50722]= -2130817471;
assign addr[50723]= -2125724211;
assign addr[50724]= -2119956737;
assign addr[50725]= -2113516878;
assign addr[50726]= -2106406677;
assign addr[50727]= -2098628387;
assign addr[50728]= -2090184478;
assign addr[50729]= -2081077626;
assign addr[50730]= -2071310720;
assign addr[50731]= -2060886858;
assign addr[50732]= -2049809346;
assign addr[50733]= -2038081698;
assign addr[50734]= -2025707632;
assign addr[50735]= -2012691075;
assign addr[50736]= -1999036154;
assign addr[50737]= -1984747199;
assign addr[50738]= -1969828744;
assign addr[50739]= -1954285520;
assign addr[50740]= -1938122457;
assign addr[50741]= -1921344681;
assign addr[50742]= -1903957513;
assign addr[50743]= -1885966468;
assign addr[50744]= -1867377253;
assign addr[50745]= -1848195763;
assign addr[50746]= -1828428082;
assign addr[50747]= -1808080480;
assign addr[50748]= -1787159411;
assign addr[50749]= -1765671509;
assign addr[50750]= -1743623590;
assign addr[50751]= -1721022648;
assign addr[50752]= -1697875851;
assign addr[50753]= -1674190539;
assign addr[50754]= -1649974225;
assign addr[50755]= -1625234591;
assign addr[50756]= -1599979481;
assign addr[50757]= -1574216908;
assign addr[50758]= -1547955041;
assign addr[50759]= -1521202211;
assign addr[50760]= -1493966902;
assign addr[50761]= -1466257752;
assign addr[50762]= -1438083551;
assign addr[50763]= -1409453233;
assign addr[50764]= -1380375881;
assign addr[50765]= -1350860716;
assign addr[50766]= -1320917099;
assign addr[50767]= -1290554528;
assign addr[50768]= -1259782632;
assign addr[50769]= -1228611172;
assign addr[50770]= -1197050035;
assign addr[50771]= -1165109230;
assign addr[50772]= -1132798888;
assign addr[50773]= -1100129257;
assign addr[50774]= -1067110699;
assign addr[50775]= -1033753687;
assign addr[50776]= -1000068799;
assign addr[50777]= -966066720;
assign addr[50778]= -931758235;
assign addr[50779]= -897154224;
assign addr[50780]= -862265664;
assign addr[50781]= -827103620;
assign addr[50782]= -791679244;
assign addr[50783]= -756003771;
assign addr[50784]= -720088517;
assign addr[50785]= -683944874;
assign addr[50786]= -647584304;
assign addr[50787]= -611018340;
assign addr[50788]= -574258580;
assign addr[50789]= -537316682;
assign addr[50790]= -500204365;
assign addr[50791]= -462933398;
assign addr[50792]= -425515602;
assign addr[50793]= -387962847;
assign addr[50794]= -350287041;
assign addr[50795]= -312500135;
assign addr[50796]= -274614114;
assign addr[50797]= -236640993;
assign addr[50798]= -198592817;
assign addr[50799]= -160481654;
assign addr[50800]= -122319591;
assign addr[50801]= -84118732;
assign addr[50802]= -45891193;
assign addr[50803]= -7649098;
assign addr[50804]= 30595422;
assign addr[50805]= 68830239;
assign addr[50806]= 107043224;
assign addr[50807]= 145222259;
assign addr[50808]= 183355234;
assign addr[50809]= 221430054;
assign addr[50810]= 259434643;
assign addr[50811]= 297356948;
assign addr[50812]= 335184940;
assign addr[50813]= 372906622;
assign addr[50814]= 410510029;
assign addr[50815]= 447983235;
assign addr[50816]= 485314355;
assign addr[50817]= 522491548;
assign addr[50818]= 559503022;
assign addr[50819]= 596337040;
assign addr[50820]= 632981917;
assign addr[50821]= 669426032;
assign addr[50822]= 705657826;
assign addr[50823]= 741665807;
assign addr[50824]= 777438554;
assign addr[50825]= 812964722;
assign addr[50826]= 848233042;
assign addr[50827]= 883232329;
assign addr[50828]= 917951481;
assign addr[50829]= 952379488;
assign addr[50830]= 986505429;
assign addr[50831]= 1020318481;
assign addr[50832]= 1053807919;
assign addr[50833]= 1086963121;
assign addr[50834]= 1119773573;
assign addr[50835]= 1152228866;
assign addr[50836]= 1184318708;
assign addr[50837]= 1216032921;
assign addr[50838]= 1247361445;
assign addr[50839]= 1278294345;
assign addr[50840]= 1308821808;
assign addr[50841]= 1338934154;
assign addr[50842]= 1368621831;
assign addr[50843]= 1397875423;
assign addr[50844]= 1426685652;
assign addr[50845]= 1455043381;
assign addr[50846]= 1482939614;
assign addr[50847]= 1510365504;
assign addr[50848]= 1537312353;
assign addr[50849]= 1563771613;
assign addr[50850]= 1589734894;
assign addr[50851]= 1615193959;
assign addr[50852]= 1640140734;
assign addr[50853]= 1664567307;
assign addr[50854]= 1688465931;
assign addr[50855]= 1711829025;
assign addr[50856]= 1734649179;
assign addr[50857]= 1756919156;
assign addr[50858]= 1778631892;
assign addr[50859]= 1799780501;
assign addr[50860]= 1820358275;
assign addr[50861]= 1840358687;
assign addr[50862]= 1859775393;
assign addr[50863]= 1878602237;
assign addr[50864]= 1896833245;
assign addr[50865]= 1914462636;
assign addr[50866]= 1931484818;
assign addr[50867]= 1947894393;
assign addr[50868]= 1963686155;
assign addr[50869]= 1978855097;
assign addr[50870]= 1993396407;
assign addr[50871]= 2007305472;
assign addr[50872]= 2020577882;
assign addr[50873]= 2033209426;
assign addr[50874]= 2045196100;
assign addr[50875]= 2056534099;
assign addr[50876]= 2067219829;
assign addr[50877]= 2077249901;
assign addr[50878]= 2086621133;
assign addr[50879]= 2095330553;
assign addr[50880]= 2103375398;
assign addr[50881]= 2110753117;
assign addr[50882]= 2117461370;
assign addr[50883]= 2123498030;
assign addr[50884]= 2128861181;
assign addr[50885]= 2133549123;
assign addr[50886]= 2137560369;
assign addr[50887]= 2140893646;
assign addr[50888]= 2143547897;
assign addr[50889]= 2145522281;
assign addr[50890]= 2146816171;
assign addr[50891]= 2147429158;
assign addr[50892]= 2147361045;
assign addr[50893]= 2146611856;
assign addr[50894]= 2145181827;
assign addr[50895]= 2143071413;
assign addr[50896]= 2140281282;
assign addr[50897]= 2136812319;
assign addr[50898]= 2132665626;
assign addr[50899]= 2127842516;
assign addr[50900]= 2122344521;
assign addr[50901]= 2116173382;
assign addr[50902]= 2109331059;
assign addr[50903]= 2101819720;
assign addr[50904]= 2093641749;
assign addr[50905]= 2084799740;
assign addr[50906]= 2075296495;
assign addr[50907]= 2065135031;
assign addr[50908]= 2054318569;
assign addr[50909]= 2042850540;
assign addr[50910]= 2030734582;
assign addr[50911]= 2017974537;
assign addr[50912]= 2004574453;
assign addr[50913]= 1990538579;
assign addr[50914]= 1975871368;
assign addr[50915]= 1960577471;
assign addr[50916]= 1944661739;
assign addr[50917]= 1928129220;
assign addr[50918]= 1910985158;
assign addr[50919]= 1893234990;
assign addr[50920]= 1874884346;
assign addr[50921]= 1855939047;
assign addr[50922]= 1836405100;
assign addr[50923]= 1816288703;
assign addr[50924]= 1795596234;
assign addr[50925]= 1774334257;
assign addr[50926]= 1752509516;
assign addr[50927]= 1730128933;
assign addr[50928]= 1707199606;
assign addr[50929]= 1683728808;
assign addr[50930]= 1659723983;
assign addr[50931]= 1635192744;
assign addr[50932]= 1610142873;
assign addr[50933]= 1584582314;
assign addr[50934]= 1558519173;
assign addr[50935]= 1531961719;
assign addr[50936]= 1504918373;
assign addr[50937]= 1477397714;
assign addr[50938]= 1449408469;
assign addr[50939]= 1420959516;
assign addr[50940]= 1392059879;
assign addr[50941]= 1362718723;
assign addr[50942]= 1332945355;
assign addr[50943]= 1302749217;
assign addr[50944]= 1272139887;
assign addr[50945]= 1241127074;
assign addr[50946]= 1209720613;
assign addr[50947]= 1177930466;
assign addr[50948]= 1145766716;
assign addr[50949]= 1113239564;
assign addr[50950]= 1080359326;
assign addr[50951]= 1047136432;
assign addr[50952]= 1013581418;
assign addr[50953]= 979704927;
assign addr[50954]= 945517704;
assign addr[50955]= 911030591;
assign addr[50956]= 876254528;
assign addr[50957]= 841200544;
assign addr[50958]= 805879757;
assign addr[50959]= 770303369;
assign addr[50960]= 734482665;
assign addr[50961]= 698429006;
assign addr[50962]= 662153826;
assign addr[50963]= 625668632;
assign addr[50964]= 588984994;
assign addr[50965]= 552114549;
assign addr[50966]= 515068990;
assign addr[50967]= 477860067;
assign addr[50968]= 440499581;
assign addr[50969]= 402999383;
assign addr[50970]= 365371365;
assign addr[50971]= 327627463;
assign addr[50972]= 289779648;
assign addr[50973]= 251839923;
assign addr[50974]= 213820322;
assign addr[50975]= 175732905;
assign addr[50976]= 137589750;
assign addr[50977]= 99402956;
assign addr[50978]= 61184634;
assign addr[50979]= 22946906;
assign addr[50980]= -15298099;
assign addr[50981]= -53538253;
assign addr[50982]= -91761426;
assign addr[50983]= -129955495;
assign addr[50984]= -168108346;
assign addr[50985]= -206207878;
assign addr[50986]= -244242007;
assign addr[50987]= -282198671;
assign addr[50988]= -320065829;
assign addr[50989]= -357831473;
assign addr[50990]= -395483624;
assign addr[50991]= -433010339;
assign addr[50992]= -470399716;
assign addr[50993]= -507639898;
assign addr[50994]= -544719071;
assign addr[50995]= -581625477;
assign addr[50996]= -618347408;
assign addr[50997]= -654873219;
assign addr[50998]= -691191324;
assign addr[50999]= -727290205;
assign addr[51000]= -763158411;
assign addr[51001]= -798784567;
assign addr[51002]= -834157373;
assign addr[51003]= -869265610;
assign addr[51004]= -904098143;
assign addr[51005]= -938643924;
assign addr[51006]= -972891995;
assign addr[51007]= -1006831495;
assign addr[51008]= -1040451659;
assign addr[51009]= -1073741824;
assign addr[51010]= -1106691431;
assign addr[51011]= -1139290029;
assign addr[51012]= -1171527280;
assign addr[51013]= -1203392958;
assign addr[51014]= -1234876957;
assign addr[51015]= -1265969291;
assign addr[51016]= -1296660098;
assign addr[51017]= -1326939644;
assign addr[51018]= -1356798326;
assign addr[51019]= -1386226674;
assign addr[51020]= -1415215352;
assign addr[51021]= -1443755168;
assign addr[51022]= -1471837070;
assign addr[51023]= -1499452149;
assign addr[51024]= -1526591649;
assign addr[51025]= -1553246960;
assign addr[51026]= -1579409630;
assign addr[51027]= -1605071359;
assign addr[51028]= -1630224009;
assign addr[51029]= -1654859602;
assign addr[51030]= -1678970324;
assign addr[51031]= -1702548529;
assign addr[51032]= -1725586737;
assign addr[51033]= -1748077642;
assign addr[51034]= -1770014111;
assign addr[51035]= -1791389186;
assign addr[51036]= -1812196087;
assign addr[51037]= -1832428215;
assign addr[51038]= -1852079154;
assign addr[51039]= -1871142669;
assign addr[51040]= -1889612716;
assign addr[51041]= -1907483436;
assign addr[51042]= -1924749160;
assign addr[51043]= -1941404413;
assign addr[51044]= -1957443913;
assign addr[51045]= -1972862571;
assign addr[51046]= -1987655498;
assign addr[51047]= -2001818002;
assign addr[51048]= -2015345591;
assign addr[51049]= -2028233973;
assign addr[51050]= -2040479063;
assign addr[51051]= -2052076975;
assign addr[51052]= -2063024031;
assign addr[51053]= -2073316760;
assign addr[51054]= -2082951896;
assign addr[51055]= -2091926384;
assign addr[51056]= -2100237377;
assign addr[51057]= -2107882239;
assign addr[51058]= -2114858546;
assign addr[51059]= -2121164085;
assign addr[51060]= -2126796855;
assign addr[51061]= -2131755071;
assign addr[51062]= -2136037160;
assign addr[51063]= -2139641764;
assign addr[51064]= -2142567738;
assign addr[51065]= -2144814157;
assign addr[51066]= -2146380306;
assign addr[51067]= -2147265689;
assign addr[51068]= -2147470025;
assign addr[51069]= -2146993250;
assign addr[51070]= -2145835515;
assign addr[51071]= -2143997187;
assign addr[51072]= -2141478848;
assign addr[51073]= -2138281298;
assign addr[51074]= -2134405552;
assign addr[51075]= -2129852837;
assign addr[51076]= -2124624598;
assign addr[51077]= -2118722494;
assign addr[51078]= -2112148396;
assign addr[51079]= -2104904390;
assign addr[51080]= -2096992772;
assign addr[51081]= -2088416053;
assign addr[51082]= -2079176953;
assign addr[51083]= -2069278401;
assign addr[51084]= -2058723538;
assign addr[51085]= -2047515711;
assign addr[51086]= -2035658475;
assign addr[51087]= -2023155591;
assign addr[51088]= -2010011024;
assign addr[51089]= -1996228943;
assign addr[51090]= -1981813720;
assign addr[51091]= -1966769926;
assign addr[51092]= -1951102334;
assign addr[51093]= -1934815911;
assign addr[51094]= -1917915825;
assign addr[51095]= -1900407434;
assign addr[51096]= -1882296293;
assign addr[51097]= -1863588145;
assign addr[51098]= -1844288924;
assign addr[51099]= -1824404752;
assign addr[51100]= -1803941934;
assign addr[51101]= -1782906961;
assign addr[51102]= -1761306505;
assign addr[51103]= -1739147417;
assign addr[51104]= -1716436725;
assign addr[51105]= -1693181631;
assign addr[51106]= -1669389513;
assign addr[51107]= -1645067915;
assign addr[51108]= -1620224553;
assign addr[51109]= -1594867305;
assign addr[51110]= -1569004214;
assign addr[51111]= -1542643483;
assign addr[51112]= -1515793473;
assign addr[51113]= -1488462700;
assign addr[51114]= -1460659832;
assign addr[51115]= -1432393688;
assign addr[51116]= -1403673233;
assign addr[51117]= -1374507575;
assign addr[51118]= -1344905966;
assign addr[51119]= -1314877795;
assign addr[51120]= -1284432584;
assign addr[51121]= -1253579991;
assign addr[51122]= -1222329801;
assign addr[51123]= -1190691925;
assign addr[51124]= -1158676398;
assign addr[51125]= -1126293375;
assign addr[51126]= -1093553126;
assign addr[51127]= -1060466036;
assign addr[51128]= -1027042599;
assign addr[51129]= -993293415;
assign addr[51130]= -959229189;
assign addr[51131]= -924860725;
assign addr[51132]= -890198924;
assign addr[51133]= -855254778;
assign addr[51134]= -820039373;
assign addr[51135]= -784563876;
assign addr[51136]= -748839539;
assign addr[51137]= -712877694;
assign addr[51138]= -676689746;
assign addr[51139]= -640287172;
assign addr[51140]= -603681519;
assign addr[51141]= -566884397;
assign addr[51142]= -529907477;
assign addr[51143]= -492762486;
assign addr[51144]= -455461206;
assign addr[51145]= -418015468;
assign addr[51146]= -380437148;
assign addr[51147]= -342738165;
assign addr[51148]= -304930476;
assign addr[51149]= -267026072;
assign addr[51150]= -229036977;
assign addr[51151]= -190975237;
assign addr[51152]= -152852926;
assign addr[51153]= -114682135;
assign addr[51154]= -76474970;
assign addr[51155]= -38243550;
assign addr[51156]= 0;
assign addr[51157]= 38243550;
assign addr[51158]= 76474970;
assign addr[51159]= 114682135;
assign addr[51160]= 152852926;
assign addr[51161]= 190975237;
assign addr[51162]= 229036977;
assign addr[51163]= 267026072;
assign addr[51164]= 304930476;
assign addr[51165]= 342738165;
assign addr[51166]= 380437148;
assign addr[51167]= 418015468;
assign addr[51168]= 455461206;
assign addr[51169]= 492762486;
assign addr[51170]= 529907477;
assign addr[51171]= 566884397;
assign addr[51172]= 603681519;
assign addr[51173]= 640287172;
assign addr[51174]= 676689746;
assign addr[51175]= 712877694;
assign addr[51176]= 748839539;
assign addr[51177]= 784563876;
assign addr[51178]= 820039373;
assign addr[51179]= 855254778;
assign addr[51180]= 890198924;
assign addr[51181]= 924860725;
assign addr[51182]= 959229189;
assign addr[51183]= 993293415;
assign addr[51184]= 1027042599;
assign addr[51185]= 1060466036;
assign addr[51186]= 1093553126;
assign addr[51187]= 1126293375;
assign addr[51188]= 1158676398;
assign addr[51189]= 1190691925;
assign addr[51190]= 1222329801;
assign addr[51191]= 1253579991;
assign addr[51192]= 1284432584;
assign addr[51193]= 1314877795;
assign addr[51194]= 1344905966;
assign addr[51195]= 1374507575;
assign addr[51196]= 1403673233;
assign addr[51197]= 1432393688;
assign addr[51198]= 1460659832;
assign addr[51199]= 1488462700;
assign addr[51200]= 1515793473;
assign addr[51201]= 1542643483;
assign addr[51202]= 1569004214;
assign addr[51203]= 1594867305;
assign addr[51204]= 1620224553;
assign addr[51205]= 1645067915;
assign addr[51206]= 1669389513;
assign addr[51207]= 1693181631;
assign addr[51208]= 1716436725;
assign addr[51209]= 1739147417;
assign addr[51210]= 1761306505;
assign addr[51211]= 1782906961;
assign addr[51212]= 1803941934;
assign addr[51213]= 1824404752;
assign addr[51214]= 1844288924;
assign addr[51215]= 1863588145;
assign addr[51216]= 1882296293;
assign addr[51217]= 1900407434;
assign addr[51218]= 1917915825;
assign addr[51219]= 1934815911;
assign addr[51220]= 1951102334;
assign addr[51221]= 1966769926;
assign addr[51222]= 1981813720;
assign addr[51223]= 1996228943;
assign addr[51224]= 2010011024;
assign addr[51225]= 2023155591;
assign addr[51226]= 2035658475;
assign addr[51227]= 2047515711;
assign addr[51228]= 2058723538;
assign addr[51229]= 2069278401;
assign addr[51230]= 2079176953;
assign addr[51231]= 2088416053;
assign addr[51232]= 2096992772;
assign addr[51233]= 2104904390;
assign addr[51234]= 2112148396;
assign addr[51235]= 2118722494;
assign addr[51236]= 2124624598;
assign addr[51237]= 2129852837;
assign addr[51238]= 2134405552;
assign addr[51239]= 2138281298;
assign addr[51240]= 2141478848;
assign addr[51241]= 2143997187;
assign addr[51242]= 2145835515;
assign addr[51243]= 2146993250;
assign addr[51244]= 2147470025;
assign addr[51245]= 2147265689;
assign addr[51246]= 2146380306;
assign addr[51247]= 2144814157;
assign addr[51248]= 2142567738;
assign addr[51249]= 2139641764;
assign addr[51250]= 2136037160;
assign addr[51251]= 2131755071;
assign addr[51252]= 2126796855;
assign addr[51253]= 2121164085;
assign addr[51254]= 2114858546;
assign addr[51255]= 2107882239;
assign addr[51256]= 2100237377;
assign addr[51257]= 2091926384;
assign addr[51258]= 2082951896;
assign addr[51259]= 2073316760;
assign addr[51260]= 2063024031;
assign addr[51261]= 2052076975;
assign addr[51262]= 2040479063;
assign addr[51263]= 2028233973;
assign addr[51264]= 2015345591;
assign addr[51265]= 2001818002;
assign addr[51266]= 1987655498;
assign addr[51267]= 1972862571;
assign addr[51268]= 1957443913;
assign addr[51269]= 1941404413;
assign addr[51270]= 1924749160;
assign addr[51271]= 1907483436;
assign addr[51272]= 1889612716;
assign addr[51273]= 1871142669;
assign addr[51274]= 1852079154;
assign addr[51275]= 1832428215;
assign addr[51276]= 1812196087;
assign addr[51277]= 1791389186;
assign addr[51278]= 1770014111;
assign addr[51279]= 1748077642;
assign addr[51280]= 1725586737;
assign addr[51281]= 1702548529;
assign addr[51282]= 1678970324;
assign addr[51283]= 1654859602;
assign addr[51284]= 1630224009;
assign addr[51285]= 1605071359;
assign addr[51286]= 1579409630;
assign addr[51287]= 1553246960;
assign addr[51288]= 1526591649;
assign addr[51289]= 1499452149;
assign addr[51290]= 1471837070;
assign addr[51291]= 1443755168;
assign addr[51292]= 1415215352;
assign addr[51293]= 1386226674;
assign addr[51294]= 1356798326;
assign addr[51295]= 1326939644;
assign addr[51296]= 1296660098;
assign addr[51297]= 1265969291;
assign addr[51298]= 1234876957;
assign addr[51299]= 1203392958;
assign addr[51300]= 1171527280;
assign addr[51301]= 1139290029;
assign addr[51302]= 1106691431;
assign addr[51303]= 1073741824;
assign addr[51304]= 1040451659;
assign addr[51305]= 1006831495;
assign addr[51306]= 972891995;
assign addr[51307]= 938643924;
assign addr[51308]= 904098143;
assign addr[51309]= 869265610;
assign addr[51310]= 834157373;
assign addr[51311]= 798784567;
assign addr[51312]= 763158411;
assign addr[51313]= 727290205;
assign addr[51314]= 691191324;
assign addr[51315]= 654873219;
assign addr[51316]= 618347408;
assign addr[51317]= 581625477;
assign addr[51318]= 544719071;
assign addr[51319]= 507639898;
assign addr[51320]= 470399716;
assign addr[51321]= 433010339;
assign addr[51322]= 395483624;
assign addr[51323]= 357831473;
assign addr[51324]= 320065829;
assign addr[51325]= 282198671;
assign addr[51326]= 244242007;
assign addr[51327]= 206207878;
assign addr[51328]= 168108346;
assign addr[51329]= 129955495;
assign addr[51330]= 91761426;
assign addr[51331]= 53538253;
assign addr[51332]= 15298099;
assign addr[51333]= -22946906;
assign addr[51334]= -61184634;
assign addr[51335]= -99402956;
assign addr[51336]= -137589750;
assign addr[51337]= -175732905;
assign addr[51338]= -213820322;
assign addr[51339]= -251839923;
assign addr[51340]= -289779648;
assign addr[51341]= -327627463;
assign addr[51342]= -365371365;
assign addr[51343]= -402999383;
assign addr[51344]= -440499581;
assign addr[51345]= -477860067;
assign addr[51346]= -515068990;
assign addr[51347]= -552114549;
assign addr[51348]= -588984994;
assign addr[51349]= -625668632;
assign addr[51350]= -662153826;
assign addr[51351]= -698429006;
assign addr[51352]= -734482665;
assign addr[51353]= -770303369;
assign addr[51354]= -805879757;
assign addr[51355]= -841200544;
assign addr[51356]= -876254528;
assign addr[51357]= -911030591;
assign addr[51358]= -945517704;
assign addr[51359]= -979704927;
assign addr[51360]= -1013581418;
assign addr[51361]= -1047136432;
assign addr[51362]= -1080359326;
assign addr[51363]= -1113239564;
assign addr[51364]= -1145766716;
assign addr[51365]= -1177930466;
assign addr[51366]= -1209720613;
assign addr[51367]= -1241127074;
assign addr[51368]= -1272139887;
assign addr[51369]= -1302749217;
assign addr[51370]= -1332945355;
assign addr[51371]= -1362718723;
assign addr[51372]= -1392059879;
assign addr[51373]= -1420959516;
assign addr[51374]= -1449408469;
assign addr[51375]= -1477397714;
assign addr[51376]= -1504918373;
assign addr[51377]= -1531961719;
assign addr[51378]= -1558519173;
assign addr[51379]= -1584582314;
assign addr[51380]= -1610142873;
assign addr[51381]= -1635192744;
assign addr[51382]= -1659723983;
assign addr[51383]= -1683728808;
assign addr[51384]= -1707199606;
assign addr[51385]= -1730128933;
assign addr[51386]= -1752509516;
assign addr[51387]= -1774334257;
assign addr[51388]= -1795596234;
assign addr[51389]= -1816288703;
assign addr[51390]= -1836405100;
assign addr[51391]= -1855939047;
assign addr[51392]= -1874884346;
assign addr[51393]= -1893234990;
assign addr[51394]= -1910985158;
assign addr[51395]= -1928129220;
assign addr[51396]= -1944661739;
assign addr[51397]= -1960577471;
assign addr[51398]= -1975871368;
assign addr[51399]= -1990538579;
assign addr[51400]= -2004574453;
assign addr[51401]= -2017974537;
assign addr[51402]= -2030734582;
assign addr[51403]= -2042850540;
assign addr[51404]= -2054318569;
assign addr[51405]= -2065135031;
assign addr[51406]= -2075296495;
assign addr[51407]= -2084799740;
assign addr[51408]= -2093641749;
assign addr[51409]= -2101819720;
assign addr[51410]= -2109331059;
assign addr[51411]= -2116173382;
assign addr[51412]= -2122344521;
assign addr[51413]= -2127842516;
assign addr[51414]= -2132665626;
assign addr[51415]= -2136812319;
assign addr[51416]= -2140281282;
assign addr[51417]= -2143071413;
assign addr[51418]= -2145181827;
assign addr[51419]= -2146611856;
assign addr[51420]= -2147361045;
assign addr[51421]= -2147429158;
assign addr[51422]= -2146816171;
assign addr[51423]= -2145522281;
assign addr[51424]= -2143547897;
assign addr[51425]= -2140893646;
assign addr[51426]= -2137560369;
assign addr[51427]= -2133549123;
assign addr[51428]= -2128861181;
assign addr[51429]= -2123498030;
assign addr[51430]= -2117461370;
assign addr[51431]= -2110753117;
assign addr[51432]= -2103375398;
assign addr[51433]= -2095330553;
assign addr[51434]= -2086621133;
assign addr[51435]= -2077249901;
assign addr[51436]= -2067219829;
assign addr[51437]= -2056534099;
assign addr[51438]= -2045196100;
assign addr[51439]= -2033209426;
assign addr[51440]= -2020577882;
assign addr[51441]= -2007305472;
assign addr[51442]= -1993396407;
assign addr[51443]= -1978855097;
assign addr[51444]= -1963686155;
assign addr[51445]= -1947894393;
assign addr[51446]= -1931484818;
assign addr[51447]= -1914462636;
assign addr[51448]= -1896833245;
assign addr[51449]= -1878602237;
assign addr[51450]= -1859775393;
assign addr[51451]= -1840358687;
assign addr[51452]= -1820358275;
assign addr[51453]= -1799780501;
assign addr[51454]= -1778631892;
assign addr[51455]= -1756919156;
assign addr[51456]= -1734649179;
assign addr[51457]= -1711829025;
assign addr[51458]= -1688465931;
assign addr[51459]= -1664567307;
assign addr[51460]= -1640140734;
assign addr[51461]= -1615193959;
assign addr[51462]= -1589734894;
assign addr[51463]= -1563771613;
assign addr[51464]= -1537312353;
assign addr[51465]= -1510365504;
assign addr[51466]= -1482939614;
assign addr[51467]= -1455043381;
assign addr[51468]= -1426685652;
assign addr[51469]= -1397875423;
assign addr[51470]= -1368621831;
assign addr[51471]= -1338934154;
assign addr[51472]= -1308821808;
assign addr[51473]= -1278294345;
assign addr[51474]= -1247361445;
assign addr[51475]= -1216032921;
assign addr[51476]= -1184318708;
assign addr[51477]= -1152228866;
assign addr[51478]= -1119773573;
assign addr[51479]= -1086963121;
assign addr[51480]= -1053807919;
assign addr[51481]= -1020318481;
assign addr[51482]= -986505429;
assign addr[51483]= -952379488;
assign addr[51484]= -917951481;
assign addr[51485]= -883232329;
assign addr[51486]= -848233042;
assign addr[51487]= -812964722;
assign addr[51488]= -777438554;
assign addr[51489]= -741665807;
assign addr[51490]= -705657826;
assign addr[51491]= -669426032;
assign addr[51492]= -632981917;
assign addr[51493]= -596337040;
assign addr[51494]= -559503022;
assign addr[51495]= -522491548;
assign addr[51496]= -485314355;
assign addr[51497]= -447983235;
assign addr[51498]= -410510029;
assign addr[51499]= -372906622;
assign addr[51500]= -335184940;
assign addr[51501]= -297356948;
assign addr[51502]= -259434643;
assign addr[51503]= -221430054;
assign addr[51504]= -183355234;
assign addr[51505]= -145222259;
assign addr[51506]= -107043224;
assign addr[51507]= -68830239;
assign addr[51508]= -30595422;
assign addr[51509]= 7649098;
assign addr[51510]= 45891193;
assign addr[51511]= 84118732;
assign addr[51512]= 122319591;
assign addr[51513]= 160481654;
assign addr[51514]= 198592817;
assign addr[51515]= 236640993;
assign addr[51516]= 274614114;
assign addr[51517]= 312500135;
assign addr[51518]= 350287041;
assign addr[51519]= 387962847;
assign addr[51520]= 425515602;
assign addr[51521]= 462933398;
assign addr[51522]= 500204365;
assign addr[51523]= 537316682;
assign addr[51524]= 574258580;
assign addr[51525]= 611018340;
assign addr[51526]= 647584304;
assign addr[51527]= 683944874;
assign addr[51528]= 720088517;
assign addr[51529]= 756003771;
assign addr[51530]= 791679244;
assign addr[51531]= 827103620;
assign addr[51532]= 862265664;
assign addr[51533]= 897154224;
assign addr[51534]= 931758235;
assign addr[51535]= 966066720;
assign addr[51536]= 1000068799;
assign addr[51537]= 1033753687;
assign addr[51538]= 1067110699;
assign addr[51539]= 1100129257;
assign addr[51540]= 1132798888;
assign addr[51541]= 1165109230;
assign addr[51542]= 1197050035;
assign addr[51543]= 1228611172;
assign addr[51544]= 1259782632;
assign addr[51545]= 1290554528;
assign addr[51546]= 1320917099;
assign addr[51547]= 1350860716;
assign addr[51548]= 1380375881;
assign addr[51549]= 1409453233;
assign addr[51550]= 1438083551;
assign addr[51551]= 1466257752;
assign addr[51552]= 1493966902;
assign addr[51553]= 1521202211;
assign addr[51554]= 1547955041;
assign addr[51555]= 1574216908;
assign addr[51556]= 1599979481;
assign addr[51557]= 1625234591;
assign addr[51558]= 1649974225;
assign addr[51559]= 1674190539;
assign addr[51560]= 1697875851;
assign addr[51561]= 1721022648;
assign addr[51562]= 1743623590;
assign addr[51563]= 1765671509;
assign addr[51564]= 1787159411;
assign addr[51565]= 1808080480;
assign addr[51566]= 1828428082;
assign addr[51567]= 1848195763;
assign addr[51568]= 1867377253;
assign addr[51569]= 1885966468;
assign addr[51570]= 1903957513;
assign addr[51571]= 1921344681;
assign addr[51572]= 1938122457;
assign addr[51573]= 1954285520;
assign addr[51574]= 1969828744;
assign addr[51575]= 1984747199;
assign addr[51576]= 1999036154;
assign addr[51577]= 2012691075;
assign addr[51578]= 2025707632;
assign addr[51579]= 2038081698;
assign addr[51580]= 2049809346;
assign addr[51581]= 2060886858;
assign addr[51582]= 2071310720;
assign addr[51583]= 2081077626;
assign addr[51584]= 2090184478;
assign addr[51585]= 2098628387;
assign addr[51586]= 2106406677;
assign addr[51587]= 2113516878;
assign addr[51588]= 2119956737;
assign addr[51589]= 2125724211;
assign addr[51590]= 2130817471;
assign addr[51591]= 2135234901;
assign addr[51592]= 2138975100;
assign addr[51593]= 2142036881;
assign addr[51594]= 2144419275;
assign addr[51595]= 2146121524;
assign addr[51596]= 2147143090;
assign addr[51597]= 2147483648;
assign addr[51598]= 2147143090;
assign addr[51599]= 2146121524;
assign addr[51600]= 2144419275;
assign addr[51601]= 2142036881;
assign addr[51602]= 2138975100;
assign addr[51603]= 2135234901;
assign addr[51604]= 2130817471;
assign addr[51605]= 2125724211;
assign addr[51606]= 2119956737;
assign addr[51607]= 2113516878;
assign addr[51608]= 2106406677;
assign addr[51609]= 2098628387;
assign addr[51610]= 2090184478;
assign addr[51611]= 2081077626;
assign addr[51612]= 2071310720;
assign addr[51613]= 2060886858;
assign addr[51614]= 2049809346;
assign addr[51615]= 2038081698;
assign addr[51616]= 2025707632;
assign addr[51617]= 2012691075;
assign addr[51618]= 1999036154;
assign addr[51619]= 1984747199;
assign addr[51620]= 1969828744;
assign addr[51621]= 1954285520;
assign addr[51622]= 1938122457;
assign addr[51623]= 1921344681;
assign addr[51624]= 1903957513;
assign addr[51625]= 1885966468;
assign addr[51626]= 1867377253;
assign addr[51627]= 1848195763;
assign addr[51628]= 1828428082;
assign addr[51629]= 1808080480;
assign addr[51630]= 1787159411;
assign addr[51631]= 1765671509;
assign addr[51632]= 1743623590;
assign addr[51633]= 1721022648;
assign addr[51634]= 1697875851;
assign addr[51635]= 1674190539;
assign addr[51636]= 1649974225;
assign addr[51637]= 1625234591;
assign addr[51638]= 1599979481;
assign addr[51639]= 1574216908;
assign addr[51640]= 1547955041;
assign addr[51641]= 1521202211;
assign addr[51642]= 1493966902;
assign addr[51643]= 1466257752;
assign addr[51644]= 1438083551;
assign addr[51645]= 1409453233;
assign addr[51646]= 1380375881;
assign addr[51647]= 1350860716;
assign addr[51648]= 1320917099;
assign addr[51649]= 1290554528;
assign addr[51650]= 1259782632;
assign addr[51651]= 1228611172;
assign addr[51652]= 1197050035;
assign addr[51653]= 1165109230;
assign addr[51654]= 1132798888;
assign addr[51655]= 1100129257;
assign addr[51656]= 1067110699;
assign addr[51657]= 1033753687;
assign addr[51658]= 1000068799;
assign addr[51659]= 966066720;
assign addr[51660]= 931758235;
assign addr[51661]= 897154224;
assign addr[51662]= 862265664;
assign addr[51663]= 827103620;
assign addr[51664]= 791679244;
assign addr[51665]= 756003771;
assign addr[51666]= 720088517;
assign addr[51667]= 683944874;
assign addr[51668]= 647584304;
assign addr[51669]= 611018340;
assign addr[51670]= 574258580;
assign addr[51671]= 537316682;
assign addr[51672]= 500204365;
assign addr[51673]= 462933398;
assign addr[51674]= 425515602;
assign addr[51675]= 387962847;
assign addr[51676]= 350287041;
assign addr[51677]= 312500135;
assign addr[51678]= 274614114;
assign addr[51679]= 236640993;
assign addr[51680]= 198592817;
assign addr[51681]= 160481654;
assign addr[51682]= 122319591;
assign addr[51683]= 84118732;
assign addr[51684]= 45891193;
assign addr[51685]= 7649098;
assign addr[51686]= -30595422;
assign addr[51687]= -68830239;
assign addr[51688]= -107043224;
assign addr[51689]= -145222259;
assign addr[51690]= -183355234;
assign addr[51691]= -221430054;
assign addr[51692]= -259434643;
assign addr[51693]= -297356948;
assign addr[51694]= -335184940;
assign addr[51695]= -372906622;
assign addr[51696]= -410510029;
assign addr[51697]= -447983235;
assign addr[51698]= -485314355;
assign addr[51699]= -522491548;
assign addr[51700]= -559503022;
assign addr[51701]= -596337040;
assign addr[51702]= -632981917;
assign addr[51703]= -669426032;
assign addr[51704]= -705657826;
assign addr[51705]= -741665807;
assign addr[51706]= -777438554;
assign addr[51707]= -812964722;
assign addr[51708]= -848233042;
assign addr[51709]= -883232329;
assign addr[51710]= -917951481;
assign addr[51711]= -952379488;
assign addr[51712]= -986505429;
assign addr[51713]= -1020318481;
assign addr[51714]= -1053807919;
assign addr[51715]= -1086963121;
assign addr[51716]= -1119773573;
assign addr[51717]= -1152228866;
assign addr[51718]= -1184318708;
assign addr[51719]= -1216032921;
assign addr[51720]= -1247361445;
assign addr[51721]= -1278294345;
assign addr[51722]= -1308821808;
assign addr[51723]= -1338934154;
assign addr[51724]= -1368621831;
assign addr[51725]= -1397875423;
assign addr[51726]= -1426685652;
assign addr[51727]= -1455043381;
assign addr[51728]= -1482939614;
assign addr[51729]= -1510365504;
assign addr[51730]= -1537312353;
assign addr[51731]= -1563771613;
assign addr[51732]= -1589734894;
assign addr[51733]= -1615193959;
assign addr[51734]= -1640140734;
assign addr[51735]= -1664567307;
assign addr[51736]= -1688465931;
assign addr[51737]= -1711829025;
assign addr[51738]= -1734649179;
assign addr[51739]= -1756919156;
assign addr[51740]= -1778631892;
assign addr[51741]= -1799780501;
assign addr[51742]= -1820358275;
assign addr[51743]= -1840358687;
assign addr[51744]= -1859775393;
assign addr[51745]= -1878602237;
assign addr[51746]= -1896833245;
assign addr[51747]= -1914462636;
assign addr[51748]= -1931484818;
assign addr[51749]= -1947894393;
assign addr[51750]= -1963686155;
assign addr[51751]= -1978855097;
assign addr[51752]= -1993396407;
assign addr[51753]= -2007305472;
assign addr[51754]= -2020577882;
assign addr[51755]= -2033209426;
assign addr[51756]= -2045196100;
assign addr[51757]= -2056534099;
assign addr[51758]= -2067219829;
assign addr[51759]= -2077249901;
assign addr[51760]= -2086621133;
assign addr[51761]= -2095330553;
assign addr[51762]= -2103375398;
assign addr[51763]= -2110753117;
assign addr[51764]= -2117461370;
assign addr[51765]= -2123498030;
assign addr[51766]= -2128861181;
assign addr[51767]= -2133549123;
assign addr[51768]= -2137560369;
assign addr[51769]= -2140893646;
assign addr[51770]= -2143547897;
assign addr[51771]= -2145522281;
assign addr[51772]= -2146816171;
assign addr[51773]= -2147429158;
assign addr[51774]= -2147361045;
assign addr[51775]= -2146611856;
assign addr[51776]= -2145181827;
assign addr[51777]= -2143071413;
assign addr[51778]= -2140281282;
assign addr[51779]= -2136812319;
assign addr[51780]= -2132665626;
assign addr[51781]= -2127842516;
assign addr[51782]= -2122344521;
assign addr[51783]= -2116173382;
assign addr[51784]= -2109331059;
assign addr[51785]= -2101819720;
assign addr[51786]= -2093641749;
assign addr[51787]= -2084799740;
assign addr[51788]= -2075296495;
assign addr[51789]= -2065135031;
assign addr[51790]= -2054318569;
assign addr[51791]= -2042850540;
assign addr[51792]= -2030734582;
assign addr[51793]= -2017974537;
assign addr[51794]= -2004574453;
assign addr[51795]= -1990538579;
assign addr[51796]= -1975871368;
assign addr[51797]= -1960577471;
assign addr[51798]= -1944661739;
assign addr[51799]= -1928129220;
assign addr[51800]= -1910985158;
assign addr[51801]= -1893234990;
assign addr[51802]= -1874884346;
assign addr[51803]= -1855939047;
assign addr[51804]= -1836405100;
assign addr[51805]= -1816288703;
assign addr[51806]= -1795596234;
assign addr[51807]= -1774334257;
assign addr[51808]= -1752509516;
assign addr[51809]= -1730128933;
assign addr[51810]= -1707199606;
assign addr[51811]= -1683728808;
assign addr[51812]= -1659723983;
assign addr[51813]= -1635192744;
assign addr[51814]= -1610142873;
assign addr[51815]= -1584582314;
assign addr[51816]= -1558519173;
assign addr[51817]= -1531961719;
assign addr[51818]= -1504918373;
assign addr[51819]= -1477397714;
assign addr[51820]= -1449408469;
assign addr[51821]= -1420959516;
assign addr[51822]= -1392059879;
assign addr[51823]= -1362718723;
assign addr[51824]= -1332945355;
assign addr[51825]= -1302749217;
assign addr[51826]= -1272139887;
assign addr[51827]= -1241127074;
assign addr[51828]= -1209720613;
assign addr[51829]= -1177930466;
assign addr[51830]= -1145766716;
assign addr[51831]= -1113239564;
assign addr[51832]= -1080359326;
assign addr[51833]= -1047136432;
assign addr[51834]= -1013581418;
assign addr[51835]= -979704927;
assign addr[51836]= -945517704;
assign addr[51837]= -911030591;
assign addr[51838]= -876254528;
assign addr[51839]= -841200544;
assign addr[51840]= -805879757;
assign addr[51841]= -770303369;
assign addr[51842]= -734482665;
assign addr[51843]= -698429006;
assign addr[51844]= -662153826;
assign addr[51845]= -625668632;
assign addr[51846]= -588984994;
assign addr[51847]= -552114549;
assign addr[51848]= -515068990;
assign addr[51849]= -477860067;
assign addr[51850]= -440499581;
assign addr[51851]= -402999383;
assign addr[51852]= -365371365;
assign addr[51853]= -327627463;
assign addr[51854]= -289779648;
assign addr[51855]= -251839923;
assign addr[51856]= -213820322;
assign addr[51857]= -175732905;
assign addr[51858]= -137589750;
assign addr[51859]= -99402956;
assign addr[51860]= -61184634;
assign addr[51861]= -22946906;
assign addr[51862]= 15298099;
assign addr[51863]= 53538253;
assign addr[51864]= 91761426;
assign addr[51865]= 129955495;
assign addr[51866]= 168108346;
assign addr[51867]= 206207878;
assign addr[51868]= 244242007;
assign addr[51869]= 282198671;
assign addr[51870]= 320065829;
assign addr[51871]= 357831473;
assign addr[51872]= 395483624;
assign addr[51873]= 433010339;
assign addr[51874]= 470399716;
assign addr[51875]= 507639898;
assign addr[51876]= 544719071;
assign addr[51877]= 581625477;
assign addr[51878]= 618347408;
assign addr[51879]= 654873219;
assign addr[51880]= 691191324;
assign addr[51881]= 727290205;
assign addr[51882]= 763158411;
assign addr[51883]= 798784567;
assign addr[51884]= 834157373;
assign addr[51885]= 869265610;
assign addr[51886]= 904098143;
assign addr[51887]= 938643924;
assign addr[51888]= 972891995;
assign addr[51889]= 1006831495;
assign addr[51890]= 1040451659;
assign addr[51891]= 1073741824;
assign addr[51892]= 1106691431;
assign addr[51893]= 1139290029;
assign addr[51894]= 1171527280;
assign addr[51895]= 1203392958;
assign addr[51896]= 1234876957;
assign addr[51897]= 1265969291;
assign addr[51898]= 1296660098;
assign addr[51899]= 1326939644;
assign addr[51900]= 1356798326;
assign addr[51901]= 1386226674;
assign addr[51902]= 1415215352;
assign addr[51903]= 1443755168;
assign addr[51904]= 1471837070;
assign addr[51905]= 1499452149;
assign addr[51906]= 1526591649;
assign addr[51907]= 1553246960;
assign addr[51908]= 1579409630;
assign addr[51909]= 1605071359;
assign addr[51910]= 1630224009;
assign addr[51911]= 1654859602;
assign addr[51912]= 1678970324;
assign addr[51913]= 1702548529;
assign addr[51914]= 1725586737;
assign addr[51915]= 1748077642;
assign addr[51916]= 1770014111;
assign addr[51917]= 1791389186;
assign addr[51918]= 1812196087;
assign addr[51919]= 1832428215;
assign addr[51920]= 1852079154;
assign addr[51921]= 1871142669;
assign addr[51922]= 1889612716;
assign addr[51923]= 1907483436;
assign addr[51924]= 1924749160;
assign addr[51925]= 1941404413;
assign addr[51926]= 1957443913;
assign addr[51927]= 1972862571;
assign addr[51928]= 1987655498;
assign addr[51929]= 2001818002;
assign addr[51930]= 2015345591;
assign addr[51931]= 2028233973;
assign addr[51932]= 2040479063;
assign addr[51933]= 2052076975;
assign addr[51934]= 2063024031;
assign addr[51935]= 2073316760;
assign addr[51936]= 2082951896;
assign addr[51937]= 2091926384;
assign addr[51938]= 2100237377;
assign addr[51939]= 2107882239;
assign addr[51940]= 2114858546;
assign addr[51941]= 2121164085;
assign addr[51942]= 2126796855;
assign addr[51943]= 2131755071;
assign addr[51944]= 2136037160;
assign addr[51945]= 2139641764;
assign addr[51946]= 2142567738;
assign addr[51947]= 2144814157;
assign addr[51948]= 2146380306;
assign addr[51949]= 2147265689;
assign addr[51950]= 2147470025;
assign addr[51951]= 2146993250;
assign addr[51952]= 2145835515;
assign addr[51953]= 2143997187;
assign addr[51954]= 2141478848;
assign addr[51955]= 2138281298;
assign addr[51956]= 2134405552;
assign addr[51957]= 2129852837;
assign addr[51958]= 2124624598;
assign addr[51959]= 2118722494;
assign addr[51960]= 2112148396;
assign addr[51961]= 2104904390;
assign addr[51962]= 2096992772;
assign addr[51963]= 2088416053;
assign addr[51964]= 2079176953;
assign addr[51965]= 2069278401;
assign addr[51966]= 2058723538;
assign addr[51967]= 2047515711;
assign addr[51968]= 2035658475;
assign addr[51969]= 2023155591;
assign addr[51970]= 2010011024;
assign addr[51971]= 1996228943;
assign addr[51972]= 1981813720;
assign addr[51973]= 1966769926;
assign addr[51974]= 1951102334;
assign addr[51975]= 1934815911;
assign addr[51976]= 1917915825;
assign addr[51977]= 1900407434;
assign addr[51978]= 1882296293;
assign addr[51979]= 1863588145;
assign addr[51980]= 1844288924;
assign addr[51981]= 1824404752;
assign addr[51982]= 1803941934;
assign addr[51983]= 1782906961;
assign addr[51984]= 1761306505;
assign addr[51985]= 1739147417;
assign addr[51986]= 1716436725;
assign addr[51987]= 1693181631;
assign addr[51988]= 1669389513;
assign addr[51989]= 1645067915;
assign addr[51990]= 1620224553;
assign addr[51991]= 1594867305;
assign addr[51992]= 1569004214;
assign addr[51993]= 1542643483;
assign addr[51994]= 1515793473;
assign addr[51995]= 1488462700;
assign addr[51996]= 1460659832;
assign addr[51997]= 1432393688;
assign addr[51998]= 1403673233;
assign addr[51999]= 1374507575;
assign addr[52000]= 1344905966;
assign addr[52001]= 1314877795;
assign addr[52002]= 1284432584;
assign addr[52003]= 1253579991;
assign addr[52004]= 1222329801;
assign addr[52005]= 1190691925;
assign addr[52006]= 1158676398;
assign addr[52007]= 1126293375;
assign addr[52008]= 1093553126;
assign addr[52009]= 1060466036;
assign addr[52010]= 1027042599;
assign addr[52011]= 993293415;
assign addr[52012]= 959229189;
assign addr[52013]= 924860725;
assign addr[52014]= 890198924;
assign addr[52015]= 855254778;
assign addr[52016]= 820039373;
assign addr[52017]= 784563876;
assign addr[52018]= 748839539;
assign addr[52019]= 712877694;
assign addr[52020]= 676689746;
assign addr[52021]= 640287172;
assign addr[52022]= 603681519;
assign addr[52023]= 566884397;
assign addr[52024]= 529907477;
assign addr[52025]= 492762486;
assign addr[52026]= 455461206;
assign addr[52027]= 418015468;
assign addr[52028]= 380437148;
assign addr[52029]= 342738165;
assign addr[52030]= 304930476;
assign addr[52031]= 267026072;
assign addr[52032]= 229036977;
assign addr[52033]= 190975237;
assign addr[52034]= 152852926;
assign addr[52035]= 114682135;
assign addr[52036]= 76474970;
assign addr[52037]= 38243550;
assign addr[52038]= 0;
assign addr[52039]= -38243550;
assign addr[52040]= -76474970;
assign addr[52041]= -114682135;
assign addr[52042]= -152852926;
assign addr[52043]= -190975237;
assign addr[52044]= -229036977;
assign addr[52045]= -267026072;
assign addr[52046]= -304930476;
assign addr[52047]= -342738165;
assign addr[52048]= -380437148;
assign addr[52049]= -418015468;
assign addr[52050]= -455461206;
assign addr[52051]= -492762486;
assign addr[52052]= -529907477;
assign addr[52053]= -566884397;
assign addr[52054]= -603681519;
assign addr[52055]= -640287172;
assign addr[52056]= -676689746;
assign addr[52057]= -712877694;
assign addr[52058]= -748839539;
assign addr[52059]= -784563876;
assign addr[52060]= -820039373;
assign addr[52061]= -855254778;
assign addr[52062]= -890198924;
assign addr[52063]= -924860725;
assign addr[52064]= -959229189;
assign addr[52065]= -993293415;
assign addr[52066]= -1027042599;
assign addr[52067]= -1060466036;
assign addr[52068]= -1093553126;
assign addr[52069]= -1126293375;
assign addr[52070]= -1158676398;
assign addr[52071]= -1190691925;
assign addr[52072]= -1222329801;
assign addr[52073]= -1253579991;
assign addr[52074]= -1284432584;
assign addr[52075]= -1314877795;
assign addr[52076]= -1344905966;
assign addr[52077]= -1374507575;
assign addr[52078]= -1403673233;
assign addr[52079]= -1432393688;
assign addr[52080]= -1460659832;
assign addr[52081]= -1488462700;
assign addr[52082]= -1515793473;
assign addr[52083]= -1542643483;
assign addr[52084]= -1569004214;
assign addr[52085]= -1594867305;
assign addr[52086]= -1620224553;
assign addr[52087]= -1645067915;
assign addr[52088]= -1669389513;
assign addr[52089]= -1693181631;
assign addr[52090]= -1716436725;
assign addr[52091]= -1739147417;
assign addr[52092]= -1761306505;
assign addr[52093]= -1782906961;
assign addr[52094]= -1803941934;
assign addr[52095]= -1824404752;
assign addr[52096]= -1844288924;
assign addr[52097]= -1863588145;
assign addr[52098]= -1882296293;
assign addr[52099]= -1900407434;
assign addr[52100]= -1917915825;
assign addr[52101]= -1934815911;
assign addr[52102]= -1951102334;
assign addr[52103]= -1966769926;
assign addr[52104]= -1981813720;
assign addr[52105]= -1996228943;
assign addr[52106]= -2010011024;
assign addr[52107]= -2023155591;
assign addr[52108]= -2035658475;
assign addr[52109]= -2047515711;
assign addr[52110]= -2058723538;
assign addr[52111]= -2069278401;
assign addr[52112]= -2079176953;
assign addr[52113]= -2088416053;
assign addr[52114]= -2096992772;
assign addr[52115]= -2104904390;
assign addr[52116]= -2112148396;
assign addr[52117]= -2118722494;
assign addr[52118]= -2124624598;
assign addr[52119]= -2129852837;
assign addr[52120]= -2134405552;
assign addr[52121]= -2138281298;
assign addr[52122]= -2141478848;
assign addr[52123]= -2143997187;
assign addr[52124]= -2145835515;
assign addr[52125]= -2146993250;
assign addr[52126]= -2147470025;
assign addr[52127]= -2147265689;
assign addr[52128]= -2146380306;
assign addr[52129]= -2144814157;
assign addr[52130]= -2142567738;
assign addr[52131]= -2139641764;
assign addr[52132]= -2136037160;
assign addr[52133]= -2131755071;
assign addr[52134]= -2126796855;
assign addr[52135]= -2121164085;
assign addr[52136]= -2114858546;
assign addr[52137]= -2107882239;
assign addr[52138]= -2100237377;
assign addr[52139]= -2091926384;
assign addr[52140]= -2082951896;
assign addr[52141]= -2073316760;
assign addr[52142]= -2063024031;
assign addr[52143]= -2052076975;
assign addr[52144]= -2040479063;
assign addr[52145]= -2028233973;
assign addr[52146]= -2015345591;
assign addr[52147]= -2001818002;
assign addr[52148]= -1987655498;
assign addr[52149]= -1972862571;
assign addr[52150]= -1957443913;
assign addr[52151]= -1941404413;
assign addr[52152]= -1924749160;
assign addr[52153]= -1907483436;
assign addr[52154]= -1889612716;
assign addr[52155]= -1871142669;
assign addr[52156]= -1852079154;
assign addr[52157]= -1832428215;
assign addr[52158]= -1812196087;
assign addr[52159]= -1791389186;
assign addr[52160]= -1770014111;
assign addr[52161]= -1748077642;
assign addr[52162]= -1725586737;
assign addr[52163]= -1702548529;
assign addr[52164]= -1678970324;
assign addr[52165]= -1654859602;
assign addr[52166]= -1630224009;
assign addr[52167]= -1605071359;
assign addr[52168]= -1579409630;
assign addr[52169]= -1553246960;
assign addr[52170]= -1526591649;
assign addr[52171]= -1499452149;
assign addr[52172]= -1471837070;
assign addr[52173]= -1443755168;
assign addr[52174]= -1415215352;
assign addr[52175]= -1386226674;
assign addr[52176]= -1356798326;
assign addr[52177]= -1326939644;
assign addr[52178]= -1296660098;
assign addr[52179]= -1265969291;
assign addr[52180]= -1234876957;
assign addr[52181]= -1203392958;
assign addr[52182]= -1171527280;
assign addr[52183]= -1139290029;
assign addr[52184]= -1106691431;
assign addr[52185]= -1073741824;
assign addr[52186]= -1040451659;
assign addr[52187]= -1006831495;
assign addr[52188]= -972891995;
assign addr[52189]= -938643924;
assign addr[52190]= -904098143;
assign addr[52191]= -869265610;
assign addr[52192]= -834157373;
assign addr[52193]= -798784567;
assign addr[52194]= -763158411;
assign addr[52195]= -727290205;
assign addr[52196]= -691191324;
assign addr[52197]= -654873219;
assign addr[52198]= -618347408;
assign addr[52199]= -581625477;
assign addr[52200]= -544719071;
assign addr[52201]= -507639898;
assign addr[52202]= -470399716;
assign addr[52203]= -433010339;
assign addr[52204]= -395483624;
assign addr[52205]= -357831473;
assign addr[52206]= -320065829;
assign addr[52207]= -282198671;
assign addr[52208]= -244242007;
assign addr[52209]= -206207878;
assign addr[52210]= -168108346;
assign addr[52211]= -129955495;
assign addr[52212]= -91761426;
assign addr[52213]= -53538253;
assign addr[52214]= -15298099;
assign addr[52215]= 22946906;
assign addr[52216]= 61184634;
assign addr[52217]= 99402956;
assign addr[52218]= 137589750;
assign addr[52219]= 175732905;
assign addr[52220]= 213820322;
assign addr[52221]= 251839923;
assign addr[52222]= 289779648;
assign addr[52223]= 327627463;
assign addr[52224]= 365371365;
assign addr[52225]= 402999383;
assign addr[52226]= 440499581;
assign addr[52227]= 477860067;
assign addr[52228]= 515068990;
assign addr[52229]= 552114549;
assign addr[52230]= 588984994;
assign addr[52231]= 625668632;
assign addr[52232]= 662153826;
assign addr[52233]= 698429006;
assign addr[52234]= 734482665;
assign addr[52235]= 770303369;
assign addr[52236]= 805879757;
assign addr[52237]= 841200544;
assign addr[52238]= 876254528;
assign addr[52239]= 911030591;
assign addr[52240]= 945517704;
assign addr[52241]= 979704927;
assign addr[52242]= 1013581418;
assign addr[52243]= 1047136432;
assign addr[52244]= 1080359326;
assign addr[52245]= 1113239564;
assign addr[52246]= 1145766716;
assign addr[52247]= 1177930466;
assign addr[52248]= 1209720613;
assign addr[52249]= 1241127074;
assign addr[52250]= 1272139887;
assign addr[52251]= 1302749217;
assign addr[52252]= 1332945355;
assign addr[52253]= 1362718723;
assign addr[52254]= 1392059879;
assign addr[52255]= 1420959516;
assign addr[52256]= 1449408469;
assign addr[52257]= 1477397714;
assign addr[52258]= 1504918373;
assign addr[52259]= 1531961719;
assign addr[52260]= 1558519173;
assign addr[52261]= 1584582314;
assign addr[52262]= 1610142873;
assign addr[52263]= 1635192744;
assign addr[52264]= 1659723983;
assign addr[52265]= 1683728808;
assign addr[52266]= 1707199606;
assign addr[52267]= 1730128933;
assign addr[52268]= 1752509516;
assign addr[52269]= 1774334257;
assign addr[52270]= 1795596234;
assign addr[52271]= 1816288703;
assign addr[52272]= 1836405100;
assign addr[52273]= 1855939047;
assign addr[52274]= 1874884346;
assign addr[52275]= 1893234990;
assign addr[52276]= 1910985158;
assign addr[52277]= 1928129220;
assign addr[52278]= 1944661739;
assign addr[52279]= 1960577471;
assign addr[52280]= 1975871368;
assign addr[52281]= 1990538579;
assign addr[52282]= 2004574453;
assign addr[52283]= 2017974537;
assign addr[52284]= 2030734582;
assign addr[52285]= 2042850540;
assign addr[52286]= 2054318569;
assign addr[52287]= 2065135031;
assign addr[52288]= 2075296495;
assign addr[52289]= 2084799740;
assign addr[52290]= 2093641749;
assign addr[52291]= 2101819720;
assign addr[52292]= 2109331059;
assign addr[52293]= 2116173382;
assign addr[52294]= 2122344521;
assign addr[52295]= 2127842516;
assign addr[52296]= 2132665626;
assign addr[52297]= 2136812319;
assign addr[52298]= 2140281282;
assign addr[52299]= 2143071413;
assign addr[52300]= 2145181827;
assign addr[52301]= 2146611856;
assign addr[52302]= 2147361045;
assign addr[52303]= 2147429158;
assign addr[52304]= 2146816171;
assign addr[52305]= 2145522281;
assign addr[52306]= 2143547897;
assign addr[52307]= 2140893646;
assign addr[52308]= 2137560369;
assign addr[52309]= 2133549123;
assign addr[52310]= 2128861181;
assign addr[52311]= 2123498030;
assign addr[52312]= 2117461370;
assign addr[52313]= 2110753117;
assign addr[52314]= 2103375398;
assign addr[52315]= 2095330553;
assign addr[52316]= 2086621133;
assign addr[52317]= 2077249901;
assign addr[52318]= 2067219829;
assign addr[52319]= 2056534099;
assign addr[52320]= 2045196100;
assign addr[52321]= 2033209426;
assign addr[52322]= 2020577882;
assign addr[52323]= 2007305472;
assign addr[52324]= 1993396407;
assign addr[52325]= 1978855097;
assign addr[52326]= 1963686155;
assign addr[52327]= 1947894393;
assign addr[52328]= 1931484818;
assign addr[52329]= 1914462636;
assign addr[52330]= 1896833245;
assign addr[52331]= 1878602237;
assign addr[52332]= 1859775393;
assign addr[52333]= 1840358687;
assign addr[52334]= 1820358275;
assign addr[52335]= 1799780501;
assign addr[52336]= 1778631892;
assign addr[52337]= 1756919156;
assign addr[52338]= 1734649179;
assign addr[52339]= 1711829025;
assign addr[52340]= 1688465931;
assign addr[52341]= 1664567307;
assign addr[52342]= 1640140734;
assign addr[52343]= 1615193959;
assign addr[52344]= 1589734894;
assign addr[52345]= 1563771613;
assign addr[52346]= 1537312353;
assign addr[52347]= 1510365504;
assign addr[52348]= 1482939614;
assign addr[52349]= 1455043381;
assign addr[52350]= 1426685652;
assign addr[52351]= 1397875423;
assign addr[52352]= 1368621831;
assign addr[52353]= 1338934154;
assign addr[52354]= 1308821808;
assign addr[52355]= 1278294345;
assign addr[52356]= 1247361445;
assign addr[52357]= 1216032921;
assign addr[52358]= 1184318708;
assign addr[52359]= 1152228866;
assign addr[52360]= 1119773573;
assign addr[52361]= 1086963121;
assign addr[52362]= 1053807919;
assign addr[52363]= 1020318481;
assign addr[52364]= 986505429;
assign addr[52365]= 952379488;
assign addr[52366]= 917951481;
assign addr[52367]= 883232329;
assign addr[52368]= 848233042;
assign addr[52369]= 812964722;
assign addr[52370]= 777438554;
assign addr[52371]= 741665807;
assign addr[52372]= 705657826;
assign addr[52373]= 669426032;
assign addr[52374]= 632981917;
assign addr[52375]= 596337040;
assign addr[52376]= 559503022;
assign addr[52377]= 522491548;
assign addr[52378]= 485314355;
assign addr[52379]= 447983235;
assign addr[52380]= 410510029;
assign addr[52381]= 372906622;
assign addr[52382]= 335184940;
assign addr[52383]= 297356948;
assign addr[52384]= 259434643;
assign addr[52385]= 221430054;
assign addr[52386]= 183355234;
assign addr[52387]= 145222259;
assign addr[52388]= 107043224;
assign addr[52389]= 68830239;
assign addr[52390]= 30595422;
assign addr[52391]= -7649098;
assign addr[52392]= -45891193;
assign addr[52393]= -84118732;
assign addr[52394]= -122319591;
assign addr[52395]= -160481654;
assign addr[52396]= -198592817;
assign addr[52397]= -236640993;
assign addr[52398]= -274614114;
assign addr[52399]= -312500135;
assign addr[52400]= -350287041;
assign addr[52401]= -387962847;
assign addr[52402]= -425515602;
assign addr[52403]= -462933398;
assign addr[52404]= -500204365;
assign addr[52405]= -537316682;
assign addr[52406]= -574258580;
assign addr[52407]= -611018340;
assign addr[52408]= -647584304;
assign addr[52409]= -683944874;
assign addr[52410]= -720088517;
assign addr[52411]= -756003771;
assign addr[52412]= -791679244;
assign addr[52413]= -827103620;
assign addr[52414]= -862265664;
assign addr[52415]= -897154224;
assign addr[52416]= -931758235;
assign addr[52417]= -966066720;
assign addr[52418]= -1000068799;
assign addr[52419]= -1033753687;
assign addr[52420]= -1067110699;
assign addr[52421]= -1100129257;
assign addr[52422]= -1132798888;
assign addr[52423]= -1165109230;
assign addr[52424]= -1197050035;
assign addr[52425]= -1228611172;
assign addr[52426]= -1259782632;
assign addr[52427]= -1290554528;
assign addr[52428]= -1320917099;
assign addr[52429]= -1350860716;
assign addr[52430]= -1380375881;
assign addr[52431]= -1409453233;
assign addr[52432]= -1438083551;
assign addr[52433]= -1466257752;
assign addr[52434]= -1493966902;
assign addr[52435]= -1521202211;
assign addr[52436]= -1547955041;
assign addr[52437]= -1574216908;
assign addr[52438]= -1599979481;
assign addr[52439]= -1625234591;
assign addr[52440]= -1649974225;
assign addr[52441]= -1674190539;
assign addr[52442]= -1697875851;
assign addr[52443]= -1721022648;
assign addr[52444]= -1743623590;
assign addr[52445]= -1765671509;
assign addr[52446]= -1787159411;
assign addr[52447]= -1808080480;
assign addr[52448]= -1828428082;
assign addr[52449]= -1848195763;
assign addr[52450]= -1867377253;
assign addr[52451]= -1885966468;
assign addr[52452]= -1903957513;
assign addr[52453]= -1921344681;
assign addr[52454]= -1938122457;
assign addr[52455]= -1954285520;
assign addr[52456]= -1969828744;
assign addr[52457]= -1984747199;
assign addr[52458]= -1999036154;
assign addr[52459]= -2012691075;
assign addr[52460]= -2025707632;
assign addr[52461]= -2038081698;
assign addr[52462]= -2049809346;
assign addr[52463]= -2060886858;
assign addr[52464]= -2071310720;
assign addr[52465]= -2081077626;
assign addr[52466]= -2090184478;
assign addr[52467]= -2098628387;
assign addr[52468]= -2106406677;
assign addr[52469]= -2113516878;
assign addr[52470]= -2119956737;
assign addr[52471]= -2125724211;
assign addr[52472]= -2130817471;
assign addr[52473]= -2135234901;
assign addr[52474]= -2138975100;
assign addr[52475]= -2142036881;
assign addr[52476]= -2144419275;
assign addr[52477]= -2146121524;
assign addr[52478]= -2147143090;
assign addr[52479]= -2147483648;
assign addr[52480]= -2147143090;
assign addr[52481]= -2146121524;
assign addr[52482]= -2144419275;
assign addr[52483]= -2142036881;
assign addr[52484]= -2138975100;
assign addr[52485]= -2135234901;
assign addr[52486]= -2130817471;
assign addr[52487]= -2125724211;
assign addr[52488]= -2119956737;
assign addr[52489]= -2113516878;
assign addr[52490]= -2106406677;
assign addr[52491]= -2098628387;
assign addr[52492]= -2090184478;
assign addr[52493]= -2081077626;
assign addr[52494]= -2071310720;
assign addr[52495]= -2060886858;
assign addr[52496]= -2049809346;
assign addr[52497]= -2038081698;
assign addr[52498]= -2025707632;
assign addr[52499]= -2012691075;
assign addr[52500]= -1999036154;
assign addr[52501]= -1984747199;
assign addr[52502]= -1969828744;
assign addr[52503]= -1954285520;
assign addr[52504]= -1938122457;
assign addr[52505]= -1921344681;
assign addr[52506]= -1903957513;
assign addr[52507]= -1885966468;
assign addr[52508]= -1867377253;
assign addr[52509]= -1848195763;
assign addr[52510]= -1828428082;
assign addr[52511]= -1808080480;
assign addr[52512]= -1787159411;
assign addr[52513]= -1765671509;
assign addr[52514]= -1743623590;
assign addr[52515]= -1721022648;
assign addr[52516]= -1697875851;
assign addr[52517]= -1674190539;
assign addr[52518]= -1649974225;
assign addr[52519]= -1625234591;
assign addr[52520]= -1599979481;
assign addr[52521]= -1574216908;
assign addr[52522]= -1547955041;
assign addr[52523]= -1521202211;
assign addr[52524]= -1493966902;
assign addr[52525]= -1466257752;
assign addr[52526]= -1438083551;
assign addr[52527]= -1409453233;
assign addr[52528]= -1380375881;
assign addr[52529]= -1350860716;
assign addr[52530]= -1320917099;
assign addr[52531]= -1290554528;
assign addr[52532]= -1259782632;
assign addr[52533]= -1228611172;
assign addr[52534]= -1197050035;
assign addr[52535]= -1165109230;
assign addr[52536]= -1132798888;
assign addr[52537]= -1100129257;
assign addr[52538]= -1067110699;
assign addr[52539]= -1033753687;
assign addr[52540]= -1000068799;
assign addr[52541]= -966066720;
assign addr[52542]= -931758235;
assign addr[52543]= -897154224;
assign addr[52544]= -862265664;
assign addr[52545]= -827103620;
assign addr[52546]= -791679244;
assign addr[52547]= -756003771;
assign addr[52548]= -720088517;
assign addr[52549]= -683944874;
assign addr[52550]= -647584304;
assign addr[52551]= -611018340;
assign addr[52552]= -574258580;
assign addr[52553]= -537316682;
assign addr[52554]= -500204365;
assign addr[52555]= -462933398;
assign addr[52556]= -425515602;
assign addr[52557]= -387962847;
assign addr[52558]= -350287041;
assign addr[52559]= -312500135;
assign addr[52560]= -274614114;
assign addr[52561]= -236640993;
assign addr[52562]= -198592817;
assign addr[52563]= -160481654;
assign addr[52564]= -122319591;
assign addr[52565]= -84118732;
assign addr[52566]= -45891193;
assign addr[52567]= -7649098;
assign addr[52568]= 30595422;
assign addr[52569]= 68830239;
assign addr[52570]= 107043224;
assign addr[52571]= 145222259;
assign addr[52572]= 183355234;
assign addr[52573]= 221430054;
assign addr[52574]= 259434643;
assign addr[52575]= 297356948;
assign addr[52576]= 335184940;
assign addr[52577]= 372906622;
assign addr[52578]= 410510029;
assign addr[52579]= 447983235;
assign addr[52580]= 485314355;
assign addr[52581]= 522491548;
assign addr[52582]= 559503022;
assign addr[52583]= 596337040;
assign addr[52584]= 632981917;
assign addr[52585]= 669426032;
assign addr[52586]= 705657826;
assign addr[52587]= 741665807;
assign addr[52588]= 777438554;
assign addr[52589]= 812964722;
assign addr[52590]= 848233042;
assign addr[52591]= 883232329;
assign addr[52592]= 917951481;
assign addr[52593]= 952379488;
assign addr[52594]= 986505429;
assign addr[52595]= 1020318481;
assign addr[52596]= 1053807919;
assign addr[52597]= 1086963121;
assign addr[52598]= 1119773573;
assign addr[52599]= 1152228866;
assign addr[52600]= 1184318708;
assign addr[52601]= 1216032921;
assign addr[52602]= 1247361445;
assign addr[52603]= 1278294345;
assign addr[52604]= 1308821808;
assign addr[52605]= 1338934154;
assign addr[52606]= 1368621831;
assign addr[52607]= 1397875423;
assign addr[52608]= 1426685652;
assign addr[52609]= 1455043381;
assign addr[52610]= 1482939614;
assign addr[52611]= 1510365504;
assign addr[52612]= 1537312353;
assign addr[52613]= 1563771613;
assign addr[52614]= 1589734894;
assign addr[52615]= 1615193959;
assign addr[52616]= 1640140734;
assign addr[52617]= 1664567307;
assign addr[52618]= 1688465931;
assign addr[52619]= 1711829025;
assign addr[52620]= 1734649179;
assign addr[52621]= 1756919156;
assign addr[52622]= 1778631892;
assign addr[52623]= 1799780501;
assign addr[52624]= 1820358275;
assign addr[52625]= 1840358687;
assign addr[52626]= 1859775393;
assign addr[52627]= 1878602237;
assign addr[52628]= 1896833245;
assign addr[52629]= 1914462636;
assign addr[52630]= 1931484818;
assign addr[52631]= 1947894393;
assign addr[52632]= 1963686155;
assign addr[52633]= 1978855097;
assign addr[52634]= 1993396407;
assign addr[52635]= 2007305472;
assign addr[52636]= 2020577882;
assign addr[52637]= 2033209426;
assign addr[52638]= 2045196100;
assign addr[52639]= 2056534099;
assign addr[52640]= 2067219829;
assign addr[52641]= 2077249901;
assign addr[52642]= 2086621133;
assign addr[52643]= 2095330553;
assign addr[52644]= 2103375398;
assign addr[52645]= 2110753117;
assign addr[52646]= 2117461370;
assign addr[52647]= 2123498030;
assign addr[52648]= 2128861181;
assign addr[52649]= 2133549123;
assign addr[52650]= 2137560369;
assign addr[52651]= 2140893646;
assign addr[52652]= 2143547897;
assign addr[52653]= 2145522281;
assign addr[52654]= 2146816171;
assign addr[52655]= 2147429158;
assign addr[52656]= 2147361045;
assign addr[52657]= 2146611856;
assign addr[52658]= 2145181827;
assign addr[52659]= 2143071413;
assign addr[52660]= 2140281282;
assign addr[52661]= 2136812319;
assign addr[52662]= 2132665626;
assign addr[52663]= 2127842516;
assign addr[52664]= 2122344521;
assign addr[52665]= 2116173382;
assign addr[52666]= 2109331059;
assign addr[52667]= 2101819720;
assign addr[52668]= 2093641749;
assign addr[52669]= 2084799740;
assign addr[52670]= 2075296495;
assign addr[52671]= 2065135031;
assign addr[52672]= 2054318569;
assign addr[52673]= 2042850540;
assign addr[52674]= 2030734582;
assign addr[52675]= 2017974537;
assign addr[52676]= 2004574453;
assign addr[52677]= 1990538579;
assign addr[52678]= 1975871368;
assign addr[52679]= 1960577471;
assign addr[52680]= 1944661739;
assign addr[52681]= 1928129220;
assign addr[52682]= 1910985158;
assign addr[52683]= 1893234990;
assign addr[52684]= 1874884346;
assign addr[52685]= 1855939047;
assign addr[52686]= 1836405100;
assign addr[52687]= 1816288703;
assign addr[52688]= 1795596234;
assign addr[52689]= 1774334257;
assign addr[52690]= 1752509516;
assign addr[52691]= 1730128933;
assign addr[52692]= 1707199606;
assign addr[52693]= 1683728808;
assign addr[52694]= 1659723983;
assign addr[52695]= 1635192744;
assign addr[52696]= 1610142873;
assign addr[52697]= 1584582314;
assign addr[52698]= 1558519173;
assign addr[52699]= 1531961719;
assign addr[52700]= 1504918373;
assign addr[52701]= 1477397714;
assign addr[52702]= 1449408469;
assign addr[52703]= 1420959516;
assign addr[52704]= 1392059879;
assign addr[52705]= 1362718723;
assign addr[52706]= 1332945355;
assign addr[52707]= 1302749217;
assign addr[52708]= 1272139887;
assign addr[52709]= 1241127074;
assign addr[52710]= 1209720613;
assign addr[52711]= 1177930466;
assign addr[52712]= 1145766716;
assign addr[52713]= 1113239564;
assign addr[52714]= 1080359326;
assign addr[52715]= 1047136432;
assign addr[52716]= 1013581418;
assign addr[52717]= 979704927;
assign addr[52718]= 945517704;
assign addr[52719]= 911030591;
assign addr[52720]= 876254528;
assign addr[52721]= 841200544;
assign addr[52722]= 805879757;
assign addr[52723]= 770303369;
assign addr[52724]= 734482665;
assign addr[52725]= 698429006;
assign addr[52726]= 662153826;
assign addr[52727]= 625668632;
assign addr[52728]= 588984994;
assign addr[52729]= 552114549;
assign addr[52730]= 515068990;
assign addr[52731]= 477860067;
assign addr[52732]= 440499581;
assign addr[52733]= 402999383;
assign addr[52734]= 365371365;
assign addr[52735]= 327627463;
assign addr[52736]= 289779648;
assign addr[52737]= 251839923;
assign addr[52738]= 213820322;
assign addr[52739]= 175732905;
assign addr[52740]= 137589750;
assign addr[52741]= 99402956;
assign addr[52742]= 61184634;
assign addr[52743]= 22946906;
assign addr[52744]= -15298099;
assign addr[52745]= -53538253;
assign addr[52746]= -91761426;
assign addr[52747]= -129955495;
assign addr[52748]= -168108346;
assign addr[52749]= -206207878;
assign addr[52750]= -244242007;
assign addr[52751]= -282198671;
assign addr[52752]= -320065829;
assign addr[52753]= -357831473;
assign addr[52754]= -395483624;
assign addr[52755]= -433010339;
assign addr[52756]= -470399716;
assign addr[52757]= -507639898;
assign addr[52758]= -544719071;
assign addr[52759]= -581625477;
assign addr[52760]= -618347408;
assign addr[52761]= -654873219;
assign addr[52762]= -691191324;
assign addr[52763]= -727290205;
assign addr[52764]= -763158411;
assign addr[52765]= -798784567;
assign addr[52766]= -834157373;
assign addr[52767]= -869265610;
assign addr[52768]= -904098143;
assign addr[52769]= -938643924;
assign addr[52770]= -972891995;
assign addr[52771]= -1006831495;
assign addr[52772]= -1040451659;
assign addr[52773]= -1073741824;
assign addr[52774]= -1106691431;
assign addr[52775]= -1139290029;
assign addr[52776]= -1171527280;
assign addr[52777]= -1203392958;
assign addr[52778]= -1234876957;
assign addr[52779]= -1265969291;
assign addr[52780]= -1296660098;
assign addr[52781]= -1326939644;
assign addr[52782]= -1356798326;
assign addr[52783]= -1386226674;
assign addr[52784]= -1415215352;
assign addr[52785]= -1443755168;
assign addr[52786]= -1471837070;
assign addr[52787]= -1499452149;
assign addr[52788]= -1526591649;
assign addr[52789]= -1553246960;
assign addr[52790]= -1579409630;
assign addr[52791]= -1605071359;
assign addr[52792]= -1630224009;
assign addr[52793]= -1654859602;
assign addr[52794]= -1678970324;
assign addr[52795]= -1702548529;
assign addr[52796]= -1725586737;
assign addr[52797]= -1748077642;
assign addr[52798]= -1770014111;
assign addr[52799]= -1791389186;
assign addr[52800]= -1812196087;
assign addr[52801]= -1832428215;
assign addr[52802]= -1852079154;
assign addr[52803]= -1871142669;
assign addr[52804]= -1889612716;
assign addr[52805]= -1907483436;
assign addr[52806]= -1924749160;
assign addr[52807]= -1941404413;
assign addr[52808]= -1957443913;
assign addr[52809]= -1972862571;
assign addr[52810]= -1987655498;
assign addr[52811]= -2001818002;
assign addr[52812]= -2015345591;
assign addr[52813]= -2028233973;
assign addr[52814]= -2040479063;
assign addr[52815]= -2052076975;
assign addr[52816]= -2063024031;
assign addr[52817]= -2073316760;
assign addr[52818]= -2082951896;
assign addr[52819]= -2091926384;
assign addr[52820]= -2100237377;
assign addr[52821]= -2107882239;
assign addr[52822]= -2114858546;
assign addr[52823]= -2121164085;
assign addr[52824]= -2126796855;
assign addr[52825]= -2131755071;
assign addr[52826]= -2136037160;
assign addr[52827]= -2139641764;
assign addr[52828]= -2142567738;
assign addr[52829]= -2144814157;
assign addr[52830]= -2146380306;
assign addr[52831]= -2147265689;
assign addr[52832]= -2147470025;
assign addr[52833]= -2146993250;
assign addr[52834]= -2145835515;
assign addr[52835]= -2143997187;
assign addr[52836]= -2141478848;
assign addr[52837]= -2138281298;
assign addr[52838]= -2134405552;
assign addr[52839]= -2129852837;
assign addr[52840]= -2124624598;
assign addr[52841]= -2118722494;
assign addr[52842]= -2112148396;
assign addr[52843]= -2104904390;
assign addr[52844]= -2096992772;
assign addr[52845]= -2088416053;
assign addr[52846]= -2079176953;
assign addr[52847]= -2069278401;
assign addr[52848]= -2058723538;
assign addr[52849]= -2047515711;
assign addr[52850]= -2035658475;
assign addr[52851]= -2023155591;
assign addr[52852]= -2010011024;
assign addr[52853]= -1996228943;
assign addr[52854]= -1981813720;
assign addr[52855]= -1966769926;
assign addr[52856]= -1951102334;
assign addr[52857]= -1934815911;
assign addr[52858]= -1917915825;
assign addr[52859]= -1900407434;
assign addr[52860]= -1882296293;
assign addr[52861]= -1863588145;
assign addr[52862]= -1844288924;
assign addr[52863]= -1824404752;
assign addr[52864]= -1803941934;
assign addr[52865]= -1782906961;
assign addr[52866]= -1761306505;
assign addr[52867]= -1739147417;
assign addr[52868]= -1716436725;
assign addr[52869]= -1693181631;
assign addr[52870]= -1669389513;
assign addr[52871]= -1645067915;
assign addr[52872]= -1620224553;
assign addr[52873]= -1594867305;
assign addr[52874]= -1569004214;
assign addr[52875]= -1542643483;
assign addr[52876]= -1515793473;
assign addr[52877]= -1488462700;
assign addr[52878]= -1460659832;
assign addr[52879]= -1432393688;
assign addr[52880]= -1403673233;
assign addr[52881]= -1374507575;
assign addr[52882]= -1344905966;
assign addr[52883]= -1314877795;
assign addr[52884]= -1284432584;
assign addr[52885]= -1253579991;
assign addr[52886]= -1222329801;
assign addr[52887]= -1190691925;
assign addr[52888]= -1158676398;
assign addr[52889]= -1126293375;
assign addr[52890]= -1093553126;
assign addr[52891]= -1060466036;
assign addr[52892]= -1027042599;
assign addr[52893]= -993293415;
assign addr[52894]= -959229189;
assign addr[52895]= -924860725;
assign addr[52896]= -890198924;
assign addr[52897]= -855254778;
assign addr[52898]= -820039373;
assign addr[52899]= -784563876;
assign addr[52900]= -748839539;
assign addr[52901]= -712877694;
assign addr[52902]= -676689746;
assign addr[52903]= -640287172;
assign addr[52904]= -603681519;
assign addr[52905]= -566884397;
assign addr[52906]= -529907477;
assign addr[52907]= -492762486;
assign addr[52908]= -455461206;
assign addr[52909]= -418015468;
assign addr[52910]= -380437148;
assign addr[52911]= -342738165;
assign addr[52912]= -304930476;
assign addr[52913]= -267026072;
assign addr[52914]= -229036977;
assign addr[52915]= -190975237;
assign addr[52916]= -152852926;
assign addr[52917]= -114682135;
assign addr[52918]= -76474970;
assign addr[52919]= -38243550;
assign addr[52920]= 0;
assign addr[52921]= 38243550;
assign addr[52922]= 76474970;
assign addr[52923]= 114682135;
assign addr[52924]= 152852926;
assign addr[52925]= 190975237;
assign addr[52926]= 229036977;
assign addr[52927]= 267026072;
assign addr[52928]= 304930476;
assign addr[52929]= 342738165;
assign addr[52930]= 380437148;
assign addr[52931]= 418015468;
assign addr[52932]= 455461206;
assign addr[52933]= 492762486;
assign addr[52934]= 529907477;
assign addr[52935]= 566884397;
assign addr[52936]= 603681519;
assign addr[52937]= 640287172;
assign addr[52938]= 676689746;
assign addr[52939]= 712877694;
assign addr[52940]= 748839539;
assign addr[52941]= 784563876;
assign addr[52942]= 820039373;
assign addr[52943]= 855254778;
assign addr[52944]= 890198924;
assign addr[52945]= 924860725;
assign addr[52946]= 959229189;
assign addr[52947]= 993293415;
assign addr[52948]= 1027042599;
assign addr[52949]= 1060466036;
assign addr[52950]= 1093553126;
assign addr[52951]= 1126293375;
assign addr[52952]= 1158676398;
assign addr[52953]= 1190691925;
assign addr[52954]= 1222329801;
assign addr[52955]= 1253579991;
assign addr[52956]= 1284432584;
assign addr[52957]= 1314877795;
assign addr[52958]= 1344905966;
assign addr[52959]= 1374507575;
assign addr[52960]= 1403673233;
assign addr[52961]= 1432393688;
assign addr[52962]= 1460659832;
assign addr[52963]= 1488462700;
assign addr[52964]= 1515793473;
assign addr[52965]= 1542643483;
assign addr[52966]= 1569004214;
assign addr[52967]= 1594867305;
assign addr[52968]= 1620224553;
assign addr[52969]= 1645067915;
assign addr[52970]= 1669389513;
assign addr[52971]= 1693181631;
assign addr[52972]= 1716436725;
assign addr[52973]= 1739147417;
assign addr[52974]= 1761306505;
assign addr[52975]= 1782906961;
assign addr[52976]= 1803941934;
assign addr[52977]= 1824404752;
assign addr[52978]= 1844288924;
assign addr[52979]= 1863588145;
assign addr[52980]= 1882296293;
assign addr[52981]= 1900407434;
assign addr[52982]= 1917915825;
assign addr[52983]= 1934815911;
assign addr[52984]= 1951102334;
assign addr[52985]= 1966769926;
assign addr[52986]= 1981813720;
assign addr[52987]= 1996228943;
assign addr[52988]= 2010011024;
assign addr[52989]= 2023155591;
assign addr[52990]= 2035658475;
assign addr[52991]= 2047515711;
assign addr[52992]= 2058723538;
assign addr[52993]= 2069278401;
assign addr[52994]= 2079176953;
assign addr[52995]= 2088416053;
assign addr[52996]= 2096992772;
assign addr[52997]= 2104904390;
assign addr[52998]= 2112148396;
assign addr[52999]= 2118722494;
assign addr[53000]= 2124624598;
assign addr[53001]= 2129852837;
assign addr[53002]= 2134405552;
assign addr[53003]= 2138281298;
assign addr[53004]= 2141478848;
assign addr[53005]= 2143997187;
assign addr[53006]= 2145835515;
assign addr[53007]= 2146993250;
assign addr[53008]= 2147470025;
assign addr[53009]= 2147265689;
assign addr[53010]= 2146380306;
assign addr[53011]= 2144814157;
assign addr[53012]= 2142567738;
assign addr[53013]= 2139641764;
assign addr[53014]= 2136037160;
assign addr[53015]= 2131755071;
assign addr[53016]= 2126796855;
assign addr[53017]= 2121164085;
assign addr[53018]= 2114858546;
assign addr[53019]= 2107882239;
assign addr[53020]= 2100237377;
assign addr[53021]= 2091926384;
assign addr[53022]= 2082951896;
assign addr[53023]= 2073316760;
assign addr[53024]= 2063024031;
assign addr[53025]= 2052076975;
assign addr[53026]= 2040479063;
assign addr[53027]= 2028233973;
assign addr[53028]= 2015345591;
assign addr[53029]= 2001818002;
assign addr[53030]= 1987655498;
assign addr[53031]= 1972862571;
assign addr[53032]= 1957443913;
assign addr[53033]= 1941404413;
assign addr[53034]= 1924749160;
assign addr[53035]= 1907483436;
assign addr[53036]= 1889612716;
assign addr[53037]= 1871142669;
assign addr[53038]= 1852079154;
assign addr[53039]= 1832428215;
assign addr[53040]= 1812196087;
assign addr[53041]= 1791389186;
assign addr[53042]= 1770014111;
assign addr[53043]= 1748077642;
assign addr[53044]= 1725586737;
assign addr[53045]= 1702548529;
assign addr[53046]= 1678970324;
assign addr[53047]= 1654859602;
assign addr[53048]= 1630224009;
assign addr[53049]= 1605071359;
assign addr[53050]= 1579409630;
assign addr[53051]= 1553246960;
assign addr[53052]= 1526591649;
assign addr[53053]= 1499452149;
assign addr[53054]= 1471837070;
assign addr[53055]= 1443755168;
assign addr[53056]= 1415215352;
assign addr[53057]= 1386226674;
assign addr[53058]= 1356798326;
assign addr[53059]= 1326939644;
assign addr[53060]= 1296660098;
assign addr[53061]= 1265969291;
assign addr[53062]= 1234876957;
assign addr[53063]= 1203392958;
assign addr[53064]= 1171527280;
assign addr[53065]= 1139290029;
assign addr[53066]= 1106691431;
assign addr[53067]= 1073741824;
assign addr[53068]= 1040451659;
assign addr[53069]= 1006831495;
assign addr[53070]= 972891995;
assign addr[53071]= 938643924;
assign addr[53072]= 904098143;
assign addr[53073]= 869265610;
assign addr[53074]= 834157373;
assign addr[53075]= 798784567;
assign addr[53076]= 763158411;
assign addr[53077]= 727290205;
assign addr[53078]= 691191324;
assign addr[53079]= 654873219;
assign addr[53080]= 618347408;
assign addr[53081]= 581625477;
assign addr[53082]= 544719071;
assign addr[53083]= 507639898;
assign addr[53084]= 470399716;
assign addr[53085]= 433010339;
assign addr[53086]= 395483624;
assign addr[53087]= 357831473;
assign addr[53088]= 320065829;
assign addr[53089]= 282198671;
assign addr[53090]= 244242007;
assign addr[53091]= 206207878;
assign addr[53092]= 168108346;
assign addr[53093]= 129955495;
assign addr[53094]= 91761426;
assign addr[53095]= 53538253;
assign addr[53096]= 15298099;
assign addr[53097]= -22946906;
assign addr[53098]= -61184634;
assign addr[53099]= -99402956;
assign addr[53100]= -137589750;
assign addr[53101]= -175732905;
assign addr[53102]= -213820322;
assign addr[53103]= -251839923;
assign addr[53104]= -289779648;
assign addr[53105]= -327627463;
assign addr[53106]= -365371365;
assign addr[53107]= -402999383;
assign addr[53108]= -440499581;
assign addr[53109]= -477860067;
assign addr[53110]= -515068990;
assign addr[53111]= -552114549;
assign addr[53112]= -588984994;
assign addr[53113]= -625668632;
assign addr[53114]= -662153826;
assign addr[53115]= -698429006;
assign addr[53116]= -734482665;
assign addr[53117]= -770303369;
assign addr[53118]= -805879757;
assign addr[53119]= -841200544;
assign addr[53120]= -876254528;
assign addr[53121]= -911030591;
assign addr[53122]= -945517704;
assign addr[53123]= -979704927;
assign addr[53124]= -1013581418;
assign addr[53125]= -1047136432;
assign addr[53126]= -1080359326;
assign addr[53127]= -1113239564;
assign addr[53128]= -1145766716;
assign addr[53129]= -1177930466;
assign addr[53130]= -1209720613;
assign addr[53131]= -1241127074;
assign addr[53132]= -1272139887;
assign addr[53133]= -1302749217;
assign addr[53134]= -1332945355;
assign addr[53135]= -1362718723;
assign addr[53136]= -1392059879;
assign addr[53137]= -1420959516;
assign addr[53138]= -1449408469;
assign addr[53139]= -1477397714;
assign addr[53140]= -1504918373;
assign addr[53141]= -1531961719;
assign addr[53142]= -1558519173;
assign addr[53143]= -1584582314;
assign addr[53144]= -1610142873;
assign addr[53145]= -1635192744;
assign addr[53146]= -1659723983;
assign addr[53147]= -1683728808;
assign addr[53148]= -1707199606;
assign addr[53149]= -1730128933;
assign addr[53150]= -1752509516;
assign addr[53151]= -1774334257;
assign addr[53152]= -1795596234;
assign addr[53153]= -1816288703;
assign addr[53154]= -1836405100;
assign addr[53155]= -1855939047;
assign addr[53156]= -1874884346;
assign addr[53157]= -1893234990;
assign addr[53158]= -1910985158;
assign addr[53159]= -1928129220;
assign addr[53160]= -1944661739;
assign addr[53161]= -1960577471;
assign addr[53162]= -1975871368;
assign addr[53163]= -1990538579;
assign addr[53164]= -2004574453;
assign addr[53165]= -2017974537;
assign addr[53166]= -2030734582;
assign addr[53167]= -2042850540;
assign addr[53168]= -2054318569;
assign addr[53169]= -2065135031;
assign addr[53170]= -2075296495;
assign addr[53171]= -2084799740;
assign addr[53172]= -2093641749;
assign addr[53173]= -2101819720;
assign addr[53174]= -2109331059;
assign addr[53175]= -2116173382;
assign addr[53176]= -2122344521;
assign addr[53177]= -2127842516;
assign addr[53178]= -2132665626;
assign addr[53179]= -2136812319;
assign addr[53180]= -2140281282;
assign addr[53181]= -2143071413;
assign addr[53182]= -2145181827;
assign addr[53183]= -2146611856;
assign addr[53184]= -2147361045;
assign addr[53185]= -2147429158;
assign addr[53186]= -2146816171;
assign addr[53187]= -2145522281;
assign addr[53188]= -2143547897;
assign addr[53189]= -2140893646;
assign addr[53190]= -2137560369;
assign addr[53191]= -2133549123;
assign addr[53192]= -2128861181;
assign addr[53193]= -2123498030;
assign addr[53194]= -2117461370;
assign addr[53195]= -2110753117;
assign addr[53196]= -2103375398;
assign addr[53197]= -2095330553;
assign addr[53198]= -2086621133;
assign addr[53199]= -2077249901;
assign addr[53200]= -2067219829;
assign addr[53201]= -2056534099;
assign addr[53202]= -2045196100;
assign addr[53203]= -2033209426;
assign addr[53204]= -2020577882;
assign addr[53205]= -2007305472;
assign addr[53206]= -1993396407;
assign addr[53207]= -1978855097;
assign addr[53208]= -1963686155;
assign addr[53209]= -1947894393;
assign addr[53210]= -1931484818;
assign addr[53211]= -1914462636;
assign addr[53212]= -1896833245;
assign addr[53213]= -1878602237;
assign addr[53214]= -1859775393;
assign addr[53215]= -1840358687;
assign addr[53216]= -1820358275;
assign addr[53217]= -1799780501;
assign addr[53218]= -1778631892;
assign addr[53219]= -1756919156;
assign addr[53220]= -1734649179;
assign addr[53221]= -1711829025;
assign addr[53222]= -1688465931;
assign addr[53223]= -1664567307;
assign addr[53224]= -1640140734;
assign addr[53225]= -1615193959;
assign addr[53226]= -1589734894;
assign addr[53227]= -1563771613;
assign addr[53228]= -1537312353;
assign addr[53229]= -1510365504;
assign addr[53230]= -1482939614;
assign addr[53231]= -1455043381;
assign addr[53232]= -1426685652;
assign addr[53233]= -1397875423;
assign addr[53234]= -1368621831;
assign addr[53235]= -1338934154;
assign addr[53236]= -1308821808;
assign addr[53237]= -1278294345;
assign addr[53238]= -1247361445;
assign addr[53239]= -1216032921;
assign addr[53240]= -1184318708;
assign addr[53241]= -1152228866;
assign addr[53242]= -1119773573;
assign addr[53243]= -1086963121;
assign addr[53244]= -1053807919;
assign addr[53245]= -1020318481;
assign addr[53246]= -986505429;
assign addr[53247]= -952379488;
assign addr[53248]= -917951481;
assign addr[53249]= -883232329;
assign addr[53250]= -848233042;
assign addr[53251]= -812964722;
assign addr[53252]= -777438554;
assign addr[53253]= -741665807;
assign addr[53254]= -705657826;
assign addr[53255]= -669426032;
assign addr[53256]= -632981917;
assign addr[53257]= -596337040;
assign addr[53258]= -559503022;
assign addr[53259]= -522491548;
assign addr[53260]= -485314355;
assign addr[53261]= -447983235;
assign addr[53262]= -410510029;
assign addr[53263]= -372906622;
assign addr[53264]= -335184940;
assign addr[53265]= -297356948;
assign addr[53266]= -259434643;
assign addr[53267]= -221430054;
assign addr[53268]= -183355234;
assign addr[53269]= -145222259;
assign addr[53270]= -107043224;
assign addr[53271]= -68830239;
assign addr[53272]= -30595422;
assign addr[53273]= 7649098;
assign addr[53274]= 45891193;
assign addr[53275]= 84118732;
assign addr[53276]= 122319591;
assign addr[53277]= 160481654;
assign addr[53278]= 198592817;
assign addr[53279]= 236640993;
assign addr[53280]= 274614114;
assign addr[53281]= 312500135;
assign addr[53282]= 350287041;
assign addr[53283]= 387962847;
assign addr[53284]= 425515602;
assign addr[53285]= 462933398;
assign addr[53286]= 500204365;
assign addr[53287]= 537316682;
assign addr[53288]= 574258580;
assign addr[53289]= 611018340;
assign addr[53290]= 647584304;
assign addr[53291]= 683944874;
assign addr[53292]= 720088517;
assign addr[53293]= 756003771;
assign addr[53294]= 791679244;
assign addr[53295]= 827103620;
assign addr[53296]= 862265664;
assign addr[53297]= 897154224;
assign addr[53298]= 931758235;
assign addr[53299]= 966066720;
assign addr[53300]= 1000068799;
assign addr[53301]= 1033753687;
assign addr[53302]= 1067110699;
assign addr[53303]= 1100129257;
assign addr[53304]= 1132798888;
assign addr[53305]= 1165109230;
assign addr[53306]= 1197050035;
assign addr[53307]= 1228611172;
assign addr[53308]= 1259782632;
assign addr[53309]= 1290554528;
assign addr[53310]= 1320917099;
assign addr[53311]= 1350860716;
assign addr[53312]= 1380375881;
assign addr[53313]= 1409453233;
assign addr[53314]= 1438083551;
assign addr[53315]= 1466257752;
assign addr[53316]= 1493966902;
assign addr[53317]= 1521202211;
assign addr[53318]= 1547955041;
assign addr[53319]= 1574216908;
assign addr[53320]= 1599979481;
assign addr[53321]= 1625234591;
assign addr[53322]= 1649974225;
assign addr[53323]= 1674190539;
assign addr[53324]= 1697875851;
assign addr[53325]= 1721022648;
assign addr[53326]= 1743623590;
assign addr[53327]= 1765671509;
assign addr[53328]= 1787159411;
assign addr[53329]= 1808080480;
assign addr[53330]= 1828428082;
assign addr[53331]= 1848195763;
assign addr[53332]= 1867377253;
assign addr[53333]= 1885966468;
assign addr[53334]= 1903957513;
assign addr[53335]= 1921344681;
assign addr[53336]= 1938122457;
assign addr[53337]= 1954285520;
assign addr[53338]= 1969828744;
assign addr[53339]= 1984747199;
assign addr[53340]= 1999036154;
assign addr[53341]= 2012691075;
assign addr[53342]= 2025707632;
assign addr[53343]= 2038081698;
assign addr[53344]= 2049809346;
assign addr[53345]= 2060886858;
assign addr[53346]= 2071310720;
assign addr[53347]= 2081077626;
assign addr[53348]= 2090184478;
assign addr[53349]= 2098628387;
assign addr[53350]= 2106406677;
assign addr[53351]= 2113516878;
assign addr[53352]= 2119956737;
assign addr[53353]= 2125724211;
assign addr[53354]= 2130817471;
assign addr[53355]= 2135234901;
assign addr[53356]= 2138975100;
assign addr[53357]= 2142036881;
assign addr[53358]= 2144419275;
assign addr[53359]= 2146121524;
assign addr[53360]= 2147143090;
assign addr[53361]= 2147483648;
assign addr[53362]= 2147143090;
assign addr[53363]= 2146121524;
assign addr[53364]= 2144419275;
assign addr[53365]= 2142036881;
assign addr[53366]= 2138975100;
assign addr[53367]= 2135234901;
assign addr[53368]= 2130817471;
assign addr[53369]= 2125724211;
assign addr[53370]= 2119956737;
assign addr[53371]= 2113516878;
assign addr[53372]= 2106406677;
assign addr[53373]= 2098628387;
assign addr[53374]= 2090184478;
assign addr[53375]= 2081077626;
assign addr[53376]= 2071310720;
assign addr[53377]= 2060886858;
assign addr[53378]= 2049809346;
assign addr[53379]= 2038081698;
assign addr[53380]= 2025707632;
assign addr[53381]= 2012691075;
assign addr[53382]= 1999036154;
assign addr[53383]= 1984747199;
assign addr[53384]= 1969828744;
assign addr[53385]= 1954285520;
assign addr[53386]= 1938122457;
assign addr[53387]= 1921344681;
assign addr[53388]= 1903957513;
assign addr[53389]= 1885966468;
assign addr[53390]= 1867377253;
assign addr[53391]= 1848195763;
assign addr[53392]= 1828428082;
assign addr[53393]= 1808080480;
assign addr[53394]= 1787159411;
assign addr[53395]= 1765671509;
assign addr[53396]= 1743623590;
assign addr[53397]= 1721022648;
assign addr[53398]= 1697875851;
assign addr[53399]= 1674190539;
assign addr[53400]= 1649974225;
assign addr[53401]= 1625234591;
assign addr[53402]= 1599979481;
assign addr[53403]= 1574216908;
assign addr[53404]= 1547955041;
assign addr[53405]= 1521202211;
assign addr[53406]= 1493966902;
assign addr[53407]= 1466257752;
assign addr[53408]= 1438083551;
assign addr[53409]= 1409453233;
assign addr[53410]= 1380375881;
assign addr[53411]= 1350860716;
assign addr[53412]= 1320917099;
assign addr[53413]= 1290554528;
assign addr[53414]= 1259782632;
assign addr[53415]= 1228611172;
assign addr[53416]= 1197050035;
assign addr[53417]= 1165109230;
assign addr[53418]= 1132798888;
assign addr[53419]= 1100129257;
assign addr[53420]= 1067110699;
assign addr[53421]= 1033753687;
assign addr[53422]= 1000068799;
assign addr[53423]= 966066720;
assign addr[53424]= 931758235;
assign addr[53425]= 897154224;
assign addr[53426]= 862265664;
assign addr[53427]= 827103620;
assign addr[53428]= 791679244;
assign addr[53429]= 756003771;
assign addr[53430]= 720088517;
assign addr[53431]= 683944874;
assign addr[53432]= 647584304;
assign addr[53433]= 611018340;
assign addr[53434]= 574258580;
assign addr[53435]= 537316682;
assign addr[53436]= 500204365;
assign addr[53437]= 462933398;
assign addr[53438]= 425515602;
assign addr[53439]= 387962847;
assign addr[53440]= 350287041;
assign addr[53441]= 312500135;
assign addr[53442]= 274614114;
assign addr[53443]= 236640993;
assign addr[53444]= 198592817;
assign addr[53445]= 160481654;
assign addr[53446]= 122319591;
assign addr[53447]= 84118732;
assign addr[53448]= 45891193;
assign addr[53449]= 7649098;
assign addr[53450]= -30595422;
assign addr[53451]= -68830239;
assign addr[53452]= -107043224;
assign addr[53453]= -145222259;
assign addr[53454]= -183355234;
assign addr[53455]= -221430054;
assign addr[53456]= -259434643;
assign addr[53457]= -297356948;
assign addr[53458]= -335184940;
assign addr[53459]= -372906622;
assign addr[53460]= -410510029;
assign addr[53461]= -447983235;
assign addr[53462]= -485314355;
assign addr[53463]= -522491548;
assign addr[53464]= -559503022;
assign addr[53465]= -596337040;
assign addr[53466]= -632981917;
assign addr[53467]= -669426032;
assign addr[53468]= -705657826;
assign addr[53469]= -741665807;
assign addr[53470]= -777438554;
assign addr[53471]= -812964722;
assign addr[53472]= -848233042;
assign addr[53473]= -883232329;
assign addr[53474]= -917951481;
assign addr[53475]= -952379488;
assign addr[53476]= -986505429;
assign addr[53477]= -1020318481;
assign addr[53478]= -1053807919;
assign addr[53479]= -1086963121;
assign addr[53480]= -1119773573;
assign addr[53481]= -1152228866;
assign addr[53482]= -1184318708;
assign addr[53483]= -1216032921;
assign addr[53484]= -1247361445;
assign addr[53485]= -1278294345;
assign addr[53486]= -1308821808;
assign addr[53487]= -1338934154;
assign addr[53488]= -1368621831;
assign addr[53489]= -1397875423;
assign addr[53490]= -1426685652;
assign addr[53491]= -1455043381;
assign addr[53492]= -1482939614;
assign addr[53493]= -1510365504;
assign addr[53494]= -1537312353;
assign addr[53495]= -1563771613;
assign addr[53496]= -1589734894;
assign addr[53497]= -1615193959;
assign addr[53498]= -1640140734;
assign addr[53499]= -1664567307;
assign addr[53500]= -1688465931;
assign addr[53501]= -1711829025;
assign addr[53502]= -1734649179;
assign addr[53503]= -1756919156;
assign addr[53504]= -1778631892;
assign addr[53505]= -1799780501;
assign addr[53506]= -1820358275;
assign addr[53507]= -1840358687;
assign addr[53508]= -1859775393;
assign addr[53509]= -1878602237;
assign addr[53510]= -1896833245;
assign addr[53511]= -1914462636;
assign addr[53512]= -1931484818;
assign addr[53513]= -1947894393;
assign addr[53514]= -1963686155;
assign addr[53515]= -1978855097;
assign addr[53516]= -1993396407;
assign addr[53517]= -2007305472;
assign addr[53518]= -2020577882;
assign addr[53519]= -2033209426;
assign addr[53520]= -2045196100;
assign addr[53521]= -2056534099;
assign addr[53522]= -2067219829;
assign addr[53523]= -2077249901;
assign addr[53524]= -2086621133;
assign addr[53525]= -2095330553;
assign addr[53526]= -2103375398;
assign addr[53527]= -2110753117;
assign addr[53528]= -2117461370;
assign addr[53529]= -2123498030;
assign addr[53530]= -2128861181;
assign addr[53531]= -2133549123;
assign addr[53532]= -2137560369;
assign addr[53533]= -2140893646;
assign addr[53534]= -2143547897;
assign addr[53535]= -2145522281;
assign addr[53536]= -2146816171;
assign addr[53537]= -2147429158;
assign addr[53538]= -2147361045;
assign addr[53539]= -2146611856;
assign addr[53540]= -2145181827;
assign addr[53541]= -2143071413;
assign addr[53542]= -2140281282;
assign addr[53543]= -2136812319;
assign addr[53544]= -2132665626;
assign addr[53545]= -2127842516;
assign addr[53546]= -2122344521;
assign addr[53547]= -2116173382;
assign addr[53548]= -2109331059;
assign addr[53549]= -2101819720;
assign addr[53550]= -2093641749;
assign addr[53551]= -2084799740;
assign addr[53552]= -2075296495;
assign addr[53553]= -2065135031;
assign addr[53554]= -2054318569;
assign addr[53555]= -2042850540;
assign addr[53556]= -2030734582;
assign addr[53557]= -2017974537;
assign addr[53558]= -2004574453;
assign addr[53559]= -1990538579;
assign addr[53560]= -1975871368;
assign addr[53561]= -1960577471;
assign addr[53562]= -1944661739;
assign addr[53563]= -1928129220;
assign addr[53564]= -1910985158;
assign addr[53565]= -1893234990;
assign addr[53566]= -1874884346;
assign addr[53567]= -1855939047;
assign addr[53568]= -1836405100;
assign addr[53569]= -1816288703;
assign addr[53570]= -1795596234;
assign addr[53571]= -1774334257;
assign addr[53572]= -1752509516;
assign addr[53573]= -1730128933;
assign addr[53574]= -1707199606;
assign addr[53575]= -1683728808;
assign addr[53576]= -1659723983;
assign addr[53577]= -1635192744;
assign addr[53578]= -1610142873;
assign addr[53579]= -1584582314;
assign addr[53580]= -1558519173;
assign addr[53581]= -1531961719;
assign addr[53582]= -1504918373;
assign addr[53583]= -1477397714;
assign addr[53584]= -1449408469;
assign addr[53585]= -1420959516;
assign addr[53586]= -1392059879;
assign addr[53587]= -1362718723;
assign addr[53588]= -1332945355;
assign addr[53589]= -1302749217;
assign addr[53590]= -1272139887;
assign addr[53591]= -1241127074;
assign addr[53592]= -1209720613;
assign addr[53593]= -1177930466;
assign addr[53594]= -1145766716;
assign addr[53595]= -1113239564;
assign addr[53596]= -1080359326;
assign addr[53597]= -1047136432;
assign addr[53598]= -1013581418;
assign addr[53599]= -979704927;
assign addr[53600]= -945517704;
assign addr[53601]= -911030591;
assign addr[53602]= -876254528;
assign addr[53603]= -841200544;
assign addr[53604]= -805879757;
assign addr[53605]= -770303369;
assign addr[53606]= -734482665;
assign addr[53607]= -698429006;
assign addr[53608]= -662153826;
assign addr[53609]= -625668632;
assign addr[53610]= -588984994;
assign addr[53611]= -552114549;
assign addr[53612]= -515068990;
assign addr[53613]= -477860067;
assign addr[53614]= -440499581;
assign addr[53615]= -402999383;
assign addr[53616]= -365371365;
assign addr[53617]= -327627463;
assign addr[53618]= -289779648;
assign addr[53619]= -251839923;
assign addr[53620]= -213820322;
assign addr[53621]= -175732905;
assign addr[53622]= -137589750;
assign addr[53623]= -99402956;
assign addr[53624]= -61184634;
assign addr[53625]= -22946906;
assign addr[53626]= 15298099;
assign addr[53627]= 53538253;
assign addr[53628]= 91761426;
assign addr[53629]= 129955495;
assign addr[53630]= 168108346;
assign addr[53631]= 206207878;
assign addr[53632]= 244242007;
assign addr[53633]= 282198671;
assign addr[53634]= 320065829;
assign addr[53635]= 357831473;
assign addr[53636]= 395483624;
assign addr[53637]= 433010339;
assign addr[53638]= 470399716;
assign addr[53639]= 507639898;
assign addr[53640]= 544719071;
assign addr[53641]= 581625477;
assign addr[53642]= 618347408;
assign addr[53643]= 654873219;
assign addr[53644]= 691191324;
assign addr[53645]= 727290205;
assign addr[53646]= 763158411;
assign addr[53647]= 798784567;
assign addr[53648]= 834157373;
assign addr[53649]= 869265610;
assign addr[53650]= 904098143;
assign addr[53651]= 938643924;
assign addr[53652]= 972891995;
assign addr[53653]= 1006831495;
assign addr[53654]= 1040451659;
assign addr[53655]= 1073741824;
assign addr[53656]= 1106691431;
assign addr[53657]= 1139290029;
assign addr[53658]= 1171527280;
assign addr[53659]= 1203392958;
assign addr[53660]= 1234876957;
assign addr[53661]= 1265969291;
assign addr[53662]= 1296660098;
assign addr[53663]= 1326939644;
assign addr[53664]= 1356798326;
assign addr[53665]= 1386226674;
assign addr[53666]= 1415215352;
assign addr[53667]= 1443755168;
assign addr[53668]= 1471837070;
assign addr[53669]= 1499452149;
assign addr[53670]= 1526591649;
assign addr[53671]= 1553246960;
assign addr[53672]= 1579409630;
assign addr[53673]= 1605071359;
assign addr[53674]= 1630224009;
assign addr[53675]= 1654859602;
assign addr[53676]= 1678970324;
assign addr[53677]= 1702548529;
assign addr[53678]= 1725586737;
assign addr[53679]= 1748077642;
assign addr[53680]= 1770014111;
assign addr[53681]= 1791389186;
assign addr[53682]= 1812196087;
assign addr[53683]= 1832428215;
assign addr[53684]= 1852079154;
assign addr[53685]= 1871142669;
assign addr[53686]= 1889612716;
assign addr[53687]= 1907483436;
assign addr[53688]= 1924749160;
assign addr[53689]= 1941404413;
assign addr[53690]= 1957443913;
assign addr[53691]= 1972862571;
assign addr[53692]= 1987655498;
assign addr[53693]= 2001818002;
assign addr[53694]= 2015345591;
assign addr[53695]= 2028233973;
assign addr[53696]= 2040479063;
assign addr[53697]= 2052076975;
assign addr[53698]= 2063024031;
assign addr[53699]= 2073316760;
assign addr[53700]= 2082951896;
assign addr[53701]= 2091926384;
assign addr[53702]= 2100237377;
assign addr[53703]= 2107882239;
assign addr[53704]= 2114858546;
assign addr[53705]= 2121164085;
assign addr[53706]= 2126796855;
assign addr[53707]= 2131755071;
assign addr[53708]= 2136037160;
assign addr[53709]= 2139641764;
assign addr[53710]= 2142567738;
assign addr[53711]= 2144814157;
assign addr[53712]= 2146380306;
assign addr[53713]= 2147265689;
assign addr[53714]= 2147470025;
assign addr[53715]= 2146993250;
assign addr[53716]= 2145835515;
assign addr[53717]= 2143997187;
assign addr[53718]= 2141478848;
assign addr[53719]= 2138281298;
assign addr[53720]= 2134405552;
assign addr[53721]= 2129852837;
assign addr[53722]= 2124624598;
assign addr[53723]= 2118722494;
assign addr[53724]= 2112148396;
assign addr[53725]= 2104904390;
assign addr[53726]= 2096992772;
assign addr[53727]= 2088416053;
assign addr[53728]= 2079176953;
assign addr[53729]= 2069278401;
assign addr[53730]= 2058723538;
assign addr[53731]= 2047515711;
assign addr[53732]= 2035658475;
assign addr[53733]= 2023155591;
assign addr[53734]= 2010011024;
assign addr[53735]= 1996228943;
assign addr[53736]= 1981813720;
assign addr[53737]= 1966769926;
assign addr[53738]= 1951102334;
assign addr[53739]= 1934815911;
assign addr[53740]= 1917915825;
assign addr[53741]= 1900407434;
assign addr[53742]= 1882296293;
assign addr[53743]= 1863588145;
assign addr[53744]= 1844288924;
assign addr[53745]= 1824404752;
assign addr[53746]= 1803941934;
assign addr[53747]= 1782906961;
assign addr[53748]= 1761306505;
assign addr[53749]= 1739147417;
assign addr[53750]= 1716436725;
assign addr[53751]= 1693181631;
assign addr[53752]= 1669389513;
assign addr[53753]= 1645067915;
assign addr[53754]= 1620224553;
assign addr[53755]= 1594867305;
assign addr[53756]= 1569004214;
assign addr[53757]= 1542643483;
assign addr[53758]= 1515793473;
assign addr[53759]= 1488462700;
assign addr[53760]= 1460659832;
assign addr[53761]= 1432393688;
assign addr[53762]= 1403673233;
assign addr[53763]= 1374507575;
assign addr[53764]= 1344905966;
assign addr[53765]= 1314877795;
assign addr[53766]= 1284432584;
assign addr[53767]= 1253579991;
assign addr[53768]= 1222329801;
assign addr[53769]= 1190691925;
assign addr[53770]= 1158676398;
assign addr[53771]= 1126293375;
assign addr[53772]= 1093553126;
assign addr[53773]= 1060466036;
assign addr[53774]= 1027042599;
assign addr[53775]= 993293415;
assign addr[53776]= 959229189;
assign addr[53777]= 924860725;
assign addr[53778]= 890198924;
assign addr[53779]= 855254778;
assign addr[53780]= 820039373;
assign addr[53781]= 784563876;
assign addr[53782]= 748839539;
assign addr[53783]= 712877694;
assign addr[53784]= 676689746;
assign addr[53785]= 640287172;
assign addr[53786]= 603681519;
assign addr[53787]= 566884397;
assign addr[53788]= 529907477;
assign addr[53789]= 492762486;
assign addr[53790]= 455461206;
assign addr[53791]= 418015468;
assign addr[53792]= 380437148;
assign addr[53793]= 342738165;
assign addr[53794]= 304930476;
assign addr[53795]= 267026072;
assign addr[53796]= 229036977;
assign addr[53797]= 190975237;
assign addr[53798]= 152852926;
assign addr[53799]= 114682135;
assign addr[53800]= 76474970;
assign addr[53801]= 38243550;
assign addr[53802]= 0;
assign addr[53803]= -38243550;
assign addr[53804]= -76474970;
assign addr[53805]= -114682135;
assign addr[53806]= -152852926;
assign addr[53807]= -190975237;
assign addr[53808]= -229036977;
assign addr[53809]= -267026072;
assign addr[53810]= -304930476;
assign addr[53811]= -342738165;
assign addr[53812]= -380437148;
assign addr[53813]= -418015468;
assign addr[53814]= -455461206;
assign addr[53815]= -492762486;
assign addr[53816]= -529907477;
assign addr[53817]= -566884397;
assign addr[53818]= -603681519;
assign addr[53819]= -640287172;
assign addr[53820]= -676689746;
assign addr[53821]= -712877694;
assign addr[53822]= -748839539;
assign addr[53823]= -784563876;
assign addr[53824]= -820039373;
assign addr[53825]= -855254778;
assign addr[53826]= -890198924;
assign addr[53827]= -924860725;
assign addr[53828]= -959229189;
assign addr[53829]= -993293415;
assign addr[53830]= -1027042599;
assign addr[53831]= -1060466036;
assign addr[53832]= -1093553126;
assign addr[53833]= -1126293375;
assign addr[53834]= -1158676398;
assign addr[53835]= -1190691925;
assign addr[53836]= -1222329801;
assign addr[53837]= -1253579991;
assign addr[53838]= -1284432584;
assign addr[53839]= -1314877795;
assign addr[53840]= -1344905966;
assign addr[53841]= -1374507575;
assign addr[53842]= -1403673233;
assign addr[53843]= -1432393688;
assign addr[53844]= -1460659832;
assign addr[53845]= -1488462700;
assign addr[53846]= -1515793473;
assign addr[53847]= -1542643483;
assign addr[53848]= -1569004214;
assign addr[53849]= -1594867305;
assign addr[53850]= -1620224553;
assign addr[53851]= -1645067915;
assign addr[53852]= -1669389513;
assign addr[53853]= -1693181631;
assign addr[53854]= -1716436725;
assign addr[53855]= -1739147417;
assign addr[53856]= -1761306505;
assign addr[53857]= -1782906961;
assign addr[53858]= -1803941934;
assign addr[53859]= -1824404752;
assign addr[53860]= -1844288924;
assign addr[53861]= -1863588145;
assign addr[53862]= -1882296293;
assign addr[53863]= -1900407434;
assign addr[53864]= -1917915825;
assign addr[53865]= -1934815911;
assign addr[53866]= -1951102334;
assign addr[53867]= -1966769926;
assign addr[53868]= -1981813720;
assign addr[53869]= -1996228943;
assign addr[53870]= -2010011024;
assign addr[53871]= -2023155591;
assign addr[53872]= -2035658475;
assign addr[53873]= -2047515711;
assign addr[53874]= -2058723538;
assign addr[53875]= -2069278401;
assign addr[53876]= -2079176953;
assign addr[53877]= -2088416053;
assign addr[53878]= -2096992772;
assign addr[53879]= -2104904390;
assign addr[53880]= -2112148396;
assign addr[53881]= -2118722494;
assign addr[53882]= -2124624598;
assign addr[53883]= -2129852837;
assign addr[53884]= -2134405552;
assign addr[53885]= -2138281298;
assign addr[53886]= -2141478848;
assign addr[53887]= -2143997187;
assign addr[53888]= -2145835515;
assign addr[53889]= -2146993250;
assign addr[53890]= -2147470025;
assign addr[53891]= -2147265689;
assign addr[53892]= -2146380306;
assign addr[53893]= -2144814157;
assign addr[53894]= -2142567738;
assign addr[53895]= -2139641764;
assign addr[53896]= -2136037160;
assign addr[53897]= -2131755071;
assign addr[53898]= -2126796855;
assign addr[53899]= -2121164085;
assign addr[53900]= -2114858546;
assign addr[53901]= -2107882239;
assign addr[53902]= -2100237377;
assign addr[53903]= -2091926384;
assign addr[53904]= -2082951896;
assign addr[53905]= -2073316760;
assign addr[53906]= -2063024031;
assign addr[53907]= -2052076975;
assign addr[53908]= -2040479063;
assign addr[53909]= -2028233973;
assign addr[53910]= -2015345591;
assign addr[53911]= -2001818002;
assign addr[53912]= -1987655498;
assign addr[53913]= -1972862571;
assign addr[53914]= -1957443913;
assign addr[53915]= -1941404413;
assign addr[53916]= -1924749160;
assign addr[53917]= -1907483436;
assign addr[53918]= -1889612716;
assign addr[53919]= -1871142669;
assign addr[53920]= -1852079154;
assign addr[53921]= -1832428215;
assign addr[53922]= -1812196087;
assign addr[53923]= -1791389186;
assign addr[53924]= -1770014111;
assign addr[53925]= -1748077642;
assign addr[53926]= -1725586737;
assign addr[53927]= -1702548529;
assign addr[53928]= -1678970324;
assign addr[53929]= -1654859602;
assign addr[53930]= -1630224009;
assign addr[53931]= -1605071359;
assign addr[53932]= -1579409630;
assign addr[53933]= -1553246960;
assign addr[53934]= -1526591649;
assign addr[53935]= -1499452149;
assign addr[53936]= -1471837070;
assign addr[53937]= -1443755168;
assign addr[53938]= -1415215352;
assign addr[53939]= -1386226674;
assign addr[53940]= -1356798326;
assign addr[53941]= -1326939644;
assign addr[53942]= -1296660098;
assign addr[53943]= -1265969291;
assign addr[53944]= -1234876957;
assign addr[53945]= -1203392958;
assign addr[53946]= -1171527280;
assign addr[53947]= -1139290029;
assign addr[53948]= -1106691431;
assign addr[53949]= -1073741824;
assign addr[53950]= -1040451659;
assign addr[53951]= -1006831495;
assign addr[53952]= -972891995;
assign addr[53953]= -938643924;
assign addr[53954]= -904098143;
assign addr[53955]= -869265610;
assign addr[53956]= -834157373;
assign addr[53957]= -798784567;
assign addr[53958]= -763158411;
assign addr[53959]= -727290205;
assign addr[53960]= -691191324;
assign addr[53961]= -654873219;
assign addr[53962]= -618347408;
assign addr[53963]= -581625477;
assign addr[53964]= -544719071;
assign addr[53965]= -507639898;
assign addr[53966]= -470399716;
assign addr[53967]= -433010339;
assign addr[53968]= -395483624;
assign addr[53969]= -357831473;
assign addr[53970]= -320065829;
assign addr[53971]= -282198671;
assign addr[53972]= -244242007;
assign addr[53973]= -206207878;
assign addr[53974]= -168108346;
assign addr[53975]= -129955495;
assign addr[53976]= -91761426;
assign addr[53977]= -53538253;
assign addr[53978]= -15298099;
assign addr[53979]= 22946906;
assign addr[53980]= 61184634;
assign addr[53981]= 99402956;
assign addr[53982]= 137589750;
assign addr[53983]= 175732905;
assign addr[53984]= 213820322;
assign addr[53985]= 251839923;
assign addr[53986]= 289779648;
assign addr[53987]= 327627463;
assign addr[53988]= 365371365;
assign addr[53989]= 402999383;
assign addr[53990]= 440499581;
assign addr[53991]= 477860067;
assign addr[53992]= 515068990;
assign addr[53993]= 552114549;
assign addr[53994]= 588984994;
assign addr[53995]= 625668632;
assign addr[53996]= 662153826;
assign addr[53997]= 698429006;
assign addr[53998]= 734482665;
assign addr[53999]= 770303369;
assign addr[54000]= 805879757;
assign addr[54001]= 841200544;
assign addr[54002]= 876254528;
assign addr[54003]= 911030591;
assign addr[54004]= 945517704;
assign addr[54005]= 979704927;
assign addr[54006]= 1013581418;
assign addr[54007]= 1047136432;
assign addr[54008]= 1080359326;
assign addr[54009]= 1113239564;
assign addr[54010]= 1145766716;
assign addr[54011]= 1177930466;
assign addr[54012]= 1209720613;
assign addr[54013]= 1241127074;
assign addr[54014]= 1272139887;
assign addr[54015]= 1302749217;
assign addr[54016]= 1332945355;
assign addr[54017]= 1362718723;
assign addr[54018]= 1392059879;
assign addr[54019]= 1420959516;
assign addr[54020]= 1449408469;
assign addr[54021]= 1477397714;
assign addr[54022]= 1504918373;
assign addr[54023]= 1531961719;
assign addr[54024]= 1558519173;
assign addr[54025]= 1584582314;
assign addr[54026]= 1610142873;
assign addr[54027]= 1635192744;
assign addr[54028]= 1659723983;
assign addr[54029]= 1683728808;
assign addr[54030]= 1707199606;
assign addr[54031]= 1730128933;
assign addr[54032]= 1752509516;
assign addr[54033]= 1774334257;
assign addr[54034]= 1795596234;
assign addr[54035]= 1816288703;
assign addr[54036]= 1836405100;
assign addr[54037]= 1855939047;
assign addr[54038]= 1874884346;
assign addr[54039]= 1893234990;
assign addr[54040]= 1910985158;
assign addr[54041]= 1928129220;
assign addr[54042]= 1944661739;
assign addr[54043]= 1960577471;
assign addr[54044]= 1975871368;
assign addr[54045]= 1990538579;
assign addr[54046]= 2004574453;
assign addr[54047]= 2017974537;
assign addr[54048]= 2030734582;
assign addr[54049]= 2042850540;
assign addr[54050]= 2054318569;
assign addr[54051]= 2065135031;
assign addr[54052]= 2075296495;
assign addr[54053]= 2084799740;
assign addr[54054]= 2093641749;
assign addr[54055]= 2101819720;
assign addr[54056]= 2109331059;
assign addr[54057]= 2116173382;
assign addr[54058]= 2122344521;
assign addr[54059]= 2127842516;
assign addr[54060]= 2132665626;
assign addr[54061]= 2136812319;
assign addr[54062]= 2140281282;
assign addr[54063]= 2143071413;
assign addr[54064]= 2145181827;
assign addr[54065]= 2146611856;
assign addr[54066]= 2147361045;
assign addr[54067]= 2147429158;
assign addr[54068]= 2146816171;
assign addr[54069]= 2145522281;
assign addr[54070]= 2143547897;
assign addr[54071]= 2140893646;
assign addr[54072]= 2137560369;
assign addr[54073]= 2133549123;
assign addr[54074]= 2128861181;
assign addr[54075]= 2123498030;
assign addr[54076]= 2117461370;
assign addr[54077]= 2110753117;
assign addr[54078]= 2103375398;
assign addr[54079]= 2095330553;
assign addr[54080]= 2086621133;
assign addr[54081]= 2077249901;
assign addr[54082]= 2067219829;
assign addr[54083]= 2056534099;
assign addr[54084]= 2045196100;
assign addr[54085]= 2033209426;
assign addr[54086]= 2020577882;
assign addr[54087]= 2007305472;
assign addr[54088]= 1993396407;
assign addr[54089]= 1978855097;
assign addr[54090]= 1963686155;
assign addr[54091]= 1947894393;
assign addr[54092]= 1931484818;
assign addr[54093]= 1914462636;
assign addr[54094]= 1896833245;
assign addr[54095]= 1878602237;
assign addr[54096]= 1859775393;
assign addr[54097]= 1840358687;
assign addr[54098]= 1820358275;
assign addr[54099]= 1799780501;
assign addr[54100]= 1778631892;
assign addr[54101]= 1756919156;
assign addr[54102]= 1734649179;
assign addr[54103]= 1711829025;
assign addr[54104]= 1688465931;
assign addr[54105]= 1664567307;
assign addr[54106]= 1640140734;
assign addr[54107]= 1615193959;
assign addr[54108]= 1589734894;
assign addr[54109]= 1563771613;
assign addr[54110]= 1537312353;
assign addr[54111]= 1510365504;
assign addr[54112]= 1482939614;
assign addr[54113]= 1455043381;
assign addr[54114]= 1426685652;
assign addr[54115]= 1397875423;
assign addr[54116]= 1368621831;
assign addr[54117]= 1338934154;
assign addr[54118]= 1308821808;
assign addr[54119]= 1278294345;
assign addr[54120]= 1247361445;
assign addr[54121]= 1216032921;
assign addr[54122]= 1184318708;
assign addr[54123]= 1152228866;
assign addr[54124]= 1119773573;
assign addr[54125]= 1086963121;
assign addr[54126]= 1053807919;
assign addr[54127]= 1020318481;
assign addr[54128]= 986505429;
assign addr[54129]= 952379488;
assign addr[54130]= 917951481;
assign addr[54131]= 883232329;
assign addr[54132]= 848233042;
assign addr[54133]= 812964722;
assign addr[54134]= 777438554;
assign addr[54135]= 741665807;
assign addr[54136]= 705657826;
assign addr[54137]= 669426032;
assign addr[54138]= 632981917;
assign addr[54139]= 596337040;
assign addr[54140]= 559503022;
assign addr[54141]= 522491548;
assign addr[54142]= 485314355;
assign addr[54143]= 447983235;
assign addr[54144]= 410510029;
assign addr[54145]= 372906622;
assign addr[54146]= 335184940;
assign addr[54147]= 297356948;
assign addr[54148]= 259434643;
assign addr[54149]= 221430054;
assign addr[54150]= 183355234;
assign addr[54151]= 145222259;
assign addr[54152]= 107043224;
assign addr[54153]= 68830239;
assign addr[54154]= 30595422;
assign addr[54155]= -7649098;
assign addr[54156]= -45891193;
assign addr[54157]= -84118732;
assign addr[54158]= -122319591;
assign addr[54159]= -160481654;
assign addr[54160]= -198592817;
assign addr[54161]= -236640993;
assign addr[54162]= -274614114;
assign addr[54163]= -312500135;
assign addr[54164]= -350287041;
assign addr[54165]= -387962847;
assign addr[54166]= -425515602;
assign addr[54167]= -462933398;
assign addr[54168]= -500204365;
assign addr[54169]= -537316682;
assign addr[54170]= -574258580;
assign addr[54171]= -611018340;
assign addr[54172]= -647584304;
assign addr[54173]= -683944874;
assign addr[54174]= -720088517;
assign addr[54175]= -756003771;
assign addr[54176]= -791679244;
assign addr[54177]= -827103620;
assign addr[54178]= -862265664;
assign addr[54179]= -897154224;
assign addr[54180]= -931758235;
assign addr[54181]= -966066720;
assign addr[54182]= -1000068799;
assign addr[54183]= -1033753687;
assign addr[54184]= -1067110699;
assign addr[54185]= -1100129257;
assign addr[54186]= -1132798888;
assign addr[54187]= -1165109230;
assign addr[54188]= -1197050035;
assign addr[54189]= -1228611172;
assign addr[54190]= -1259782632;
assign addr[54191]= -1290554528;
assign addr[54192]= -1320917099;
assign addr[54193]= -1350860716;
assign addr[54194]= -1380375881;
assign addr[54195]= -1409453233;
assign addr[54196]= -1438083551;
assign addr[54197]= -1466257752;
assign addr[54198]= -1493966902;
assign addr[54199]= -1521202211;
assign addr[54200]= -1547955041;
assign addr[54201]= -1574216908;
assign addr[54202]= -1599979481;
assign addr[54203]= -1625234591;
assign addr[54204]= -1649974225;
assign addr[54205]= -1674190539;
assign addr[54206]= -1697875851;
assign addr[54207]= -1721022648;
assign addr[54208]= -1743623590;
assign addr[54209]= -1765671509;
assign addr[54210]= -1787159411;
assign addr[54211]= -1808080480;
assign addr[54212]= -1828428082;
assign addr[54213]= -1848195763;
assign addr[54214]= -1867377253;
assign addr[54215]= -1885966468;
assign addr[54216]= -1903957513;
assign addr[54217]= -1921344681;
assign addr[54218]= -1938122457;
assign addr[54219]= -1954285520;
assign addr[54220]= -1969828744;
assign addr[54221]= -1984747199;
assign addr[54222]= -1999036154;
assign addr[54223]= -2012691075;
assign addr[54224]= -2025707632;
assign addr[54225]= -2038081698;
assign addr[54226]= -2049809346;
assign addr[54227]= -2060886858;
assign addr[54228]= -2071310720;
assign addr[54229]= -2081077626;
assign addr[54230]= -2090184478;
assign addr[54231]= -2098628387;
assign addr[54232]= -2106406677;
assign addr[54233]= -2113516878;
assign addr[54234]= -2119956737;
assign addr[54235]= -2125724211;
assign addr[54236]= -2130817471;
assign addr[54237]= -2135234901;
assign addr[54238]= -2138975100;
assign addr[54239]= -2142036881;
assign addr[54240]= -2144419275;
assign addr[54241]= -2146121524;
assign addr[54242]= -2147143090;
assign addr[54243]= -2147483648;
assign addr[54244]= -2147143090;
assign addr[54245]= -2146121524;
assign addr[54246]= -2144419275;
assign addr[54247]= -2142036881;
assign addr[54248]= -2138975100;
assign addr[54249]= -2135234901;
assign addr[54250]= -2130817471;
assign addr[54251]= -2125724211;
assign addr[54252]= -2119956737;
assign addr[54253]= -2113516878;
assign addr[54254]= -2106406677;
assign addr[54255]= -2098628387;
assign addr[54256]= -2090184478;
assign addr[54257]= -2081077626;
assign addr[54258]= -2071310720;
assign addr[54259]= -2060886858;
assign addr[54260]= -2049809346;
assign addr[54261]= -2038081698;
assign addr[54262]= -2025707632;
assign addr[54263]= -2012691075;
assign addr[54264]= -1999036154;
assign addr[54265]= -1984747199;
assign addr[54266]= -1969828744;
assign addr[54267]= -1954285520;
assign addr[54268]= -1938122457;
assign addr[54269]= -1921344681;
assign addr[54270]= -1903957513;
assign addr[54271]= -1885966468;
assign addr[54272]= -1867377253;
assign addr[54273]= -1848195763;
assign addr[54274]= -1828428082;
assign addr[54275]= -1808080480;
assign addr[54276]= -1787159411;
assign addr[54277]= -1765671509;
assign addr[54278]= -1743623590;
assign addr[54279]= -1721022648;
assign addr[54280]= -1697875851;
assign addr[54281]= -1674190539;
assign addr[54282]= -1649974225;
assign addr[54283]= -1625234591;
assign addr[54284]= -1599979481;
assign addr[54285]= -1574216908;
assign addr[54286]= -1547955041;
assign addr[54287]= -1521202211;
assign addr[54288]= -1493966902;
assign addr[54289]= -1466257752;
assign addr[54290]= -1438083551;
assign addr[54291]= -1409453233;
assign addr[54292]= -1380375881;
assign addr[54293]= -1350860716;
assign addr[54294]= -1320917099;
assign addr[54295]= -1290554528;
assign addr[54296]= -1259782632;
assign addr[54297]= -1228611172;
assign addr[54298]= -1197050035;
assign addr[54299]= -1165109230;
assign addr[54300]= -1132798888;
assign addr[54301]= -1100129257;
assign addr[54302]= -1067110699;
assign addr[54303]= -1033753687;
assign addr[54304]= -1000068799;
assign addr[54305]= -966066720;
assign addr[54306]= -931758235;
assign addr[54307]= -897154224;
assign addr[54308]= -862265664;
assign addr[54309]= -827103620;
assign addr[54310]= -791679244;
assign addr[54311]= -756003771;
assign addr[54312]= -720088517;
assign addr[54313]= -683944874;
assign addr[54314]= -647584304;
assign addr[54315]= -611018340;
assign addr[54316]= -574258580;
assign addr[54317]= -537316682;
assign addr[54318]= -500204365;
assign addr[54319]= -462933398;
assign addr[54320]= -425515602;
assign addr[54321]= -387962847;
assign addr[54322]= -350287041;
assign addr[54323]= -312500135;
assign addr[54324]= -274614114;
assign addr[54325]= -236640993;
assign addr[54326]= -198592817;
assign addr[54327]= -160481654;
assign addr[54328]= -122319591;
assign addr[54329]= -84118732;
assign addr[54330]= -45891193;
assign addr[54331]= -7649098;
assign addr[54332]= 30595422;
assign addr[54333]= 68830239;
assign addr[54334]= 107043224;
assign addr[54335]= 145222259;
assign addr[54336]= 183355234;
assign addr[54337]= 221430054;
assign addr[54338]= 259434643;
assign addr[54339]= 297356948;
assign addr[54340]= 335184940;
assign addr[54341]= 372906622;
assign addr[54342]= 410510029;
assign addr[54343]= 447983235;
assign addr[54344]= 485314355;
assign addr[54345]= 522491548;
assign addr[54346]= 559503022;
assign addr[54347]= 596337040;
assign addr[54348]= 632981917;
assign addr[54349]= 669426032;
assign addr[54350]= 705657826;
assign addr[54351]= 741665807;
assign addr[54352]= 777438554;
assign addr[54353]= 812964722;
assign addr[54354]= 848233042;
assign addr[54355]= 883232329;
assign addr[54356]= 917951481;
assign addr[54357]= 952379488;
assign addr[54358]= 986505429;
assign addr[54359]= 1020318481;
assign addr[54360]= 1053807919;
assign addr[54361]= 1086963121;
assign addr[54362]= 1119773573;
assign addr[54363]= 1152228866;
assign addr[54364]= 1184318708;
assign addr[54365]= 1216032921;
assign addr[54366]= 1247361445;
assign addr[54367]= 1278294345;
assign addr[54368]= 1308821808;
assign addr[54369]= 1338934154;
assign addr[54370]= 1368621831;
assign addr[54371]= 1397875423;
assign addr[54372]= 1426685652;
assign addr[54373]= 1455043381;
assign addr[54374]= 1482939614;
assign addr[54375]= 1510365504;
assign addr[54376]= 1537312353;
assign addr[54377]= 1563771613;
assign addr[54378]= 1589734894;
assign addr[54379]= 1615193959;
assign addr[54380]= 1640140734;
assign addr[54381]= 1664567307;
assign addr[54382]= 1688465931;
assign addr[54383]= 1711829025;
assign addr[54384]= 1734649179;
assign addr[54385]= 1756919156;
assign addr[54386]= 1778631892;
assign addr[54387]= 1799780501;
assign addr[54388]= 1820358275;
assign addr[54389]= 1840358687;
assign addr[54390]= 1859775393;
assign addr[54391]= 1878602237;
assign addr[54392]= 1896833245;
assign addr[54393]= 1914462636;
assign addr[54394]= 1931484818;
assign addr[54395]= 1947894393;
assign addr[54396]= 1963686155;
assign addr[54397]= 1978855097;
assign addr[54398]= 1993396407;
assign addr[54399]= 2007305472;
assign addr[54400]= 2020577882;
assign addr[54401]= 2033209426;
assign addr[54402]= 2045196100;
assign addr[54403]= 2056534099;
assign addr[54404]= 2067219829;
assign addr[54405]= 2077249901;
assign addr[54406]= 2086621133;
assign addr[54407]= 2095330553;
assign addr[54408]= 2103375398;
assign addr[54409]= 2110753117;
assign addr[54410]= 2117461370;
assign addr[54411]= 2123498030;
assign addr[54412]= 2128861181;
assign addr[54413]= 2133549123;
assign addr[54414]= 2137560369;
assign addr[54415]= 2140893646;
assign addr[54416]= 2143547897;
assign addr[54417]= 2145522281;
assign addr[54418]= 2146816171;
assign addr[54419]= 2147429158;
assign addr[54420]= 2147361045;
assign addr[54421]= 2146611856;
assign addr[54422]= 2145181827;
assign addr[54423]= 2143071413;
assign addr[54424]= 2140281282;
assign addr[54425]= 2136812319;
assign addr[54426]= 2132665626;
assign addr[54427]= 2127842516;
assign addr[54428]= 2122344521;
assign addr[54429]= 2116173382;
assign addr[54430]= 2109331059;
assign addr[54431]= 2101819720;
assign addr[54432]= 2093641749;
assign addr[54433]= 2084799740;
assign addr[54434]= 2075296495;
assign addr[54435]= 2065135031;
assign addr[54436]= 2054318569;
assign addr[54437]= 2042850540;
assign addr[54438]= 2030734582;
assign addr[54439]= 2017974537;
assign addr[54440]= 2004574453;
assign addr[54441]= 1990538579;
assign addr[54442]= 1975871368;
assign addr[54443]= 1960577471;
assign addr[54444]= 1944661739;
assign addr[54445]= 1928129220;
assign addr[54446]= 1910985158;
assign addr[54447]= 1893234990;
assign addr[54448]= 1874884346;
assign addr[54449]= 1855939047;
assign addr[54450]= 1836405100;
assign addr[54451]= 1816288703;
assign addr[54452]= 1795596234;
assign addr[54453]= 1774334257;
assign addr[54454]= 1752509516;
assign addr[54455]= 1730128933;
assign addr[54456]= 1707199606;
assign addr[54457]= 1683728808;
assign addr[54458]= 1659723983;
assign addr[54459]= 1635192744;
assign addr[54460]= 1610142873;
assign addr[54461]= 1584582314;
assign addr[54462]= 1558519173;
assign addr[54463]= 1531961719;
assign addr[54464]= 1504918373;
assign addr[54465]= 1477397714;
assign addr[54466]= 1449408469;
assign addr[54467]= 1420959516;
assign addr[54468]= 1392059879;
assign addr[54469]= 1362718723;
assign addr[54470]= 1332945355;
assign addr[54471]= 1302749217;
assign addr[54472]= 1272139887;
assign addr[54473]= 1241127074;
assign addr[54474]= 1209720613;
assign addr[54475]= 1177930466;
assign addr[54476]= 1145766716;
assign addr[54477]= 1113239564;
assign addr[54478]= 1080359326;
assign addr[54479]= 1047136432;
assign addr[54480]= 1013581418;
assign addr[54481]= 979704927;
assign addr[54482]= 945517704;
assign addr[54483]= 911030591;
assign addr[54484]= 876254528;
assign addr[54485]= 841200544;
assign addr[54486]= 805879757;
assign addr[54487]= 770303369;
assign addr[54488]= 734482665;
assign addr[54489]= 698429006;
assign addr[54490]= 662153826;
assign addr[54491]= 625668632;
assign addr[54492]= 588984994;
assign addr[54493]= 552114549;
assign addr[54494]= 515068990;
assign addr[54495]= 477860067;
assign addr[54496]= 440499581;
assign addr[54497]= 402999383;
assign addr[54498]= 365371365;
assign addr[54499]= 327627463;
assign addr[54500]= 289779648;
assign addr[54501]= 251839923;
assign addr[54502]= 213820322;
assign addr[54503]= 175732905;
assign addr[54504]= 137589750;
assign addr[54505]= 99402956;
assign addr[54506]= 61184634;
assign addr[54507]= 22946906;
assign addr[54508]= -15298099;
assign addr[54509]= -53538253;
assign addr[54510]= -91761426;
assign addr[54511]= -129955495;
assign addr[54512]= -168108346;
assign addr[54513]= -206207878;
assign addr[54514]= -244242007;
assign addr[54515]= -282198671;
assign addr[54516]= -320065829;
assign addr[54517]= -357831473;
assign addr[54518]= -395483624;
assign addr[54519]= -433010339;
assign addr[54520]= -470399716;
assign addr[54521]= -507639898;
assign addr[54522]= -544719071;
assign addr[54523]= -581625477;
assign addr[54524]= -618347408;
assign addr[54525]= -654873219;
assign addr[54526]= -691191324;
assign addr[54527]= -727290205;
assign addr[54528]= -763158411;
assign addr[54529]= -798784567;
assign addr[54530]= -834157373;
assign addr[54531]= -869265610;
assign addr[54532]= -904098143;
assign addr[54533]= -938643924;
assign addr[54534]= -972891995;
assign addr[54535]= -1006831495;
assign addr[54536]= -1040451659;
assign addr[54537]= -1073741824;
assign addr[54538]= -1106691431;
assign addr[54539]= -1139290029;
assign addr[54540]= -1171527280;
assign addr[54541]= -1203392958;
assign addr[54542]= -1234876957;
assign addr[54543]= -1265969291;
assign addr[54544]= -1296660098;
assign addr[54545]= -1326939644;
assign addr[54546]= -1356798326;
assign addr[54547]= -1386226674;
assign addr[54548]= -1415215352;
assign addr[54549]= -1443755168;
assign addr[54550]= -1471837070;
assign addr[54551]= -1499452149;
assign addr[54552]= -1526591649;
assign addr[54553]= -1553246960;
assign addr[54554]= -1579409630;
assign addr[54555]= -1605071359;
assign addr[54556]= -1630224009;
assign addr[54557]= -1654859602;
assign addr[54558]= -1678970324;
assign addr[54559]= -1702548529;
assign addr[54560]= -1725586737;
assign addr[54561]= -1748077642;
assign addr[54562]= -1770014111;
assign addr[54563]= -1791389186;
assign addr[54564]= -1812196087;
assign addr[54565]= -1832428215;
assign addr[54566]= -1852079154;
assign addr[54567]= -1871142669;
assign addr[54568]= -1889612716;
assign addr[54569]= -1907483436;
assign addr[54570]= -1924749160;
assign addr[54571]= -1941404413;
assign addr[54572]= -1957443913;
assign addr[54573]= -1972862571;
assign addr[54574]= -1987655498;
assign addr[54575]= -2001818002;
assign addr[54576]= -2015345591;
assign addr[54577]= -2028233973;
assign addr[54578]= -2040479063;
assign addr[54579]= -2052076975;
assign addr[54580]= -2063024031;
assign addr[54581]= -2073316760;
assign addr[54582]= -2082951896;
assign addr[54583]= -2091926384;
assign addr[54584]= -2100237377;
assign addr[54585]= -2107882239;
assign addr[54586]= -2114858546;
assign addr[54587]= -2121164085;
assign addr[54588]= -2126796855;
assign addr[54589]= -2131755071;
assign addr[54590]= -2136037160;
assign addr[54591]= -2139641764;
assign addr[54592]= -2142567738;
assign addr[54593]= -2144814157;
assign addr[54594]= -2146380306;
assign addr[54595]= -2147265689;
assign addr[54596]= -2147470025;
assign addr[54597]= -2146993250;
assign addr[54598]= -2145835515;
assign addr[54599]= -2143997187;
assign addr[54600]= -2141478848;
assign addr[54601]= -2138281298;
assign addr[54602]= -2134405552;
assign addr[54603]= -2129852837;
assign addr[54604]= -2124624598;
assign addr[54605]= -2118722494;
assign addr[54606]= -2112148396;
assign addr[54607]= -2104904390;
assign addr[54608]= -2096992772;
assign addr[54609]= -2088416053;
assign addr[54610]= -2079176953;
assign addr[54611]= -2069278401;
assign addr[54612]= -2058723538;
assign addr[54613]= -2047515711;
assign addr[54614]= -2035658475;
assign addr[54615]= -2023155591;
assign addr[54616]= -2010011024;
assign addr[54617]= -1996228943;
assign addr[54618]= -1981813720;
assign addr[54619]= -1966769926;
assign addr[54620]= -1951102334;
assign addr[54621]= -1934815911;
assign addr[54622]= -1917915825;
assign addr[54623]= -1900407434;
assign addr[54624]= -1882296293;
assign addr[54625]= -1863588145;
assign addr[54626]= -1844288924;
assign addr[54627]= -1824404752;
assign addr[54628]= -1803941934;
assign addr[54629]= -1782906961;
assign addr[54630]= -1761306505;
assign addr[54631]= -1739147417;
assign addr[54632]= -1716436725;
assign addr[54633]= -1693181631;
assign addr[54634]= -1669389513;
assign addr[54635]= -1645067915;
assign addr[54636]= -1620224553;
assign addr[54637]= -1594867305;
assign addr[54638]= -1569004214;
assign addr[54639]= -1542643483;
assign addr[54640]= -1515793473;
assign addr[54641]= -1488462700;
assign addr[54642]= -1460659832;
assign addr[54643]= -1432393688;
assign addr[54644]= -1403673233;
assign addr[54645]= -1374507575;
assign addr[54646]= -1344905966;
assign addr[54647]= -1314877795;
assign addr[54648]= -1284432584;
assign addr[54649]= -1253579991;
assign addr[54650]= -1222329801;
assign addr[54651]= -1190691925;
assign addr[54652]= -1158676398;
assign addr[54653]= -1126293375;
assign addr[54654]= -1093553126;
assign addr[54655]= -1060466036;
assign addr[54656]= -1027042599;
assign addr[54657]= -993293415;
assign addr[54658]= -959229189;
assign addr[54659]= -924860725;
assign addr[54660]= -890198924;
assign addr[54661]= -855254778;
assign addr[54662]= -820039373;
assign addr[54663]= -784563876;
assign addr[54664]= -748839539;
assign addr[54665]= -712877694;
assign addr[54666]= -676689746;
assign addr[54667]= -640287172;
assign addr[54668]= -603681519;
assign addr[54669]= -566884397;
assign addr[54670]= -529907477;
assign addr[54671]= -492762486;
assign addr[54672]= -455461206;
assign addr[54673]= -418015468;
assign addr[54674]= -380437148;
assign addr[54675]= -342738165;
assign addr[54676]= -304930476;
assign addr[54677]= -267026072;
assign addr[54678]= -229036977;
assign addr[54679]= -190975237;
assign addr[54680]= -152852926;
assign addr[54681]= -114682135;
assign addr[54682]= -76474970;
assign addr[54683]= -38243550;
assign addr[54684]= 0;
assign addr[54685]= 38243550;
assign addr[54686]= 76474970;
assign addr[54687]= 114682135;
assign addr[54688]= 152852926;
assign addr[54689]= 190975237;
assign addr[54690]= 229036977;
assign addr[54691]= 267026072;
assign addr[54692]= 304930476;
assign addr[54693]= 342738165;
assign addr[54694]= 380437148;
assign addr[54695]= 418015468;
assign addr[54696]= 455461206;
assign addr[54697]= 492762486;
assign addr[54698]= 529907477;
assign addr[54699]= 566884397;
assign addr[54700]= 603681519;
assign addr[54701]= 640287172;
assign addr[54702]= 676689746;
assign addr[54703]= 712877694;
assign addr[54704]= 748839539;
assign addr[54705]= 784563876;
assign addr[54706]= 820039373;
assign addr[54707]= 855254778;
assign addr[54708]= 890198924;
assign addr[54709]= 924860725;
assign addr[54710]= 959229189;
assign addr[54711]= 993293415;
assign addr[54712]= 1027042599;
assign addr[54713]= 1060466036;
assign addr[54714]= 1093553126;
assign addr[54715]= 1126293375;
assign addr[54716]= 1158676398;
assign addr[54717]= 1190691925;
assign addr[54718]= 1222329801;
assign addr[54719]= 1253579991;
assign addr[54720]= 1284432584;
assign addr[54721]= 1314877795;
assign addr[54722]= 1344905966;
assign addr[54723]= 1374507575;
assign addr[54724]= 1403673233;
assign addr[54725]= 1432393688;
assign addr[54726]= 1460659832;
assign addr[54727]= 1488462700;
assign addr[54728]= 1515793473;
assign addr[54729]= 1542643483;
assign addr[54730]= 1569004214;
assign addr[54731]= 1594867305;
assign addr[54732]= 1620224553;
assign addr[54733]= 1645067915;
assign addr[54734]= 1669389513;
assign addr[54735]= 1693181631;
assign addr[54736]= 1716436725;
assign addr[54737]= 1739147417;
assign addr[54738]= 1761306505;
assign addr[54739]= 1782906961;
assign addr[54740]= 1803941934;
assign addr[54741]= 1824404752;
assign addr[54742]= 1844288924;
assign addr[54743]= 1863588145;
assign addr[54744]= 1882296293;
assign addr[54745]= 1900407434;
assign addr[54746]= 1917915825;
assign addr[54747]= 1934815911;
assign addr[54748]= 1951102334;
assign addr[54749]= 1966769926;
assign addr[54750]= 1981813720;
assign addr[54751]= 1996228943;
assign addr[54752]= 2010011024;
assign addr[54753]= 2023155591;
assign addr[54754]= 2035658475;
assign addr[54755]= 2047515711;
assign addr[54756]= 2058723538;
assign addr[54757]= 2069278401;
assign addr[54758]= 2079176953;
assign addr[54759]= 2088416053;
assign addr[54760]= 2096992772;
assign addr[54761]= 2104904390;
assign addr[54762]= 2112148396;
assign addr[54763]= 2118722494;
assign addr[54764]= 2124624598;
assign addr[54765]= 2129852837;
assign addr[54766]= 2134405552;
assign addr[54767]= 2138281298;
assign addr[54768]= 2141478848;
assign addr[54769]= 2143997187;
assign addr[54770]= 2145835515;
assign addr[54771]= 2146993250;
assign addr[54772]= 2147470025;
assign addr[54773]= 2147265689;
assign addr[54774]= 2146380306;
assign addr[54775]= 2144814157;
assign addr[54776]= 2142567738;
assign addr[54777]= 2139641764;
assign addr[54778]= 2136037160;
assign addr[54779]= 2131755071;
assign addr[54780]= 2126796855;
assign addr[54781]= 2121164085;
assign addr[54782]= 2114858546;
assign addr[54783]= 2107882239;
assign addr[54784]= 2100237377;
assign addr[54785]= 2091926384;
assign addr[54786]= 2082951896;
assign addr[54787]= 2073316760;
assign addr[54788]= 2063024031;
assign addr[54789]= 2052076975;
assign addr[54790]= 2040479063;
assign addr[54791]= 2028233973;
assign addr[54792]= 2015345591;
assign addr[54793]= 2001818002;
assign addr[54794]= 1987655498;
assign addr[54795]= 1972862571;
assign addr[54796]= 1957443913;
assign addr[54797]= 1941404413;
assign addr[54798]= 1924749160;
assign addr[54799]= 1907483436;
assign addr[54800]= 1889612716;
assign addr[54801]= 1871142669;
assign addr[54802]= 1852079154;
assign addr[54803]= 1832428215;
assign addr[54804]= 1812196087;
assign addr[54805]= 1791389186;
assign addr[54806]= 1770014111;
assign addr[54807]= 1748077642;
assign addr[54808]= 1725586737;
assign addr[54809]= 1702548529;
assign addr[54810]= 1678970324;
assign addr[54811]= 1654859602;
assign addr[54812]= 1630224009;
assign addr[54813]= 1605071359;
assign addr[54814]= 1579409630;
assign addr[54815]= 1553246960;
assign addr[54816]= 1526591649;
assign addr[54817]= 1499452149;
assign addr[54818]= 1471837070;
assign addr[54819]= 1443755168;
assign addr[54820]= 1415215352;
assign addr[54821]= 1386226674;
assign addr[54822]= 1356798326;
assign addr[54823]= 1326939644;
assign addr[54824]= 1296660098;
assign addr[54825]= 1265969291;
assign addr[54826]= 1234876957;
assign addr[54827]= 1203392958;
assign addr[54828]= 1171527280;
assign addr[54829]= 1139290029;
assign addr[54830]= 1106691431;
assign addr[54831]= 1073741824;
assign addr[54832]= 1040451659;
assign addr[54833]= 1006831495;
assign addr[54834]= 972891995;
assign addr[54835]= 938643924;
assign addr[54836]= 904098143;
assign addr[54837]= 869265610;
assign addr[54838]= 834157373;
assign addr[54839]= 798784567;
assign addr[54840]= 763158411;
assign addr[54841]= 727290205;
assign addr[54842]= 691191324;
assign addr[54843]= 654873219;
assign addr[54844]= 618347408;
assign addr[54845]= 581625477;
assign addr[54846]= 544719071;
assign addr[54847]= 507639898;
assign addr[54848]= 470399716;
assign addr[54849]= 433010339;
assign addr[54850]= 395483624;
assign addr[54851]= 357831473;
assign addr[54852]= 320065829;
assign addr[54853]= 282198671;
assign addr[54854]= 244242007;
assign addr[54855]= 206207878;
assign addr[54856]= 168108346;
assign addr[54857]= 129955495;
assign addr[54858]= 91761426;
assign addr[54859]= 53538253;
assign addr[54860]= 15298099;
assign addr[54861]= -22946906;
assign addr[54862]= -61184634;
assign addr[54863]= -99402956;
assign addr[54864]= -137589750;
assign addr[54865]= -175732905;
assign addr[54866]= -213820322;
assign addr[54867]= -251839923;
assign addr[54868]= -289779648;
assign addr[54869]= -327627463;
assign addr[54870]= -365371365;
assign addr[54871]= -402999383;
assign addr[54872]= -440499581;
assign addr[54873]= -477860067;
assign addr[54874]= -515068990;
assign addr[54875]= -552114549;
assign addr[54876]= -588984994;
assign addr[54877]= -625668632;
assign addr[54878]= -662153826;
assign addr[54879]= -698429006;
assign addr[54880]= -734482665;
assign addr[54881]= -770303369;
assign addr[54882]= -805879757;
assign addr[54883]= -841200544;
assign addr[54884]= -876254528;
assign addr[54885]= -911030591;
assign addr[54886]= -945517704;
assign addr[54887]= -979704927;
assign addr[54888]= -1013581418;
assign addr[54889]= -1047136432;
assign addr[54890]= -1080359326;
assign addr[54891]= -1113239564;
assign addr[54892]= -1145766716;
assign addr[54893]= -1177930466;
assign addr[54894]= -1209720613;
assign addr[54895]= -1241127074;
assign addr[54896]= -1272139887;
assign addr[54897]= -1302749217;
assign addr[54898]= -1332945355;
assign addr[54899]= -1362718723;
assign addr[54900]= -1392059879;
assign addr[54901]= -1420959516;
assign addr[54902]= -1449408469;
assign addr[54903]= -1477397714;
assign addr[54904]= -1504918373;
assign addr[54905]= -1531961719;
assign addr[54906]= -1558519173;
assign addr[54907]= -1584582314;
assign addr[54908]= -1610142873;
assign addr[54909]= -1635192744;
assign addr[54910]= -1659723983;
assign addr[54911]= -1683728808;
assign addr[54912]= -1707199606;
assign addr[54913]= -1730128933;
assign addr[54914]= -1752509516;
assign addr[54915]= -1774334257;
assign addr[54916]= -1795596234;
assign addr[54917]= -1816288703;
assign addr[54918]= -1836405100;
assign addr[54919]= -1855939047;
assign addr[54920]= -1874884346;
assign addr[54921]= -1893234990;
assign addr[54922]= -1910985158;
assign addr[54923]= -1928129220;
assign addr[54924]= -1944661739;
assign addr[54925]= -1960577471;
assign addr[54926]= -1975871368;
assign addr[54927]= -1990538579;
assign addr[54928]= -2004574453;
assign addr[54929]= -2017974537;
assign addr[54930]= -2030734582;
assign addr[54931]= -2042850540;
assign addr[54932]= -2054318569;
assign addr[54933]= -2065135031;
assign addr[54934]= -2075296495;
assign addr[54935]= -2084799740;
assign addr[54936]= -2093641749;
assign addr[54937]= -2101819720;
assign addr[54938]= -2109331059;
assign addr[54939]= -2116173382;
assign addr[54940]= -2122344521;
assign addr[54941]= -2127842516;
assign addr[54942]= -2132665626;
assign addr[54943]= -2136812319;
assign addr[54944]= -2140281282;
assign addr[54945]= -2143071413;
assign addr[54946]= -2145181827;
assign addr[54947]= -2146611856;
assign addr[54948]= -2147361045;
assign addr[54949]= -2147429158;
assign addr[54950]= -2146816171;
assign addr[54951]= -2145522281;
assign addr[54952]= -2143547897;
assign addr[54953]= -2140893646;
assign addr[54954]= -2137560369;
assign addr[54955]= -2133549123;
assign addr[54956]= -2128861181;
assign addr[54957]= -2123498030;
assign addr[54958]= -2117461370;
assign addr[54959]= -2110753117;
assign addr[54960]= -2103375398;
assign addr[54961]= -2095330553;
assign addr[54962]= -2086621133;
assign addr[54963]= -2077249901;
assign addr[54964]= -2067219829;
assign addr[54965]= -2056534099;
assign addr[54966]= -2045196100;
assign addr[54967]= -2033209426;
assign addr[54968]= -2020577882;
assign addr[54969]= -2007305472;
assign addr[54970]= -1993396407;
assign addr[54971]= -1978855097;
assign addr[54972]= -1963686155;
assign addr[54973]= -1947894393;
assign addr[54974]= -1931484818;
assign addr[54975]= -1914462636;
assign addr[54976]= -1896833245;
assign addr[54977]= -1878602237;
assign addr[54978]= -1859775393;
assign addr[54979]= -1840358687;
assign addr[54980]= -1820358275;
assign addr[54981]= -1799780501;
assign addr[54982]= -1778631892;
assign addr[54983]= -1756919156;
assign addr[54984]= -1734649179;
assign addr[54985]= -1711829025;
assign addr[54986]= -1688465931;
assign addr[54987]= -1664567307;
assign addr[54988]= -1640140734;
assign addr[54989]= -1615193959;
assign addr[54990]= -1589734894;
assign addr[54991]= -1563771613;
assign addr[54992]= -1537312353;
assign addr[54993]= -1510365504;
assign addr[54994]= -1482939614;
assign addr[54995]= -1455043381;
assign addr[54996]= -1426685652;
assign addr[54997]= -1397875423;
assign addr[54998]= -1368621831;
assign addr[54999]= -1338934154;
assign addr[55000]= -1308821808;
assign addr[55001]= -1278294345;
assign addr[55002]= -1247361445;
assign addr[55003]= -1216032921;
assign addr[55004]= -1184318708;
assign addr[55005]= -1152228866;
assign addr[55006]= -1119773573;
assign addr[55007]= -1086963121;
assign addr[55008]= -1053807919;
assign addr[55009]= -1020318481;
assign addr[55010]= -986505429;
assign addr[55011]= -952379488;
assign addr[55012]= -917951481;
assign addr[55013]= -883232329;
assign addr[55014]= -848233042;
assign addr[55015]= -812964722;
assign addr[55016]= -777438554;
assign addr[55017]= -741665807;
assign addr[55018]= -705657826;
assign addr[55019]= -669426032;
assign addr[55020]= -632981917;
assign addr[55021]= -596337040;
assign addr[55022]= -559503022;
assign addr[55023]= -522491548;
assign addr[55024]= -485314355;
assign addr[55025]= -447983235;
assign addr[55026]= -410510029;
assign addr[55027]= -372906622;
assign addr[55028]= -335184940;
assign addr[55029]= -297356948;
assign addr[55030]= -259434643;
assign addr[55031]= -221430054;
assign addr[55032]= -183355234;
assign addr[55033]= -145222259;
assign addr[55034]= -107043224;
assign addr[55035]= -68830239;
assign addr[55036]= -30595422;
assign addr[55037]= 7649098;
assign addr[55038]= 45891193;
assign addr[55039]= 84118732;
assign addr[55040]= 122319591;
assign addr[55041]= 160481654;
assign addr[55042]= 198592817;
assign addr[55043]= 236640993;
assign addr[55044]= 274614114;
assign addr[55045]= 312500135;
assign addr[55046]= 350287041;
assign addr[55047]= 387962847;
assign addr[55048]= 425515602;
assign addr[55049]= 462933398;
assign addr[55050]= 500204365;
assign addr[55051]= 537316682;
assign addr[55052]= 574258580;
assign addr[55053]= 611018340;
assign addr[55054]= 647584304;
assign addr[55055]= 683944874;
assign addr[55056]= 720088517;
assign addr[55057]= 756003771;
assign addr[55058]= 791679244;
assign addr[55059]= 827103620;
assign addr[55060]= 862265664;
assign addr[55061]= 897154224;
assign addr[55062]= 931758235;
assign addr[55063]= 966066720;
assign addr[55064]= 1000068799;
assign addr[55065]= 1033753687;
assign addr[55066]= 1067110699;
assign addr[55067]= 1100129257;
assign addr[55068]= 1132798888;
assign addr[55069]= 1165109230;
assign addr[55070]= 1197050035;
assign addr[55071]= 1228611172;
assign addr[55072]= 1259782632;
assign addr[55073]= 1290554528;
assign addr[55074]= 1320917099;
assign addr[55075]= 1350860716;
assign addr[55076]= 1380375881;
assign addr[55077]= 1409453233;
assign addr[55078]= 1438083551;
assign addr[55079]= 1466257752;
assign addr[55080]= 1493966902;
assign addr[55081]= 1521202211;
assign addr[55082]= 1547955041;
assign addr[55083]= 1574216908;
assign addr[55084]= 1599979481;
assign addr[55085]= 1625234591;
assign addr[55086]= 1649974225;
assign addr[55087]= 1674190539;
assign addr[55088]= 1697875851;
assign addr[55089]= 1721022648;
assign addr[55090]= 1743623590;
assign addr[55091]= 1765671509;
assign addr[55092]= 1787159411;
assign addr[55093]= 1808080480;
assign addr[55094]= 1828428082;
assign addr[55095]= 1848195763;
assign addr[55096]= 1867377253;
assign addr[55097]= 1885966468;
assign addr[55098]= 1903957513;
assign addr[55099]= 1921344681;
assign addr[55100]= 1938122457;
assign addr[55101]= 1954285520;
assign addr[55102]= 1969828744;
assign addr[55103]= 1984747199;
assign addr[55104]= 1999036154;
assign addr[55105]= 2012691075;
assign addr[55106]= 2025707632;
assign addr[55107]= 2038081698;
assign addr[55108]= 2049809346;
assign addr[55109]= 2060886858;
assign addr[55110]= 2071310720;
assign addr[55111]= 2081077626;
assign addr[55112]= 2090184478;
assign addr[55113]= 2098628387;
assign addr[55114]= 2106406677;
assign addr[55115]= 2113516878;
assign addr[55116]= 2119956737;
assign addr[55117]= 2125724211;
assign addr[55118]= 2130817471;
assign addr[55119]= 2135234901;
assign addr[55120]= 2138975100;
assign addr[55121]= 2142036881;
assign addr[55122]= 2144419275;
assign addr[55123]= 2146121524;
assign addr[55124]= 2147143090;
assign addr[55125]= 2147483648;
assign addr[55126]= 2147143090;
assign addr[55127]= 2146121524;
assign addr[55128]= 2144419275;
assign addr[55129]= 2142036881;
assign addr[55130]= 2138975100;
assign addr[55131]= 2135234901;
assign addr[55132]= 2130817471;
assign addr[55133]= 2125724211;
assign addr[55134]= 2119956737;
assign addr[55135]= 2113516878;
assign addr[55136]= 2106406677;
assign addr[55137]= 2098628387;
assign addr[55138]= 2090184478;
assign addr[55139]= 2081077626;
assign addr[55140]= 2071310720;
assign addr[55141]= 2060886858;
assign addr[55142]= 2049809346;
assign addr[55143]= 2038081698;
assign addr[55144]= 2025707632;
assign addr[55145]= 2012691075;
assign addr[55146]= 1999036154;
assign addr[55147]= 1984747199;
assign addr[55148]= 1969828744;
assign addr[55149]= 1954285520;
assign addr[55150]= 1938122457;
assign addr[55151]= 1921344681;
assign addr[55152]= 1903957513;
assign addr[55153]= 1885966468;
assign addr[55154]= 1867377253;
assign addr[55155]= 1848195763;
assign addr[55156]= 1828428082;
assign addr[55157]= 1808080480;
assign addr[55158]= 1787159411;
assign addr[55159]= 1765671509;
assign addr[55160]= 1743623590;
assign addr[55161]= 1721022648;
assign addr[55162]= 1697875851;
assign addr[55163]= 1674190539;
assign addr[55164]= 1649974225;
assign addr[55165]= 1625234591;
assign addr[55166]= 1599979481;
assign addr[55167]= 1574216908;
assign addr[55168]= 1547955041;
assign addr[55169]= 1521202211;
assign addr[55170]= 1493966902;
assign addr[55171]= 1466257752;
assign addr[55172]= 1438083551;
assign addr[55173]= 1409453233;
assign addr[55174]= 1380375881;
assign addr[55175]= 1350860716;
assign addr[55176]= 1320917099;
assign addr[55177]= 1290554528;
assign addr[55178]= 1259782632;
assign addr[55179]= 1228611172;
assign addr[55180]= 1197050035;
assign addr[55181]= 1165109230;
assign addr[55182]= 1132798888;
assign addr[55183]= 1100129257;
assign addr[55184]= 1067110699;
assign addr[55185]= 1033753687;
assign addr[55186]= 1000068799;
assign addr[55187]= 966066720;
assign addr[55188]= 931758235;
assign addr[55189]= 897154224;
assign addr[55190]= 862265664;
assign addr[55191]= 827103620;
assign addr[55192]= 791679244;
assign addr[55193]= 756003771;
assign addr[55194]= 720088517;
assign addr[55195]= 683944874;
assign addr[55196]= 647584304;
assign addr[55197]= 611018340;
assign addr[55198]= 574258580;
assign addr[55199]= 537316682;
assign addr[55200]= 500204365;
assign addr[55201]= 462933398;
assign addr[55202]= 425515602;
assign addr[55203]= 387962847;
assign addr[55204]= 350287041;
assign addr[55205]= 312500135;
assign addr[55206]= 274614114;
assign addr[55207]= 236640993;
assign addr[55208]= 198592817;
assign addr[55209]= 160481654;
assign addr[55210]= 122319591;
assign addr[55211]= 84118732;
assign addr[55212]= 45891193;
assign addr[55213]= 7649098;
assign addr[55214]= -30595422;
assign addr[55215]= -68830239;
assign addr[55216]= -107043224;
assign addr[55217]= -145222259;
assign addr[55218]= -183355234;
assign addr[55219]= -221430054;
assign addr[55220]= -259434643;
assign addr[55221]= -297356948;
assign addr[55222]= -335184940;
assign addr[55223]= -372906622;
assign addr[55224]= -410510029;
assign addr[55225]= -447983235;
assign addr[55226]= -485314355;
assign addr[55227]= -522491548;
assign addr[55228]= -559503022;
assign addr[55229]= -596337040;
assign addr[55230]= -632981917;
assign addr[55231]= -669426032;
assign addr[55232]= -705657826;
assign addr[55233]= -741665807;
assign addr[55234]= -777438554;
assign addr[55235]= -812964722;
assign addr[55236]= -848233042;
assign addr[55237]= -883232329;
assign addr[55238]= -917951481;
assign addr[55239]= -952379488;
assign addr[55240]= -986505429;
assign addr[55241]= -1020318481;
assign addr[55242]= -1053807919;
assign addr[55243]= -1086963121;
assign addr[55244]= -1119773573;
assign addr[55245]= -1152228866;
assign addr[55246]= -1184318708;
assign addr[55247]= -1216032921;
assign addr[55248]= -1247361445;
assign addr[55249]= -1278294345;
assign addr[55250]= -1308821808;
assign addr[55251]= -1338934154;
assign addr[55252]= -1368621831;
assign addr[55253]= -1397875423;
assign addr[55254]= -1426685652;
assign addr[55255]= -1455043381;
assign addr[55256]= -1482939614;
assign addr[55257]= -1510365504;
assign addr[55258]= -1537312353;
assign addr[55259]= -1563771613;
assign addr[55260]= -1589734894;
assign addr[55261]= -1615193959;
assign addr[55262]= -1640140734;
assign addr[55263]= -1664567307;
assign addr[55264]= -1688465931;
assign addr[55265]= -1711829025;
assign addr[55266]= -1734649179;
assign addr[55267]= -1756919156;
assign addr[55268]= -1778631892;
assign addr[55269]= -1799780501;
assign addr[55270]= -1820358275;
assign addr[55271]= -1840358687;
assign addr[55272]= -1859775393;
assign addr[55273]= -1878602237;
assign addr[55274]= -1896833245;
assign addr[55275]= -1914462636;
assign addr[55276]= -1931484818;
assign addr[55277]= -1947894393;
assign addr[55278]= -1963686155;
assign addr[55279]= -1978855097;
assign addr[55280]= -1993396407;
assign addr[55281]= -2007305472;
assign addr[55282]= -2020577882;
assign addr[55283]= -2033209426;
assign addr[55284]= -2045196100;
assign addr[55285]= -2056534099;
assign addr[55286]= -2067219829;
assign addr[55287]= -2077249901;
assign addr[55288]= -2086621133;
assign addr[55289]= -2095330553;
assign addr[55290]= -2103375398;
assign addr[55291]= -2110753117;
assign addr[55292]= -2117461370;
assign addr[55293]= -2123498030;
assign addr[55294]= -2128861181;
assign addr[55295]= -2133549123;
assign addr[55296]= -2137560369;
assign addr[55297]= -2140893646;
assign addr[55298]= -2143547897;
assign addr[55299]= -2145522281;
assign addr[55300]= -2146816171;
assign addr[55301]= -2147429158;
assign addr[55302]= -2147361045;
assign addr[55303]= -2146611856;
assign addr[55304]= -2145181827;
assign addr[55305]= -2143071413;
assign addr[55306]= -2140281282;
assign addr[55307]= -2136812319;
assign addr[55308]= -2132665626;
assign addr[55309]= -2127842516;
assign addr[55310]= -2122344521;
assign addr[55311]= -2116173382;
assign addr[55312]= -2109331059;
assign addr[55313]= -2101819720;
assign addr[55314]= -2093641749;
assign addr[55315]= -2084799740;
assign addr[55316]= -2075296495;
assign addr[55317]= -2065135031;
assign addr[55318]= -2054318569;
assign addr[55319]= -2042850540;
assign addr[55320]= -2030734582;
assign addr[55321]= -2017974537;
assign addr[55322]= -2004574453;
assign addr[55323]= -1990538579;
assign addr[55324]= -1975871368;
assign addr[55325]= -1960577471;
assign addr[55326]= -1944661739;
assign addr[55327]= -1928129220;
assign addr[55328]= -1910985158;
assign addr[55329]= -1893234990;
assign addr[55330]= -1874884346;
assign addr[55331]= -1855939047;
assign addr[55332]= -1836405100;
assign addr[55333]= -1816288703;
assign addr[55334]= -1795596234;
assign addr[55335]= -1774334257;
assign addr[55336]= -1752509516;
assign addr[55337]= -1730128933;
assign addr[55338]= -1707199606;
assign addr[55339]= -1683728808;
assign addr[55340]= -1659723983;
assign addr[55341]= -1635192744;
assign addr[55342]= -1610142873;
assign addr[55343]= -1584582314;
assign addr[55344]= -1558519173;
assign addr[55345]= -1531961719;
assign addr[55346]= -1504918373;
assign addr[55347]= -1477397714;
assign addr[55348]= -1449408469;
assign addr[55349]= -1420959516;
assign addr[55350]= -1392059879;
assign addr[55351]= -1362718723;
assign addr[55352]= -1332945355;
assign addr[55353]= -1302749217;
assign addr[55354]= -1272139887;
assign addr[55355]= -1241127074;
assign addr[55356]= -1209720613;
assign addr[55357]= -1177930466;
assign addr[55358]= -1145766716;
assign addr[55359]= -1113239564;
assign addr[55360]= -1080359326;
assign addr[55361]= -1047136432;
assign addr[55362]= -1013581418;
assign addr[55363]= -979704927;
assign addr[55364]= -945517704;
assign addr[55365]= -911030591;
assign addr[55366]= -876254528;
assign addr[55367]= -841200544;
assign addr[55368]= -805879757;
assign addr[55369]= -770303369;
assign addr[55370]= -734482665;
assign addr[55371]= -698429006;
assign addr[55372]= -662153826;
assign addr[55373]= -625668632;
assign addr[55374]= -588984994;
assign addr[55375]= -552114549;
assign addr[55376]= -515068990;
assign addr[55377]= -477860067;
assign addr[55378]= -440499581;
assign addr[55379]= -402999383;
assign addr[55380]= -365371365;
assign addr[55381]= -327627463;
assign addr[55382]= -289779648;
assign addr[55383]= -251839923;
assign addr[55384]= -213820322;
assign addr[55385]= -175732905;
assign addr[55386]= -137589750;
assign addr[55387]= -99402956;
assign addr[55388]= -61184634;
assign addr[55389]= -22946906;
assign addr[55390]= 15298099;
assign addr[55391]= 53538253;
assign addr[55392]= 91761426;
assign addr[55393]= 129955495;
assign addr[55394]= 168108346;
assign addr[55395]= 206207878;
assign addr[55396]= 244242007;
assign addr[55397]= 282198671;
assign addr[55398]= 320065829;
assign addr[55399]= 357831473;
assign addr[55400]= 395483624;
assign addr[55401]= 433010339;
assign addr[55402]= 470399716;
assign addr[55403]= 507639898;
assign addr[55404]= 544719071;
assign addr[55405]= 581625477;
assign addr[55406]= 618347408;
assign addr[55407]= 654873219;
assign addr[55408]= 691191324;
assign addr[55409]= 727290205;
assign addr[55410]= 763158411;
assign addr[55411]= 798784567;
assign addr[55412]= 834157373;
assign addr[55413]= 869265610;
assign addr[55414]= 904098143;
assign addr[55415]= 938643924;
assign addr[55416]= 972891995;
assign addr[55417]= 1006831495;
assign addr[55418]= 1040451659;
assign addr[55419]= 1073741824;
assign addr[55420]= 1106691431;
assign addr[55421]= 1139290029;
assign addr[55422]= 1171527280;
assign addr[55423]= 1203392958;
assign addr[55424]= 1234876957;
assign addr[55425]= 1265969291;
assign addr[55426]= 1296660098;
assign addr[55427]= 1326939644;
assign addr[55428]= 1356798326;
assign addr[55429]= 1386226674;
assign addr[55430]= 1415215352;
assign addr[55431]= 1443755168;
assign addr[55432]= 1471837070;
assign addr[55433]= 1499452149;
assign addr[55434]= 1526591649;
assign addr[55435]= 1553246960;
assign addr[55436]= 1579409630;
assign addr[55437]= 1605071359;
assign addr[55438]= 1630224009;
assign addr[55439]= 1654859602;
assign addr[55440]= 1678970324;
assign addr[55441]= 1702548529;
assign addr[55442]= 1725586737;
assign addr[55443]= 1748077642;
assign addr[55444]= 1770014111;
assign addr[55445]= 1791389186;
assign addr[55446]= 1812196087;
assign addr[55447]= 1832428215;
assign addr[55448]= 1852079154;
assign addr[55449]= 1871142669;
assign addr[55450]= 1889612716;
assign addr[55451]= 1907483436;
assign addr[55452]= 1924749160;
assign addr[55453]= 1941404413;
assign addr[55454]= 1957443913;
assign addr[55455]= 1972862571;
assign addr[55456]= 1987655498;
assign addr[55457]= 2001818002;
assign addr[55458]= 2015345591;
assign addr[55459]= 2028233973;
assign addr[55460]= 2040479063;
assign addr[55461]= 2052076975;
assign addr[55462]= 2063024031;
assign addr[55463]= 2073316760;
assign addr[55464]= 2082951896;
assign addr[55465]= 2091926384;
assign addr[55466]= 2100237377;
assign addr[55467]= 2107882239;
assign addr[55468]= 2114858546;
assign addr[55469]= 2121164085;
assign addr[55470]= 2126796855;
assign addr[55471]= 2131755071;
assign addr[55472]= 2136037160;
assign addr[55473]= 2139641764;
assign addr[55474]= 2142567738;
assign addr[55475]= 2144814157;
assign addr[55476]= 2146380306;
assign addr[55477]= 2147265689;
assign addr[55478]= 2147470025;
assign addr[55479]= 2146993250;
assign addr[55480]= 2145835515;
assign addr[55481]= 2143997187;
assign addr[55482]= 2141478848;
assign addr[55483]= 2138281298;
assign addr[55484]= 2134405552;
assign addr[55485]= 2129852837;
assign addr[55486]= 2124624598;
assign addr[55487]= 2118722494;
assign addr[55488]= 2112148396;
assign addr[55489]= 2104904390;
assign addr[55490]= 2096992772;
assign addr[55491]= 2088416053;
assign addr[55492]= 2079176953;
assign addr[55493]= 2069278401;
assign addr[55494]= 2058723538;
assign addr[55495]= 2047515711;
assign addr[55496]= 2035658475;
assign addr[55497]= 2023155591;
assign addr[55498]= 2010011024;
assign addr[55499]= 1996228943;
assign addr[55500]= 1981813720;
assign addr[55501]= 1966769926;
assign addr[55502]= 1951102334;
assign addr[55503]= 1934815911;
assign addr[55504]= 1917915825;
assign addr[55505]= 1900407434;
assign addr[55506]= 1882296293;
assign addr[55507]= 1863588145;
assign addr[55508]= 1844288924;
assign addr[55509]= 1824404752;
assign addr[55510]= 1803941934;
assign addr[55511]= 1782906961;
assign addr[55512]= 1761306505;
assign addr[55513]= 1739147417;
assign addr[55514]= 1716436725;
assign addr[55515]= 1693181631;
assign addr[55516]= 1669389513;
assign addr[55517]= 1645067915;
assign addr[55518]= 1620224553;
assign addr[55519]= 1594867305;
assign addr[55520]= 1569004214;
assign addr[55521]= 1542643483;
assign addr[55522]= 1515793473;
assign addr[55523]= 1488462700;
assign addr[55524]= 1460659832;
assign addr[55525]= 1432393688;
assign addr[55526]= 1403673233;
assign addr[55527]= 1374507575;
assign addr[55528]= 1344905966;
assign addr[55529]= 1314877795;
assign addr[55530]= 1284432584;
assign addr[55531]= 1253579991;
assign addr[55532]= 1222329801;
assign addr[55533]= 1190691925;
assign addr[55534]= 1158676398;
assign addr[55535]= 1126293375;
assign addr[55536]= 1093553126;
assign addr[55537]= 1060466036;
assign addr[55538]= 1027042599;
assign addr[55539]= 993293415;
assign addr[55540]= 959229189;
assign addr[55541]= 924860725;
assign addr[55542]= 890198924;
assign addr[55543]= 855254778;
assign addr[55544]= 820039373;
assign addr[55545]= 784563876;
assign addr[55546]= 748839539;
assign addr[55547]= 712877694;
assign addr[55548]= 676689746;
assign addr[55549]= 640287172;
assign addr[55550]= 603681519;
assign addr[55551]= 566884397;
assign addr[55552]= 529907477;
assign addr[55553]= 492762486;
assign addr[55554]= 455461206;
assign addr[55555]= 418015468;
assign addr[55556]= 380437148;
assign addr[55557]= 342738165;
assign addr[55558]= 304930476;
assign addr[55559]= 267026072;
assign addr[55560]= 229036977;
assign addr[55561]= 190975237;
assign addr[55562]= 152852926;
assign addr[55563]= 114682135;
assign addr[55564]= 76474970;
assign addr[55565]= 38243550;
assign addr[55566]= 0;
assign addr[55567]= -38243550;
assign addr[55568]= -76474970;
assign addr[55569]= -114682135;
assign addr[55570]= -152852926;
assign addr[55571]= -190975237;
assign addr[55572]= -229036977;
assign addr[55573]= -267026072;
assign addr[55574]= -304930476;
assign addr[55575]= -342738165;
assign addr[55576]= -380437148;
assign addr[55577]= -418015468;
assign addr[55578]= -455461206;
assign addr[55579]= -492762486;
assign addr[55580]= -529907477;
assign addr[55581]= -566884397;
assign addr[55582]= -603681519;
assign addr[55583]= -640287172;
assign addr[55584]= -676689746;
assign addr[55585]= -712877694;
assign addr[55586]= -748839539;
assign addr[55587]= -784563876;
assign addr[55588]= -820039373;
assign addr[55589]= -855254778;
assign addr[55590]= -890198924;
assign addr[55591]= -924860725;
assign addr[55592]= -959229189;
assign addr[55593]= -993293415;
assign addr[55594]= -1027042599;
assign addr[55595]= -1060466036;
assign addr[55596]= -1093553126;
assign addr[55597]= -1126293375;
assign addr[55598]= -1158676398;
assign addr[55599]= -1190691925;
assign addr[55600]= -1222329801;
assign addr[55601]= -1253579991;
assign addr[55602]= -1284432584;
assign addr[55603]= -1314877795;
assign addr[55604]= -1344905966;
assign addr[55605]= -1374507575;
assign addr[55606]= -1403673233;
assign addr[55607]= -1432393688;
assign addr[55608]= -1460659832;
assign addr[55609]= -1488462700;
assign addr[55610]= -1515793473;
assign addr[55611]= -1542643483;
assign addr[55612]= -1569004214;
assign addr[55613]= -1594867305;
assign addr[55614]= -1620224553;
assign addr[55615]= -1645067915;
assign addr[55616]= -1669389513;
assign addr[55617]= -1693181631;
assign addr[55618]= -1716436725;
assign addr[55619]= -1739147417;
assign addr[55620]= -1761306505;
assign addr[55621]= -1782906961;
assign addr[55622]= -1803941934;
assign addr[55623]= -1824404752;
assign addr[55624]= -1844288924;
assign addr[55625]= -1863588145;
assign addr[55626]= -1882296293;
assign addr[55627]= -1900407434;
assign addr[55628]= -1917915825;
assign addr[55629]= -1934815911;
assign addr[55630]= -1951102334;
assign addr[55631]= -1966769926;
assign addr[55632]= -1981813720;
assign addr[55633]= -1996228943;
assign addr[55634]= -2010011024;
assign addr[55635]= -2023155591;
assign addr[55636]= -2035658475;
assign addr[55637]= -2047515711;
assign addr[55638]= -2058723538;
assign addr[55639]= -2069278401;
assign addr[55640]= -2079176953;
assign addr[55641]= -2088416053;
assign addr[55642]= -2096992772;
assign addr[55643]= -2104904390;
assign addr[55644]= -2112148396;
assign addr[55645]= -2118722494;
assign addr[55646]= -2124624598;
assign addr[55647]= -2129852837;
assign addr[55648]= -2134405552;
assign addr[55649]= -2138281298;
assign addr[55650]= -2141478848;
assign addr[55651]= -2143997187;
assign addr[55652]= -2145835515;
assign addr[55653]= -2146993250;
assign addr[55654]= -2147470025;
assign addr[55655]= -2147265689;
assign addr[55656]= -2146380306;
assign addr[55657]= -2144814157;
assign addr[55658]= -2142567738;
assign addr[55659]= -2139641764;
assign addr[55660]= -2136037160;
assign addr[55661]= -2131755071;
assign addr[55662]= -2126796855;
assign addr[55663]= -2121164085;
assign addr[55664]= -2114858546;
assign addr[55665]= -2107882239;
assign addr[55666]= -2100237377;
assign addr[55667]= -2091926384;
assign addr[55668]= -2082951896;
assign addr[55669]= -2073316760;
assign addr[55670]= -2063024031;
assign addr[55671]= -2052076975;
assign addr[55672]= -2040479063;
assign addr[55673]= -2028233973;
assign addr[55674]= -2015345591;
assign addr[55675]= -2001818002;
assign addr[55676]= -1987655498;
assign addr[55677]= -1972862571;
assign addr[55678]= -1957443913;
assign addr[55679]= -1941404413;
assign addr[55680]= -1924749160;
assign addr[55681]= -1907483436;
assign addr[55682]= -1889612716;
assign addr[55683]= -1871142669;
assign addr[55684]= -1852079154;
assign addr[55685]= -1832428215;
assign addr[55686]= -1812196087;
assign addr[55687]= -1791389186;
assign addr[55688]= -1770014111;
assign addr[55689]= -1748077642;
assign addr[55690]= -1725586737;
assign addr[55691]= -1702548529;
assign addr[55692]= -1678970324;
assign addr[55693]= -1654859602;
assign addr[55694]= -1630224009;
assign addr[55695]= -1605071359;
assign addr[55696]= -1579409630;
assign addr[55697]= -1553246960;
assign addr[55698]= -1526591649;
assign addr[55699]= -1499452149;
assign addr[55700]= -1471837070;
assign addr[55701]= -1443755168;
assign addr[55702]= -1415215352;
assign addr[55703]= -1386226674;
assign addr[55704]= -1356798326;
assign addr[55705]= -1326939644;
assign addr[55706]= -1296660098;
assign addr[55707]= -1265969291;
assign addr[55708]= -1234876957;
assign addr[55709]= -1203392958;
assign addr[55710]= -1171527280;
assign addr[55711]= -1139290029;
assign addr[55712]= -1106691431;
assign addr[55713]= -1073741824;
assign addr[55714]= -1040451659;
assign addr[55715]= -1006831495;
assign addr[55716]= -972891995;
assign addr[55717]= -938643924;
assign addr[55718]= -904098143;
assign addr[55719]= -869265610;
assign addr[55720]= -834157373;
assign addr[55721]= -798784567;
assign addr[55722]= -763158411;
assign addr[55723]= -727290205;
assign addr[55724]= -691191324;
assign addr[55725]= -654873219;
assign addr[55726]= -618347408;
assign addr[55727]= -581625477;
assign addr[55728]= -544719071;
assign addr[55729]= -507639898;
assign addr[55730]= -470399716;
assign addr[55731]= -433010339;
assign addr[55732]= -395483624;
assign addr[55733]= -357831473;
assign addr[55734]= -320065829;
assign addr[55735]= -282198671;
assign addr[55736]= -244242007;
assign addr[55737]= -206207878;
assign addr[55738]= -168108346;
assign addr[55739]= -129955495;
assign addr[55740]= -91761426;
assign addr[55741]= -53538253;
assign addr[55742]= -15298099;
assign addr[55743]= 22946906;
assign addr[55744]= 61184634;
assign addr[55745]= 99402956;
assign addr[55746]= 137589750;
assign addr[55747]= 175732905;
assign addr[55748]= 213820322;
assign addr[55749]= 251839923;
assign addr[55750]= 289779648;
assign addr[55751]= 327627463;
assign addr[55752]= 365371365;
assign addr[55753]= 402999383;
assign addr[55754]= 440499581;
assign addr[55755]= 477860067;
assign addr[55756]= 515068990;
assign addr[55757]= 552114549;
assign addr[55758]= 588984994;
assign addr[55759]= 625668632;
assign addr[55760]= 662153826;
assign addr[55761]= 698429006;
assign addr[55762]= 734482665;
assign addr[55763]= 770303369;
assign addr[55764]= 805879757;
assign addr[55765]= 841200544;
assign addr[55766]= 876254528;
assign addr[55767]= 911030591;
assign addr[55768]= 945517704;
assign addr[55769]= 979704927;
assign addr[55770]= 1013581418;
assign addr[55771]= 1047136432;
assign addr[55772]= 1080359326;
assign addr[55773]= 1113239564;
assign addr[55774]= 1145766716;
assign addr[55775]= 1177930466;
assign addr[55776]= 1209720613;
assign addr[55777]= 1241127074;
assign addr[55778]= 1272139887;
assign addr[55779]= 1302749217;
assign addr[55780]= 1332945355;
assign addr[55781]= 1362718723;
assign addr[55782]= 1392059879;
assign addr[55783]= 1420959516;
assign addr[55784]= 1449408469;
assign addr[55785]= 1477397714;
assign addr[55786]= 1504918373;
assign addr[55787]= 1531961719;
assign addr[55788]= 1558519173;
assign addr[55789]= 1584582314;
assign addr[55790]= 1610142873;
assign addr[55791]= 1635192744;
assign addr[55792]= 1659723983;
assign addr[55793]= 1683728808;
assign addr[55794]= 1707199606;
assign addr[55795]= 1730128933;
assign addr[55796]= 1752509516;
assign addr[55797]= 1774334257;
assign addr[55798]= 1795596234;
assign addr[55799]= 1816288703;
assign addr[55800]= 1836405100;
assign addr[55801]= 1855939047;
assign addr[55802]= 1874884346;
assign addr[55803]= 1893234990;
assign addr[55804]= 1910985158;
assign addr[55805]= 1928129220;
assign addr[55806]= 1944661739;
assign addr[55807]= 1960577471;
assign addr[55808]= 1975871368;
assign addr[55809]= 1990538579;
assign addr[55810]= 2004574453;
assign addr[55811]= 2017974537;
assign addr[55812]= 2030734582;
assign addr[55813]= 2042850540;
assign addr[55814]= 2054318569;
assign addr[55815]= 2065135031;
assign addr[55816]= 2075296495;
assign addr[55817]= 2084799740;
assign addr[55818]= 2093641749;
assign addr[55819]= 2101819720;
assign addr[55820]= 2109331059;
assign addr[55821]= 2116173382;
assign addr[55822]= 2122344521;
assign addr[55823]= 2127842516;
assign addr[55824]= 2132665626;
assign addr[55825]= 2136812319;
assign addr[55826]= 2140281282;
assign addr[55827]= 2143071413;
assign addr[55828]= 2145181827;
assign addr[55829]= 2146611856;
assign addr[55830]= 2147361045;
assign addr[55831]= 2147429158;
assign addr[55832]= 2146816171;
assign addr[55833]= 2145522281;
assign addr[55834]= 2143547897;
assign addr[55835]= 2140893646;
assign addr[55836]= 2137560369;
assign addr[55837]= 2133549123;
assign addr[55838]= 2128861181;
assign addr[55839]= 2123498030;
assign addr[55840]= 2117461370;
assign addr[55841]= 2110753117;
assign addr[55842]= 2103375398;
assign addr[55843]= 2095330553;
assign addr[55844]= 2086621133;
assign addr[55845]= 2077249901;
assign addr[55846]= 2067219829;
assign addr[55847]= 2056534099;
assign addr[55848]= 2045196100;
assign addr[55849]= 2033209426;
assign addr[55850]= 2020577882;
assign addr[55851]= 2007305472;
assign addr[55852]= 1993396407;
assign addr[55853]= 1978855097;
assign addr[55854]= 1963686155;
assign addr[55855]= 1947894393;
assign addr[55856]= 1931484818;
assign addr[55857]= 1914462636;
assign addr[55858]= 1896833245;
assign addr[55859]= 1878602237;
assign addr[55860]= 1859775393;
assign addr[55861]= 1840358687;
assign addr[55862]= 1820358275;
assign addr[55863]= 1799780501;
assign addr[55864]= 1778631892;
assign addr[55865]= 1756919156;
assign addr[55866]= 1734649179;
assign addr[55867]= 1711829025;
assign addr[55868]= 1688465931;
assign addr[55869]= 1664567307;
assign addr[55870]= 1640140734;
assign addr[55871]= 1615193959;
assign addr[55872]= 1589734894;
assign addr[55873]= 1563771613;
assign addr[55874]= 1537312353;
assign addr[55875]= 1510365504;
assign addr[55876]= 1482939614;
assign addr[55877]= 1455043381;
assign addr[55878]= 1426685652;
assign addr[55879]= 1397875423;
assign addr[55880]= 1368621831;
assign addr[55881]= 1338934154;
assign addr[55882]= 1308821808;
assign addr[55883]= 1278294345;
assign addr[55884]= 1247361445;
assign addr[55885]= 1216032921;
assign addr[55886]= 1184318708;
assign addr[55887]= 1152228866;
assign addr[55888]= 1119773573;
assign addr[55889]= 1086963121;
assign addr[55890]= 1053807919;
assign addr[55891]= 1020318481;
assign addr[55892]= 986505429;
assign addr[55893]= 952379488;
assign addr[55894]= 917951481;
assign addr[55895]= 883232329;
assign addr[55896]= 848233042;
assign addr[55897]= 812964722;
assign addr[55898]= 777438554;
assign addr[55899]= 741665807;
assign addr[55900]= 705657826;
assign addr[55901]= 669426032;
assign addr[55902]= 632981917;
assign addr[55903]= 596337040;
assign addr[55904]= 559503022;
assign addr[55905]= 522491548;
assign addr[55906]= 485314355;
assign addr[55907]= 447983235;
assign addr[55908]= 410510029;
assign addr[55909]= 372906622;
assign addr[55910]= 335184940;
assign addr[55911]= 297356948;
assign addr[55912]= 259434643;
assign addr[55913]= 221430054;
assign addr[55914]= 183355234;
assign addr[55915]= 145222259;
assign addr[55916]= 107043224;
assign addr[55917]= 68830239;
assign addr[55918]= 30595422;
assign addr[55919]= -7649098;
assign addr[55920]= -45891193;
assign addr[55921]= -84118732;
assign addr[55922]= -122319591;
assign addr[55923]= -160481654;
assign addr[55924]= -198592817;
assign addr[55925]= -236640993;
assign addr[55926]= -274614114;
assign addr[55927]= -312500135;
assign addr[55928]= -350287041;
assign addr[55929]= -387962847;
assign addr[55930]= -425515602;
assign addr[55931]= -462933398;
assign addr[55932]= -500204365;
assign addr[55933]= -537316682;
assign addr[55934]= -574258580;
assign addr[55935]= -611018340;
assign addr[55936]= -647584304;
assign addr[55937]= -683944874;
assign addr[55938]= -720088517;
assign addr[55939]= -756003771;
assign addr[55940]= -791679244;
assign addr[55941]= -827103620;
assign addr[55942]= -862265664;
assign addr[55943]= -897154224;
assign addr[55944]= -931758235;
assign addr[55945]= -966066720;
assign addr[55946]= -1000068799;
assign addr[55947]= -1033753687;
assign addr[55948]= -1067110699;
assign addr[55949]= -1100129257;
assign addr[55950]= -1132798888;
assign addr[55951]= -1165109230;
assign addr[55952]= -1197050035;
assign addr[55953]= -1228611172;
assign addr[55954]= -1259782632;
assign addr[55955]= -1290554528;
assign addr[55956]= -1320917099;
assign addr[55957]= -1350860716;
assign addr[55958]= -1380375881;
assign addr[55959]= -1409453233;
assign addr[55960]= -1438083551;
assign addr[55961]= -1466257752;
assign addr[55962]= -1493966902;
assign addr[55963]= -1521202211;
assign addr[55964]= -1547955041;
assign addr[55965]= -1574216908;
assign addr[55966]= -1599979481;
assign addr[55967]= -1625234591;
assign addr[55968]= -1649974225;
assign addr[55969]= -1674190539;
assign addr[55970]= -1697875851;
assign addr[55971]= -1721022648;
assign addr[55972]= -1743623590;
assign addr[55973]= -1765671509;
assign addr[55974]= -1787159411;
assign addr[55975]= -1808080480;
assign addr[55976]= -1828428082;
assign addr[55977]= -1848195763;
assign addr[55978]= -1867377253;
assign addr[55979]= -1885966468;
assign addr[55980]= -1903957513;
assign addr[55981]= -1921344681;
assign addr[55982]= -1938122457;
assign addr[55983]= -1954285520;
assign addr[55984]= -1969828744;
assign addr[55985]= -1984747199;
assign addr[55986]= -1999036154;
assign addr[55987]= -2012691075;
assign addr[55988]= -2025707632;
assign addr[55989]= -2038081698;
assign addr[55990]= -2049809346;
assign addr[55991]= -2060886858;
assign addr[55992]= -2071310720;
assign addr[55993]= -2081077626;
assign addr[55994]= -2090184478;
assign addr[55995]= -2098628387;
assign addr[55996]= -2106406677;
assign addr[55997]= -2113516878;
assign addr[55998]= -2119956737;
assign addr[55999]= -2125724211;
assign addr[56000]= -2130817471;
assign addr[56001]= -2135234901;
assign addr[56002]= -2138975100;
assign addr[56003]= -2142036881;
assign addr[56004]= -2144419275;
assign addr[56005]= -2146121524;
assign addr[56006]= -2147143090;
assign addr[56007]= -2147483648;
assign addr[56008]= -2147143090;
assign addr[56009]= -2146121524;
assign addr[56010]= -2144419275;
assign addr[56011]= -2142036881;
assign addr[56012]= -2138975100;
assign addr[56013]= -2135234901;
assign addr[56014]= -2130817471;
assign addr[56015]= -2125724211;
assign addr[56016]= -2119956737;
assign addr[56017]= -2113516878;
assign addr[56018]= -2106406677;
assign addr[56019]= -2098628387;
assign addr[56020]= -2090184478;
assign addr[56021]= -2081077626;
assign addr[56022]= -2071310720;
assign addr[56023]= -2060886858;
assign addr[56024]= -2049809346;
assign addr[56025]= -2038081698;
assign addr[56026]= -2025707632;
assign addr[56027]= -2012691075;
assign addr[56028]= -1999036154;
assign addr[56029]= -1984747199;
assign addr[56030]= -1969828744;
assign addr[56031]= -1954285520;
assign addr[56032]= -1938122457;
assign addr[56033]= -1921344681;
assign addr[56034]= -1903957513;
assign addr[56035]= -1885966468;
assign addr[56036]= -1867377253;
assign addr[56037]= -1848195763;
assign addr[56038]= -1828428082;
assign addr[56039]= -1808080480;
assign addr[56040]= -1787159411;
assign addr[56041]= -1765671509;
assign addr[56042]= -1743623590;
assign addr[56043]= -1721022648;
assign addr[56044]= -1697875851;
assign addr[56045]= -1674190539;
assign addr[56046]= -1649974225;
assign addr[56047]= -1625234591;
assign addr[56048]= -1599979481;
assign addr[56049]= -1574216908;
assign addr[56050]= -1547955041;
assign addr[56051]= -1521202211;
assign addr[56052]= -1493966902;
assign addr[56053]= -1466257752;
assign addr[56054]= -1438083551;
assign addr[56055]= -1409453233;
assign addr[56056]= -1380375881;
assign addr[56057]= -1350860716;
assign addr[56058]= -1320917099;
assign addr[56059]= -1290554528;
assign addr[56060]= -1259782632;
assign addr[56061]= -1228611172;
assign addr[56062]= -1197050035;
assign addr[56063]= -1165109230;
assign addr[56064]= -1132798888;
assign addr[56065]= -1100129257;
assign addr[56066]= -1067110699;
assign addr[56067]= -1033753687;
assign addr[56068]= -1000068799;
assign addr[56069]= -966066720;
assign addr[56070]= -931758235;
assign addr[56071]= -897154224;
assign addr[56072]= -862265664;
assign addr[56073]= -827103620;
assign addr[56074]= -791679244;
assign addr[56075]= -756003771;
assign addr[56076]= -720088517;
assign addr[56077]= -683944874;
assign addr[56078]= -647584304;
assign addr[56079]= -611018340;
assign addr[56080]= -574258580;
assign addr[56081]= -537316682;
assign addr[56082]= -500204365;
assign addr[56083]= -462933398;
assign addr[56084]= -425515602;
assign addr[56085]= -387962847;
assign addr[56086]= -350287041;
assign addr[56087]= -312500135;
assign addr[56088]= -274614114;
assign addr[56089]= -236640993;
assign addr[56090]= -198592817;
assign addr[56091]= -160481654;
assign addr[56092]= -122319591;
assign addr[56093]= -84118732;
assign addr[56094]= -45891193;
assign addr[56095]= -7649098;
assign addr[56096]= 30595422;
assign addr[56097]= 68830239;
assign addr[56098]= 107043224;
assign addr[56099]= 145222259;
assign addr[56100]= 183355234;
assign addr[56101]= 221430054;
assign addr[56102]= 259434643;
assign addr[56103]= 297356948;
assign addr[56104]= 335184940;
assign addr[56105]= 372906622;
assign addr[56106]= 410510029;
assign addr[56107]= 447983235;
assign addr[56108]= 485314355;
assign addr[56109]= 522491548;
assign addr[56110]= 559503022;
assign addr[56111]= 596337040;
assign addr[56112]= 632981917;
assign addr[56113]= 669426032;
assign addr[56114]= 705657826;
assign addr[56115]= 741665807;
assign addr[56116]= 777438554;
assign addr[56117]= 812964722;
assign addr[56118]= 848233042;
assign addr[56119]= 883232329;
assign addr[56120]= 917951481;
assign addr[56121]= 952379488;
assign addr[56122]= 986505429;
assign addr[56123]= 1020318481;
assign addr[56124]= 1053807919;
assign addr[56125]= 1086963121;
assign addr[56126]= 1119773573;
assign addr[56127]= 1152228866;
assign addr[56128]= 1184318708;
assign addr[56129]= 1216032921;
assign addr[56130]= 1247361445;
assign addr[56131]= 1278294345;
assign addr[56132]= 1308821808;
assign addr[56133]= 1338934154;
assign addr[56134]= 1368621831;
assign addr[56135]= 1397875423;
assign addr[56136]= 1426685652;
assign addr[56137]= 1455043381;
assign addr[56138]= 1482939614;
assign addr[56139]= 1510365504;
assign addr[56140]= 1537312353;
assign addr[56141]= 1563771613;
assign addr[56142]= 1589734894;
assign addr[56143]= 1615193959;
assign addr[56144]= 1640140734;
assign addr[56145]= 1664567307;
assign addr[56146]= 1688465931;
assign addr[56147]= 1711829025;
assign addr[56148]= 1734649179;
assign addr[56149]= 1756919156;
assign addr[56150]= 1778631892;
assign addr[56151]= 1799780501;
assign addr[56152]= 1820358275;
assign addr[56153]= 1840358687;
assign addr[56154]= 1859775393;
assign addr[56155]= 1878602237;
assign addr[56156]= 1896833245;
assign addr[56157]= 1914462636;
assign addr[56158]= 1931484818;
assign addr[56159]= 1947894393;
assign addr[56160]= 1963686155;
assign addr[56161]= 1978855097;
assign addr[56162]= 1993396407;
assign addr[56163]= 2007305472;
assign addr[56164]= 2020577882;
assign addr[56165]= 2033209426;
assign addr[56166]= 2045196100;
assign addr[56167]= 2056534099;
assign addr[56168]= 2067219829;
assign addr[56169]= 2077249901;
assign addr[56170]= 2086621133;
assign addr[56171]= 2095330553;
assign addr[56172]= 2103375398;
assign addr[56173]= 2110753117;
assign addr[56174]= 2117461370;
assign addr[56175]= 2123498030;
assign addr[56176]= 2128861181;
assign addr[56177]= 2133549123;
assign addr[56178]= 2137560369;
assign addr[56179]= 2140893646;
assign addr[56180]= 2143547897;
assign addr[56181]= 2145522281;
assign addr[56182]= 2146816171;
assign addr[56183]= 2147429158;
assign addr[56184]= 2147361045;
assign addr[56185]= 2146611856;
assign addr[56186]= 2145181827;
assign addr[56187]= 2143071413;
assign addr[56188]= 2140281282;
assign addr[56189]= 2136812319;
assign addr[56190]= 2132665626;
assign addr[56191]= 2127842516;
assign addr[56192]= 2122344521;
assign addr[56193]= 2116173382;
assign addr[56194]= 2109331059;
assign addr[56195]= 2101819720;
assign addr[56196]= 2093641749;
assign addr[56197]= 2084799740;
assign addr[56198]= 2075296495;
assign addr[56199]= 2065135031;
assign addr[56200]= 2054318569;
assign addr[56201]= 2042850540;
assign addr[56202]= 2030734582;
assign addr[56203]= 2017974537;
assign addr[56204]= 2004574453;
assign addr[56205]= 1990538579;
assign addr[56206]= 1975871368;
assign addr[56207]= 1960577471;
assign addr[56208]= 1944661739;
assign addr[56209]= 1928129220;
assign addr[56210]= 1910985158;
assign addr[56211]= 1893234990;
assign addr[56212]= 1874884346;
assign addr[56213]= 1855939047;
assign addr[56214]= 1836405100;
assign addr[56215]= 1816288703;
assign addr[56216]= 1795596234;
assign addr[56217]= 1774334257;
assign addr[56218]= 1752509516;
assign addr[56219]= 1730128933;
assign addr[56220]= 1707199606;
assign addr[56221]= 1683728808;
assign addr[56222]= 1659723983;
assign addr[56223]= 1635192744;
assign addr[56224]= 1610142873;
assign addr[56225]= 1584582314;
assign addr[56226]= 1558519173;
assign addr[56227]= 1531961719;
assign addr[56228]= 1504918373;
assign addr[56229]= 1477397714;
assign addr[56230]= 1449408469;
assign addr[56231]= 1420959516;
assign addr[56232]= 1392059879;
assign addr[56233]= 1362718723;
assign addr[56234]= 1332945355;
assign addr[56235]= 1302749217;
assign addr[56236]= 1272139887;
assign addr[56237]= 1241127074;
assign addr[56238]= 1209720613;
assign addr[56239]= 1177930466;
assign addr[56240]= 1145766716;
assign addr[56241]= 1113239564;
assign addr[56242]= 1080359326;
assign addr[56243]= 1047136432;
assign addr[56244]= 1013581418;
assign addr[56245]= 979704927;
assign addr[56246]= 945517704;
assign addr[56247]= 911030591;
assign addr[56248]= 876254528;
assign addr[56249]= 841200544;
assign addr[56250]= 805879757;
assign addr[56251]= 770303369;
assign addr[56252]= 734482665;
assign addr[56253]= 698429006;
assign addr[56254]= 662153826;
assign addr[56255]= 625668632;
assign addr[56256]= 588984994;
assign addr[56257]= 552114549;
assign addr[56258]= 515068990;
assign addr[56259]= 477860067;
assign addr[56260]= 440499581;
assign addr[56261]= 402999383;
assign addr[56262]= 365371365;
assign addr[56263]= 327627463;
assign addr[56264]= 289779648;
assign addr[56265]= 251839923;
assign addr[56266]= 213820322;
assign addr[56267]= 175732905;
assign addr[56268]= 137589750;
assign addr[56269]= 99402956;
assign addr[56270]= 61184634;
assign addr[56271]= 22946906;
assign addr[56272]= -15298099;
assign addr[56273]= -53538253;
assign addr[56274]= -91761426;
assign addr[56275]= -129955495;
assign addr[56276]= -168108346;
assign addr[56277]= -206207878;
assign addr[56278]= -244242007;
assign addr[56279]= -282198671;
assign addr[56280]= -320065829;
assign addr[56281]= -357831473;
assign addr[56282]= -395483624;
assign addr[56283]= -433010339;
assign addr[56284]= -470399716;
assign addr[56285]= -507639898;
assign addr[56286]= -544719071;
assign addr[56287]= -581625477;
assign addr[56288]= -618347408;
assign addr[56289]= -654873219;
assign addr[56290]= -691191324;
assign addr[56291]= -727290205;
assign addr[56292]= -763158411;
assign addr[56293]= -798784567;
assign addr[56294]= -834157373;
assign addr[56295]= -869265610;
assign addr[56296]= -904098143;
assign addr[56297]= -938643924;
assign addr[56298]= -972891995;
assign addr[56299]= -1006831495;
assign addr[56300]= -1040451659;
assign addr[56301]= -1073741824;
assign addr[56302]= -1106691431;
assign addr[56303]= -1139290029;
assign addr[56304]= -1171527280;
assign addr[56305]= -1203392958;
assign addr[56306]= -1234876957;
assign addr[56307]= -1265969291;
assign addr[56308]= -1296660098;
assign addr[56309]= -1326939644;
assign addr[56310]= -1356798326;
assign addr[56311]= -1386226674;
assign addr[56312]= -1415215352;
assign addr[56313]= -1443755168;
assign addr[56314]= -1471837070;
assign addr[56315]= -1499452149;
assign addr[56316]= -1526591649;
assign addr[56317]= -1553246960;
assign addr[56318]= -1579409630;
assign addr[56319]= -1605071359;
assign addr[56320]= -1630224009;
assign addr[56321]= -1654859602;
assign addr[56322]= -1678970324;
assign addr[56323]= -1702548529;
assign addr[56324]= -1725586737;
assign addr[56325]= -1748077642;
assign addr[56326]= -1770014111;
assign addr[56327]= -1791389186;
assign addr[56328]= -1812196087;
assign addr[56329]= -1832428215;
assign addr[56330]= -1852079154;
assign addr[56331]= -1871142669;
assign addr[56332]= -1889612716;
assign addr[56333]= -1907483436;
assign addr[56334]= -1924749160;
assign addr[56335]= -1941404413;
assign addr[56336]= -1957443913;
assign addr[56337]= -1972862571;
assign addr[56338]= -1987655498;
assign addr[56339]= -2001818002;
assign addr[56340]= -2015345591;
assign addr[56341]= -2028233973;
assign addr[56342]= -2040479063;
assign addr[56343]= -2052076975;
assign addr[56344]= -2063024031;
assign addr[56345]= -2073316760;
assign addr[56346]= -2082951896;
assign addr[56347]= -2091926384;
assign addr[56348]= -2100237377;
assign addr[56349]= -2107882239;
assign addr[56350]= -2114858546;
assign addr[56351]= -2121164085;
assign addr[56352]= -2126796855;
assign addr[56353]= -2131755071;
assign addr[56354]= -2136037160;
assign addr[56355]= -2139641764;
assign addr[56356]= -2142567738;
assign addr[56357]= -2144814157;
assign addr[56358]= -2146380306;
assign addr[56359]= -2147265689;
assign addr[56360]= -2147470025;
assign addr[56361]= -2146993250;
assign addr[56362]= -2145835515;
assign addr[56363]= -2143997187;
assign addr[56364]= -2141478848;
assign addr[56365]= -2138281298;
assign addr[56366]= -2134405552;
assign addr[56367]= -2129852837;
assign addr[56368]= -2124624598;
assign addr[56369]= -2118722494;
assign addr[56370]= -2112148396;
assign addr[56371]= -2104904390;
assign addr[56372]= -2096992772;
assign addr[56373]= -2088416053;
assign addr[56374]= -2079176953;
assign addr[56375]= -2069278401;
assign addr[56376]= -2058723538;
assign addr[56377]= -2047515711;
assign addr[56378]= -2035658475;
assign addr[56379]= -2023155591;
assign addr[56380]= -2010011024;
assign addr[56381]= -1996228943;
assign addr[56382]= -1981813720;
assign addr[56383]= -1966769926;
assign addr[56384]= -1951102334;
assign addr[56385]= -1934815911;
assign addr[56386]= -1917915825;
assign addr[56387]= -1900407434;
assign addr[56388]= -1882296293;
assign addr[56389]= -1863588145;
assign addr[56390]= -1844288924;
assign addr[56391]= -1824404752;
assign addr[56392]= -1803941934;
assign addr[56393]= -1782906961;
assign addr[56394]= -1761306505;
assign addr[56395]= -1739147417;
assign addr[56396]= -1716436725;
assign addr[56397]= -1693181631;
assign addr[56398]= -1669389513;
assign addr[56399]= -1645067915;
assign addr[56400]= -1620224553;
assign addr[56401]= -1594867305;
assign addr[56402]= -1569004214;
assign addr[56403]= -1542643483;
assign addr[56404]= -1515793473;
assign addr[56405]= -1488462700;
assign addr[56406]= -1460659832;
assign addr[56407]= -1432393688;
assign addr[56408]= -1403673233;
assign addr[56409]= -1374507575;
assign addr[56410]= -1344905966;
assign addr[56411]= -1314877795;
assign addr[56412]= -1284432584;
assign addr[56413]= -1253579991;
assign addr[56414]= -1222329801;
assign addr[56415]= -1190691925;
assign addr[56416]= -1158676398;
assign addr[56417]= -1126293375;
assign addr[56418]= -1093553126;
assign addr[56419]= -1060466036;
assign addr[56420]= -1027042599;
assign addr[56421]= -993293415;
assign addr[56422]= -959229189;
assign addr[56423]= -924860725;
assign addr[56424]= -890198924;
assign addr[56425]= -855254778;
assign addr[56426]= -820039373;
assign addr[56427]= -784563876;
assign addr[56428]= -748839539;
assign addr[56429]= -712877694;
assign addr[56430]= -676689746;
assign addr[56431]= -640287172;
assign addr[56432]= -603681519;
assign addr[56433]= -566884397;
assign addr[56434]= -529907477;
assign addr[56435]= -492762486;
assign addr[56436]= -455461206;
assign addr[56437]= -418015468;
assign addr[56438]= -380437148;
assign addr[56439]= -342738165;
assign addr[56440]= -304930476;
assign addr[56441]= -267026072;
assign addr[56442]= -229036977;
assign addr[56443]= -190975237;
assign addr[56444]= -152852926;
assign addr[56445]= -114682135;
assign addr[56446]= -76474970;
assign addr[56447]= -38243550;
assign addr[56448]= 0;
assign addr[56449]= 38243550;
assign addr[56450]= 76474970;
assign addr[56451]= 114682135;
assign addr[56452]= 152852926;
assign addr[56453]= 190975237;
assign addr[56454]= 229036977;
assign addr[56455]= 267026072;
assign addr[56456]= 304930476;
assign addr[56457]= 342738165;
assign addr[56458]= 380437148;
assign addr[56459]= 418015468;
assign addr[56460]= 455461206;
assign addr[56461]= 492762486;
assign addr[56462]= 529907477;
assign addr[56463]= 566884397;
assign addr[56464]= 603681519;
assign addr[56465]= 640287172;
assign addr[56466]= 676689746;
assign addr[56467]= 712877694;
assign addr[56468]= 748839539;
assign addr[56469]= 784563876;
assign addr[56470]= 820039373;
assign addr[56471]= 855254778;
assign addr[56472]= 890198924;
assign addr[56473]= 924860725;
assign addr[56474]= 959229189;
assign addr[56475]= 993293415;
assign addr[56476]= 1027042599;
assign addr[56477]= 1060466036;
assign addr[56478]= 1093553126;
assign addr[56479]= 1126293375;
assign addr[56480]= 1158676398;
assign addr[56481]= 1190691925;
assign addr[56482]= 1222329801;
assign addr[56483]= 1253579991;
assign addr[56484]= 1284432584;
assign addr[56485]= 1314877795;
assign addr[56486]= 1344905966;
assign addr[56487]= 1374507575;
assign addr[56488]= 1403673233;
assign addr[56489]= 1432393688;
assign addr[56490]= 1460659832;
assign addr[56491]= 1488462700;
assign addr[56492]= 1515793473;
assign addr[56493]= 1542643483;
assign addr[56494]= 1569004214;
assign addr[56495]= 1594867305;
assign addr[56496]= 1620224553;
assign addr[56497]= 1645067915;
assign addr[56498]= 1669389513;
assign addr[56499]= 1693181631;
assign addr[56500]= 1716436725;
assign addr[56501]= 1739147417;
assign addr[56502]= 1761306505;
assign addr[56503]= 1782906961;
assign addr[56504]= 1803941934;
assign addr[56505]= 1824404752;
assign addr[56506]= 1844288924;
assign addr[56507]= 1863588145;
assign addr[56508]= 1882296293;
assign addr[56509]= 1900407434;
assign addr[56510]= 1917915825;
assign addr[56511]= 1934815911;
assign addr[56512]= 1951102334;
assign addr[56513]= 1966769926;
assign addr[56514]= 1981813720;
assign addr[56515]= 1996228943;
assign addr[56516]= 2010011024;
assign addr[56517]= 2023155591;
assign addr[56518]= 2035658475;
assign addr[56519]= 2047515711;
assign addr[56520]= 2058723538;
assign addr[56521]= 2069278401;
assign addr[56522]= 2079176953;
assign addr[56523]= 2088416053;
assign addr[56524]= 2096992772;
assign addr[56525]= 2104904390;
assign addr[56526]= 2112148396;
assign addr[56527]= 2118722494;
assign addr[56528]= 2124624598;
assign addr[56529]= 2129852837;
assign addr[56530]= 2134405552;
assign addr[56531]= 2138281298;
assign addr[56532]= 2141478848;
assign addr[56533]= 2143997187;
assign addr[56534]= 2145835515;
assign addr[56535]= 2146993250;
assign addr[56536]= 2147470025;
assign addr[56537]= 2147265689;
assign addr[56538]= 2146380306;
assign addr[56539]= 2144814157;
assign addr[56540]= 2142567738;
assign addr[56541]= 2139641764;
assign addr[56542]= 2136037160;
assign addr[56543]= 2131755071;
assign addr[56544]= 2126796855;
assign addr[56545]= 2121164085;
assign addr[56546]= 2114858546;
assign addr[56547]= 2107882239;
assign addr[56548]= 2100237377;
assign addr[56549]= 2091926384;
assign addr[56550]= 2082951896;
assign addr[56551]= 2073316760;
assign addr[56552]= 2063024031;
assign addr[56553]= 2052076975;
assign addr[56554]= 2040479063;
assign addr[56555]= 2028233973;
assign addr[56556]= 2015345591;
assign addr[56557]= 2001818002;
assign addr[56558]= 1987655498;
assign addr[56559]= 1972862571;
assign addr[56560]= 1957443913;
assign addr[56561]= 1941404413;
assign addr[56562]= 1924749160;
assign addr[56563]= 1907483436;
assign addr[56564]= 1889612716;
assign addr[56565]= 1871142669;
assign addr[56566]= 1852079154;
assign addr[56567]= 1832428215;
assign addr[56568]= 1812196087;
assign addr[56569]= 1791389186;
assign addr[56570]= 1770014111;
assign addr[56571]= 1748077642;
assign addr[56572]= 1725586737;
assign addr[56573]= 1702548529;
assign addr[56574]= 1678970324;
assign addr[56575]= 1654859602;
assign addr[56576]= 1630224009;
assign addr[56577]= 1605071359;
assign addr[56578]= 1579409630;
assign addr[56579]= 1553246960;
assign addr[56580]= 1526591649;
assign addr[56581]= 1499452149;
assign addr[56582]= 1471837070;
assign addr[56583]= 1443755168;
assign addr[56584]= 1415215352;
assign addr[56585]= 1386226674;
assign addr[56586]= 1356798326;
assign addr[56587]= 1326939644;
assign addr[56588]= 1296660098;
assign addr[56589]= 1265969291;
assign addr[56590]= 1234876957;
assign addr[56591]= 1203392958;
assign addr[56592]= 1171527280;
assign addr[56593]= 1139290029;
assign addr[56594]= 1106691431;
assign addr[56595]= 1073741824;
assign addr[56596]= 1040451659;
assign addr[56597]= 1006831495;
assign addr[56598]= 972891995;
assign addr[56599]= 938643924;
assign addr[56600]= 904098143;
assign addr[56601]= 869265610;
assign addr[56602]= 834157373;
assign addr[56603]= 798784567;
assign addr[56604]= 763158411;
assign addr[56605]= 727290205;
assign addr[56606]= 691191324;
assign addr[56607]= 654873219;
assign addr[56608]= 618347408;
assign addr[56609]= 581625477;
assign addr[56610]= 544719071;
assign addr[56611]= 507639898;
assign addr[56612]= 470399716;
assign addr[56613]= 433010339;
assign addr[56614]= 395483624;
assign addr[56615]= 357831473;
assign addr[56616]= 320065829;
assign addr[56617]= 282198671;
assign addr[56618]= 244242007;
assign addr[56619]= 206207878;
assign addr[56620]= 168108346;
assign addr[56621]= 129955495;
assign addr[56622]= 91761426;
assign addr[56623]= 53538253;
assign addr[56624]= 15298099;
assign addr[56625]= -22946906;
assign addr[56626]= -61184634;
assign addr[56627]= -99402956;
assign addr[56628]= -137589750;
assign addr[56629]= -175732905;
assign addr[56630]= -213820322;
assign addr[56631]= -251839923;
assign addr[56632]= -289779648;
assign addr[56633]= -327627463;
assign addr[56634]= -365371365;
assign addr[56635]= -402999383;
assign addr[56636]= -440499581;
assign addr[56637]= -477860067;
assign addr[56638]= -515068990;
assign addr[56639]= -552114549;
assign addr[56640]= -588984994;
assign addr[56641]= -625668632;
assign addr[56642]= -662153826;
assign addr[56643]= -698429006;
assign addr[56644]= -734482665;
assign addr[56645]= -770303369;
assign addr[56646]= -805879757;
assign addr[56647]= -841200544;
assign addr[56648]= -876254528;
assign addr[56649]= -911030591;
assign addr[56650]= -945517704;
assign addr[56651]= -979704927;
assign addr[56652]= -1013581418;
assign addr[56653]= -1047136432;
assign addr[56654]= -1080359326;
assign addr[56655]= -1113239564;
assign addr[56656]= -1145766716;
assign addr[56657]= -1177930466;
assign addr[56658]= -1209720613;
assign addr[56659]= -1241127074;
assign addr[56660]= -1272139887;
assign addr[56661]= -1302749217;
assign addr[56662]= -1332945355;
assign addr[56663]= -1362718723;
assign addr[56664]= -1392059879;
assign addr[56665]= -1420959516;
assign addr[56666]= -1449408469;
assign addr[56667]= -1477397714;
assign addr[56668]= -1504918373;
assign addr[56669]= -1531961719;
assign addr[56670]= -1558519173;
assign addr[56671]= -1584582314;
assign addr[56672]= -1610142873;
assign addr[56673]= -1635192744;
assign addr[56674]= -1659723983;
assign addr[56675]= -1683728808;
assign addr[56676]= -1707199606;
assign addr[56677]= -1730128933;
assign addr[56678]= -1752509516;
assign addr[56679]= -1774334257;
assign addr[56680]= -1795596234;
assign addr[56681]= -1816288703;
assign addr[56682]= -1836405100;
assign addr[56683]= -1855939047;
assign addr[56684]= -1874884346;
assign addr[56685]= -1893234990;
assign addr[56686]= -1910985158;
assign addr[56687]= -1928129220;
assign addr[56688]= -1944661739;
assign addr[56689]= -1960577471;
assign addr[56690]= -1975871368;
assign addr[56691]= -1990538579;
assign addr[56692]= -2004574453;
assign addr[56693]= -2017974537;
assign addr[56694]= -2030734582;
assign addr[56695]= -2042850540;
assign addr[56696]= -2054318569;
assign addr[56697]= -2065135031;
assign addr[56698]= -2075296495;
assign addr[56699]= -2084799740;
assign addr[56700]= -2093641749;
assign addr[56701]= -2101819720;
assign addr[56702]= -2109331059;
assign addr[56703]= -2116173382;
assign addr[56704]= -2122344521;
assign addr[56705]= -2127842516;
assign addr[56706]= -2132665626;
assign addr[56707]= -2136812319;
assign addr[56708]= -2140281282;
assign addr[56709]= -2143071413;
assign addr[56710]= -2145181827;
assign addr[56711]= -2146611856;
assign addr[56712]= -2147361045;
assign addr[56713]= -2147429158;
assign addr[56714]= -2146816171;
assign addr[56715]= -2145522281;
assign addr[56716]= -2143547897;
assign addr[56717]= -2140893646;
assign addr[56718]= -2137560369;
assign addr[56719]= -2133549123;
assign addr[56720]= -2128861181;
assign addr[56721]= -2123498030;
assign addr[56722]= -2117461370;
assign addr[56723]= -2110753117;
assign addr[56724]= -2103375398;
assign addr[56725]= -2095330553;
assign addr[56726]= -2086621133;
assign addr[56727]= -2077249901;
assign addr[56728]= -2067219829;
assign addr[56729]= -2056534099;
assign addr[56730]= -2045196100;
assign addr[56731]= -2033209426;
assign addr[56732]= -2020577882;
assign addr[56733]= -2007305472;
assign addr[56734]= -1993396407;
assign addr[56735]= -1978855097;
assign addr[56736]= -1963686155;
assign addr[56737]= -1947894393;
assign addr[56738]= -1931484818;
assign addr[56739]= -1914462636;
assign addr[56740]= -1896833245;
assign addr[56741]= -1878602237;
assign addr[56742]= -1859775393;
assign addr[56743]= -1840358687;
assign addr[56744]= -1820358275;
assign addr[56745]= -1799780501;
assign addr[56746]= -1778631892;
assign addr[56747]= -1756919156;
assign addr[56748]= -1734649179;
assign addr[56749]= -1711829025;
assign addr[56750]= -1688465931;
assign addr[56751]= -1664567307;
assign addr[56752]= -1640140734;
assign addr[56753]= -1615193959;
assign addr[56754]= -1589734894;
assign addr[56755]= -1563771613;
assign addr[56756]= -1537312353;
assign addr[56757]= -1510365504;
assign addr[56758]= -1482939614;
assign addr[56759]= -1455043381;
assign addr[56760]= -1426685652;
assign addr[56761]= -1397875423;
assign addr[56762]= -1368621831;
assign addr[56763]= -1338934154;
assign addr[56764]= -1308821808;
assign addr[56765]= -1278294345;
assign addr[56766]= -1247361445;
assign addr[56767]= -1216032921;
assign addr[56768]= -1184318708;
assign addr[56769]= -1152228866;
assign addr[56770]= -1119773573;
assign addr[56771]= -1086963121;
assign addr[56772]= -1053807919;
assign addr[56773]= -1020318481;
assign addr[56774]= -986505429;
assign addr[56775]= -952379488;
assign addr[56776]= -917951481;
assign addr[56777]= -883232329;
assign addr[56778]= -848233042;
assign addr[56779]= -812964722;
assign addr[56780]= -777438554;
assign addr[56781]= -741665807;
assign addr[56782]= -705657826;
assign addr[56783]= -669426032;
assign addr[56784]= -632981917;
assign addr[56785]= -596337040;
assign addr[56786]= -559503022;
assign addr[56787]= -522491548;
assign addr[56788]= -485314355;
assign addr[56789]= -447983235;
assign addr[56790]= -410510029;
assign addr[56791]= -372906622;
assign addr[56792]= -335184940;
assign addr[56793]= -297356948;
assign addr[56794]= -259434643;
assign addr[56795]= -221430054;
assign addr[56796]= -183355234;
assign addr[56797]= -145222259;
assign addr[56798]= -107043224;
assign addr[56799]= -68830239;
assign addr[56800]= -30595422;
assign addr[56801]= 7649098;
assign addr[56802]= 45891193;
assign addr[56803]= 84118732;
assign addr[56804]= 122319591;
assign addr[56805]= 160481654;
assign addr[56806]= 198592817;
assign addr[56807]= 236640993;
assign addr[56808]= 274614114;
assign addr[56809]= 312500135;
assign addr[56810]= 350287041;
assign addr[56811]= 387962847;
assign addr[56812]= 425515602;
assign addr[56813]= 462933398;
assign addr[56814]= 500204365;
assign addr[56815]= 537316682;
assign addr[56816]= 574258580;
assign addr[56817]= 611018340;
assign addr[56818]= 647584304;
assign addr[56819]= 683944874;
assign addr[56820]= 720088517;
assign addr[56821]= 756003771;
assign addr[56822]= 791679244;
assign addr[56823]= 827103620;
assign addr[56824]= 862265664;
assign addr[56825]= 897154224;
assign addr[56826]= 931758235;
assign addr[56827]= 966066720;
assign addr[56828]= 1000068799;
assign addr[56829]= 1033753687;
assign addr[56830]= 1067110699;
assign addr[56831]= 1100129257;
assign addr[56832]= 1132798888;
assign addr[56833]= 1165109230;
assign addr[56834]= 1197050035;
assign addr[56835]= 1228611172;
assign addr[56836]= 1259782632;
assign addr[56837]= 1290554528;
assign addr[56838]= 1320917099;
assign addr[56839]= 1350860716;
assign addr[56840]= 1380375881;
assign addr[56841]= 1409453233;
assign addr[56842]= 1438083551;
assign addr[56843]= 1466257752;
assign addr[56844]= 1493966902;
assign addr[56845]= 1521202211;
assign addr[56846]= 1547955041;
assign addr[56847]= 1574216908;
assign addr[56848]= 1599979481;
assign addr[56849]= 1625234591;
assign addr[56850]= 1649974225;
assign addr[56851]= 1674190539;
assign addr[56852]= 1697875851;
assign addr[56853]= 1721022648;
assign addr[56854]= 1743623590;
assign addr[56855]= 1765671509;
assign addr[56856]= 1787159411;
assign addr[56857]= 1808080480;
assign addr[56858]= 1828428082;
assign addr[56859]= 1848195763;
assign addr[56860]= 1867377253;
assign addr[56861]= 1885966468;
assign addr[56862]= 1903957513;
assign addr[56863]= 1921344681;
assign addr[56864]= 1938122457;
assign addr[56865]= 1954285520;
assign addr[56866]= 1969828744;
assign addr[56867]= 1984747199;
assign addr[56868]= 1999036154;
assign addr[56869]= 2012691075;
assign addr[56870]= 2025707632;
assign addr[56871]= 2038081698;
assign addr[56872]= 2049809346;
assign addr[56873]= 2060886858;
assign addr[56874]= 2071310720;
assign addr[56875]= 2081077626;
assign addr[56876]= 2090184478;
assign addr[56877]= 2098628387;
assign addr[56878]= 2106406677;
assign addr[56879]= 2113516878;
assign addr[56880]= 2119956737;
assign addr[56881]= 2125724211;
assign addr[56882]= 2130817471;
assign addr[56883]= 2135234901;
assign addr[56884]= 2138975100;
assign addr[56885]= 2142036881;
assign addr[56886]= 2144419275;
assign addr[56887]= 2146121524;
assign addr[56888]= 2147143090;
assign addr[56889]= 2147483648;
assign addr[56890]= 2147143090;
assign addr[56891]= 2146121524;
assign addr[56892]= 2144419275;
assign addr[56893]= 2142036881;
assign addr[56894]= 2138975100;
assign addr[56895]= 2135234901;
assign addr[56896]= 2130817471;
assign addr[56897]= 2125724211;
assign addr[56898]= 2119956737;
assign addr[56899]= 2113516878;
assign addr[56900]= 2106406677;
assign addr[56901]= 2098628387;
assign addr[56902]= 2090184478;
assign addr[56903]= 2081077626;
assign addr[56904]= 2071310720;
assign addr[56905]= 2060886858;
assign addr[56906]= 2049809346;
assign addr[56907]= 2038081698;
assign addr[56908]= 2025707632;
assign addr[56909]= 2012691075;
assign addr[56910]= 1999036154;
assign addr[56911]= 1984747199;
assign addr[56912]= 1969828744;
assign addr[56913]= 1954285520;
assign addr[56914]= 1938122457;
assign addr[56915]= 1921344681;
assign addr[56916]= 1903957513;
assign addr[56917]= 1885966468;
assign addr[56918]= 1867377253;
assign addr[56919]= 1848195763;
assign addr[56920]= 1828428082;
assign addr[56921]= 1808080480;
assign addr[56922]= 1787159411;
assign addr[56923]= 1765671509;
assign addr[56924]= 1743623590;
assign addr[56925]= 1721022648;
assign addr[56926]= 1697875851;
assign addr[56927]= 1674190539;
assign addr[56928]= 1649974225;
assign addr[56929]= 1625234591;
assign addr[56930]= 1599979481;
assign addr[56931]= 1574216908;
assign addr[56932]= 1547955041;
assign addr[56933]= 1521202211;
assign addr[56934]= 1493966902;
assign addr[56935]= 1466257752;
assign addr[56936]= 1438083551;
assign addr[56937]= 1409453233;
assign addr[56938]= 1380375881;
assign addr[56939]= 1350860716;
assign addr[56940]= 1320917099;
assign addr[56941]= 1290554528;
assign addr[56942]= 1259782632;
assign addr[56943]= 1228611172;
assign addr[56944]= 1197050035;
assign addr[56945]= 1165109230;
assign addr[56946]= 1132798888;
assign addr[56947]= 1100129257;
assign addr[56948]= 1067110699;
assign addr[56949]= 1033753687;
assign addr[56950]= 1000068799;
assign addr[56951]= 966066720;
assign addr[56952]= 931758235;
assign addr[56953]= 897154224;
assign addr[56954]= 862265664;
assign addr[56955]= 827103620;
assign addr[56956]= 791679244;
assign addr[56957]= 756003771;
assign addr[56958]= 720088517;
assign addr[56959]= 683944874;
assign addr[56960]= 647584304;
assign addr[56961]= 611018340;
assign addr[56962]= 574258580;
assign addr[56963]= 537316682;
assign addr[56964]= 500204365;
assign addr[56965]= 462933398;
assign addr[56966]= 425515602;
assign addr[56967]= 387962847;
assign addr[56968]= 350287041;
assign addr[56969]= 312500135;
assign addr[56970]= 274614114;
assign addr[56971]= 236640993;
assign addr[56972]= 198592817;
assign addr[56973]= 160481654;
assign addr[56974]= 122319591;
assign addr[56975]= 84118732;
assign addr[56976]= 45891193;
assign addr[56977]= 7649098;
assign addr[56978]= -30595422;
assign addr[56979]= -68830239;
assign addr[56980]= -107043224;
assign addr[56981]= -145222259;
assign addr[56982]= -183355234;
assign addr[56983]= -221430054;
assign addr[56984]= -259434643;
assign addr[56985]= -297356948;
assign addr[56986]= -335184940;
assign addr[56987]= -372906622;
assign addr[56988]= -410510029;
assign addr[56989]= -447983235;
assign addr[56990]= -485314355;
assign addr[56991]= -522491548;
assign addr[56992]= -559503022;
assign addr[56993]= -596337040;
assign addr[56994]= -632981917;
assign addr[56995]= -669426032;
assign addr[56996]= -705657826;
assign addr[56997]= -741665807;
assign addr[56998]= -777438554;
assign addr[56999]= -812964722;
assign addr[57000]= -848233042;
assign addr[57001]= -883232329;
assign addr[57002]= -917951481;
assign addr[57003]= -952379488;
assign addr[57004]= -986505429;
assign addr[57005]= -1020318481;
assign addr[57006]= -1053807919;
assign addr[57007]= -1086963121;
assign addr[57008]= -1119773573;
assign addr[57009]= -1152228866;
assign addr[57010]= -1184318708;
assign addr[57011]= -1216032921;
assign addr[57012]= -1247361445;
assign addr[57013]= -1278294345;
assign addr[57014]= -1308821808;
assign addr[57015]= -1338934154;
assign addr[57016]= -1368621831;
assign addr[57017]= -1397875423;
assign addr[57018]= -1426685652;
assign addr[57019]= -1455043381;
assign addr[57020]= -1482939614;
assign addr[57021]= -1510365504;
assign addr[57022]= -1537312353;
assign addr[57023]= -1563771613;
assign addr[57024]= -1589734894;
assign addr[57025]= -1615193959;
assign addr[57026]= -1640140734;
assign addr[57027]= -1664567307;
assign addr[57028]= -1688465931;
assign addr[57029]= -1711829025;
assign addr[57030]= -1734649179;
assign addr[57031]= -1756919156;
assign addr[57032]= -1778631892;
assign addr[57033]= -1799780501;
assign addr[57034]= -1820358275;
assign addr[57035]= -1840358687;
assign addr[57036]= -1859775393;
assign addr[57037]= -1878602237;
assign addr[57038]= -1896833245;
assign addr[57039]= -1914462636;
assign addr[57040]= -1931484818;
assign addr[57041]= -1947894393;
assign addr[57042]= -1963686155;
assign addr[57043]= -1978855097;
assign addr[57044]= -1993396407;
assign addr[57045]= -2007305472;
assign addr[57046]= -2020577882;
assign addr[57047]= -2033209426;
assign addr[57048]= -2045196100;
assign addr[57049]= -2056534099;
assign addr[57050]= -2067219829;
assign addr[57051]= -2077249901;
assign addr[57052]= -2086621133;
assign addr[57053]= -2095330553;
assign addr[57054]= -2103375398;
assign addr[57055]= -2110753117;
assign addr[57056]= -2117461370;
assign addr[57057]= -2123498030;
assign addr[57058]= -2128861181;
assign addr[57059]= -2133549123;
assign addr[57060]= -2137560369;
assign addr[57061]= -2140893646;
assign addr[57062]= -2143547897;
assign addr[57063]= -2145522281;
assign addr[57064]= -2146816171;
assign addr[57065]= -2147429158;
assign addr[57066]= -2147361045;
assign addr[57067]= -2146611856;
assign addr[57068]= -2145181827;
assign addr[57069]= -2143071413;
assign addr[57070]= -2140281282;
assign addr[57071]= -2136812319;
assign addr[57072]= -2132665626;
assign addr[57073]= -2127842516;
assign addr[57074]= -2122344521;
assign addr[57075]= -2116173382;
assign addr[57076]= -2109331059;
assign addr[57077]= -2101819720;
assign addr[57078]= -2093641749;
assign addr[57079]= -2084799740;
assign addr[57080]= -2075296495;
assign addr[57081]= -2065135031;
assign addr[57082]= -2054318569;
assign addr[57083]= -2042850540;
assign addr[57084]= -2030734582;
assign addr[57085]= -2017974537;
assign addr[57086]= -2004574453;
assign addr[57087]= -1990538579;
assign addr[57088]= -1975871368;
assign addr[57089]= -1960577471;
assign addr[57090]= -1944661739;
assign addr[57091]= -1928129220;
assign addr[57092]= -1910985158;
assign addr[57093]= -1893234990;
assign addr[57094]= -1874884346;
assign addr[57095]= -1855939047;
assign addr[57096]= -1836405100;
assign addr[57097]= -1816288703;
assign addr[57098]= -1795596234;
assign addr[57099]= -1774334257;
assign addr[57100]= -1752509516;
assign addr[57101]= -1730128933;
assign addr[57102]= -1707199606;
assign addr[57103]= -1683728808;
assign addr[57104]= -1659723983;
assign addr[57105]= -1635192744;
assign addr[57106]= -1610142873;
assign addr[57107]= -1584582314;
assign addr[57108]= -1558519173;
assign addr[57109]= -1531961719;
assign addr[57110]= -1504918373;
assign addr[57111]= -1477397714;
assign addr[57112]= -1449408469;
assign addr[57113]= -1420959516;
assign addr[57114]= -1392059879;
assign addr[57115]= -1362718723;
assign addr[57116]= -1332945355;
assign addr[57117]= -1302749217;
assign addr[57118]= -1272139887;
assign addr[57119]= -1241127074;
assign addr[57120]= -1209720613;
assign addr[57121]= -1177930466;
assign addr[57122]= -1145766716;
assign addr[57123]= -1113239564;
assign addr[57124]= -1080359326;
assign addr[57125]= -1047136432;
assign addr[57126]= -1013581418;
assign addr[57127]= -979704927;
assign addr[57128]= -945517704;
assign addr[57129]= -911030591;
assign addr[57130]= -876254528;
assign addr[57131]= -841200544;
assign addr[57132]= -805879757;
assign addr[57133]= -770303369;
assign addr[57134]= -734482665;
assign addr[57135]= -698429006;
assign addr[57136]= -662153826;
assign addr[57137]= -625668632;
assign addr[57138]= -588984994;
assign addr[57139]= -552114549;
assign addr[57140]= -515068990;
assign addr[57141]= -477860067;
assign addr[57142]= -440499581;
assign addr[57143]= -402999383;
assign addr[57144]= -365371365;
assign addr[57145]= -327627463;
assign addr[57146]= -289779648;
assign addr[57147]= -251839923;
assign addr[57148]= -213820322;
assign addr[57149]= -175732905;
assign addr[57150]= -137589750;
assign addr[57151]= -99402956;
assign addr[57152]= -61184634;
assign addr[57153]= -22946906;
assign addr[57154]= 15298099;
assign addr[57155]= 53538253;
assign addr[57156]= 91761426;
assign addr[57157]= 129955495;
assign addr[57158]= 168108346;
assign addr[57159]= 206207878;
assign addr[57160]= 244242007;
assign addr[57161]= 282198671;
assign addr[57162]= 320065829;
assign addr[57163]= 357831473;
assign addr[57164]= 395483624;
assign addr[57165]= 433010339;
assign addr[57166]= 470399716;
assign addr[57167]= 507639898;
assign addr[57168]= 544719071;
assign addr[57169]= 581625477;
assign addr[57170]= 618347408;
assign addr[57171]= 654873219;
assign addr[57172]= 691191324;
assign addr[57173]= 727290205;
assign addr[57174]= 763158411;
assign addr[57175]= 798784567;
assign addr[57176]= 834157373;
assign addr[57177]= 869265610;
assign addr[57178]= 904098143;
assign addr[57179]= 938643924;
assign addr[57180]= 972891995;
assign addr[57181]= 1006831495;
assign addr[57182]= 1040451659;
assign addr[57183]= 1073741824;
assign addr[57184]= 1106691431;
assign addr[57185]= 1139290029;
assign addr[57186]= 1171527280;
assign addr[57187]= 1203392958;
assign addr[57188]= 1234876957;
assign addr[57189]= 1265969291;
assign addr[57190]= 1296660098;
assign addr[57191]= 1326939644;
assign addr[57192]= 1356798326;
assign addr[57193]= 1386226674;
assign addr[57194]= 1415215352;
assign addr[57195]= 1443755168;
assign addr[57196]= 1471837070;
assign addr[57197]= 1499452149;
assign addr[57198]= 1526591649;
assign addr[57199]= 1553246960;
assign addr[57200]= 1579409630;
assign addr[57201]= 1605071359;
assign addr[57202]= 1630224009;
assign addr[57203]= 1654859602;
assign addr[57204]= 1678970324;
assign addr[57205]= 1702548529;
assign addr[57206]= 1725586737;
assign addr[57207]= 1748077642;
assign addr[57208]= 1770014111;
assign addr[57209]= 1791389186;
assign addr[57210]= 1812196087;
assign addr[57211]= 1832428215;
assign addr[57212]= 1852079154;
assign addr[57213]= 1871142669;
assign addr[57214]= 1889612716;
assign addr[57215]= 1907483436;
assign addr[57216]= 1924749160;
assign addr[57217]= 1941404413;
assign addr[57218]= 1957443913;
assign addr[57219]= 1972862571;
assign addr[57220]= 1987655498;
assign addr[57221]= 2001818002;
assign addr[57222]= 2015345591;
assign addr[57223]= 2028233973;
assign addr[57224]= 2040479063;
assign addr[57225]= 2052076975;
assign addr[57226]= 2063024031;
assign addr[57227]= 2073316760;
assign addr[57228]= 2082951896;
assign addr[57229]= 2091926384;
assign addr[57230]= 2100237377;
assign addr[57231]= 2107882239;
assign addr[57232]= 2114858546;
assign addr[57233]= 2121164085;
assign addr[57234]= 2126796855;
assign addr[57235]= 2131755071;
assign addr[57236]= 2136037160;
assign addr[57237]= 2139641764;
assign addr[57238]= 2142567738;
assign addr[57239]= 2144814157;
assign addr[57240]= 2146380306;
assign addr[57241]= 2147265689;
assign addr[57242]= 2147470025;
assign addr[57243]= 2146993250;
assign addr[57244]= 2145835515;
assign addr[57245]= 2143997187;
assign addr[57246]= 2141478848;
assign addr[57247]= 2138281298;
assign addr[57248]= 2134405552;
assign addr[57249]= 2129852837;
assign addr[57250]= 2124624598;
assign addr[57251]= 2118722494;
assign addr[57252]= 2112148396;
assign addr[57253]= 2104904390;
assign addr[57254]= 2096992772;
assign addr[57255]= 2088416053;
assign addr[57256]= 2079176953;
assign addr[57257]= 2069278401;
assign addr[57258]= 2058723538;
assign addr[57259]= 2047515711;
assign addr[57260]= 2035658475;
assign addr[57261]= 2023155591;
assign addr[57262]= 2010011024;
assign addr[57263]= 1996228943;
assign addr[57264]= 1981813720;
assign addr[57265]= 1966769926;
assign addr[57266]= 1951102334;
assign addr[57267]= 1934815911;
assign addr[57268]= 1917915825;
assign addr[57269]= 1900407434;
assign addr[57270]= 1882296293;
assign addr[57271]= 1863588145;
assign addr[57272]= 1844288924;
assign addr[57273]= 1824404752;
assign addr[57274]= 1803941934;
assign addr[57275]= 1782906961;
assign addr[57276]= 1761306505;
assign addr[57277]= 1739147417;
assign addr[57278]= 1716436725;
assign addr[57279]= 1693181631;
assign addr[57280]= 1669389513;
assign addr[57281]= 1645067915;
assign addr[57282]= 1620224553;
assign addr[57283]= 1594867305;
assign addr[57284]= 1569004214;
assign addr[57285]= 1542643483;
assign addr[57286]= 1515793473;
assign addr[57287]= 1488462700;
assign addr[57288]= 1460659832;
assign addr[57289]= 1432393688;
assign addr[57290]= 1403673233;
assign addr[57291]= 1374507575;
assign addr[57292]= 1344905966;
assign addr[57293]= 1314877795;
assign addr[57294]= 1284432584;
assign addr[57295]= 1253579991;
assign addr[57296]= 1222329801;
assign addr[57297]= 1190691925;
assign addr[57298]= 1158676398;
assign addr[57299]= 1126293375;
assign addr[57300]= 1093553126;
assign addr[57301]= 1060466036;
assign addr[57302]= 1027042599;
assign addr[57303]= 993293415;
assign addr[57304]= 959229189;
assign addr[57305]= 924860725;
assign addr[57306]= 890198924;
assign addr[57307]= 855254778;
assign addr[57308]= 820039373;
assign addr[57309]= 784563876;
assign addr[57310]= 748839539;
assign addr[57311]= 712877694;
assign addr[57312]= 676689746;
assign addr[57313]= 640287172;
assign addr[57314]= 603681519;
assign addr[57315]= 566884397;
assign addr[57316]= 529907477;
assign addr[57317]= 492762486;
assign addr[57318]= 455461206;
assign addr[57319]= 418015468;
assign addr[57320]= 380437148;
assign addr[57321]= 342738165;
assign addr[57322]= 304930476;
assign addr[57323]= 267026072;
assign addr[57324]= 229036977;
assign addr[57325]= 190975237;
assign addr[57326]= 152852926;
assign addr[57327]= 114682135;
assign addr[57328]= 76474970;
assign addr[57329]= 38243550;
assign addr[57330]= 0;
assign addr[57331]= -38243550;
assign addr[57332]= -76474970;
assign addr[57333]= -114682135;
assign addr[57334]= -152852926;
assign addr[57335]= -190975237;
assign addr[57336]= -229036977;
assign addr[57337]= -267026072;
assign addr[57338]= -304930476;
assign addr[57339]= -342738165;
assign addr[57340]= -380437148;
assign addr[57341]= -418015468;
assign addr[57342]= -455461206;
assign addr[57343]= -492762486;
assign addr[57344]= -529907477;
assign addr[57345]= -566884397;
assign addr[57346]= -603681519;
assign addr[57347]= -640287172;
assign addr[57348]= -676689746;
assign addr[57349]= -712877694;
assign addr[57350]= -748839539;
assign addr[57351]= -784563876;
assign addr[57352]= -820039373;
assign addr[57353]= -855254778;
assign addr[57354]= -890198924;
assign addr[57355]= -924860725;
assign addr[57356]= -959229189;
assign addr[57357]= -993293415;
assign addr[57358]= -1027042599;
assign addr[57359]= -1060466036;
assign addr[57360]= -1093553126;
assign addr[57361]= -1126293375;
assign addr[57362]= -1158676398;
assign addr[57363]= -1190691925;
assign addr[57364]= -1222329801;
assign addr[57365]= -1253579991;
assign addr[57366]= -1284432584;
assign addr[57367]= -1314877795;
assign addr[57368]= -1344905966;
assign addr[57369]= -1374507575;
assign addr[57370]= -1403673233;
assign addr[57371]= -1432393688;
assign addr[57372]= -1460659832;
assign addr[57373]= -1488462700;
assign addr[57374]= -1515793473;
assign addr[57375]= -1542643483;
assign addr[57376]= -1569004214;
assign addr[57377]= -1594867305;
assign addr[57378]= -1620224553;
assign addr[57379]= -1645067915;
assign addr[57380]= -1669389513;
assign addr[57381]= -1693181631;
assign addr[57382]= -1716436725;
assign addr[57383]= -1739147417;
assign addr[57384]= -1761306505;
assign addr[57385]= -1782906961;
assign addr[57386]= -1803941934;
assign addr[57387]= -1824404752;
assign addr[57388]= -1844288924;
assign addr[57389]= -1863588145;
assign addr[57390]= -1882296293;
assign addr[57391]= -1900407434;
assign addr[57392]= -1917915825;
assign addr[57393]= -1934815911;
assign addr[57394]= -1951102334;
assign addr[57395]= -1966769926;
assign addr[57396]= -1981813720;
assign addr[57397]= -1996228943;
assign addr[57398]= -2010011024;
assign addr[57399]= -2023155591;
assign addr[57400]= -2035658475;
assign addr[57401]= -2047515711;
assign addr[57402]= -2058723538;
assign addr[57403]= -2069278401;
assign addr[57404]= -2079176953;
assign addr[57405]= -2088416053;
assign addr[57406]= -2096992772;
assign addr[57407]= -2104904390;
assign addr[57408]= -2112148396;
assign addr[57409]= -2118722494;
assign addr[57410]= -2124624598;
assign addr[57411]= -2129852837;
assign addr[57412]= -2134405552;
assign addr[57413]= -2138281298;
assign addr[57414]= -2141478848;
assign addr[57415]= -2143997187;
assign addr[57416]= -2145835515;
assign addr[57417]= -2146993250;
assign addr[57418]= -2147470025;
assign addr[57419]= -2147265689;
assign addr[57420]= -2146380306;
assign addr[57421]= -2144814157;
assign addr[57422]= -2142567738;
assign addr[57423]= -2139641764;
assign addr[57424]= -2136037160;
assign addr[57425]= -2131755071;
assign addr[57426]= -2126796855;
assign addr[57427]= -2121164085;
assign addr[57428]= -2114858546;
assign addr[57429]= -2107882239;
assign addr[57430]= -2100237377;
assign addr[57431]= -2091926384;
assign addr[57432]= -2082951896;
assign addr[57433]= -2073316760;
assign addr[57434]= -2063024031;
assign addr[57435]= -2052076975;
assign addr[57436]= -2040479063;
assign addr[57437]= -2028233973;
assign addr[57438]= -2015345591;
assign addr[57439]= -2001818002;
assign addr[57440]= -1987655498;
assign addr[57441]= -1972862571;
assign addr[57442]= -1957443913;
assign addr[57443]= -1941404413;
assign addr[57444]= -1924749160;
assign addr[57445]= -1907483436;
assign addr[57446]= -1889612716;
assign addr[57447]= -1871142669;
assign addr[57448]= -1852079154;
assign addr[57449]= -1832428215;
assign addr[57450]= -1812196087;
assign addr[57451]= -1791389186;
assign addr[57452]= -1770014111;
assign addr[57453]= -1748077642;
assign addr[57454]= -1725586737;
assign addr[57455]= -1702548529;
assign addr[57456]= -1678970324;
assign addr[57457]= -1654859602;
assign addr[57458]= -1630224009;
assign addr[57459]= -1605071359;
assign addr[57460]= -1579409630;
assign addr[57461]= -1553246960;
assign addr[57462]= -1526591649;
assign addr[57463]= -1499452149;
assign addr[57464]= -1471837070;
assign addr[57465]= -1443755168;
assign addr[57466]= -1415215352;
assign addr[57467]= -1386226674;
assign addr[57468]= -1356798326;
assign addr[57469]= -1326939644;
assign addr[57470]= -1296660098;
assign addr[57471]= -1265969291;
assign addr[57472]= -1234876957;
assign addr[57473]= -1203392958;
assign addr[57474]= -1171527280;
assign addr[57475]= -1139290029;
assign addr[57476]= -1106691431;
assign addr[57477]= -1073741824;
assign addr[57478]= -1040451659;
assign addr[57479]= -1006831495;
assign addr[57480]= -972891995;
assign addr[57481]= -938643924;
assign addr[57482]= -904098143;
assign addr[57483]= -869265610;
assign addr[57484]= -834157373;
assign addr[57485]= -798784567;
assign addr[57486]= -763158411;
assign addr[57487]= -727290205;
assign addr[57488]= -691191324;
assign addr[57489]= -654873219;
assign addr[57490]= -618347408;
assign addr[57491]= -581625477;
assign addr[57492]= -544719071;
assign addr[57493]= -507639898;
assign addr[57494]= -470399716;
assign addr[57495]= -433010339;
assign addr[57496]= -395483624;
assign addr[57497]= -357831473;
assign addr[57498]= -320065829;
assign addr[57499]= -282198671;
assign addr[57500]= -244242007;
assign addr[57501]= -206207878;
assign addr[57502]= -168108346;
assign addr[57503]= -129955495;
assign addr[57504]= -91761426;
assign addr[57505]= -53538253;
assign addr[57506]= -15298099;
assign addr[57507]= 22946906;
assign addr[57508]= 61184634;
assign addr[57509]= 99402956;
assign addr[57510]= 137589750;
assign addr[57511]= 175732905;
assign addr[57512]= 213820322;
assign addr[57513]= 251839923;
assign addr[57514]= 289779648;
assign addr[57515]= 327627463;
assign addr[57516]= 365371365;
assign addr[57517]= 402999383;
assign addr[57518]= 440499581;
assign addr[57519]= 477860067;
assign addr[57520]= 515068990;
assign addr[57521]= 552114549;
assign addr[57522]= 588984994;
assign addr[57523]= 625668632;
assign addr[57524]= 662153826;
assign addr[57525]= 698429006;
assign addr[57526]= 734482665;
assign addr[57527]= 770303369;
assign addr[57528]= 805879757;
assign addr[57529]= 841200544;
assign addr[57530]= 876254528;
assign addr[57531]= 911030591;
assign addr[57532]= 945517704;
assign addr[57533]= 979704927;
assign addr[57534]= 1013581418;
assign addr[57535]= 1047136432;
assign addr[57536]= 1080359326;
assign addr[57537]= 1113239564;
assign addr[57538]= 1145766716;
assign addr[57539]= 1177930466;
assign addr[57540]= 1209720613;
assign addr[57541]= 1241127074;
assign addr[57542]= 1272139887;
assign addr[57543]= 1302749217;
assign addr[57544]= 1332945355;
assign addr[57545]= 1362718723;
assign addr[57546]= 1392059879;
assign addr[57547]= 1420959516;
assign addr[57548]= 1449408469;
assign addr[57549]= 1477397714;
assign addr[57550]= 1504918373;
assign addr[57551]= 1531961719;
assign addr[57552]= 1558519173;
assign addr[57553]= 1584582314;
assign addr[57554]= 1610142873;
assign addr[57555]= 1635192744;
assign addr[57556]= 1659723983;
assign addr[57557]= 1683728808;
assign addr[57558]= 1707199606;
assign addr[57559]= 1730128933;
assign addr[57560]= 1752509516;
assign addr[57561]= 1774334257;
assign addr[57562]= 1795596234;
assign addr[57563]= 1816288703;
assign addr[57564]= 1836405100;
assign addr[57565]= 1855939047;
assign addr[57566]= 1874884346;
assign addr[57567]= 1893234990;
assign addr[57568]= 1910985158;
assign addr[57569]= 1928129220;
assign addr[57570]= 1944661739;
assign addr[57571]= 1960577471;
assign addr[57572]= 1975871368;
assign addr[57573]= 1990538579;
assign addr[57574]= 2004574453;
assign addr[57575]= 2017974537;
assign addr[57576]= 2030734582;
assign addr[57577]= 2042850540;
assign addr[57578]= 2054318569;
assign addr[57579]= 2065135031;
assign addr[57580]= 2075296495;
assign addr[57581]= 2084799740;
assign addr[57582]= 2093641749;
assign addr[57583]= 2101819720;
assign addr[57584]= 2109331059;
assign addr[57585]= 2116173382;
assign addr[57586]= 2122344521;
assign addr[57587]= 2127842516;
assign addr[57588]= 2132665626;
assign addr[57589]= 2136812319;
assign addr[57590]= 2140281282;
assign addr[57591]= 2143071413;
assign addr[57592]= 2145181827;
assign addr[57593]= 2146611856;
assign addr[57594]= 2147361045;
assign addr[57595]= 2147429158;
assign addr[57596]= 2146816171;
assign addr[57597]= 2145522281;
assign addr[57598]= 2143547897;
assign addr[57599]= 2140893646;
assign addr[57600]= 2137560369;
assign addr[57601]= 2133549123;
assign addr[57602]= 2128861181;
assign addr[57603]= 2123498030;
assign addr[57604]= 2117461370;
assign addr[57605]= 2110753117;
assign addr[57606]= 2103375398;
assign addr[57607]= 2095330553;
assign addr[57608]= 2086621133;
assign addr[57609]= 2077249901;
assign addr[57610]= 2067219829;
assign addr[57611]= 2056534099;
assign addr[57612]= 2045196100;
assign addr[57613]= 2033209426;
assign addr[57614]= 2020577882;
assign addr[57615]= 2007305472;
assign addr[57616]= 1993396407;
assign addr[57617]= 1978855097;
assign addr[57618]= 1963686155;
assign addr[57619]= 1947894393;
assign addr[57620]= 1931484818;
assign addr[57621]= 1914462636;
assign addr[57622]= 1896833245;
assign addr[57623]= 1878602237;
assign addr[57624]= 1859775393;
assign addr[57625]= 1840358687;
assign addr[57626]= 1820358275;
assign addr[57627]= 1799780501;
assign addr[57628]= 1778631892;
assign addr[57629]= 1756919156;
assign addr[57630]= 1734649179;
assign addr[57631]= 1711829025;
assign addr[57632]= 1688465931;
assign addr[57633]= 1664567307;
assign addr[57634]= 1640140734;
assign addr[57635]= 1615193959;
assign addr[57636]= 1589734894;
assign addr[57637]= 1563771613;
assign addr[57638]= 1537312353;
assign addr[57639]= 1510365504;
assign addr[57640]= 1482939614;
assign addr[57641]= 1455043381;
assign addr[57642]= 1426685652;
assign addr[57643]= 1397875423;
assign addr[57644]= 1368621831;
assign addr[57645]= 1338934154;
assign addr[57646]= 1308821808;
assign addr[57647]= 1278294345;
assign addr[57648]= 1247361445;
assign addr[57649]= 1216032921;
assign addr[57650]= 1184318708;
assign addr[57651]= 1152228866;
assign addr[57652]= 1119773573;
assign addr[57653]= 1086963121;
assign addr[57654]= 1053807919;
assign addr[57655]= 1020318481;
assign addr[57656]= 986505429;
assign addr[57657]= 952379488;
assign addr[57658]= 917951481;
assign addr[57659]= 883232329;
assign addr[57660]= 848233042;
assign addr[57661]= 812964722;
assign addr[57662]= 777438554;
assign addr[57663]= 741665807;
assign addr[57664]= 705657826;
assign addr[57665]= 669426032;
assign addr[57666]= 632981917;
assign addr[57667]= 596337040;
assign addr[57668]= 559503022;
assign addr[57669]= 522491548;
assign addr[57670]= 485314355;
assign addr[57671]= 447983235;
assign addr[57672]= 410510029;
assign addr[57673]= 372906622;
assign addr[57674]= 335184940;
assign addr[57675]= 297356948;
assign addr[57676]= 259434643;
assign addr[57677]= 221430054;
assign addr[57678]= 183355234;
assign addr[57679]= 145222259;
assign addr[57680]= 107043224;
assign addr[57681]= 68830239;
assign addr[57682]= 30595422;
assign addr[57683]= -7649098;
assign addr[57684]= -45891193;
assign addr[57685]= -84118732;
assign addr[57686]= -122319591;
assign addr[57687]= -160481654;
assign addr[57688]= -198592817;
assign addr[57689]= -236640993;
assign addr[57690]= -274614114;
assign addr[57691]= -312500135;
assign addr[57692]= -350287041;
assign addr[57693]= -387962847;
assign addr[57694]= -425515602;
assign addr[57695]= -462933398;
assign addr[57696]= -500204365;
assign addr[57697]= -537316682;
assign addr[57698]= -574258580;
assign addr[57699]= -611018340;
assign addr[57700]= -647584304;
assign addr[57701]= -683944874;
assign addr[57702]= -720088517;
assign addr[57703]= -756003771;
assign addr[57704]= -791679244;
assign addr[57705]= -827103620;
assign addr[57706]= -862265664;
assign addr[57707]= -897154224;
assign addr[57708]= -931758235;
assign addr[57709]= -966066720;
assign addr[57710]= -1000068799;
assign addr[57711]= -1033753687;
assign addr[57712]= -1067110699;
assign addr[57713]= -1100129257;
assign addr[57714]= -1132798888;
assign addr[57715]= -1165109230;
assign addr[57716]= -1197050035;
assign addr[57717]= -1228611172;
assign addr[57718]= -1259782632;
assign addr[57719]= -1290554528;
assign addr[57720]= -1320917099;
assign addr[57721]= -1350860716;
assign addr[57722]= -1380375881;
assign addr[57723]= -1409453233;
assign addr[57724]= -1438083551;
assign addr[57725]= -1466257752;
assign addr[57726]= -1493966902;
assign addr[57727]= -1521202211;
assign addr[57728]= -1547955041;
assign addr[57729]= -1574216908;
assign addr[57730]= -1599979481;
assign addr[57731]= -1625234591;
assign addr[57732]= -1649974225;
assign addr[57733]= -1674190539;
assign addr[57734]= -1697875851;
assign addr[57735]= -1721022648;
assign addr[57736]= -1743623590;
assign addr[57737]= -1765671509;
assign addr[57738]= -1787159411;
assign addr[57739]= -1808080480;
assign addr[57740]= -1828428082;
assign addr[57741]= -1848195763;
assign addr[57742]= -1867377253;
assign addr[57743]= -1885966468;
assign addr[57744]= -1903957513;
assign addr[57745]= -1921344681;
assign addr[57746]= -1938122457;
assign addr[57747]= -1954285520;
assign addr[57748]= -1969828744;
assign addr[57749]= -1984747199;
assign addr[57750]= -1999036154;
assign addr[57751]= -2012691075;
assign addr[57752]= -2025707632;
assign addr[57753]= -2038081698;
assign addr[57754]= -2049809346;
assign addr[57755]= -2060886858;
assign addr[57756]= -2071310720;
assign addr[57757]= -2081077626;
assign addr[57758]= -2090184478;
assign addr[57759]= -2098628387;
assign addr[57760]= -2106406677;
assign addr[57761]= -2113516878;
assign addr[57762]= -2119956737;
assign addr[57763]= -2125724211;
assign addr[57764]= -2130817471;
assign addr[57765]= -2135234901;
assign addr[57766]= -2138975100;
assign addr[57767]= -2142036881;
assign addr[57768]= -2144419275;
assign addr[57769]= -2146121524;
assign addr[57770]= -2147143090;
assign addr[57771]= -2147483648;
assign addr[57772]= -2147143090;
assign addr[57773]= -2146121524;
assign addr[57774]= -2144419275;
assign addr[57775]= -2142036881;
assign addr[57776]= -2138975100;
assign addr[57777]= -2135234901;
assign addr[57778]= -2130817471;
assign addr[57779]= -2125724211;
assign addr[57780]= -2119956737;
assign addr[57781]= -2113516878;
assign addr[57782]= -2106406677;
assign addr[57783]= -2098628387;
assign addr[57784]= -2090184478;
assign addr[57785]= -2081077626;
assign addr[57786]= -2071310720;
assign addr[57787]= -2060886858;
assign addr[57788]= -2049809346;
assign addr[57789]= -2038081698;
assign addr[57790]= -2025707632;
assign addr[57791]= -2012691075;
assign addr[57792]= -1999036154;
assign addr[57793]= -1984747199;
assign addr[57794]= -1969828744;
assign addr[57795]= -1954285520;
assign addr[57796]= -1938122457;
assign addr[57797]= -1921344681;
assign addr[57798]= -1903957513;
assign addr[57799]= -1885966468;
assign addr[57800]= -1867377253;
assign addr[57801]= -1848195763;
assign addr[57802]= -1828428082;
assign addr[57803]= -1808080480;
assign addr[57804]= -1787159411;
assign addr[57805]= -1765671509;
assign addr[57806]= -1743623590;
assign addr[57807]= -1721022648;
assign addr[57808]= -1697875851;
assign addr[57809]= -1674190539;
assign addr[57810]= -1649974225;
assign addr[57811]= -1625234591;
assign addr[57812]= -1599979481;
assign addr[57813]= -1574216908;
assign addr[57814]= -1547955041;
assign addr[57815]= -1521202211;
assign addr[57816]= -1493966902;
assign addr[57817]= -1466257752;
assign addr[57818]= -1438083551;
assign addr[57819]= -1409453233;
assign addr[57820]= -1380375881;
assign addr[57821]= -1350860716;
assign addr[57822]= -1320917099;
assign addr[57823]= -1290554528;
assign addr[57824]= -1259782632;
assign addr[57825]= -1228611172;
assign addr[57826]= -1197050035;
assign addr[57827]= -1165109230;
assign addr[57828]= -1132798888;
assign addr[57829]= -1100129257;
assign addr[57830]= -1067110699;
assign addr[57831]= -1033753687;
assign addr[57832]= -1000068799;
assign addr[57833]= -966066720;
assign addr[57834]= -931758235;
assign addr[57835]= -897154224;
assign addr[57836]= -862265664;
assign addr[57837]= -827103620;
assign addr[57838]= -791679244;
assign addr[57839]= -756003771;
assign addr[57840]= -720088517;
assign addr[57841]= -683944874;
assign addr[57842]= -647584304;
assign addr[57843]= -611018340;
assign addr[57844]= -574258580;
assign addr[57845]= -537316682;
assign addr[57846]= -500204365;
assign addr[57847]= -462933398;
assign addr[57848]= -425515602;
assign addr[57849]= -387962847;
assign addr[57850]= -350287041;
assign addr[57851]= -312500135;
assign addr[57852]= -274614114;
assign addr[57853]= -236640993;
assign addr[57854]= -198592817;
assign addr[57855]= -160481654;
assign addr[57856]= -122319591;
assign addr[57857]= -84118732;
assign addr[57858]= -45891193;
assign addr[57859]= -7649098;
assign addr[57860]= 30595422;
assign addr[57861]= 68830239;
assign addr[57862]= 107043224;
assign addr[57863]= 145222259;
assign addr[57864]= 183355234;
assign addr[57865]= 221430054;
assign addr[57866]= 259434643;
assign addr[57867]= 297356948;
assign addr[57868]= 335184940;
assign addr[57869]= 372906622;
assign addr[57870]= 410510029;
assign addr[57871]= 447983235;
assign addr[57872]= 485314355;
assign addr[57873]= 522491548;
assign addr[57874]= 559503022;
assign addr[57875]= 596337040;
assign addr[57876]= 632981917;
assign addr[57877]= 669426032;
assign addr[57878]= 705657826;
assign addr[57879]= 741665807;
assign addr[57880]= 777438554;
assign addr[57881]= 812964722;
assign addr[57882]= 848233042;
assign addr[57883]= 883232329;
assign addr[57884]= 917951481;
assign addr[57885]= 952379488;
assign addr[57886]= 986505429;
assign addr[57887]= 1020318481;
assign addr[57888]= 1053807919;
assign addr[57889]= 1086963121;
assign addr[57890]= 1119773573;
assign addr[57891]= 1152228866;
assign addr[57892]= 1184318708;
assign addr[57893]= 1216032921;
assign addr[57894]= 1247361445;
assign addr[57895]= 1278294345;
assign addr[57896]= 1308821808;
assign addr[57897]= 1338934154;
assign addr[57898]= 1368621831;
assign addr[57899]= 1397875423;
assign addr[57900]= 1426685652;
assign addr[57901]= 1455043381;
assign addr[57902]= 1482939614;
assign addr[57903]= 1510365504;
assign addr[57904]= 1537312353;
assign addr[57905]= 1563771613;
assign addr[57906]= 1589734894;
assign addr[57907]= 1615193959;
assign addr[57908]= 1640140734;
assign addr[57909]= 1664567307;
assign addr[57910]= 1688465931;
assign addr[57911]= 1711829025;
assign addr[57912]= 1734649179;
assign addr[57913]= 1756919156;
assign addr[57914]= 1778631892;
assign addr[57915]= 1799780501;
assign addr[57916]= 1820358275;
assign addr[57917]= 1840358687;
assign addr[57918]= 1859775393;
assign addr[57919]= 1878602237;
assign addr[57920]= 1896833245;
assign addr[57921]= 1914462636;
assign addr[57922]= 1931484818;
assign addr[57923]= 1947894393;
assign addr[57924]= 1963686155;
assign addr[57925]= 1978855097;
assign addr[57926]= 1993396407;
assign addr[57927]= 2007305472;
assign addr[57928]= 2020577882;
assign addr[57929]= 2033209426;
assign addr[57930]= 2045196100;
assign addr[57931]= 2056534099;
assign addr[57932]= 2067219829;
assign addr[57933]= 2077249901;
assign addr[57934]= 2086621133;
assign addr[57935]= 2095330553;
assign addr[57936]= 2103375398;
assign addr[57937]= 2110753117;
assign addr[57938]= 2117461370;
assign addr[57939]= 2123498030;
assign addr[57940]= 2128861181;
assign addr[57941]= 2133549123;
assign addr[57942]= 2137560369;
assign addr[57943]= 2140893646;
assign addr[57944]= 2143547897;
assign addr[57945]= 2145522281;
assign addr[57946]= 2146816171;
assign addr[57947]= 2147429158;
assign addr[57948]= 2147361045;
assign addr[57949]= 2146611856;
assign addr[57950]= 2145181827;
assign addr[57951]= 2143071413;
assign addr[57952]= 2140281282;
assign addr[57953]= 2136812319;
assign addr[57954]= 2132665626;
assign addr[57955]= 2127842516;
assign addr[57956]= 2122344521;
assign addr[57957]= 2116173382;
assign addr[57958]= 2109331059;
assign addr[57959]= 2101819720;
assign addr[57960]= 2093641749;
assign addr[57961]= 2084799740;
assign addr[57962]= 2075296495;
assign addr[57963]= 2065135031;
assign addr[57964]= 2054318569;
assign addr[57965]= 2042850540;
assign addr[57966]= 2030734582;
assign addr[57967]= 2017974537;
assign addr[57968]= 2004574453;
assign addr[57969]= 1990538579;
assign addr[57970]= 1975871368;
assign addr[57971]= 1960577471;
assign addr[57972]= 1944661739;
assign addr[57973]= 1928129220;
assign addr[57974]= 1910985158;
assign addr[57975]= 1893234990;
assign addr[57976]= 1874884346;
assign addr[57977]= 1855939047;
assign addr[57978]= 1836405100;
assign addr[57979]= 1816288703;
assign addr[57980]= 1795596234;
assign addr[57981]= 1774334257;
assign addr[57982]= 1752509516;
assign addr[57983]= 1730128933;
assign addr[57984]= 1707199606;
assign addr[57985]= 1683728808;
assign addr[57986]= 1659723983;
assign addr[57987]= 1635192744;
assign addr[57988]= 1610142873;
assign addr[57989]= 1584582314;
assign addr[57990]= 1558519173;
assign addr[57991]= 1531961719;
assign addr[57992]= 1504918373;
assign addr[57993]= 1477397714;
assign addr[57994]= 1449408469;
assign addr[57995]= 1420959516;
assign addr[57996]= 1392059879;
assign addr[57997]= 1362718723;
assign addr[57998]= 1332945355;
assign addr[57999]= 1302749217;
assign addr[58000]= 1272139887;
assign addr[58001]= 1241127074;
assign addr[58002]= 1209720613;
assign addr[58003]= 1177930466;
assign addr[58004]= 1145766716;
assign addr[58005]= 1113239564;
assign addr[58006]= 1080359326;
assign addr[58007]= 1047136432;
assign addr[58008]= 1013581418;
assign addr[58009]= 979704927;
assign addr[58010]= 945517704;
assign addr[58011]= 911030591;
assign addr[58012]= 876254528;
assign addr[58013]= 841200544;
assign addr[58014]= 805879757;
assign addr[58015]= 770303369;
assign addr[58016]= 734482665;
assign addr[58017]= 698429006;
assign addr[58018]= 662153826;
assign addr[58019]= 625668632;
assign addr[58020]= 588984994;
assign addr[58021]= 552114549;
assign addr[58022]= 515068990;
assign addr[58023]= 477860067;
assign addr[58024]= 440499581;
assign addr[58025]= 402999383;
assign addr[58026]= 365371365;
assign addr[58027]= 327627463;
assign addr[58028]= 289779648;
assign addr[58029]= 251839923;
assign addr[58030]= 213820322;
assign addr[58031]= 175732905;
assign addr[58032]= 137589750;
assign addr[58033]= 99402956;
assign addr[58034]= 61184634;
assign addr[58035]= 22946906;
assign addr[58036]= -15298099;
assign addr[58037]= -53538253;
assign addr[58038]= -91761426;
assign addr[58039]= -129955495;
assign addr[58040]= -168108346;
assign addr[58041]= -206207878;
assign addr[58042]= -244242007;
assign addr[58043]= -282198671;
assign addr[58044]= -320065829;
assign addr[58045]= -357831473;
assign addr[58046]= -395483624;
assign addr[58047]= -433010339;
assign addr[58048]= -470399716;
assign addr[58049]= -507639898;
assign addr[58050]= -544719071;
assign addr[58051]= -581625477;
assign addr[58052]= -618347408;
assign addr[58053]= -654873219;
assign addr[58054]= -691191324;
assign addr[58055]= -727290205;
assign addr[58056]= -763158411;
assign addr[58057]= -798784567;
assign addr[58058]= -834157373;
assign addr[58059]= -869265610;
assign addr[58060]= -904098143;
assign addr[58061]= -938643924;
assign addr[58062]= -972891995;
assign addr[58063]= -1006831495;
assign addr[58064]= -1040451659;
assign addr[58065]= -1073741824;
assign addr[58066]= -1106691431;
assign addr[58067]= -1139290029;
assign addr[58068]= -1171527280;
assign addr[58069]= -1203392958;
assign addr[58070]= -1234876957;
assign addr[58071]= -1265969291;
assign addr[58072]= -1296660098;
assign addr[58073]= -1326939644;
assign addr[58074]= -1356798326;
assign addr[58075]= -1386226674;
assign addr[58076]= -1415215352;
assign addr[58077]= -1443755168;
assign addr[58078]= -1471837070;
assign addr[58079]= -1499452149;
assign addr[58080]= -1526591649;
assign addr[58081]= -1553246960;
assign addr[58082]= -1579409630;
assign addr[58083]= -1605071359;
assign addr[58084]= -1630224009;
assign addr[58085]= -1654859602;
assign addr[58086]= -1678970324;
assign addr[58087]= -1702548529;
assign addr[58088]= -1725586737;
assign addr[58089]= -1748077642;
assign addr[58090]= -1770014111;
assign addr[58091]= -1791389186;
assign addr[58092]= -1812196087;
assign addr[58093]= -1832428215;
assign addr[58094]= -1852079154;
assign addr[58095]= -1871142669;
assign addr[58096]= -1889612716;
assign addr[58097]= -1907483436;
assign addr[58098]= -1924749160;
assign addr[58099]= -1941404413;
assign addr[58100]= -1957443913;
assign addr[58101]= -1972862571;
assign addr[58102]= -1987655498;
assign addr[58103]= -2001818002;
assign addr[58104]= -2015345591;
assign addr[58105]= -2028233973;
assign addr[58106]= -2040479063;
assign addr[58107]= -2052076975;
assign addr[58108]= -2063024031;
assign addr[58109]= -2073316760;
assign addr[58110]= -2082951896;
assign addr[58111]= -2091926384;
assign addr[58112]= -2100237377;
assign addr[58113]= -2107882239;
assign addr[58114]= -2114858546;
assign addr[58115]= -2121164085;
assign addr[58116]= -2126796855;
assign addr[58117]= -2131755071;
assign addr[58118]= -2136037160;
assign addr[58119]= -2139641764;
assign addr[58120]= -2142567738;
assign addr[58121]= -2144814157;
assign addr[58122]= -2146380306;
assign addr[58123]= -2147265689;
assign addr[58124]= -2147470025;
assign addr[58125]= -2146993250;
assign addr[58126]= -2145835515;
assign addr[58127]= -2143997187;
assign addr[58128]= -2141478848;
assign addr[58129]= -2138281298;
assign addr[58130]= -2134405552;
assign addr[58131]= -2129852837;
assign addr[58132]= -2124624598;
assign addr[58133]= -2118722494;
assign addr[58134]= -2112148396;
assign addr[58135]= -2104904390;
assign addr[58136]= -2096992772;
assign addr[58137]= -2088416053;
assign addr[58138]= -2079176953;
assign addr[58139]= -2069278401;
assign addr[58140]= -2058723538;
assign addr[58141]= -2047515711;
assign addr[58142]= -2035658475;
assign addr[58143]= -2023155591;
assign addr[58144]= -2010011024;
assign addr[58145]= -1996228943;
assign addr[58146]= -1981813720;
assign addr[58147]= -1966769926;
assign addr[58148]= -1951102334;
assign addr[58149]= -1934815911;
assign addr[58150]= -1917915825;
assign addr[58151]= -1900407434;
assign addr[58152]= -1882296293;
assign addr[58153]= -1863588145;
assign addr[58154]= -1844288924;
assign addr[58155]= -1824404752;
assign addr[58156]= -1803941934;
assign addr[58157]= -1782906961;
assign addr[58158]= -1761306505;
assign addr[58159]= -1739147417;
assign addr[58160]= -1716436725;
assign addr[58161]= -1693181631;
assign addr[58162]= -1669389513;
assign addr[58163]= -1645067915;
assign addr[58164]= -1620224553;
assign addr[58165]= -1594867305;
assign addr[58166]= -1569004214;
assign addr[58167]= -1542643483;
assign addr[58168]= -1515793473;
assign addr[58169]= -1488462700;
assign addr[58170]= -1460659832;
assign addr[58171]= -1432393688;
assign addr[58172]= -1403673233;
assign addr[58173]= -1374507575;
assign addr[58174]= -1344905966;
assign addr[58175]= -1314877795;
assign addr[58176]= -1284432584;
assign addr[58177]= -1253579991;
assign addr[58178]= -1222329801;
assign addr[58179]= -1190691925;
assign addr[58180]= -1158676398;
assign addr[58181]= -1126293375;
assign addr[58182]= -1093553126;
assign addr[58183]= -1060466036;
assign addr[58184]= -1027042599;
assign addr[58185]= -993293415;
assign addr[58186]= -959229189;
assign addr[58187]= -924860725;
assign addr[58188]= -890198924;
assign addr[58189]= -855254778;
assign addr[58190]= -820039373;
assign addr[58191]= -784563876;
assign addr[58192]= -748839539;
assign addr[58193]= -712877694;
assign addr[58194]= -676689746;
assign addr[58195]= -640287172;
assign addr[58196]= -603681519;
assign addr[58197]= -566884397;
assign addr[58198]= -529907477;
assign addr[58199]= -492762486;
assign addr[58200]= -455461206;
assign addr[58201]= -418015468;
assign addr[58202]= -380437148;
assign addr[58203]= -342738165;
assign addr[58204]= -304930476;
assign addr[58205]= -267026072;
assign addr[58206]= -229036977;
assign addr[58207]= -190975237;
assign addr[58208]= -152852926;
assign addr[58209]= -114682135;
assign addr[58210]= -76474970;
assign addr[58211]= -38243550;
assign addr[58212]= 0;
assign addr[58213]= 38243550;
assign addr[58214]= 76474970;
assign addr[58215]= 114682135;
assign addr[58216]= 152852926;
assign addr[58217]= 190975237;
assign addr[58218]= 229036977;
assign addr[58219]= 267026072;
assign addr[58220]= 304930476;
assign addr[58221]= 342738165;
assign addr[58222]= 380437148;
assign addr[58223]= 418015468;
assign addr[58224]= 455461206;
assign addr[58225]= 492762486;
assign addr[58226]= 529907477;
assign addr[58227]= 566884397;
assign addr[58228]= 603681519;
assign addr[58229]= 640287172;
assign addr[58230]= 676689746;
assign addr[58231]= 712877694;
assign addr[58232]= 748839539;
assign addr[58233]= 784563876;
assign addr[58234]= 820039373;
assign addr[58235]= 855254778;
assign addr[58236]= 890198924;
assign addr[58237]= 924860725;
assign addr[58238]= 959229189;
assign addr[58239]= 993293415;
assign addr[58240]= 1027042599;
assign addr[58241]= 1060466036;
assign addr[58242]= 1093553126;
assign addr[58243]= 1126293375;
assign addr[58244]= 1158676398;
assign addr[58245]= 1190691925;
assign addr[58246]= 1222329801;
assign addr[58247]= 1253579991;
assign addr[58248]= 1284432584;
assign addr[58249]= 1314877795;
assign addr[58250]= 1344905966;
assign addr[58251]= 1374507575;
assign addr[58252]= 1403673233;
assign addr[58253]= 1432393688;
assign addr[58254]= 1460659832;
assign addr[58255]= 1488462700;
assign addr[58256]= 1515793473;
assign addr[58257]= 1542643483;
assign addr[58258]= 1569004214;
assign addr[58259]= 1594867305;
assign addr[58260]= 1620224553;
assign addr[58261]= 1645067915;
assign addr[58262]= 1669389513;
assign addr[58263]= 1693181631;
assign addr[58264]= 1716436725;
assign addr[58265]= 1739147417;
assign addr[58266]= 1761306505;
assign addr[58267]= 1782906961;
assign addr[58268]= 1803941934;
assign addr[58269]= 1824404752;
assign addr[58270]= 1844288924;
assign addr[58271]= 1863588145;
assign addr[58272]= 1882296293;
assign addr[58273]= 1900407434;
assign addr[58274]= 1917915825;
assign addr[58275]= 1934815911;
assign addr[58276]= 1951102334;
assign addr[58277]= 1966769926;
assign addr[58278]= 1981813720;
assign addr[58279]= 1996228943;
assign addr[58280]= 2010011024;
assign addr[58281]= 2023155591;
assign addr[58282]= 2035658475;
assign addr[58283]= 2047515711;
assign addr[58284]= 2058723538;
assign addr[58285]= 2069278401;
assign addr[58286]= 2079176953;
assign addr[58287]= 2088416053;
assign addr[58288]= 2096992772;
assign addr[58289]= 2104904390;
assign addr[58290]= 2112148396;
assign addr[58291]= 2118722494;
assign addr[58292]= 2124624598;
assign addr[58293]= 2129852837;
assign addr[58294]= 2134405552;
assign addr[58295]= 2138281298;
assign addr[58296]= 2141478848;
assign addr[58297]= 2143997187;
assign addr[58298]= 2145835515;
assign addr[58299]= 2146993250;
assign addr[58300]= 2147470025;
assign addr[58301]= 2147265689;
assign addr[58302]= 2146380306;
assign addr[58303]= 2144814157;
assign addr[58304]= 2142567738;
assign addr[58305]= 2139641764;
assign addr[58306]= 2136037160;
assign addr[58307]= 2131755071;
assign addr[58308]= 2126796855;
assign addr[58309]= 2121164085;
assign addr[58310]= 2114858546;
assign addr[58311]= 2107882239;
assign addr[58312]= 2100237377;
assign addr[58313]= 2091926384;
assign addr[58314]= 2082951896;
assign addr[58315]= 2073316760;
assign addr[58316]= 2063024031;
assign addr[58317]= 2052076975;
assign addr[58318]= 2040479063;
assign addr[58319]= 2028233973;
assign addr[58320]= 2015345591;
assign addr[58321]= 2001818002;
assign addr[58322]= 1987655498;
assign addr[58323]= 1972862571;
assign addr[58324]= 1957443913;
assign addr[58325]= 1941404413;
assign addr[58326]= 1924749160;
assign addr[58327]= 1907483436;
assign addr[58328]= 1889612716;
assign addr[58329]= 1871142669;
assign addr[58330]= 1852079154;
assign addr[58331]= 1832428215;
assign addr[58332]= 1812196087;
assign addr[58333]= 1791389186;
assign addr[58334]= 1770014111;
assign addr[58335]= 1748077642;
assign addr[58336]= 1725586737;
assign addr[58337]= 1702548529;
assign addr[58338]= 1678970324;
assign addr[58339]= 1654859602;
assign addr[58340]= 1630224009;
assign addr[58341]= 1605071359;
assign addr[58342]= 1579409630;
assign addr[58343]= 1553246960;
assign addr[58344]= 1526591649;
assign addr[58345]= 1499452149;
assign addr[58346]= 1471837070;
assign addr[58347]= 1443755168;
assign addr[58348]= 1415215352;
assign addr[58349]= 1386226674;
assign addr[58350]= 1356798326;
assign addr[58351]= 1326939644;
assign addr[58352]= 1296660098;
assign addr[58353]= 1265969291;
assign addr[58354]= 1234876957;
assign addr[58355]= 1203392958;
assign addr[58356]= 1171527280;
assign addr[58357]= 1139290029;
assign addr[58358]= 1106691431;
assign addr[58359]= 1073741824;
assign addr[58360]= 1040451659;
assign addr[58361]= 1006831495;
assign addr[58362]= 972891995;
assign addr[58363]= 938643924;
assign addr[58364]= 904098143;
assign addr[58365]= 869265610;
assign addr[58366]= 834157373;
assign addr[58367]= 798784567;
assign addr[58368]= 763158411;
assign addr[58369]= 727290205;
assign addr[58370]= 691191324;
assign addr[58371]= 654873219;
assign addr[58372]= 618347408;
assign addr[58373]= 581625477;
assign addr[58374]= 544719071;
assign addr[58375]= 507639898;
assign addr[58376]= 470399716;
assign addr[58377]= 433010339;
assign addr[58378]= 395483624;
assign addr[58379]= 357831473;
assign addr[58380]= 320065829;
assign addr[58381]= 282198671;
assign addr[58382]= 244242007;
assign addr[58383]= 206207878;
assign addr[58384]= 168108346;
assign addr[58385]= 129955495;
assign addr[58386]= 91761426;
assign addr[58387]= 53538253;
assign addr[58388]= 15298099;
assign addr[58389]= -22946906;
assign addr[58390]= -61184634;
assign addr[58391]= -99402956;
assign addr[58392]= -137589750;
assign addr[58393]= -175732905;
assign addr[58394]= -213820322;
assign addr[58395]= -251839923;
assign addr[58396]= -289779648;
assign addr[58397]= -327627463;
assign addr[58398]= -365371365;
assign addr[58399]= -402999383;
assign addr[58400]= -440499581;
assign addr[58401]= -477860067;
assign addr[58402]= -515068990;
assign addr[58403]= -552114549;
assign addr[58404]= -588984994;
assign addr[58405]= -625668632;
assign addr[58406]= -662153826;
assign addr[58407]= -698429006;
assign addr[58408]= -734482665;
assign addr[58409]= -770303369;
assign addr[58410]= -805879757;
assign addr[58411]= -841200544;
assign addr[58412]= -876254528;
assign addr[58413]= -911030591;
assign addr[58414]= -945517704;
assign addr[58415]= -979704927;
assign addr[58416]= -1013581418;
assign addr[58417]= -1047136432;
assign addr[58418]= -1080359326;
assign addr[58419]= -1113239564;
assign addr[58420]= -1145766716;
assign addr[58421]= -1177930466;
assign addr[58422]= -1209720613;
assign addr[58423]= -1241127074;
assign addr[58424]= -1272139887;
assign addr[58425]= -1302749217;
assign addr[58426]= -1332945355;
assign addr[58427]= -1362718723;
assign addr[58428]= -1392059879;
assign addr[58429]= -1420959516;
assign addr[58430]= -1449408469;
assign addr[58431]= -1477397714;
assign addr[58432]= -1504918373;
assign addr[58433]= -1531961719;
assign addr[58434]= -1558519173;
assign addr[58435]= -1584582314;
assign addr[58436]= -1610142873;
assign addr[58437]= -1635192744;
assign addr[58438]= -1659723983;
assign addr[58439]= -1683728808;
assign addr[58440]= -1707199606;
assign addr[58441]= -1730128933;
assign addr[58442]= -1752509516;
assign addr[58443]= -1774334257;
assign addr[58444]= -1795596234;
assign addr[58445]= -1816288703;
assign addr[58446]= -1836405100;
assign addr[58447]= -1855939047;
assign addr[58448]= -1874884346;
assign addr[58449]= -1893234990;
assign addr[58450]= -1910985158;
assign addr[58451]= -1928129220;
assign addr[58452]= -1944661739;
assign addr[58453]= -1960577471;
assign addr[58454]= -1975871368;
assign addr[58455]= -1990538579;
assign addr[58456]= -2004574453;
assign addr[58457]= -2017974537;
assign addr[58458]= -2030734582;
assign addr[58459]= -2042850540;
assign addr[58460]= -2054318569;
assign addr[58461]= -2065135031;
assign addr[58462]= -2075296495;
assign addr[58463]= -2084799740;
assign addr[58464]= -2093641749;
assign addr[58465]= -2101819720;
assign addr[58466]= -2109331059;
assign addr[58467]= -2116173382;
assign addr[58468]= -2122344521;
assign addr[58469]= -2127842516;
assign addr[58470]= -2132665626;
assign addr[58471]= -2136812319;
assign addr[58472]= -2140281282;
assign addr[58473]= -2143071413;
assign addr[58474]= -2145181827;
assign addr[58475]= -2146611856;
assign addr[58476]= -2147361045;
assign addr[58477]= -2147429158;
assign addr[58478]= -2146816171;
assign addr[58479]= -2145522281;
assign addr[58480]= -2143547897;
assign addr[58481]= -2140893646;
assign addr[58482]= -2137560369;
assign addr[58483]= -2133549123;
assign addr[58484]= -2128861181;
assign addr[58485]= -2123498030;
assign addr[58486]= -2117461370;
assign addr[58487]= -2110753117;
assign addr[58488]= -2103375398;
assign addr[58489]= -2095330553;
assign addr[58490]= -2086621133;
assign addr[58491]= -2077249901;
assign addr[58492]= -2067219829;
assign addr[58493]= -2056534099;
assign addr[58494]= -2045196100;
assign addr[58495]= -2033209426;
assign addr[58496]= -2020577882;
assign addr[58497]= -2007305472;
assign addr[58498]= -1993396407;
assign addr[58499]= -1978855097;
assign addr[58500]= -1963686155;
assign addr[58501]= -1947894393;
assign addr[58502]= -1931484818;
assign addr[58503]= -1914462636;
assign addr[58504]= -1896833245;
assign addr[58505]= -1878602237;
assign addr[58506]= -1859775393;
assign addr[58507]= -1840358687;
assign addr[58508]= -1820358275;
assign addr[58509]= -1799780501;
assign addr[58510]= -1778631892;
assign addr[58511]= -1756919156;
assign addr[58512]= -1734649179;
assign addr[58513]= -1711829025;
assign addr[58514]= -1688465931;
assign addr[58515]= -1664567307;
assign addr[58516]= -1640140734;
assign addr[58517]= -1615193959;
assign addr[58518]= -1589734894;
assign addr[58519]= -1563771613;
assign addr[58520]= -1537312353;
assign addr[58521]= -1510365504;
assign addr[58522]= -1482939614;
assign addr[58523]= -1455043381;
assign addr[58524]= -1426685652;
assign addr[58525]= -1397875423;
assign addr[58526]= -1368621831;
assign addr[58527]= -1338934154;
assign addr[58528]= -1308821808;
assign addr[58529]= -1278294345;
assign addr[58530]= -1247361445;
assign addr[58531]= -1216032921;
assign addr[58532]= -1184318708;
assign addr[58533]= -1152228866;
assign addr[58534]= -1119773573;
assign addr[58535]= -1086963121;
assign addr[58536]= -1053807919;
assign addr[58537]= -1020318481;
assign addr[58538]= -986505429;
assign addr[58539]= -952379488;
assign addr[58540]= -917951481;
assign addr[58541]= -883232329;
assign addr[58542]= -848233042;
assign addr[58543]= -812964722;
assign addr[58544]= -777438554;
assign addr[58545]= -741665807;
assign addr[58546]= -705657826;
assign addr[58547]= -669426032;
assign addr[58548]= -632981917;
assign addr[58549]= -596337040;
assign addr[58550]= -559503022;
assign addr[58551]= -522491548;
assign addr[58552]= -485314355;
assign addr[58553]= -447983235;
assign addr[58554]= -410510029;
assign addr[58555]= -372906622;
assign addr[58556]= -335184940;
assign addr[58557]= -297356948;
assign addr[58558]= -259434643;
assign addr[58559]= -221430054;
assign addr[58560]= -183355234;
assign addr[58561]= -145222259;
assign addr[58562]= -107043224;
assign addr[58563]= -68830239;
assign addr[58564]= -30595422;
assign addr[58565]= 7649098;
assign addr[58566]= 45891193;
assign addr[58567]= 84118732;
assign addr[58568]= 122319591;
assign addr[58569]= 160481654;
assign addr[58570]= 198592817;
assign addr[58571]= 236640993;
assign addr[58572]= 274614114;
assign addr[58573]= 312500135;
assign addr[58574]= 350287041;
assign addr[58575]= 387962847;
assign addr[58576]= 425515602;
assign addr[58577]= 462933398;
assign addr[58578]= 500204365;
assign addr[58579]= 537316682;
assign addr[58580]= 574258580;
assign addr[58581]= 611018340;
assign addr[58582]= 647584304;
assign addr[58583]= 683944874;
assign addr[58584]= 720088517;
assign addr[58585]= 756003771;
assign addr[58586]= 791679244;
assign addr[58587]= 827103620;
assign addr[58588]= 862265664;
assign addr[58589]= 897154224;
assign addr[58590]= 931758235;
assign addr[58591]= 966066720;
assign addr[58592]= 1000068799;
assign addr[58593]= 1033753687;
assign addr[58594]= 1067110699;
assign addr[58595]= 1100129257;
assign addr[58596]= 1132798888;
assign addr[58597]= 1165109230;
assign addr[58598]= 1197050035;
assign addr[58599]= 1228611172;
assign addr[58600]= 1259782632;
assign addr[58601]= 1290554528;
assign addr[58602]= 1320917099;
assign addr[58603]= 1350860716;
assign addr[58604]= 1380375881;
assign addr[58605]= 1409453233;
assign addr[58606]= 1438083551;
assign addr[58607]= 1466257752;
assign addr[58608]= 1493966902;
assign addr[58609]= 1521202211;
assign addr[58610]= 1547955041;
assign addr[58611]= 1574216908;
assign addr[58612]= 1599979481;
assign addr[58613]= 1625234591;
assign addr[58614]= 1649974225;
assign addr[58615]= 1674190539;
assign addr[58616]= 1697875851;
assign addr[58617]= 1721022648;
assign addr[58618]= 1743623590;
assign addr[58619]= 1765671509;
assign addr[58620]= 1787159411;
assign addr[58621]= 1808080480;
assign addr[58622]= 1828428082;
assign addr[58623]= 1848195763;
assign addr[58624]= 1867377253;
assign addr[58625]= 1885966468;
assign addr[58626]= 1903957513;
assign addr[58627]= 1921344681;
assign addr[58628]= 1938122457;
assign addr[58629]= 1954285520;
assign addr[58630]= 1969828744;
assign addr[58631]= 1984747199;
assign addr[58632]= 1999036154;
assign addr[58633]= 2012691075;
assign addr[58634]= 2025707632;
assign addr[58635]= 2038081698;
assign addr[58636]= 2049809346;
assign addr[58637]= 2060886858;
assign addr[58638]= 2071310720;
assign addr[58639]= 2081077626;
assign addr[58640]= 2090184478;
assign addr[58641]= 2098628387;
assign addr[58642]= 2106406677;
assign addr[58643]= 2113516878;
assign addr[58644]= 2119956737;
assign addr[58645]= 2125724211;
assign addr[58646]= 2130817471;
assign addr[58647]= 2135234901;
assign addr[58648]= 2138975100;
assign addr[58649]= 2142036881;
assign addr[58650]= 2144419275;
assign addr[58651]= 2146121524;
assign addr[58652]= 2147143090;
assign addr[58653]= 2147483648;
assign addr[58654]= 2147143090;
assign addr[58655]= 2146121524;
assign addr[58656]= 2144419275;
assign addr[58657]= 2142036881;
assign addr[58658]= 2138975100;
assign addr[58659]= 2135234901;
assign addr[58660]= 2130817471;
assign addr[58661]= 2125724211;
assign addr[58662]= 2119956737;
assign addr[58663]= 2113516878;
assign addr[58664]= 2106406677;
assign addr[58665]= 2098628387;
assign addr[58666]= 2090184478;
assign addr[58667]= 2081077626;
assign addr[58668]= 2071310720;
assign addr[58669]= 2060886858;
assign addr[58670]= 2049809346;
assign addr[58671]= 2038081698;
assign addr[58672]= 2025707632;
assign addr[58673]= 2012691075;
assign addr[58674]= 1999036154;
assign addr[58675]= 1984747199;
assign addr[58676]= 1969828744;
assign addr[58677]= 1954285520;
assign addr[58678]= 1938122457;
assign addr[58679]= 1921344681;
assign addr[58680]= 1903957513;
assign addr[58681]= 1885966468;
assign addr[58682]= 1867377253;
assign addr[58683]= 1848195763;
assign addr[58684]= 1828428082;
assign addr[58685]= 1808080480;
assign addr[58686]= 1787159411;
assign addr[58687]= 1765671509;
assign addr[58688]= 1743623590;
assign addr[58689]= 1721022648;
assign addr[58690]= 1697875851;
assign addr[58691]= 1674190539;
assign addr[58692]= 1649974225;
assign addr[58693]= 1625234591;
assign addr[58694]= 1599979481;
assign addr[58695]= 1574216908;
assign addr[58696]= 1547955041;
assign addr[58697]= 1521202211;
assign addr[58698]= 1493966902;
assign addr[58699]= 1466257752;
assign addr[58700]= 1438083551;
assign addr[58701]= 1409453233;
assign addr[58702]= 1380375881;
assign addr[58703]= 1350860716;
assign addr[58704]= 1320917099;
assign addr[58705]= 1290554528;
assign addr[58706]= 1259782632;
assign addr[58707]= 1228611172;
assign addr[58708]= 1197050035;
assign addr[58709]= 1165109230;
assign addr[58710]= 1132798888;
assign addr[58711]= 1100129257;
assign addr[58712]= 1067110699;
assign addr[58713]= 1033753687;
assign addr[58714]= 1000068799;
assign addr[58715]= 966066720;
assign addr[58716]= 931758235;
assign addr[58717]= 897154224;
assign addr[58718]= 862265664;
assign addr[58719]= 827103620;
assign addr[58720]= 791679244;
assign addr[58721]= 756003771;
assign addr[58722]= 720088517;
assign addr[58723]= 683944874;
assign addr[58724]= 647584304;
assign addr[58725]= 611018340;
assign addr[58726]= 574258580;
assign addr[58727]= 537316682;
assign addr[58728]= 500204365;
assign addr[58729]= 462933398;
assign addr[58730]= 425515602;
assign addr[58731]= 387962847;
assign addr[58732]= 350287041;
assign addr[58733]= 312500135;
assign addr[58734]= 274614114;
assign addr[58735]= 236640993;
assign addr[58736]= 198592817;
assign addr[58737]= 160481654;
assign addr[58738]= 122319591;
assign addr[58739]= 84118732;
assign addr[58740]= 45891193;
assign addr[58741]= 7649098;
assign addr[58742]= -30595422;
assign addr[58743]= -68830239;
assign addr[58744]= -107043224;
assign addr[58745]= -145222259;
assign addr[58746]= -183355234;
assign addr[58747]= -221430054;
assign addr[58748]= -259434643;
assign addr[58749]= -297356948;
assign addr[58750]= -335184940;
assign addr[58751]= -372906622;
assign addr[58752]= -410510029;
assign addr[58753]= -447983235;
assign addr[58754]= -485314355;
assign addr[58755]= -522491548;
assign addr[58756]= -559503022;
assign addr[58757]= -596337040;
assign addr[58758]= -632981917;
assign addr[58759]= -669426032;
assign addr[58760]= -705657826;
assign addr[58761]= -741665807;
assign addr[58762]= -777438554;
assign addr[58763]= -812964722;
assign addr[58764]= -848233042;
assign addr[58765]= -883232329;
assign addr[58766]= -917951481;
assign addr[58767]= -952379488;
assign addr[58768]= -986505429;
assign addr[58769]= -1020318481;
assign addr[58770]= -1053807919;
assign addr[58771]= -1086963121;
assign addr[58772]= -1119773573;
assign addr[58773]= -1152228866;
assign addr[58774]= -1184318708;
assign addr[58775]= -1216032921;
assign addr[58776]= -1247361445;
assign addr[58777]= -1278294345;
assign addr[58778]= -1308821808;
assign addr[58779]= -1338934154;
assign addr[58780]= -1368621831;
assign addr[58781]= -1397875423;
assign addr[58782]= -1426685652;
assign addr[58783]= -1455043381;
assign addr[58784]= -1482939614;
assign addr[58785]= -1510365504;
assign addr[58786]= -1537312353;
assign addr[58787]= -1563771613;
assign addr[58788]= -1589734894;
assign addr[58789]= -1615193959;
assign addr[58790]= -1640140734;
assign addr[58791]= -1664567307;
assign addr[58792]= -1688465931;
assign addr[58793]= -1711829025;
assign addr[58794]= -1734649179;
assign addr[58795]= -1756919156;
assign addr[58796]= -1778631892;
assign addr[58797]= -1799780501;
assign addr[58798]= -1820358275;
assign addr[58799]= -1840358687;
assign addr[58800]= -1859775393;
assign addr[58801]= -1878602237;
assign addr[58802]= -1896833245;
assign addr[58803]= -1914462636;
assign addr[58804]= -1931484818;
assign addr[58805]= -1947894393;
assign addr[58806]= -1963686155;
assign addr[58807]= -1978855097;
assign addr[58808]= -1993396407;
assign addr[58809]= -2007305472;
assign addr[58810]= -2020577882;
assign addr[58811]= -2033209426;
assign addr[58812]= -2045196100;
assign addr[58813]= -2056534099;
assign addr[58814]= -2067219829;
assign addr[58815]= -2077249901;
assign addr[58816]= -2086621133;
assign addr[58817]= -2095330553;
assign addr[58818]= -2103375398;
assign addr[58819]= -2110753117;
assign addr[58820]= -2117461370;
assign addr[58821]= -2123498030;
assign addr[58822]= -2128861181;
assign addr[58823]= -2133549123;
assign addr[58824]= -2137560369;
assign addr[58825]= -2140893646;
assign addr[58826]= -2143547897;
assign addr[58827]= -2145522281;
assign addr[58828]= -2146816171;
assign addr[58829]= -2147429158;
assign addr[58830]= -2147361045;
assign addr[58831]= -2146611856;
assign addr[58832]= -2145181827;
assign addr[58833]= -2143071413;
assign addr[58834]= -2140281282;
assign addr[58835]= -2136812319;
assign addr[58836]= -2132665626;
assign addr[58837]= -2127842516;
assign addr[58838]= -2122344521;
assign addr[58839]= -2116173382;
assign addr[58840]= -2109331059;
assign addr[58841]= -2101819720;
assign addr[58842]= -2093641749;
assign addr[58843]= -2084799740;
assign addr[58844]= -2075296495;
assign addr[58845]= -2065135031;
assign addr[58846]= -2054318569;
assign addr[58847]= -2042850540;
assign addr[58848]= -2030734582;
assign addr[58849]= -2017974537;
assign addr[58850]= -2004574453;
assign addr[58851]= -1990538579;
assign addr[58852]= -1975871368;
assign addr[58853]= -1960577471;
assign addr[58854]= -1944661739;
assign addr[58855]= -1928129220;
assign addr[58856]= -1910985158;
assign addr[58857]= -1893234990;
assign addr[58858]= -1874884346;
assign addr[58859]= -1855939047;
assign addr[58860]= -1836405100;
assign addr[58861]= -1816288703;
assign addr[58862]= -1795596234;
assign addr[58863]= -1774334257;
assign addr[58864]= -1752509516;
assign addr[58865]= -1730128933;
assign addr[58866]= -1707199606;
assign addr[58867]= -1683728808;
assign addr[58868]= -1659723983;
assign addr[58869]= -1635192744;
assign addr[58870]= -1610142873;
assign addr[58871]= -1584582314;
assign addr[58872]= -1558519173;
assign addr[58873]= -1531961719;
assign addr[58874]= -1504918373;
assign addr[58875]= -1477397714;
assign addr[58876]= -1449408469;
assign addr[58877]= -1420959516;
assign addr[58878]= -1392059879;
assign addr[58879]= -1362718723;
assign addr[58880]= -1332945355;
assign addr[58881]= -1302749217;
assign addr[58882]= -1272139887;
assign addr[58883]= -1241127074;
assign addr[58884]= -1209720613;
assign addr[58885]= -1177930466;
assign addr[58886]= -1145766716;
assign addr[58887]= -1113239564;
assign addr[58888]= -1080359326;
assign addr[58889]= -1047136432;
assign addr[58890]= -1013581418;
assign addr[58891]= -979704927;
assign addr[58892]= -945517704;
assign addr[58893]= -911030591;
assign addr[58894]= -876254528;
assign addr[58895]= -841200544;
assign addr[58896]= -805879757;
assign addr[58897]= -770303369;
assign addr[58898]= -734482665;
assign addr[58899]= -698429006;
assign addr[58900]= -662153826;
assign addr[58901]= -625668632;
assign addr[58902]= -588984994;
assign addr[58903]= -552114549;
assign addr[58904]= -515068990;
assign addr[58905]= -477860067;
assign addr[58906]= -440499581;
assign addr[58907]= -402999383;
assign addr[58908]= -365371365;
assign addr[58909]= -327627463;
assign addr[58910]= -289779648;
assign addr[58911]= -251839923;
assign addr[58912]= -213820322;
assign addr[58913]= -175732905;
assign addr[58914]= -137589750;
assign addr[58915]= -99402956;
assign addr[58916]= -61184634;
assign addr[58917]= -22946906;
assign addr[58918]= 15298099;
assign addr[58919]= 53538253;
assign addr[58920]= 91761426;
assign addr[58921]= 129955495;
assign addr[58922]= 168108346;
assign addr[58923]= 206207878;
assign addr[58924]= 244242007;
assign addr[58925]= 282198671;
assign addr[58926]= 320065829;
assign addr[58927]= 357831473;
assign addr[58928]= 395483624;
assign addr[58929]= 433010339;
assign addr[58930]= 470399716;
assign addr[58931]= 507639898;
assign addr[58932]= 544719071;
assign addr[58933]= 581625477;
assign addr[58934]= 618347408;
assign addr[58935]= 654873219;
assign addr[58936]= 691191324;
assign addr[58937]= 727290205;
assign addr[58938]= 763158411;
assign addr[58939]= 798784567;
assign addr[58940]= 834157373;
assign addr[58941]= 869265610;
assign addr[58942]= 904098143;
assign addr[58943]= 938643924;
assign addr[58944]= 972891995;
assign addr[58945]= 1006831495;
assign addr[58946]= 1040451659;
assign addr[58947]= 1073741824;
assign addr[58948]= 1106691431;
assign addr[58949]= 1139290029;
assign addr[58950]= 1171527280;
assign addr[58951]= 1203392958;
assign addr[58952]= 1234876957;
assign addr[58953]= 1265969291;
assign addr[58954]= 1296660098;
assign addr[58955]= 1326939644;
assign addr[58956]= 1356798326;
assign addr[58957]= 1386226674;
assign addr[58958]= 1415215352;
assign addr[58959]= 1443755168;
assign addr[58960]= 1471837070;
assign addr[58961]= 1499452149;
assign addr[58962]= 1526591649;
assign addr[58963]= 1553246960;
assign addr[58964]= 1579409630;
assign addr[58965]= 1605071359;
assign addr[58966]= 1630224009;
assign addr[58967]= 1654859602;
assign addr[58968]= 1678970324;
assign addr[58969]= 1702548529;
assign addr[58970]= 1725586737;
assign addr[58971]= 1748077642;
assign addr[58972]= 1770014111;
assign addr[58973]= 1791389186;
assign addr[58974]= 1812196087;
assign addr[58975]= 1832428215;
assign addr[58976]= 1852079154;
assign addr[58977]= 1871142669;
assign addr[58978]= 1889612716;
assign addr[58979]= 1907483436;
assign addr[58980]= 1924749160;
assign addr[58981]= 1941404413;
assign addr[58982]= 1957443913;
assign addr[58983]= 1972862571;
assign addr[58984]= 1987655498;
assign addr[58985]= 2001818002;
assign addr[58986]= 2015345591;
assign addr[58987]= 2028233973;
assign addr[58988]= 2040479063;
assign addr[58989]= 2052076975;
assign addr[58990]= 2063024031;
assign addr[58991]= 2073316760;
assign addr[58992]= 2082951896;
assign addr[58993]= 2091926384;
assign addr[58994]= 2100237377;
assign addr[58995]= 2107882239;
assign addr[58996]= 2114858546;
assign addr[58997]= 2121164085;
assign addr[58998]= 2126796855;
assign addr[58999]= 2131755071;
assign addr[59000]= 2136037160;
assign addr[59001]= 2139641764;
assign addr[59002]= 2142567738;
assign addr[59003]= 2144814157;
assign addr[59004]= 2146380306;
assign addr[59005]= 2147265689;
assign addr[59006]= 2147470025;
assign addr[59007]= 2146993250;
assign addr[59008]= 2145835515;
assign addr[59009]= 2143997187;
assign addr[59010]= 2141478848;
assign addr[59011]= 2138281298;
assign addr[59012]= 2134405552;
assign addr[59013]= 2129852837;
assign addr[59014]= 2124624598;
assign addr[59015]= 2118722494;
assign addr[59016]= 2112148396;
assign addr[59017]= 2104904390;
assign addr[59018]= 2096992772;
assign addr[59019]= 2088416053;
assign addr[59020]= 2079176953;
assign addr[59021]= 2069278401;
assign addr[59022]= 2058723538;
assign addr[59023]= 2047515711;
assign addr[59024]= 2035658475;
assign addr[59025]= 2023155591;
assign addr[59026]= 2010011024;
assign addr[59027]= 1996228943;
assign addr[59028]= 1981813720;
assign addr[59029]= 1966769926;
assign addr[59030]= 1951102334;
assign addr[59031]= 1934815911;
assign addr[59032]= 1917915825;
assign addr[59033]= 1900407434;
assign addr[59034]= 1882296293;
assign addr[59035]= 1863588145;
assign addr[59036]= 1844288924;
assign addr[59037]= 1824404752;
assign addr[59038]= 1803941934;
assign addr[59039]= 1782906961;
assign addr[59040]= 1761306505;
assign addr[59041]= 1739147417;
assign addr[59042]= 1716436725;
assign addr[59043]= 1693181631;
assign addr[59044]= 1669389513;
assign addr[59045]= 1645067915;
assign addr[59046]= 1620224553;
assign addr[59047]= 1594867305;
assign addr[59048]= 1569004214;
assign addr[59049]= 1542643483;
assign addr[59050]= 1515793473;
assign addr[59051]= 1488462700;
assign addr[59052]= 1460659832;
assign addr[59053]= 1432393688;
assign addr[59054]= 1403673233;
assign addr[59055]= 1374507575;
assign addr[59056]= 1344905966;
assign addr[59057]= 1314877795;
assign addr[59058]= 1284432584;
assign addr[59059]= 1253579991;
assign addr[59060]= 1222329801;
assign addr[59061]= 1190691925;
assign addr[59062]= 1158676398;
assign addr[59063]= 1126293375;
assign addr[59064]= 1093553126;
assign addr[59065]= 1060466036;
assign addr[59066]= 1027042599;
assign addr[59067]= 993293415;
assign addr[59068]= 959229189;
assign addr[59069]= 924860725;
assign addr[59070]= 890198924;
assign addr[59071]= 855254778;
assign addr[59072]= 820039373;
assign addr[59073]= 784563876;
assign addr[59074]= 748839539;
assign addr[59075]= 712877694;
assign addr[59076]= 676689746;
assign addr[59077]= 640287172;
assign addr[59078]= 603681519;
assign addr[59079]= 566884397;
assign addr[59080]= 529907477;
assign addr[59081]= 492762486;
assign addr[59082]= 455461206;
assign addr[59083]= 418015468;
assign addr[59084]= 380437148;
assign addr[59085]= 342738165;
assign addr[59086]= 304930476;
assign addr[59087]= 267026072;
assign addr[59088]= 229036977;
assign addr[59089]= 190975237;
assign addr[59090]= 152852926;
assign addr[59091]= 114682135;
assign addr[59092]= 76474970;
assign addr[59093]= 38243550;
assign addr[59094]= 0;
assign addr[59095]= -38243550;
assign addr[59096]= -76474970;
assign addr[59097]= -114682135;
assign addr[59098]= -152852926;
assign addr[59099]= -190975237;
assign addr[59100]= -229036977;
assign addr[59101]= -267026072;
assign addr[59102]= -304930476;
assign addr[59103]= -342738165;
assign addr[59104]= -380437148;
assign addr[59105]= -418015468;
assign addr[59106]= -455461206;
assign addr[59107]= -492762486;
assign addr[59108]= -529907477;
assign addr[59109]= -566884397;
assign addr[59110]= -603681519;
assign addr[59111]= -640287172;
assign addr[59112]= -676689746;
assign addr[59113]= -712877694;
assign addr[59114]= -748839539;
assign addr[59115]= -784563876;
assign addr[59116]= -820039373;
assign addr[59117]= -855254778;
assign addr[59118]= -890198924;
assign addr[59119]= -924860725;
assign addr[59120]= -959229189;
assign addr[59121]= -993293415;
assign addr[59122]= -1027042599;
assign addr[59123]= -1060466036;
assign addr[59124]= -1093553126;
assign addr[59125]= -1126293375;
assign addr[59126]= -1158676398;
assign addr[59127]= -1190691925;
assign addr[59128]= -1222329801;
assign addr[59129]= -1253579991;
assign addr[59130]= -1284432584;
assign addr[59131]= -1314877795;
assign addr[59132]= -1344905966;
assign addr[59133]= -1374507575;
assign addr[59134]= -1403673233;
assign addr[59135]= -1432393688;
assign addr[59136]= -1460659832;
assign addr[59137]= -1488462700;
assign addr[59138]= -1515793473;
assign addr[59139]= -1542643483;
assign addr[59140]= -1569004214;
assign addr[59141]= -1594867305;
assign addr[59142]= -1620224553;
assign addr[59143]= -1645067915;
assign addr[59144]= -1669389513;
assign addr[59145]= -1693181631;
assign addr[59146]= -1716436725;
assign addr[59147]= -1739147417;
assign addr[59148]= -1761306505;
assign addr[59149]= -1782906961;
assign addr[59150]= -1803941934;
assign addr[59151]= -1824404752;
assign addr[59152]= -1844288924;
assign addr[59153]= -1863588145;
assign addr[59154]= -1882296293;
assign addr[59155]= -1900407434;
assign addr[59156]= -1917915825;
assign addr[59157]= -1934815911;
assign addr[59158]= -1951102334;
assign addr[59159]= -1966769926;
assign addr[59160]= -1981813720;
assign addr[59161]= -1996228943;
assign addr[59162]= -2010011024;
assign addr[59163]= -2023155591;
assign addr[59164]= -2035658475;
assign addr[59165]= -2047515711;
assign addr[59166]= -2058723538;
assign addr[59167]= -2069278401;
assign addr[59168]= -2079176953;
assign addr[59169]= -2088416053;
assign addr[59170]= -2096992772;
assign addr[59171]= -2104904390;
assign addr[59172]= -2112148396;
assign addr[59173]= -2118722494;
assign addr[59174]= -2124624598;
assign addr[59175]= -2129852837;
assign addr[59176]= -2134405552;
assign addr[59177]= -2138281298;
assign addr[59178]= -2141478848;
assign addr[59179]= -2143997187;
assign addr[59180]= -2145835515;
assign addr[59181]= -2146993250;
assign addr[59182]= -2147470025;
assign addr[59183]= -2147265689;
assign addr[59184]= -2146380306;
assign addr[59185]= -2144814157;
assign addr[59186]= -2142567738;
assign addr[59187]= -2139641764;
assign addr[59188]= -2136037160;
assign addr[59189]= -2131755071;
assign addr[59190]= -2126796855;
assign addr[59191]= -2121164085;
assign addr[59192]= -2114858546;
assign addr[59193]= -2107882239;
assign addr[59194]= -2100237377;
assign addr[59195]= -2091926384;
assign addr[59196]= -2082951896;
assign addr[59197]= -2073316760;
assign addr[59198]= -2063024031;
assign addr[59199]= -2052076975;
assign addr[59200]= -2040479063;
assign addr[59201]= -2028233973;
assign addr[59202]= -2015345591;
assign addr[59203]= -2001818002;
assign addr[59204]= -1987655498;
assign addr[59205]= -1972862571;
assign addr[59206]= -1957443913;
assign addr[59207]= -1941404413;
assign addr[59208]= -1924749160;
assign addr[59209]= -1907483436;
assign addr[59210]= -1889612716;
assign addr[59211]= -1871142669;
assign addr[59212]= -1852079154;
assign addr[59213]= -1832428215;
assign addr[59214]= -1812196087;
assign addr[59215]= -1791389186;
assign addr[59216]= -1770014111;
assign addr[59217]= -1748077642;
assign addr[59218]= -1725586737;
assign addr[59219]= -1702548529;
assign addr[59220]= -1678970324;
assign addr[59221]= -1654859602;
assign addr[59222]= -1630224009;
assign addr[59223]= -1605071359;
assign addr[59224]= -1579409630;
assign addr[59225]= -1553246960;
assign addr[59226]= -1526591649;
assign addr[59227]= -1499452149;
assign addr[59228]= -1471837070;
assign addr[59229]= -1443755168;
assign addr[59230]= -1415215352;
assign addr[59231]= -1386226674;
assign addr[59232]= -1356798326;
assign addr[59233]= -1326939644;
assign addr[59234]= -1296660098;
assign addr[59235]= -1265969291;
assign addr[59236]= -1234876957;
assign addr[59237]= -1203392958;
assign addr[59238]= -1171527280;
assign addr[59239]= -1139290029;
assign addr[59240]= -1106691431;
assign addr[59241]= -1073741824;
assign addr[59242]= -1040451659;
assign addr[59243]= -1006831495;
assign addr[59244]= -972891995;
assign addr[59245]= -938643924;
assign addr[59246]= -904098143;
assign addr[59247]= -869265610;
assign addr[59248]= -834157373;
assign addr[59249]= -798784567;
assign addr[59250]= -763158411;
assign addr[59251]= -727290205;
assign addr[59252]= -691191324;
assign addr[59253]= -654873219;
assign addr[59254]= -618347408;
assign addr[59255]= -581625477;
assign addr[59256]= -544719071;
assign addr[59257]= -507639898;
assign addr[59258]= -470399716;
assign addr[59259]= -433010339;
assign addr[59260]= -395483624;
assign addr[59261]= -357831473;
assign addr[59262]= -320065829;
assign addr[59263]= -282198671;
assign addr[59264]= -244242007;
assign addr[59265]= -206207878;
assign addr[59266]= -168108346;
assign addr[59267]= -129955495;
assign addr[59268]= -91761426;
assign addr[59269]= -53538253;
assign addr[59270]= -15298099;
assign addr[59271]= 22946906;
assign addr[59272]= 61184634;
assign addr[59273]= 99402956;
assign addr[59274]= 137589750;
assign addr[59275]= 175732905;
assign addr[59276]= 213820322;
assign addr[59277]= 251839923;
assign addr[59278]= 289779648;
assign addr[59279]= 327627463;
assign addr[59280]= 365371365;
assign addr[59281]= 402999383;
assign addr[59282]= 440499581;
assign addr[59283]= 477860067;
assign addr[59284]= 515068990;
assign addr[59285]= 552114549;
assign addr[59286]= 588984994;
assign addr[59287]= 625668632;
assign addr[59288]= 662153826;
assign addr[59289]= 698429006;
assign addr[59290]= 734482665;
assign addr[59291]= 770303369;
assign addr[59292]= 805879757;
assign addr[59293]= 841200544;
assign addr[59294]= 876254528;
assign addr[59295]= 911030591;
assign addr[59296]= 945517704;
assign addr[59297]= 979704927;
assign addr[59298]= 1013581418;
assign addr[59299]= 1047136432;
assign addr[59300]= 1080359326;
assign addr[59301]= 1113239564;
assign addr[59302]= 1145766716;
assign addr[59303]= 1177930466;
assign addr[59304]= 1209720613;
assign addr[59305]= 1241127074;
assign addr[59306]= 1272139887;
assign addr[59307]= 1302749217;
assign addr[59308]= 1332945355;
assign addr[59309]= 1362718723;
assign addr[59310]= 1392059879;
assign addr[59311]= 1420959516;
assign addr[59312]= 1449408469;
assign addr[59313]= 1477397714;
assign addr[59314]= 1504918373;
assign addr[59315]= 1531961719;
assign addr[59316]= 1558519173;
assign addr[59317]= 1584582314;
assign addr[59318]= 1610142873;
assign addr[59319]= 1635192744;
assign addr[59320]= 1659723983;
assign addr[59321]= 1683728808;
assign addr[59322]= 1707199606;
assign addr[59323]= 1730128933;
assign addr[59324]= 1752509516;
assign addr[59325]= 1774334257;
assign addr[59326]= 1795596234;
assign addr[59327]= 1816288703;
assign addr[59328]= 1836405100;
assign addr[59329]= 1855939047;
assign addr[59330]= 1874884346;
assign addr[59331]= 1893234990;
assign addr[59332]= 1910985158;
assign addr[59333]= 1928129220;
assign addr[59334]= 1944661739;
assign addr[59335]= 1960577471;
assign addr[59336]= 1975871368;
assign addr[59337]= 1990538579;
assign addr[59338]= 2004574453;
assign addr[59339]= 2017974537;
assign addr[59340]= 2030734582;
assign addr[59341]= 2042850540;
assign addr[59342]= 2054318569;
assign addr[59343]= 2065135031;
assign addr[59344]= 2075296495;
assign addr[59345]= 2084799740;
assign addr[59346]= 2093641749;
assign addr[59347]= 2101819720;
assign addr[59348]= 2109331059;
assign addr[59349]= 2116173382;
assign addr[59350]= 2122344521;
assign addr[59351]= 2127842516;
assign addr[59352]= 2132665626;
assign addr[59353]= 2136812319;
assign addr[59354]= 2140281282;
assign addr[59355]= 2143071413;
assign addr[59356]= 2145181827;
assign addr[59357]= 2146611856;
assign addr[59358]= 2147361045;
assign addr[59359]= 2147429158;
assign addr[59360]= 2146816171;
assign addr[59361]= 2145522281;
assign addr[59362]= 2143547897;
assign addr[59363]= 2140893646;
assign addr[59364]= 2137560369;
assign addr[59365]= 2133549123;
assign addr[59366]= 2128861181;
assign addr[59367]= 2123498030;
assign addr[59368]= 2117461370;
assign addr[59369]= 2110753117;
assign addr[59370]= 2103375398;
assign addr[59371]= 2095330553;
assign addr[59372]= 2086621133;
assign addr[59373]= 2077249901;
assign addr[59374]= 2067219829;
assign addr[59375]= 2056534099;
assign addr[59376]= 2045196100;
assign addr[59377]= 2033209426;
assign addr[59378]= 2020577882;
assign addr[59379]= 2007305472;
assign addr[59380]= 1993396407;
assign addr[59381]= 1978855097;
assign addr[59382]= 1963686155;
assign addr[59383]= 1947894393;
assign addr[59384]= 1931484818;
assign addr[59385]= 1914462636;
assign addr[59386]= 1896833245;
assign addr[59387]= 1878602237;
assign addr[59388]= 1859775393;
assign addr[59389]= 1840358687;
assign addr[59390]= 1820358275;
assign addr[59391]= 1799780501;
assign addr[59392]= 1778631892;
assign addr[59393]= 1756919156;
assign addr[59394]= 1734649179;
assign addr[59395]= 1711829025;
assign addr[59396]= 1688465931;
assign addr[59397]= 1664567307;
assign addr[59398]= 1640140734;
assign addr[59399]= 1615193959;
assign addr[59400]= 1589734894;
assign addr[59401]= 1563771613;
assign addr[59402]= 1537312353;
assign addr[59403]= 1510365504;
assign addr[59404]= 1482939614;
assign addr[59405]= 1455043381;
assign addr[59406]= 1426685652;
assign addr[59407]= 1397875423;
assign addr[59408]= 1368621831;
assign addr[59409]= 1338934154;
assign addr[59410]= 1308821808;
assign addr[59411]= 1278294345;
assign addr[59412]= 1247361445;
assign addr[59413]= 1216032921;
assign addr[59414]= 1184318708;
assign addr[59415]= 1152228866;
assign addr[59416]= 1119773573;
assign addr[59417]= 1086963121;
assign addr[59418]= 1053807919;
assign addr[59419]= 1020318481;
assign addr[59420]= 986505429;
assign addr[59421]= 952379488;
assign addr[59422]= 917951481;
assign addr[59423]= 883232329;
assign addr[59424]= 848233042;
assign addr[59425]= 812964722;
assign addr[59426]= 777438554;
assign addr[59427]= 741665807;
assign addr[59428]= 705657826;
assign addr[59429]= 669426032;
assign addr[59430]= 632981917;
assign addr[59431]= 596337040;
assign addr[59432]= 559503022;
assign addr[59433]= 522491548;
assign addr[59434]= 485314355;
assign addr[59435]= 447983235;
assign addr[59436]= 410510029;
assign addr[59437]= 372906622;
assign addr[59438]= 335184940;
assign addr[59439]= 297356948;
assign addr[59440]= 259434643;
assign addr[59441]= 221430054;
assign addr[59442]= 183355234;
assign addr[59443]= 145222259;
assign addr[59444]= 107043224;
assign addr[59445]= 68830239;
assign addr[59446]= 30595422;
assign addr[59447]= -7649098;
assign addr[59448]= -45891193;
assign addr[59449]= -84118732;
assign addr[59450]= -122319591;
assign addr[59451]= -160481654;
assign addr[59452]= -198592817;
assign addr[59453]= -236640993;
assign addr[59454]= -274614114;
assign addr[59455]= -312500135;
assign addr[59456]= -350287041;
assign addr[59457]= -387962847;
assign addr[59458]= -425515602;
assign addr[59459]= -462933398;
assign addr[59460]= -500204365;
assign addr[59461]= -537316682;
assign addr[59462]= -574258580;
assign addr[59463]= -611018340;
assign addr[59464]= -647584304;
assign addr[59465]= -683944874;
assign addr[59466]= -720088517;
assign addr[59467]= -756003771;
assign addr[59468]= -791679244;
assign addr[59469]= -827103620;
assign addr[59470]= -862265664;
assign addr[59471]= -897154224;
assign addr[59472]= -931758235;
assign addr[59473]= -966066720;
assign addr[59474]= -1000068799;
assign addr[59475]= -1033753687;
assign addr[59476]= -1067110699;
assign addr[59477]= -1100129257;
assign addr[59478]= -1132798888;
assign addr[59479]= -1165109230;
assign addr[59480]= -1197050035;
assign addr[59481]= -1228611172;
assign addr[59482]= -1259782632;
assign addr[59483]= -1290554528;
assign addr[59484]= -1320917099;
assign addr[59485]= -1350860716;
assign addr[59486]= -1380375881;
assign addr[59487]= -1409453233;
assign addr[59488]= -1438083551;
assign addr[59489]= -1466257752;
assign addr[59490]= -1493966902;
assign addr[59491]= -1521202211;
assign addr[59492]= -1547955041;
assign addr[59493]= -1574216908;
assign addr[59494]= -1599979481;
assign addr[59495]= -1625234591;
assign addr[59496]= -1649974225;
assign addr[59497]= -1674190539;
assign addr[59498]= -1697875851;
assign addr[59499]= -1721022648;
assign addr[59500]= -1743623590;
assign addr[59501]= -1765671509;
assign addr[59502]= -1787159411;
assign addr[59503]= -1808080480;
assign addr[59504]= -1828428082;
assign addr[59505]= -1848195763;
assign addr[59506]= -1867377253;
assign addr[59507]= -1885966468;
assign addr[59508]= -1903957513;
assign addr[59509]= -1921344681;
assign addr[59510]= -1938122457;
assign addr[59511]= -1954285520;
assign addr[59512]= -1969828744;
assign addr[59513]= -1984747199;
assign addr[59514]= -1999036154;
assign addr[59515]= -2012691075;
assign addr[59516]= -2025707632;
assign addr[59517]= -2038081698;
assign addr[59518]= -2049809346;
assign addr[59519]= -2060886858;
assign addr[59520]= -2071310720;
assign addr[59521]= -2081077626;
assign addr[59522]= -2090184478;
assign addr[59523]= -2098628387;
assign addr[59524]= -2106406677;
assign addr[59525]= -2113516878;
assign addr[59526]= -2119956737;
assign addr[59527]= -2125724211;
assign addr[59528]= -2130817471;
assign addr[59529]= -2135234901;
assign addr[59530]= -2138975100;
assign addr[59531]= -2142036881;
assign addr[59532]= -2144419275;
assign addr[59533]= -2146121524;
assign addr[59534]= -2147143090;
assign addr[59535]= -2147483648;
assign addr[59536]= -2147143090;
assign addr[59537]= -2146121524;
assign addr[59538]= -2144419275;
assign addr[59539]= -2142036881;
assign addr[59540]= -2138975100;
assign addr[59541]= -2135234901;
assign addr[59542]= -2130817471;
assign addr[59543]= -2125724211;
assign addr[59544]= -2119956737;
assign addr[59545]= -2113516878;
assign addr[59546]= -2106406677;
assign addr[59547]= -2098628387;
assign addr[59548]= -2090184478;
assign addr[59549]= -2081077626;
assign addr[59550]= -2071310720;
assign addr[59551]= -2060886858;
assign addr[59552]= -2049809346;
assign addr[59553]= -2038081698;
assign addr[59554]= -2025707632;
assign addr[59555]= -2012691075;
assign addr[59556]= -1999036154;
assign addr[59557]= -1984747199;
assign addr[59558]= -1969828744;
assign addr[59559]= -1954285520;
assign addr[59560]= -1938122457;
assign addr[59561]= -1921344681;
assign addr[59562]= -1903957513;
assign addr[59563]= -1885966468;
assign addr[59564]= -1867377253;
assign addr[59565]= -1848195763;
assign addr[59566]= -1828428082;
assign addr[59567]= -1808080480;
assign addr[59568]= -1787159411;
assign addr[59569]= -1765671509;
assign addr[59570]= -1743623590;
assign addr[59571]= -1721022648;
assign addr[59572]= -1697875851;
assign addr[59573]= -1674190539;
assign addr[59574]= -1649974225;
assign addr[59575]= -1625234591;
assign addr[59576]= -1599979481;
assign addr[59577]= -1574216908;
assign addr[59578]= -1547955041;
assign addr[59579]= -1521202211;
assign addr[59580]= -1493966902;
assign addr[59581]= -1466257752;
assign addr[59582]= -1438083551;
assign addr[59583]= -1409453233;
assign addr[59584]= -1380375881;
assign addr[59585]= -1350860716;
assign addr[59586]= -1320917099;
assign addr[59587]= -1290554528;
assign addr[59588]= -1259782632;
assign addr[59589]= -1228611172;
assign addr[59590]= -1197050035;
assign addr[59591]= -1165109230;
assign addr[59592]= -1132798888;
assign addr[59593]= -1100129257;
assign addr[59594]= -1067110699;
assign addr[59595]= -1033753687;
assign addr[59596]= -1000068799;
assign addr[59597]= -966066720;
assign addr[59598]= -931758235;
assign addr[59599]= -897154224;
assign addr[59600]= -862265664;
assign addr[59601]= -827103620;
assign addr[59602]= -791679244;
assign addr[59603]= -756003771;
assign addr[59604]= -720088517;
assign addr[59605]= -683944874;
assign addr[59606]= -647584304;
assign addr[59607]= -611018340;
assign addr[59608]= -574258580;
assign addr[59609]= -537316682;
assign addr[59610]= -500204365;
assign addr[59611]= -462933398;
assign addr[59612]= -425515602;
assign addr[59613]= -387962847;
assign addr[59614]= -350287041;
assign addr[59615]= -312500135;
assign addr[59616]= -274614114;
assign addr[59617]= -236640993;
assign addr[59618]= -198592817;
assign addr[59619]= -160481654;
assign addr[59620]= -122319591;
assign addr[59621]= -84118732;
assign addr[59622]= -45891193;
assign addr[59623]= -7649098;
assign addr[59624]= 30595422;
assign addr[59625]= 68830239;
assign addr[59626]= 107043224;
assign addr[59627]= 145222259;
assign addr[59628]= 183355234;
assign addr[59629]= 221430054;
assign addr[59630]= 259434643;
assign addr[59631]= 297356948;
assign addr[59632]= 335184940;
assign addr[59633]= 372906622;
assign addr[59634]= 410510029;
assign addr[59635]= 447983235;
assign addr[59636]= 485314355;
assign addr[59637]= 522491548;
assign addr[59638]= 559503022;
assign addr[59639]= 596337040;
assign addr[59640]= 632981917;
assign addr[59641]= 669426032;
assign addr[59642]= 705657826;
assign addr[59643]= 741665807;
assign addr[59644]= 777438554;
assign addr[59645]= 812964722;
assign addr[59646]= 848233042;
assign addr[59647]= 883232329;
assign addr[59648]= 917951481;
assign addr[59649]= 952379488;
assign addr[59650]= 986505429;
assign addr[59651]= 1020318481;
assign addr[59652]= 1053807919;
assign addr[59653]= 1086963121;
assign addr[59654]= 1119773573;
assign addr[59655]= 1152228866;
assign addr[59656]= 1184318708;
assign addr[59657]= 1216032921;
assign addr[59658]= 1247361445;
assign addr[59659]= 1278294345;
assign addr[59660]= 1308821808;
assign addr[59661]= 1338934154;
assign addr[59662]= 1368621831;
assign addr[59663]= 1397875423;
assign addr[59664]= 1426685652;
assign addr[59665]= 1455043381;
assign addr[59666]= 1482939614;
assign addr[59667]= 1510365504;
assign addr[59668]= 1537312353;
assign addr[59669]= 1563771613;
assign addr[59670]= 1589734894;
assign addr[59671]= 1615193959;
assign addr[59672]= 1640140734;
assign addr[59673]= 1664567307;
assign addr[59674]= 1688465931;
assign addr[59675]= 1711829025;
assign addr[59676]= 1734649179;
assign addr[59677]= 1756919156;
assign addr[59678]= 1778631892;
assign addr[59679]= 1799780501;
assign addr[59680]= 1820358275;
assign addr[59681]= 1840358687;
assign addr[59682]= 1859775393;
assign addr[59683]= 1878602237;
assign addr[59684]= 1896833245;
assign addr[59685]= 1914462636;
assign addr[59686]= 1931484818;
assign addr[59687]= 1947894393;
assign addr[59688]= 1963686155;
assign addr[59689]= 1978855097;
assign addr[59690]= 1993396407;
assign addr[59691]= 2007305472;
assign addr[59692]= 2020577882;
assign addr[59693]= 2033209426;
assign addr[59694]= 2045196100;
assign addr[59695]= 2056534099;
assign addr[59696]= 2067219829;
assign addr[59697]= 2077249901;
assign addr[59698]= 2086621133;
assign addr[59699]= 2095330553;
assign addr[59700]= 2103375398;
assign addr[59701]= 2110753117;
assign addr[59702]= 2117461370;
assign addr[59703]= 2123498030;
assign addr[59704]= 2128861181;
assign addr[59705]= 2133549123;
assign addr[59706]= 2137560369;
assign addr[59707]= 2140893646;
assign addr[59708]= 2143547897;
assign addr[59709]= 2145522281;
assign addr[59710]= 2146816171;
assign addr[59711]= 2147429158;
assign addr[59712]= 2147361045;
assign addr[59713]= 2146611856;
assign addr[59714]= 2145181827;
assign addr[59715]= 2143071413;
assign addr[59716]= 2140281282;
assign addr[59717]= 2136812319;
assign addr[59718]= 2132665626;
assign addr[59719]= 2127842516;
assign addr[59720]= 2122344521;
assign addr[59721]= 2116173382;
assign addr[59722]= 2109331059;
assign addr[59723]= 2101819720;
assign addr[59724]= 2093641749;
assign addr[59725]= 2084799740;
assign addr[59726]= 2075296495;
assign addr[59727]= 2065135031;
assign addr[59728]= 2054318569;
assign addr[59729]= 2042850540;
assign addr[59730]= 2030734582;
assign addr[59731]= 2017974537;
assign addr[59732]= 2004574453;
assign addr[59733]= 1990538579;
assign addr[59734]= 1975871368;
assign addr[59735]= 1960577471;
assign addr[59736]= 1944661739;
assign addr[59737]= 1928129220;
assign addr[59738]= 1910985158;
assign addr[59739]= 1893234990;
assign addr[59740]= 1874884346;
assign addr[59741]= 1855939047;
assign addr[59742]= 1836405100;
assign addr[59743]= 1816288703;
assign addr[59744]= 1795596234;
assign addr[59745]= 1774334257;
assign addr[59746]= 1752509516;
assign addr[59747]= 1730128933;
assign addr[59748]= 1707199606;
assign addr[59749]= 1683728808;
assign addr[59750]= 1659723983;
assign addr[59751]= 1635192744;
assign addr[59752]= 1610142873;
assign addr[59753]= 1584582314;
assign addr[59754]= 1558519173;
assign addr[59755]= 1531961719;
assign addr[59756]= 1504918373;
assign addr[59757]= 1477397714;
assign addr[59758]= 1449408469;
assign addr[59759]= 1420959516;
assign addr[59760]= 1392059879;
assign addr[59761]= 1362718723;
assign addr[59762]= 1332945355;
assign addr[59763]= 1302749217;
assign addr[59764]= 1272139887;
assign addr[59765]= 1241127074;
assign addr[59766]= 1209720613;
assign addr[59767]= 1177930466;
assign addr[59768]= 1145766716;
assign addr[59769]= 1113239564;
assign addr[59770]= 1080359326;
assign addr[59771]= 1047136432;
assign addr[59772]= 1013581418;
assign addr[59773]= 979704927;
assign addr[59774]= 945517704;
assign addr[59775]= 911030591;
assign addr[59776]= 876254528;
assign addr[59777]= 841200544;
assign addr[59778]= 805879757;
assign addr[59779]= 770303369;
assign addr[59780]= 734482665;
assign addr[59781]= 698429006;
assign addr[59782]= 662153826;
assign addr[59783]= 625668632;
assign addr[59784]= 588984994;
assign addr[59785]= 552114549;
assign addr[59786]= 515068990;
assign addr[59787]= 477860067;
assign addr[59788]= 440499581;
assign addr[59789]= 402999383;
assign addr[59790]= 365371365;
assign addr[59791]= 327627463;
assign addr[59792]= 289779648;
assign addr[59793]= 251839923;
assign addr[59794]= 213820322;
assign addr[59795]= 175732905;
assign addr[59796]= 137589750;
assign addr[59797]= 99402956;
assign addr[59798]= 61184634;
assign addr[59799]= 22946906;
assign addr[59800]= -15298099;
assign addr[59801]= -53538253;
assign addr[59802]= -91761426;
assign addr[59803]= -129955495;
assign addr[59804]= -168108346;
assign addr[59805]= -206207878;
assign addr[59806]= -244242007;
assign addr[59807]= -282198671;
assign addr[59808]= -320065829;
assign addr[59809]= -357831473;
assign addr[59810]= -395483624;
assign addr[59811]= -433010339;
assign addr[59812]= -470399716;
assign addr[59813]= -507639898;
assign addr[59814]= -544719071;
assign addr[59815]= -581625477;
assign addr[59816]= -618347408;
assign addr[59817]= -654873219;
assign addr[59818]= -691191324;
assign addr[59819]= -727290205;
assign addr[59820]= -763158411;
assign addr[59821]= -798784567;
assign addr[59822]= -834157373;
assign addr[59823]= -869265610;
assign addr[59824]= -904098143;
assign addr[59825]= -938643924;
assign addr[59826]= -972891995;
assign addr[59827]= -1006831495;
assign addr[59828]= -1040451659;
assign addr[59829]= -1073741824;
assign addr[59830]= -1106691431;
assign addr[59831]= -1139290029;
assign addr[59832]= -1171527280;
assign addr[59833]= -1203392958;
assign addr[59834]= -1234876957;
assign addr[59835]= -1265969291;
assign addr[59836]= -1296660098;
assign addr[59837]= -1326939644;
assign addr[59838]= -1356798326;
assign addr[59839]= -1386226674;
assign addr[59840]= -1415215352;
assign addr[59841]= -1443755168;
assign addr[59842]= -1471837070;
assign addr[59843]= -1499452149;
assign addr[59844]= -1526591649;
assign addr[59845]= -1553246960;
assign addr[59846]= -1579409630;
assign addr[59847]= -1605071359;
assign addr[59848]= -1630224009;
assign addr[59849]= -1654859602;
assign addr[59850]= -1678970324;
assign addr[59851]= -1702548529;
assign addr[59852]= -1725586737;
assign addr[59853]= -1748077642;
assign addr[59854]= -1770014111;
assign addr[59855]= -1791389186;
assign addr[59856]= -1812196087;
assign addr[59857]= -1832428215;
assign addr[59858]= -1852079154;
assign addr[59859]= -1871142669;
assign addr[59860]= -1889612716;
assign addr[59861]= -1907483436;
assign addr[59862]= -1924749160;
assign addr[59863]= -1941404413;
assign addr[59864]= -1957443913;
assign addr[59865]= -1972862571;
assign addr[59866]= -1987655498;
assign addr[59867]= -2001818002;
assign addr[59868]= -2015345591;
assign addr[59869]= -2028233973;
assign addr[59870]= -2040479063;
assign addr[59871]= -2052076975;
assign addr[59872]= -2063024031;
assign addr[59873]= -2073316760;
assign addr[59874]= -2082951896;
assign addr[59875]= -2091926384;
assign addr[59876]= -2100237377;
assign addr[59877]= -2107882239;
assign addr[59878]= -2114858546;
assign addr[59879]= -2121164085;
assign addr[59880]= -2126796855;
assign addr[59881]= -2131755071;
assign addr[59882]= -2136037160;
assign addr[59883]= -2139641764;
assign addr[59884]= -2142567738;
assign addr[59885]= -2144814157;
assign addr[59886]= -2146380306;
assign addr[59887]= -2147265689;
assign addr[59888]= -2147470025;
assign addr[59889]= -2146993250;
assign addr[59890]= -2145835515;
assign addr[59891]= -2143997187;
assign addr[59892]= -2141478848;
assign addr[59893]= -2138281298;
assign addr[59894]= -2134405552;
assign addr[59895]= -2129852837;
assign addr[59896]= -2124624598;
assign addr[59897]= -2118722494;
assign addr[59898]= -2112148396;
assign addr[59899]= -2104904390;
assign addr[59900]= -2096992772;
assign addr[59901]= -2088416053;
assign addr[59902]= -2079176953;
assign addr[59903]= -2069278401;
assign addr[59904]= -2058723538;
assign addr[59905]= -2047515711;
assign addr[59906]= -2035658475;
assign addr[59907]= -2023155591;
assign addr[59908]= -2010011024;
assign addr[59909]= -1996228943;
assign addr[59910]= -1981813720;
assign addr[59911]= -1966769926;
assign addr[59912]= -1951102334;
assign addr[59913]= -1934815911;
assign addr[59914]= -1917915825;
assign addr[59915]= -1900407434;
assign addr[59916]= -1882296293;
assign addr[59917]= -1863588145;
assign addr[59918]= -1844288924;
assign addr[59919]= -1824404752;
assign addr[59920]= -1803941934;
assign addr[59921]= -1782906961;
assign addr[59922]= -1761306505;
assign addr[59923]= -1739147417;
assign addr[59924]= -1716436725;
assign addr[59925]= -1693181631;
assign addr[59926]= -1669389513;
assign addr[59927]= -1645067915;
assign addr[59928]= -1620224553;
assign addr[59929]= -1594867305;
assign addr[59930]= -1569004214;
assign addr[59931]= -1542643483;
assign addr[59932]= -1515793473;
assign addr[59933]= -1488462700;
assign addr[59934]= -1460659832;
assign addr[59935]= -1432393688;
assign addr[59936]= -1403673233;
assign addr[59937]= -1374507575;
assign addr[59938]= -1344905966;
assign addr[59939]= -1314877795;
assign addr[59940]= -1284432584;
assign addr[59941]= -1253579991;
assign addr[59942]= -1222329801;
assign addr[59943]= -1190691925;
assign addr[59944]= -1158676398;
assign addr[59945]= -1126293375;
assign addr[59946]= -1093553126;
assign addr[59947]= -1060466036;
assign addr[59948]= -1027042599;
assign addr[59949]= -993293415;
assign addr[59950]= -959229189;
assign addr[59951]= -924860725;
assign addr[59952]= -890198924;
assign addr[59953]= -855254778;
assign addr[59954]= -820039373;
assign addr[59955]= -784563876;
assign addr[59956]= -748839539;
assign addr[59957]= -712877694;
assign addr[59958]= -676689746;
assign addr[59959]= -640287172;
assign addr[59960]= -603681519;
assign addr[59961]= -566884397;
assign addr[59962]= -529907477;
assign addr[59963]= -492762486;
assign addr[59964]= -455461206;
assign addr[59965]= -418015468;
assign addr[59966]= -380437148;
assign addr[59967]= -342738165;
assign addr[59968]= -304930476;
assign addr[59969]= -267026072;
assign addr[59970]= -229036977;
assign addr[59971]= -190975237;
assign addr[59972]= -152852926;
assign addr[59973]= -114682135;
assign addr[59974]= -76474970;
assign addr[59975]= -38243550;
assign addr[59976]= 0;
assign addr[59977]= 38243550;
assign addr[59978]= 76474970;
assign addr[59979]= 114682135;
assign addr[59980]= 152852926;
assign addr[59981]= 190975237;
assign addr[59982]= 229036977;
assign addr[59983]= 267026072;
assign addr[59984]= 304930476;
assign addr[59985]= 342738165;
assign addr[59986]= 380437148;
assign addr[59987]= 418015468;
assign addr[59988]= 455461206;
assign addr[59989]= 492762486;
assign addr[59990]= 529907477;
assign addr[59991]= 566884397;
assign addr[59992]= 603681519;
assign addr[59993]= 640287172;
assign addr[59994]= 676689746;
assign addr[59995]= 712877694;
assign addr[59996]= 748839539;
assign addr[59997]= 784563876;
assign addr[59998]= 820039373;
assign addr[59999]= 855254778;
assign addr[60000]= 890198924;
assign addr[60001]= 924860725;
assign addr[60002]= 959229189;
assign addr[60003]= 993293415;
assign addr[60004]= 1027042599;
assign addr[60005]= 1060466036;
assign addr[60006]= 1093553126;
assign addr[60007]= 1126293375;
assign addr[60008]= 1158676398;
assign addr[60009]= 1190691925;
assign addr[60010]= 1222329801;
assign addr[60011]= 1253579991;
assign addr[60012]= 1284432584;
assign addr[60013]= 1314877795;
assign addr[60014]= 1344905966;
assign addr[60015]= 1374507575;
assign addr[60016]= 1403673233;
assign addr[60017]= 1432393688;
assign addr[60018]= 1460659832;
assign addr[60019]= 1488462700;
assign addr[60020]= 1515793473;
assign addr[60021]= 1542643483;
assign addr[60022]= 1569004214;
assign addr[60023]= 1594867305;
assign addr[60024]= 1620224553;
assign addr[60025]= 1645067915;
assign addr[60026]= 1669389513;
assign addr[60027]= 1693181631;
assign addr[60028]= 1716436725;
assign addr[60029]= 1739147417;
assign addr[60030]= 1761306505;
assign addr[60031]= 1782906961;
assign addr[60032]= 1803941934;
assign addr[60033]= 1824404752;
assign addr[60034]= 1844288924;
assign addr[60035]= 1863588145;
assign addr[60036]= 1882296293;
assign addr[60037]= 1900407434;
assign addr[60038]= 1917915825;
assign addr[60039]= 1934815911;
assign addr[60040]= 1951102334;
assign addr[60041]= 1966769926;
assign addr[60042]= 1981813720;
assign addr[60043]= 1996228943;
assign addr[60044]= 2010011024;
assign addr[60045]= 2023155591;
assign addr[60046]= 2035658475;
assign addr[60047]= 2047515711;
assign addr[60048]= 2058723538;
assign addr[60049]= 2069278401;
assign addr[60050]= 2079176953;
assign addr[60051]= 2088416053;
assign addr[60052]= 2096992772;
assign addr[60053]= 2104904390;
assign addr[60054]= 2112148396;
assign addr[60055]= 2118722494;
assign addr[60056]= 2124624598;
assign addr[60057]= 2129852837;
assign addr[60058]= 2134405552;
assign addr[60059]= 2138281298;
assign addr[60060]= 2141478848;
assign addr[60061]= 2143997187;
assign addr[60062]= 2145835515;
assign addr[60063]= 2146993250;
assign addr[60064]= 2147470025;
assign addr[60065]= 2147265689;
assign addr[60066]= 2146380306;
assign addr[60067]= 2144814157;
assign addr[60068]= 2142567738;
assign addr[60069]= 2139641764;
assign addr[60070]= 2136037160;
assign addr[60071]= 2131755071;
assign addr[60072]= 2126796855;
assign addr[60073]= 2121164085;
assign addr[60074]= 2114858546;
assign addr[60075]= 2107882239;
assign addr[60076]= 2100237377;
assign addr[60077]= 2091926384;
assign addr[60078]= 2082951896;
assign addr[60079]= 2073316760;
assign addr[60080]= 2063024031;
assign addr[60081]= 2052076975;
assign addr[60082]= 2040479063;
assign addr[60083]= 2028233973;
assign addr[60084]= 2015345591;
assign addr[60085]= 2001818002;
assign addr[60086]= 1987655498;
assign addr[60087]= 1972862571;
assign addr[60088]= 1957443913;
assign addr[60089]= 1941404413;
assign addr[60090]= 1924749160;
assign addr[60091]= 1907483436;
assign addr[60092]= 1889612716;
assign addr[60093]= 1871142669;
assign addr[60094]= 1852079154;
assign addr[60095]= 1832428215;
assign addr[60096]= 1812196087;
assign addr[60097]= 1791389186;
assign addr[60098]= 1770014111;
assign addr[60099]= 1748077642;
assign addr[60100]= 1725586737;
assign addr[60101]= 1702548529;
assign addr[60102]= 1678970324;
assign addr[60103]= 1654859602;
assign addr[60104]= 1630224009;
assign addr[60105]= 1605071359;
assign addr[60106]= 1579409630;
assign addr[60107]= 1553246960;
assign addr[60108]= 1526591649;
assign addr[60109]= 1499452149;
assign addr[60110]= 1471837070;
assign addr[60111]= 1443755168;
assign addr[60112]= 1415215352;
assign addr[60113]= 1386226674;
assign addr[60114]= 1356798326;
assign addr[60115]= 1326939644;
assign addr[60116]= 1296660098;
assign addr[60117]= 1265969291;
assign addr[60118]= 1234876957;
assign addr[60119]= 1203392958;
assign addr[60120]= 1171527280;
assign addr[60121]= 1139290029;
assign addr[60122]= 1106691431;
assign addr[60123]= 1073741824;
assign addr[60124]= 1040451659;
assign addr[60125]= 1006831495;
assign addr[60126]= 972891995;
assign addr[60127]= 938643924;
assign addr[60128]= 904098143;
assign addr[60129]= 869265610;
assign addr[60130]= 834157373;
assign addr[60131]= 798784567;
assign addr[60132]= 763158411;
assign addr[60133]= 727290205;
assign addr[60134]= 691191324;
assign addr[60135]= 654873219;
assign addr[60136]= 618347408;
assign addr[60137]= 581625477;
assign addr[60138]= 544719071;
assign addr[60139]= 507639898;
assign addr[60140]= 470399716;
assign addr[60141]= 433010339;
assign addr[60142]= 395483624;
assign addr[60143]= 357831473;
assign addr[60144]= 320065829;
assign addr[60145]= 282198671;
assign addr[60146]= 244242007;
assign addr[60147]= 206207878;
assign addr[60148]= 168108346;
assign addr[60149]= 129955495;
assign addr[60150]= 91761426;
assign addr[60151]= 53538253;
assign addr[60152]= 15298099;
assign addr[60153]= -22946906;
assign addr[60154]= -61184634;
assign addr[60155]= -99402956;
assign addr[60156]= -137589750;
assign addr[60157]= -175732905;
assign addr[60158]= -213820322;
assign addr[60159]= -251839923;
assign addr[60160]= -289779648;
assign addr[60161]= -327627463;
assign addr[60162]= -365371365;
assign addr[60163]= -402999383;
assign addr[60164]= -440499581;
assign addr[60165]= -477860067;
assign addr[60166]= -515068990;
assign addr[60167]= -552114549;
assign addr[60168]= -588984994;
assign addr[60169]= -625668632;
assign addr[60170]= -662153826;
assign addr[60171]= -698429006;
assign addr[60172]= -734482665;
assign addr[60173]= -770303369;
assign addr[60174]= -805879757;
assign addr[60175]= -841200544;
assign addr[60176]= -876254528;
assign addr[60177]= -911030591;
assign addr[60178]= -945517704;
assign addr[60179]= -979704927;
assign addr[60180]= -1013581418;
assign addr[60181]= -1047136432;
assign addr[60182]= -1080359326;
assign addr[60183]= -1113239564;
assign addr[60184]= -1145766716;
assign addr[60185]= -1177930466;
assign addr[60186]= -1209720613;
assign addr[60187]= -1241127074;
assign addr[60188]= -1272139887;
assign addr[60189]= -1302749217;
assign addr[60190]= -1332945355;
assign addr[60191]= -1362718723;
assign addr[60192]= -1392059879;
assign addr[60193]= -1420959516;
assign addr[60194]= -1449408469;
assign addr[60195]= -1477397714;
assign addr[60196]= -1504918373;
assign addr[60197]= -1531961719;
assign addr[60198]= -1558519173;
assign addr[60199]= -1584582314;
assign addr[60200]= -1610142873;
assign addr[60201]= -1635192744;
assign addr[60202]= -1659723983;
assign addr[60203]= -1683728808;
assign addr[60204]= -1707199606;
assign addr[60205]= -1730128933;
assign addr[60206]= -1752509516;
assign addr[60207]= -1774334257;
assign addr[60208]= -1795596234;
assign addr[60209]= -1816288703;
assign addr[60210]= -1836405100;
assign addr[60211]= -1855939047;
assign addr[60212]= -1874884346;
assign addr[60213]= -1893234990;
assign addr[60214]= -1910985158;
assign addr[60215]= -1928129220;
assign addr[60216]= -1944661739;
assign addr[60217]= -1960577471;
assign addr[60218]= -1975871368;
assign addr[60219]= -1990538579;
assign addr[60220]= -2004574453;
assign addr[60221]= -2017974537;
assign addr[60222]= -2030734582;
assign addr[60223]= -2042850540;
assign addr[60224]= -2054318569;
assign addr[60225]= -2065135031;
assign addr[60226]= -2075296495;
assign addr[60227]= -2084799740;
assign addr[60228]= -2093641749;
assign addr[60229]= -2101819720;
assign addr[60230]= -2109331059;
assign addr[60231]= -2116173382;
assign addr[60232]= -2122344521;
assign addr[60233]= -2127842516;
assign addr[60234]= -2132665626;
assign addr[60235]= -2136812319;
assign addr[60236]= -2140281282;
assign addr[60237]= -2143071413;
assign addr[60238]= -2145181827;
assign addr[60239]= -2146611856;
assign addr[60240]= -2147361045;
assign addr[60241]= -2147429158;
assign addr[60242]= -2146816171;
assign addr[60243]= -2145522281;
assign addr[60244]= -2143547897;
assign addr[60245]= -2140893646;
assign addr[60246]= -2137560369;
assign addr[60247]= -2133549123;
assign addr[60248]= -2128861181;
assign addr[60249]= -2123498030;
assign addr[60250]= -2117461370;
assign addr[60251]= -2110753117;
assign addr[60252]= -2103375398;
assign addr[60253]= -2095330553;
assign addr[60254]= -2086621133;
assign addr[60255]= -2077249901;
assign addr[60256]= -2067219829;
assign addr[60257]= -2056534099;
assign addr[60258]= -2045196100;
assign addr[60259]= -2033209426;
assign addr[60260]= -2020577882;
assign addr[60261]= -2007305472;
assign addr[60262]= -1993396407;
assign addr[60263]= -1978855097;
assign addr[60264]= -1963686155;
assign addr[60265]= -1947894393;
assign addr[60266]= -1931484818;
assign addr[60267]= -1914462636;
assign addr[60268]= -1896833245;
assign addr[60269]= -1878602237;
assign addr[60270]= -1859775393;
assign addr[60271]= -1840358687;
assign addr[60272]= -1820358275;
assign addr[60273]= -1799780501;
assign addr[60274]= -1778631892;
assign addr[60275]= -1756919156;
assign addr[60276]= -1734649179;
assign addr[60277]= -1711829025;
assign addr[60278]= -1688465931;
assign addr[60279]= -1664567307;
assign addr[60280]= -1640140734;
assign addr[60281]= -1615193959;
assign addr[60282]= -1589734894;
assign addr[60283]= -1563771613;
assign addr[60284]= -1537312353;
assign addr[60285]= -1510365504;
assign addr[60286]= -1482939614;
assign addr[60287]= -1455043381;
assign addr[60288]= -1426685652;
assign addr[60289]= -1397875423;
assign addr[60290]= -1368621831;
assign addr[60291]= -1338934154;
assign addr[60292]= -1308821808;
assign addr[60293]= -1278294345;
assign addr[60294]= -1247361445;
assign addr[60295]= -1216032921;
assign addr[60296]= -1184318708;
assign addr[60297]= -1152228866;
assign addr[60298]= -1119773573;
assign addr[60299]= -1086963121;
assign addr[60300]= -1053807919;
assign addr[60301]= -1020318481;
assign addr[60302]= -986505429;
assign addr[60303]= -952379488;
assign addr[60304]= -917951481;
assign addr[60305]= -883232329;
assign addr[60306]= -848233042;
assign addr[60307]= -812964722;
assign addr[60308]= -777438554;
assign addr[60309]= -741665807;
assign addr[60310]= -705657826;
assign addr[60311]= -669426032;
assign addr[60312]= -632981917;
assign addr[60313]= -596337040;
assign addr[60314]= -559503022;
assign addr[60315]= -522491548;
assign addr[60316]= -485314355;
assign addr[60317]= -447983235;
assign addr[60318]= -410510029;
assign addr[60319]= -372906622;
assign addr[60320]= -335184940;
assign addr[60321]= -297356948;
assign addr[60322]= -259434643;
assign addr[60323]= -221430054;
assign addr[60324]= -183355234;
assign addr[60325]= -145222259;
assign addr[60326]= -107043224;
assign addr[60327]= -68830239;
assign addr[60328]= -30595422;
assign addr[60329]= 7649098;
assign addr[60330]= 45891193;
assign addr[60331]= 84118732;
assign addr[60332]= 122319591;
assign addr[60333]= 160481654;
assign addr[60334]= 198592817;
assign addr[60335]= 236640993;
assign addr[60336]= 274614114;
assign addr[60337]= 312500135;
assign addr[60338]= 350287041;
assign addr[60339]= 387962847;
assign addr[60340]= 425515602;
assign addr[60341]= 462933398;
assign addr[60342]= 500204365;
assign addr[60343]= 537316682;
assign addr[60344]= 574258580;
assign addr[60345]= 611018340;
assign addr[60346]= 647584304;
assign addr[60347]= 683944874;
assign addr[60348]= 720088517;
assign addr[60349]= 756003771;
assign addr[60350]= 791679244;
assign addr[60351]= 827103620;
assign addr[60352]= 862265664;
assign addr[60353]= 897154224;
assign addr[60354]= 931758235;
assign addr[60355]= 966066720;
assign addr[60356]= 1000068799;
assign addr[60357]= 1033753687;
assign addr[60358]= 1067110699;
assign addr[60359]= 1100129257;
assign addr[60360]= 1132798888;
assign addr[60361]= 1165109230;
assign addr[60362]= 1197050035;
assign addr[60363]= 1228611172;
assign addr[60364]= 1259782632;
assign addr[60365]= 1290554528;
assign addr[60366]= 1320917099;
assign addr[60367]= 1350860716;
assign addr[60368]= 1380375881;
assign addr[60369]= 1409453233;
assign addr[60370]= 1438083551;
assign addr[60371]= 1466257752;
assign addr[60372]= 1493966902;
assign addr[60373]= 1521202211;
assign addr[60374]= 1547955041;
assign addr[60375]= 1574216908;
assign addr[60376]= 1599979481;
assign addr[60377]= 1625234591;
assign addr[60378]= 1649974225;
assign addr[60379]= 1674190539;
assign addr[60380]= 1697875851;
assign addr[60381]= 1721022648;
assign addr[60382]= 1743623590;
assign addr[60383]= 1765671509;
assign addr[60384]= 1787159411;
assign addr[60385]= 1808080480;
assign addr[60386]= 1828428082;
assign addr[60387]= 1848195763;
assign addr[60388]= 1867377253;
assign addr[60389]= 1885966468;
assign addr[60390]= 1903957513;
assign addr[60391]= 1921344681;
assign addr[60392]= 1938122457;
assign addr[60393]= 1954285520;
assign addr[60394]= 1969828744;
assign addr[60395]= 1984747199;
assign addr[60396]= 1999036154;
assign addr[60397]= 2012691075;
assign addr[60398]= 2025707632;
assign addr[60399]= 2038081698;
assign addr[60400]= 2049809346;
assign addr[60401]= 2060886858;
assign addr[60402]= 2071310720;
assign addr[60403]= 2081077626;
assign addr[60404]= 2090184478;
assign addr[60405]= 2098628387;
assign addr[60406]= 2106406677;
assign addr[60407]= 2113516878;
assign addr[60408]= 2119956737;
assign addr[60409]= 2125724211;
assign addr[60410]= 2130817471;
assign addr[60411]= 2135234901;
assign addr[60412]= 2138975100;
assign addr[60413]= 2142036881;
assign addr[60414]= 2144419275;
assign addr[60415]= 2146121524;
assign addr[60416]= 2147143090;
assign addr[60417]= 2147483648;
assign addr[60418]= 2147143090;
assign addr[60419]= 2146121524;
assign addr[60420]= 2144419275;
assign addr[60421]= 2142036881;
assign addr[60422]= 2138975100;
assign addr[60423]= 2135234901;
assign addr[60424]= 2130817471;
assign addr[60425]= 2125724211;
assign addr[60426]= 2119956737;
assign addr[60427]= 2113516878;
assign addr[60428]= 2106406677;
assign addr[60429]= 2098628387;
assign addr[60430]= 2090184478;
assign addr[60431]= 2081077626;
assign addr[60432]= 2071310720;
assign addr[60433]= 2060886858;
assign addr[60434]= 2049809346;
assign addr[60435]= 2038081698;
assign addr[60436]= 2025707632;
assign addr[60437]= 2012691075;
assign addr[60438]= 1999036154;
assign addr[60439]= 1984747199;
assign addr[60440]= 1969828744;
assign addr[60441]= 1954285520;
assign addr[60442]= 1938122457;
assign addr[60443]= 1921344681;
assign addr[60444]= 1903957513;
assign addr[60445]= 1885966468;
assign addr[60446]= 1867377253;
assign addr[60447]= 1848195763;
assign addr[60448]= 1828428082;
assign addr[60449]= 1808080480;
assign addr[60450]= 1787159411;
assign addr[60451]= 1765671509;
assign addr[60452]= 1743623590;
assign addr[60453]= 1721022648;
assign addr[60454]= 1697875851;
assign addr[60455]= 1674190539;
assign addr[60456]= 1649974225;
assign addr[60457]= 1625234591;
assign addr[60458]= 1599979481;
assign addr[60459]= 1574216908;
assign addr[60460]= 1547955041;
assign addr[60461]= 1521202211;
assign addr[60462]= 1493966902;
assign addr[60463]= 1466257752;
assign addr[60464]= 1438083551;
assign addr[60465]= 1409453233;
assign addr[60466]= 1380375881;
assign addr[60467]= 1350860716;
assign addr[60468]= 1320917099;
assign addr[60469]= 1290554528;
assign addr[60470]= 1259782632;
assign addr[60471]= 1228611172;
assign addr[60472]= 1197050035;
assign addr[60473]= 1165109230;
assign addr[60474]= 1132798888;
assign addr[60475]= 1100129257;
assign addr[60476]= 1067110699;
assign addr[60477]= 1033753687;
assign addr[60478]= 1000068799;
assign addr[60479]= 966066720;
assign addr[60480]= 931758235;
assign addr[60481]= 897154224;
assign addr[60482]= 862265664;
assign addr[60483]= 827103620;
assign addr[60484]= 791679244;
assign addr[60485]= 756003771;
assign addr[60486]= 720088517;
assign addr[60487]= 683944874;
assign addr[60488]= 647584304;
assign addr[60489]= 611018340;
assign addr[60490]= 574258580;
assign addr[60491]= 537316682;
assign addr[60492]= 500204365;
assign addr[60493]= 462933398;
assign addr[60494]= 425515602;
assign addr[60495]= 387962847;
assign addr[60496]= 350287041;
assign addr[60497]= 312500135;
assign addr[60498]= 274614114;
assign addr[60499]= 236640993;
assign addr[60500]= 198592817;
assign addr[60501]= 160481654;
assign addr[60502]= 122319591;
assign addr[60503]= 84118732;
assign addr[60504]= 45891193;
assign addr[60505]= 7649098;
assign addr[60506]= -30595422;
assign addr[60507]= -68830239;
assign addr[60508]= -107043224;
assign addr[60509]= -145222259;
assign addr[60510]= -183355234;
assign addr[60511]= -221430054;
assign addr[60512]= -259434643;
assign addr[60513]= -297356948;
assign addr[60514]= -335184940;
assign addr[60515]= -372906622;
assign addr[60516]= -410510029;
assign addr[60517]= -447983235;
assign addr[60518]= -485314355;
assign addr[60519]= -522491548;
assign addr[60520]= -559503022;
assign addr[60521]= -596337040;
assign addr[60522]= -632981917;
assign addr[60523]= -669426032;
assign addr[60524]= -705657826;
assign addr[60525]= -741665807;
assign addr[60526]= -777438554;
assign addr[60527]= -812964722;
assign addr[60528]= -848233042;
assign addr[60529]= -883232329;
assign addr[60530]= -917951481;
assign addr[60531]= -952379488;
assign addr[60532]= -986505429;
assign addr[60533]= -1020318481;
assign addr[60534]= -1053807919;
assign addr[60535]= -1086963121;
assign addr[60536]= -1119773573;
assign addr[60537]= -1152228866;
assign addr[60538]= -1184318708;
assign addr[60539]= -1216032921;
assign addr[60540]= -1247361445;
assign addr[60541]= -1278294345;
assign addr[60542]= -1308821808;
assign addr[60543]= -1338934154;
assign addr[60544]= -1368621831;
assign addr[60545]= -1397875423;
assign addr[60546]= -1426685652;
assign addr[60547]= -1455043381;
assign addr[60548]= -1482939614;
assign addr[60549]= -1510365504;
assign addr[60550]= -1537312353;
assign addr[60551]= -1563771613;
assign addr[60552]= -1589734894;
assign addr[60553]= -1615193959;
assign addr[60554]= -1640140734;
assign addr[60555]= -1664567307;
assign addr[60556]= -1688465931;
assign addr[60557]= -1711829025;
assign addr[60558]= -1734649179;
assign addr[60559]= -1756919156;
assign addr[60560]= -1778631892;
assign addr[60561]= -1799780501;
assign addr[60562]= -1820358275;
assign addr[60563]= -1840358687;
assign addr[60564]= -1859775393;
assign addr[60565]= -1878602237;
assign addr[60566]= -1896833245;
assign addr[60567]= -1914462636;
assign addr[60568]= -1931484818;
assign addr[60569]= -1947894393;
assign addr[60570]= -1963686155;
assign addr[60571]= -1978855097;
assign addr[60572]= -1993396407;
assign addr[60573]= -2007305472;
assign addr[60574]= -2020577882;
assign addr[60575]= -2033209426;
assign addr[60576]= -2045196100;
assign addr[60577]= -2056534099;
assign addr[60578]= -2067219829;
assign addr[60579]= -2077249901;
assign addr[60580]= -2086621133;
assign addr[60581]= -2095330553;
assign addr[60582]= -2103375398;
assign addr[60583]= -2110753117;
assign addr[60584]= -2117461370;
assign addr[60585]= -2123498030;
assign addr[60586]= -2128861181;
assign addr[60587]= -2133549123;
assign addr[60588]= -2137560369;
assign addr[60589]= -2140893646;
assign addr[60590]= -2143547897;
assign addr[60591]= -2145522281;
assign addr[60592]= -2146816171;
assign addr[60593]= -2147429158;
assign addr[60594]= -2147361045;
assign addr[60595]= -2146611856;
assign addr[60596]= -2145181827;
assign addr[60597]= -2143071413;
assign addr[60598]= -2140281282;
assign addr[60599]= -2136812319;
assign addr[60600]= -2132665626;
assign addr[60601]= -2127842516;
assign addr[60602]= -2122344521;
assign addr[60603]= -2116173382;
assign addr[60604]= -2109331059;
assign addr[60605]= -2101819720;
assign addr[60606]= -2093641749;
assign addr[60607]= -2084799740;
assign addr[60608]= -2075296495;
assign addr[60609]= -2065135031;
assign addr[60610]= -2054318569;
assign addr[60611]= -2042850540;
assign addr[60612]= -2030734582;
assign addr[60613]= -2017974537;
assign addr[60614]= -2004574453;
assign addr[60615]= -1990538579;
assign addr[60616]= -1975871368;
assign addr[60617]= -1960577471;
assign addr[60618]= -1944661739;
assign addr[60619]= -1928129220;
assign addr[60620]= -1910985158;
assign addr[60621]= -1893234990;
assign addr[60622]= -1874884346;
assign addr[60623]= -1855939047;
assign addr[60624]= -1836405100;
assign addr[60625]= -1816288703;
assign addr[60626]= -1795596234;
assign addr[60627]= -1774334257;
assign addr[60628]= -1752509516;
assign addr[60629]= -1730128933;
assign addr[60630]= -1707199606;
assign addr[60631]= -1683728808;
assign addr[60632]= -1659723983;
assign addr[60633]= -1635192744;
assign addr[60634]= -1610142873;
assign addr[60635]= -1584582314;
assign addr[60636]= -1558519173;
assign addr[60637]= -1531961719;
assign addr[60638]= -1504918373;
assign addr[60639]= -1477397714;
assign addr[60640]= -1449408469;
assign addr[60641]= -1420959516;
assign addr[60642]= -1392059879;
assign addr[60643]= -1362718723;
assign addr[60644]= -1332945355;
assign addr[60645]= -1302749217;
assign addr[60646]= -1272139887;
assign addr[60647]= -1241127074;
assign addr[60648]= -1209720613;
assign addr[60649]= -1177930466;
assign addr[60650]= -1145766716;
assign addr[60651]= -1113239564;
assign addr[60652]= -1080359326;
assign addr[60653]= -1047136432;
assign addr[60654]= -1013581418;
assign addr[60655]= -979704927;
assign addr[60656]= -945517704;
assign addr[60657]= -911030591;
assign addr[60658]= -876254528;
assign addr[60659]= -841200544;
assign addr[60660]= -805879757;
assign addr[60661]= -770303369;
assign addr[60662]= -734482665;
assign addr[60663]= -698429006;
assign addr[60664]= -662153826;
assign addr[60665]= -625668632;
assign addr[60666]= -588984994;
assign addr[60667]= -552114549;
assign addr[60668]= -515068990;
assign addr[60669]= -477860067;
assign addr[60670]= -440499581;
assign addr[60671]= -402999383;
assign addr[60672]= -365371365;
assign addr[60673]= -327627463;
assign addr[60674]= -289779648;
assign addr[60675]= -251839923;
assign addr[60676]= -213820322;
assign addr[60677]= -175732905;
assign addr[60678]= -137589750;
assign addr[60679]= -99402956;
assign addr[60680]= -61184634;
assign addr[60681]= -22946906;
assign addr[60682]= 15298099;
assign addr[60683]= 53538253;
assign addr[60684]= 91761426;
assign addr[60685]= 129955495;
assign addr[60686]= 168108346;
assign addr[60687]= 206207878;
assign addr[60688]= 244242007;
assign addr[60689]= 282198671;
assign addr[60690]= 320065829;
assign addr[60691]= 357831473;
assign addr[60692]= 395483624;
assign addr[60693]= 433010339;
assign addr[60694]= 470399716;
assign addr[60695]= 507639898;
assign addr[60696]= 544719071;
assign addr[60697]= 581625477;
assign addr[60698]= 618347408;
assign addr[60699]= 654873219;
assign addr[60700]= 691191324;
assign addr[60701]= 727290205;
assign addr[60702]= 763158411;
assign addr[60703]= 798784567;
assign addr[60704]= 834157373;
assign addr[60705]= 869265610;
assign addr[60706]= 904098143;
assign addr[60707]= 938643924;
assign addr[60708]= 972891995;
assign addr[60709]= 1006831495;
assign addr[60710]= 1040451659;
assign addr[60711]= 1073741824;
assign addr[60712]= 1106691431;
assign addr[60713]= 1139290029;
assign addr[60714]= 1171527280;
assign addr[60715]= 1203392958;
assign addr[60716]= 1234876957;
assign addr[60717]= 1265969291;
assign addr[60718]= 1296660098;
assign addr[60719]= 1326939644;
assign addr[60720]= 1356798326;
assign addr[60721]= 1386226674;
assign addr[60722]= 1415215352;
assign addr[60723]= 1443755168;
assign addr[60724]= 1471837070;
assign addr[60725]= 1499452149;
assign addr[60726]= 1526591649;
assign addr[60727]= 1553246960;
assign addr[60728]= 1579409630;
assign addr[60729]= 1605071359;
assign addr[60730]= 1630224009;
assign addr[60731]= 1654859602;
assign addr[60732]= 1678970324;
assign addr[60733]= 1702548529;
assign addr[60734]= 1725586737;
assign addr[60735]= 1748077642;
assign addr[60736]= 1770014111;
assign addr[60737]= 1791389186;
assign addr[60738]= 1812196087;
assign addr[60739]= 1832428215;
assign addr[60740]= 1852079154;
assign addr[60741]= 1871142669;
assign addr[60742]= 1889612716;
assign addr[60743]= 1907483436;
assign addr[60744]= 1924749160;
assign addr[60745]= 1941404413;
assign addr[60746]= 1957443913;
assign addr[60747]= 1972862571;
assign addr[60748]= 1987655498;
assign addr[60749]= 2001818002;
assign addr[60750]= 2015345591;
assign addr[60751]= 2028233973;
assign addr[60752]= 2040479063;
assign addr[60753]= 2052076975;
assign addr[60754]= 2063024031;
assign addr[60755]= 2073316760;
assign addr[60756]= 2082951896;
assign addr[60757]= 2091926384;
assign addr[60758]= 2100237377;
assign addr[60759]= 2107882239;
assign addr[60760]= 2114858546;
assign addr[60761]= 2121164085;
assign addr[60762]= 2126796855;
assign addr[60763]= 2131755071;
assign addr[60764]= 2136037160;
assign addr[60765]= 2139641764;
assign addr[60766]= 2142567738;
assign addr[60767]= 2144814157;
assign addr[60768]= 2146380306;
assign addr[60769]= 2147265689;
assign addr[60770]= 2147470025;
assign addr[60771]= 2146993250;
assign addr[60772]= 2145835515;
assign addr[60773]= 2143997187;
assign addr[60774]= 2141478848;
assign addr[60775]= 2138281298;
assign addr[60776]= 2134405552;
assign addr[60777]= 2129852837;
assign addr[60778]= 2124624598;
assign addr[60779]= 2118722494;
assign addr[60780]= 2112148396;
assign addr[60781]= 2104904390;
assign addr[60782]= 2096992772;
assign addr[60783]= 2088416053;
assign addr[60784]= 2079176953;
assign addr[60785]= 2069278401;
assign addr[60786]= 2058723538;
assign addr[60787]= 2047515711;
assign addr[60788]= 2035658475;
assign addr[60789]= 2023155591;
assign addr[60790]= 2010011024;
assign addr[60791]= 1996228943;
assign addr[60792]= 1981813720;
assign addr[60793]= 1966769926;
assign addr[60794]= 1951102334;
assign addr[60795]= 1934815911;
assign addr[60796]= 1917915825;
assign addr[60797]= 1900407434;
assign addr[60798]= 1882296293;
assign addr[60799]= 1863588145;
assign addr[60800]= 1844288924;
assign addr[60801]= 1824404752;
assign addr[60802]= 1803941934;
assign addr[60803]= 1782906961;
assign addr[60804]= 1761306505;
assign addr[60805]= 1739147417;
assign addr[60806]= 1716436725;
assign addr[60807]= 1693181631;
assign addr[60808]= 1669389513;
assign addr[60809]= 1645067915;
assign addr[60810]= 1620224553;
assign addr[60811]= 1594867305;
assign addr[60812]= 1569004214;
assign addr[60813]= 1542643483;
assign addr[60814]= 1515793473;
assign addr[60815]= 1488462700;
assign addr[60816]= 1460659832;
assign addr[60817]= 1432393688;
assign addr[60818]= 1403673233;
assign addr[60819]= 1374507575;
assign addr[60820]= 1344905966;
assign addr[60821]= 1314877795;
assign addr[60822]= 1284432584;
assign addr[60823]= 1253579991;
assign addr[60824]= 1222329801;
assign addr[60825]= 1190691925;
assign addr[60826]= 1158676398;
assign addr[60827]= 1126293375;
assign addr[60828]= 1093553126;
assign addr[60829]= 1060466036;
assign addr[60830]= 1027042599;
assign addr[60831]= 993293415;
assign addr[60832]= 959229189;
assign addr[60833]= 924860725;
assign addr[60834]= 890198924;
assign addr[60835]= 855254778;
assign addr[60836]= 820039373;
assign addr[60837]= 784563876;
assign addr[60838]= 748839539;
assign addr[60839]= 712877694;
assign addr[60840]= 676689746;
assign addr[60841]= 640287172;
assign addr[60842]= 603681519;
assign addr[60843]= 566884397;
assign addr[60844]= 529907477;
assign addr[60845]= 492762486;
assign addr[60846]= 455461206;
assign addr[60847]= 418015468;
assign addr[60848]= 380437148;
assign addr[60849]= 342738165;
assign addr[60850]= 304930476;
assign addr[60851]= 267026072;
assign addr[60852]= 229036977;
assign addr[60853]= 190975237;
assign addr[60854]= 152852926;
assign addr[60855]= 114682135;
assign addr[60856]= 76474970;
assign addr[60857]= 38243550;
assign addr[60858]= 0;
assign addr[60859]= -38243550;
assign addr[60860]= -76474970;
assign addr[60861]= -114682135;
assign addr[60862]= -152852926;
assign addr[60863]= -190975237;
assign addr[60864]= -229036977;
assign addr[60865]= -267026072;
assign addr[60866]= -304930476;
assign addr[60867]= -342738165;
assign addr[60868]= -380437148;
assign addr[60869]= -418015468;
assign addr[60870]= -455461206;
assign addr[60871]= -492762486;
assign addr[60872]= -529907477;
assign addr[60873]= -566884397;
assign addr[60874]= -603681519;
assign addr[60875]= -640287172;
assign addr[60876]= -676689746;
assign addr[60877]= -712877694;
assign addr[60878]= -748839539;
assign addr[60879]= -784563876;
assign addr[60880]= -820039373;
assign addr[60881]= -855254778;
assign addr[60882]= -890198924;
assign addr[60883]= -924860725;
assign addr[60884]= -959229189;
assign addr[60885]= -993293415;
assign addr[60886]= -1027042599;
assign addr[60887]= -1060466036;
assign addr[60888]= -1093553126;
assign addr[60889]= -1126293375;
assign addr[60890]= -1158676398;
assign addr[60891]= -1190691925;
assign addr[60892]= -1222329801;
assign addr[60893]= -1253579991;
assign addr[60894]= -1284432584;
assign addr[60895]= -1314877795;
assign addr[60896]= -1344905966;
assign addr[60897]= -1374507575;
assign addr[60898]= -1403673233;
assign addr[60899]= -1432393688;
assign addr[60900]= -1460659832;
assign addr[60901]= -1488462700;
assign addr[60902]= -1515793473;
assign addr[60903]= -1542643483;
assign addr[60904]= -1569004214;
assign addr[60905]= -1594867305;
assign addr[60906]= -1620224553;
assign addr[60907]= -1645067915;
assign addr[60908]= -1669389513;
assign addr[60909]= -1693181631;
assign addr[60910]= -1716436725;
assign addr[60911]= -1739147417;
assign addr[60912]= -1761306505;
assign addr[60913]= -1782906961;
assign addr[60914]= -1803941934;
assign addr[60915]= -1824404752;
assign addr[60916]= -1844288924;
assign addr[60917]= -1863588145;
assign addr[60918]= -1882296293;
assign addr[60919]= -1900407434;
assign addr[60920]= -1917915825;
assign addr[60921]= -1934815911;
assign addr[60922]= -1951102334;
assign addr[60923]= -1966769926;
assign addr[60924]= -1981813720;
assign addr[60925]= -1996228943;
assign addr[60926]= -2010011024;
assign addr[60927]= -2023155591;
assign addr[60928]= -2035658475;
assign addr[60929]= -2047515711;
assign addr[60930]= -2058723538;
assign addr[60931]= -2069278401;
assign addr[60932]= -2079176953;
assign addr[60933]= -2088416053;
assign addr[60934]= -2096992772;
assign addr[60935]= -2104904390;
assign addr[60936]= -2112148396;
assign addr[60937]= -2118722494;
assign addr[60938]= -2124624598;
assign addr[60939]= -2129852837;
assign addr[60940]= -2134405552;
assign addr[60941]= -2138281298;
assign addr[60942]= -2141478848;
assign addr[60943]= -2143997187;
assign addr[60944]= -2145835515;
assign addr[60945]= -2146993250;
assign addr[60946]= -2147470025;
assign addr[60947]= -2147265689;
assign addr[60948]= -2146380306;
assign addr[60949]= -2144814157;
assign addr[60950]= -2142567738;
assign addr[60951]= -2139641764;
assign addr[60952]= -2136037160;
assign addr[60953]= -2131755071;
assign addr[60954]= -2126796855;
assign addr[60955]= -2121164085;
assign addr[60956]= -2114858546;
assign addr[60957]= -2107882239;
assign addr[60958]= -2100237377;
assign addr[60959]= -2091926384;
assign addr[60960]= -2082951896;
assign addr[60961]= -2073316760;
assign addr[60962]= -2063024031;
assign addr[60963]= -2052076975;
assign addr[60964]= -2040479063;
assign addr[60965]= -2028233973;
assign addr[60966]= -2015345591;
assign addr[60967]= -2001818002;
assign addr[60968]= -1987655498;
assign addr[60969]= -1972862571;
assign addr[60970]= -1957443913;
assign addr[60971]= -1941404413;
assign addr[60972]= -1924749160;
assign addr[60973]= -1907483436;
assign addr[60974]= -1889612716;
assign addr[60975]= -1871142669;
assign addr[60976]= -1852079154;
assign addr[60977]= -1832428215;
assign addr[60978]= -1812196087;
assign addr[60979]= -1791389186;
assign addr[60980]= -1770014111;
assign addr[60981]= -1748077642;
assign addr[60982]= -1725586737;
assign addr[60983]= -1702548529;
assign addr[60984]= -1678970324;
assign addr[60985]= -1654859602;
assign addr[60986]= -1630224009;
assign addr[60987]= -1605071359;
assign addr[60988]= -1579409630;
assign addr[60989]= -1553246960;
assign addr[60990]= -1526591649;
assign addr[60991]= -1499452149;
assign addr[60992]= -1471837070;
assign addr[60993]= -1443755168;
assign addr[60994]= -1415215352;
assign addr[60995]= -1386226674;
assign addr[60996]= -1356798326;
assign addr[60997]= -1326939644;
assign addr[60998]= -1296660098;
assign addr[60999]= -1265969291;
assign addr[61000]= -1234876957;
assign addr[61001]= -1203392958;
assign addr[61002]= -1171527280;
assign addr[61003]= -1139290029;
assign addr[61004]= -1106691431;
assign addr[61005]= -1073741824;
assign addr[61006]= -1040451659;
assign addr[61007]= -1006831495;
assign addr[61008]= -972891995;
assign addr[61009]= -938643924;
assign addr[61010]= -904098143;
assign addr[61011]= -869265610;
assign addr[61012]= -834157373;
assign addr[61013]= -798784567;
assign addr[61014]= -763158411;
assign addr[61015]= -727290205;
assign addr[61016]= -691191324;
assign addr[61017]= -654873219;
assign addr[61018]= -618347408;
assign addr[61019]= -581625477;
assign addr[61020]= -544719071;
assign addr[61021]= -507639898;
assign addr[61022]= -470399716;
assign addr[61023]= -433010339;
assign addr[61024]= -395483624;
assign addr[61025]= -357831473;
assign addr[61026]= -320065829;
assign addr[61027]= -282198671;
assign addr[61028]= -244242007;
assign addr[61029]= -206207878;
assign addr[61030]= -168108346;
assign addr[61031]= -129955495;
assign addr[61032]= -91761426;
assign addr[61033]= -53538253;
assign addr[61034]= -15298099;
assign addr[61035]= 22946906;
assign addr[61036]= 61184634;
assign addr[61037]= 99402956;
assign addr[61038]= 137589750;
assign addr[61039]= 175732905;
assign addr[61040]= 213820322;
assign addr[61041]= 251839923;
assign addr[61042]= 289779648;
assign addr[61043]= 327627463;
assign addr[61044]= 365371365;
assign addr[61045]= 402999383;
assign addr[61046]= 440499581;
assign addr[61047]= 477860067;
assign addr[61048]= 515068990;
assign addr[61049]= 552114549;
assign addr[61050]= 588984994;
assign addr[61051]= 625668632;
assign addr[61052]= 662153826;
assign addr[61053]= 698429006;
assign addr[61054]= 734482665;
assign addr[61055]= 770303369;
assign addr[61056]= 805879757;
assign addr[61057]= 841200544;
assign addr[61058]= 876254528;
assign addr[61059]= 911030591;
assign addr[61060]= 945517704;
assign addr[61061]= 979704927;
assign addr[61062]= 1013581418;
assign addr[61063]= 1047136432;
assign addr[61064]= 1080359326;
assign addr[61065]= 1113239564;
assign addr[61066]= 1145766716;
assign addr[61067]= 1177930466;
assign addr[61068]= 1209720613;
assign addr[61069]= 1241127074;
assign addr[61070]= 1272139887;
assign addr[61071]= 1302749217;
assign addr[61072]= 1332945355;
assign addr[61073]= 1362718723;
assign addr[61074]= 1392059879;
assign addr[61075]= 1420959516;
assign addr[61076]= 1449408469;
assign addr[61077]= 1477397714;
assign addr[61078]= 1504918373;
assign addr[61079]= 1531961719;
assign addr[61080]= 1558519173;
assign addr[61081]= 1584582314;
assign addr[61082]= 1610142873;
assign addr[61083]= 1635192744;
assign addr[61084]= 1659723983;
assign addr[61085]= 1683728808;
assign addr[61086]= 1707199606;
assign addr[61087]= 1730128933;
assign addr[61088]= 1752509516;
assign addr[61089]= 1774334257;
assign addr[61090]= 1795596234;
assign addr[61091]= 1816288703;
assign addr[61092]= 1836405100;
assign addr[61093]= 1855939047;
assign addr[61094]= 1874884346;
assign addr[61095]= 1893234990;
assign addr[61096]= 1910985158;
assign addr[61097]= 1928129220;
assign addr[61098]= 1944661739;
assign addr[61099]= 1960577471;
assign addr[61100]= 1975871368;
assign addr[61101]= 1990538579;
assign addr[61102]= 2004574453;
assign addr[61103]= 2017974537;
assign addr[61104]= 2030734582;
assign addr[61105]= 2042850540;
assign addr[61106]= 2054318569;
assign addr[61107]= 2065135031;
assign addr[61108]= 2075296495;
assign addr[61109]= 2084799740;
assign addr[61110]= 2093641749;
assign addr[61111]= 2101819720;
assign addr[61112]= 2109331059;
assign addr[61113]= 2116173382;
assign addr[61114]= 2122344521;
assign addr[61115]= 2127842516;
assign addr[61116]= 2132665626;
assign addr[61117]= 2136812319;
assign addr[61118]= 2140281282;
assign addr[61119]= 2143071413;
assign addr[61120]= 2145181827;
assign addr[61121]= 2146611856;
assign addr[61122]= 2147361045;
assign addr[61123]= 2147429158;
assign addr[61124]= 2146816171;
assign addr[61125]= 2145522281;
assign addr[61126]= 2143547897;
assign addr[61127]= 2140893646;
assign addr[61128]= 2137560369;
assign addr[61129]= 2133549123;
assign addr[61130]= 2128861181;
assign addr[61131]= 2123498030;
assign addr[61132]= 2117461370;
assign addr[61133]= 2110753117;
assign addr[61134]= 2103375398;
assign addr[61135]= 2095330553;
assign addr[61136]= 2086621133;
assign addr[61137]= 2077249901;
assign addr[61138]= 2067219829;
assign addr[61139]= 2056534099;
assign addr[61140]= 2045196100;
assign addr[61141]= 2033209426;
assign addr[61142]= 2020577882;
assign addr[61143]= 2007305472;
assign addr[61144]= 1993396407;
assign addr[61145]= 1978855097;
assign addr[61146]= 1963686155;
assign addr[61147]= 1947894393;
assign addr[61148]= 1931484818;
assign addr[61149]= 1914462636;
assign addr[61150]= 1896833245;
assign addr[61151]= 1878602237;
assign addr[61152]= 1859775393;
assign addr[61153]= 1840358687;
assign addr[61154]= 1820358275;
assign addr[61155]= 1799780501;
assign addr[61156]= 1778631892;
assign addr[61157]= 1756919156;
assign addr[61158]= 1734649179;
assign addr[61159]= 1711829025;
assign addr[61160]= 1688465931;
assign addr[61161]= 1664567307;
assign addr[61162]= 1640140734;
assign addr[61163]= 1615193959;
assign addr[61164]= 1589734894;
assign addr[61165]= 1563771613;
assign addr[61166]= 1537312353;
assign addr[61167]= 1510365504;
assign addr[61168]= 1482939614;
assign addr[61169]= 1455043381;
assign addr[61170]= 1426685652;
assign addr[61171]= 1397875423;
assign addr[61172]= 1368621831;
assign addr[61173]= 1338934154;
assign addr[61174]= 1308821808;
assign addr[61175]= 1278294345;
assign addr[61176]= 1247361445;
assign addr[61177]= 1216032921;
assign addr[61178]= 1184318708;
assign addr[61179]= 1152228866;
assign addr[61180]= 1119773573;
assign addr[61181]= 1086963121;
assign addr[61182]= 1053807919;
assign addr[61183]= 1020318481;
assign addr[61184]= 986505429;
assign addr[61185]= 952379488;
assign addr[61186]= 917951481;
assign addr[61187]= 883232329;
assign addr[61188]= 848233042;
assign addr[61189]= 812964722;
assign addr[61190]= 777438554;
assign addr[61191]= 741665807;
assign addr[61192]= 705657826;
assign addr[61193]= 669426032;
assign addr[61194]= 632981917;
assign addr[61195]= 596337040;
assign addr[61196]= 559503022;
assign addr[61197]= 522491548;
assign addr[61198]= 485314355;
assign addr[61199]= 447983235;
assign addr[61200]= 410510029;
assign addr[61201]= 372906622;
assign addr[61202]= 335184940;
assign addr[61203]= 297356948;
assign addr[61204]= 259434643;
assign addr[61205]= 221430054;
assign addr[61206]= 183355234;
assign addr[61207]= 145222259;
assign addr[61208]= 107043224;
assign addr[61209]= 68830239;
assign addr[61210]= 30595422;
assign addr[61211]= -7649098;
assign addr[61212]= -45891193;
assign addr[61213]= -84118732;
assign addr[61214]= -122319591;
assign addr[61215]= -160481654;
assign addr[61216]= -198592817;
assign addr[61217]= -236640993;
assign addr[61218]= -274614114;
assign addr[61219]= -312500135;
assign addr[61220]= -350287041;
assign addr[61221]= -387962847;
assign addr[61222]= -425515602;
assign addr[61223]= -462933398;
assign addr[61224]= -500204365;
assign addr[61225]= -537316682;
assign addr[61226]= -574258580;
assign addr[61227]= -611018340;
assign addr[61228]= -647584304;
assign addr[61229]= -683944874;
assign addr[61230]= -720088517;
assign addr[61231]= -756003771;
assign addr[61232]= -791679244;
assign addr[61233]= -827103620;
assign addr[61234]= -862265664;
assign addr[61235]= -897154224;
assign addr[61236]= -931758235;
assign addr[61237]= -966066720;
assign addr[61238]= -1000068799;
assign addr[61239]= -1033753687;
assign addr[61240]= -1067110699;
assign addr[61241]= -1100129257;
assign addr[61242]= -1132798888;
assign addr[61243]= -1165109230;
assign addr[61244]= -1197050035;
assign addr[61245]= -1228611172;
assign addr[61246]= -1259782632;
assign addr[61247]= -1290554528;
assign addr[61248]= -1320917099;
assign addr[61249]= -1350860716;
assign addr[61250]= -1380375881;
assign addr[61251]= -1409453233;
assign addr[61252]= -1438083551;
assign addr[61253]= -1466257752;
assign addr[61254]= -1493966902;
assign addr[61255]= -1521202211;
assign addr[61256]= -1547955041;
assign addr[61257]= -1574216908;
assign addr[61258]= -1599979481;
assign addr[61259]= -1625234591;
assign addr[61260]= -1649974225;
assign addr[61261]= -1674190539;
assign addr[61262]= -1697875851;
assign addr[61263]= -1721022648;
assign addr[61264]= -1743623590;
assign addr[61265]= -1765671509;
assign addr[61266]= -1787159411;
assign addr[61267]= -1808080480;
assign addr[61268]= -1828428082;
assign addr[61269]= -1848195763;
assign addr[61270]= -1867377253;
assign addr[61271]= -1885966468;
assign addr[61272]= -1903957513;
assign addr[61273]= -1921344681;
assign addr[61274]= -1938122457;
assign addr[61275]= -1954285520;
assign addr[61276]= -1969828744;
assign addr[61277]= -1984747199;
assign addr[61278]= -1999036154;
assign addr[61279]= -2012691075;
assign addr[61280]= -2025707632;
assign addr[61281]= -2038081698;
assign addr[61282]= -2049809346;
assign addr[61283]= -2060886858;
assign addr[61284]= -2071310720;
assign addr[61285]= -2081077626;
assign addr[61286]= -2090184478;
assign addr[61287]= -2098628387;
assign addr[61288]= -2106406677;
assign addr[61289]= -2113516878;
assign addr[61290]= -2119956737;
assign addr[61291]= -2125724211;
assign addr[61292]= -2130817471;
assign addr[61293]= -2135234901;
assign addr[61294]= -2138975100;
assign addr[61295]= -2142036881;
assign addr[61296]= -2144419275;
assign addr[61297]= -2146121524;
assign addr[61298]= -2147143090;
assign addr[61299]= -2147483648;
assign addr[61300]= -2147143090;
assign addr[61301]= -2146121524;
assign addr[61302]= -2144419275;
assign addr[61303]= -2142036881;
assign addr[61304]= -2138975100;
assign addr[61305]= -2135234901;
assign addr[61306]= -2130817471;
assign addr[61307]= -2125724211;
assign addr[61308]= -2119956737;
assign addr[61309]= -2113516878;
assign addr[61310]= -2106406677;
assign addr[61311]= -2098628387;
assign addr[61312]= -2090184478;
assign addr[61313]= -2081077626;
assign addr[61314]= -2071310720;
assign addr[61315]= -2060886858;
assign addr[61316]= -2049809346;
assign addr[61317]= -2038081698;
assign addr[61318]= -2025707632;
assign addr[61319]= -2012691075;
assign addr[61320]= -1999036154;
assign addr[61321]= -1984747199;
assign addr[61322]= -1969828744;
assign addr[61323]= -1954285520;
assign addr[61324]= -1938122457;
assign addr[61325]= -1921344681;
assign addr[61326]= -1903957513;
assign addr[61327]= -1885966468;
assign addr[61328]= -1867377253;
assign addr[61329]= -1848195763;
assign addr[61330]= -1828428082;
assign addr[61331]= -1808080480;
assign addr[61332]= -1787159411;
assign addr[61333]= -1765671509;
assign addr[61334]= -1743623590;
assign addr[61335]= -1721022648;
assign addr[61336]= -1697875851;
assign addr[61337]= -1674190539;
assign addr[61338]= -1649974225;
assign addr[61339]= -1625234591;
assign addr[61340]= -1599979481;
assign addr[61341]= -1574216908;
assign addr[61342]= -1547955041;
assign addr[61343]= -1521202211;
assign addr[61344]= -1493966902;
assign addr[61345]= -1466257752;
assign addr[61346]= -1438083551;
assign addr[61347]= -1409453233;
assign addr[61348]= -1380375881;
assign addr[61349]= -1350860716;
assign addr[61350]= -1320917099;
assign addr[61351]= -1290554528;
assign addr[61352]= -1259782632;
assign addr[61353]= -1228611172;
assign addr[61354]= -1197050035;
assign addr[61355]= -1165109230;
assign addr[61356]= -1132798888;
assign addr[61357]= -1100129257;
assign addr[61358]= -1067110699;
assign addr[61359]= -1033753687;
assign addr[61360]= -1000068799;
assign addr[61361]= -966066720;
assign addr[61362]= -931758235;
assign addr[61363]= -897154224;
assign addr[61364]= -862265664;
assign addr[61365]= -827103620;
assign addr[61366]= -791679244;
assign addr[61367]= -756003771;
assign addr[61368]= -720088517;
assign addr[61369]= -683944874;
assign addr[61370]= -647584304;
assign addr[61371]= -611018340;
assign addr[61372]= -574258580;
assign addr[61373]= -537316682;
assign addr[61374]= -500204365;
assign addr[61375]= -462933398;
assign addr[61376]= -425515602;
assign addr[61377]= -387962847;
assign addr[61378]= -350287041;
assign addr[61379]= -312500135;
assign addr[61380]= -274614114;
assign addr[61381]= -236640993;
assign addr[61382]= -198592817;
assign addr[61383]= -160481654;
assign addr[61384]= -122319591;
assign addr[61385]= -84118732;
assign addr[61386]= -45891193;
assign addr[61387]= -7649098;
assign addr[61388]= 30595422;
assign addr[61389]= 68830239;
assign addr[61390]= 107043224;
assign addr[61391]= 145222259;
assign addr[61392]= 183355234;
assign addr[61393]= 221430054;
assign addr[61394]= 259434643;
assign addr[61395]= 297356948;
assign addr[61396]= 335184940;
assign addr[61397]= 372906622;
assign addr[61398]= 410510029;
assign addr[61399]= 447983235;
assign addr[61400]= 485314355;
assign addr[61401]= 522491548;
assign addr[61402]= 559503022;
assign addr[61403]= 596337040;
assign addr[61404]= 632981917;
assign addr[61405]= 669426032;
assign addr[61406]= 705657826;
assign addr[61407]= 741665807;
assign addr[61408]= 777438554;
assign addr[61409]= 812964722;
assign addr[61410]= 848233042;
assign addr[61411]= 883232329;
assign addr[61412]= 917951481;
assign addr[61413]= 952379488;
assign addr[61414]= 986505429;
assign addr[61415]= 1020318481;
assign addr[61416]= 1053807919;
assign addr[61417]= 1086963121;
assign addr[61418]= 1119773573;
assign addr[61419]= 1152228866;
assign addr[61420]= 1184318708;
assign addr[61421]= 1216032921;
assign addr[61422]= 1247361445;
assign addr[61423]= 1278294345;
assign addr[61424]= 1308821808;
assign addr[61425]= 1338934154;
assign addr[61426]= 1368621831;
assign addr[61427]= 1397875423;
assign addr[61428]= 1426685652;
assign addr[61429]= 1455043381;
assign addr[61430]= 1482939614;
assign addr[61431]= 1510365504;
assign addr[61432]= 1537312353;
assign addr[61433]= 1563771613;
assign addr[61434]= 1589734894;
assign addr[61435]= 1615193959;
assign addr[61436]= 1640140734;
assign addr[61437]= 1664567307;
assign addr[61438]= 1688465931;
assign addr[61439]= 1711829025;
assign addr[61440]= 1734649179;
assign addr[61441]= 1756919156;
assign addr[61442]= 1778631892;
assign addr[61443]= 1799780501;
assign addr[61444]= 1820358275;
assign addr[61445]= 1840358687;
assign addr[61446]= 1859775393;
assign addr[61447]= 1878602237;
assign addr[61448]= 1896833245;
assign addr[61449]= 1914462636;
assign addr[61450]= 1931484818;
assign addr[61451]= 1947894393;
assign addr[61452]= 1963686155;
assign addr[61453]= 1978855097;
assign addr[61454]= 1993396407;
assign addr[61455]= 2007305472;
assign addr[61456]= 2020577882;
assign addr[61457]= 2033209426;
assign addr[61458]= 2045196100;
assign addr[61459]= 2056534099;
assign addr[61460]= 2067219829;
assign addr[61461]= 2077249901;
assign addr[61462]= 2086621133;
assign addr[61463]= 2095330553;
assign addr[61464]= 2103375398;
assign addr[61465]= 2110753117;
assign addr[61466]= 2117461370;
assign addr[61467]= 2123498030;
assign addr[61468]= 2128861181;
assign addr[61469]= 2133549123;
assign addr[61470]= 2137560369;
assign addr[61471]= 2140893646;
assign addr[61472]= 2143547897;
assign addr[61473]= 2145522281;
assign addr[61474]= 2146816171;
assign addr[61475]= 2147429158;
assign addr[61476]= 2147361045;
assign addr[61477]= 2146611856;
assign addr[61478]= 2145181827;
assign addr[61479]= 2143071413;
assign addr[61480]= 2140281282;
assign addr[61481]= 2136812319;
assign addr[61482]= 2132665626;
assign addr[61483]= 2127842516;
assign addr[61484]= 2122344521;
assign addr[61485]= 2116173382;
assign addr[61486]= 2109331059;
assign addr[61487]= 2101819720;
assign addr[61488]= 2093641749;
assign addr[61489]= 2084799740;
assign addr[61490]= 2075296495;
assign addr[61491]= 2065135031;
assign addr[61492]= 2054318569;
assign addr[61493]= 2042850540;
assign addr[61494]= 2030734582;
assign addr[61495]= 2017974537;
assign addr[61496]= 2004574453;
assign addr[61497]= 1990538579;
assign addr[61498]= 1975871368;
assign addr[61499]= 1960577471;
assign addr[61500]= 1944661739;
assign addr[61501]= 1928129220;
assign addr[61502]= 1910985158;
assign addr[61503]= 1893234990;
assign addr[61504]= 1874884346;
assign addr[61505]= 1855939047;
assign addr[61506]= 1836405100;
assign addr[61507]= 1816288703;
assign addr[61508]= 1795596234;
assign addr[61509]= 1774334257;
assign addr[61510]= 1752509516;
assign addr[61511]= 1730128933;
assign addr[61512]= 1707199606;
assign addr[61513]= 1683728808;
assign addr[61514]= 1659723983;
assign addr[61515]= 1635192744;
assign addr[61516]= 1610142873;
assign addr[61517]= 1584582314;
assign addr[61518]= 1558519173;
assign addr[61519]= 1531961719;
assign addr[61520]= 1504918373;
assign addr[61521]= 1477397714;
assign addr[61522]= 1449408469;
assign addr[61523]= 1420959516;
assign addr[61524]= 1392059879;
assign addr[61525]= 1362718723;
assign addr[61526]= 1332945355;
assign addr[61527]= 1302749217;
assign addr[61528]= 1272139887;
assign addr[61529]= 1241127074;
assign addr[61530]= 1209720613;
assign addr[61531]= 1177930466;
assign addr[61532]= 1145766716;
assign addr[61533]= 1113239564;
assign addr[61534]= 1080359326;
assign addr[61535]= 1047136432;
assign addr[61536]= 1013581418;
assign addr[61537]= 979704927;
assign addr[61538]= 945517704;
assign addr[61539]= 911030591;
assign addr[61540]= 876254528;
assign addr[61541]= 841200544;
assign addr[61542]= 805879757;
assign addr[61543]= 770303369;
assign addr[61544]= 734482665;
assign addr[61545]= 698429006;
assign addr[61546]= 662153826;
assign addr[61547]= 625668632;
assign addr[61548]= 588984994;
assign addr[61549]= 552114549;
assign addr[61550]= 515068990;
assign addr[61551]= 477860067;
assign addr[61552]= 440499581;
assign addr[61553]= 402999383;
assign addr[61554]= 365371365;
assign addr[61555]= 327627463;
assign addr[61556]= 289779648;
assign addr[61557]= 251839923;
assign addr[61558]= 213820322;
assign addr[61559]= 175732905;
assign addr[61560]= 137589750;
assign addr[61561]= 99402956;
assign addr[61562]= 61184634;
assign addr[61563]= 22946906;
assign addr[61564]= -15298099;
assign addr[61565]= -53538253;
assign addr[61566]= -91761426;
assign addr[61567]= -129955495;
assign addr[61568]= -168108346;
assign addr[61569]= -206207878;
assign addr[61570]= -244242007;
assign addr[61571]= -282198671;
assign addr[61572]= -320065829;
assign addr[61573]= -357831473;
assign addr[61574]= -395483624;
assign addr[61575]= -433010339;
assign addr[61576]= -470399716;
assign addr[61577]= -507639898;
assign addr[61578]= -544719071;
assign addr[61579]= -581625477;
assign addr[61580]= -618347408;
assign addr[61581]= -654873219;
assign addr[61582]= -691191324;
assign addr[61583]= -727290205;
assign addr[61584]= -763158411;
assign addr[61585]= -798784567;
assign addr[61586]= -834157373;
assign addr[61587]= -869265610;
assign addr[61588]= -904098143;
assign addr[61589]= -938643924;
assign addr[61590]= -972891995;
assign addr[61591]= -1006831495;
assign addr[61592]= -1040451659;
assign addr[61593]= -1073741824;
assign addr[61594]= -1106691431;
assign addr[61595]= -1139290029;
assign addr[61596]= -1171527280;
assign addr[61597]= -1203392958;
assign addr[61598]= -1234876957;
assign addr[61599]= -1265969291;
assign addr[61600]= -1296660098;
assign addr[61601]= -1326939644;
assign addr[61602]= -1356798326;
assign addr[61603]= -1386226674;
assign addr[61604]= -1415215352;
assign addr[61605]= -1443755168;
assign addr[61606]= -1471837070;
assign addr[61607]= -1499452149;
assign addr[61608]= -1526591649;
assign addr[61609]= -1553246960;
assign addr[61610]= -1579409630;
assign addr[61611]= -1605071359;
assign addr[61612]= -1630224009;
assign addr[61613]= -1654859602;
assign addr[61614]= -1678970324;
assign addr[61615]= -1702548529;
assign addr[61616]= -1725586737;
assign addr[61617]= -1748077642;
assign addr[61618]= -1770014111;
assign addr[61619]= -1791389186;
assign addr[61620]= -1812196087;
assign addr[61621]= -1832428215;
assign addr[61622]= -1852079154;
assign addr[61623]= -1871142669;
assign addr[61624]= -1889612716;
assign addr[61625]= -1907483436;
assign addr[61626]= -1924749160;
assign addr[61627]= -1941404413;
assign addr[61628]= -1957443913;
assign addr[61629]= -1972862571;
assign addr[61630]= -1987655498;
assign addr[61631]= -2001818002;
assign addr[61632]= -2015345591;
assign addr[61633]= -2028233973;
assign addr[61634]= -2040479063;
assign addr[61635]= -2052076975;
assign addr[61636]= -2063024031;
assign addr[61637]= -2073316760;
assign addr[61638]= -2082951896;
assign addr[61639]= -2091926384;
assign addr[61640]= -2100237377;
assign addr[61641]= -2107882239;
assign addr[61642]= -2114858546;
assign addr[61643]= -2121164085;
assign addr[61644]= -2126796855;
assign addr[61645]= -2131755071;
assign addr[61646]= -2136037160;
assign addr[61647]= -2139641764;
assign addr[61648]= -2142567738;
assign addr[61649]= -2144814157;
assign addr[61650]= -2146380306;
assign addr[61651]= -2147265689;
assign addr[61652]= -2147470025;
assign addr[61653]= -2146993250;
assign addr[61654]= -2145835515;
assign addr[61655]= -2143997187;
assign addr[61656]= -2141478848;
assign addr[61657]= -2138281298;
assign addr[61658]= -2134405552;
assign addr[61659]= -2129852837;
assign addr[61660]= -2124624598;
assign addr[61661]= -2118722494;
assign addr[61662]= -2112148396;
assign addr[61663]= -2104904390;
assign addr[61664]= -2096992772;
assign addr[61665]= -2088416053;
assign addr[61666]= -2079176953;
assign addr[61667]= -2069278401;
assign addr[61668]= -2058723538;
assign addr[61669]= -2047515711;
assign addr[61670]= -2035658475;
assign addr[61671]= -2023155591;
assign addr[61672]= -2010011024;
assign addr[61673]= -1996228943;
assign addr[61674]= -1981813720;
assign addr[61675]= -1966769926;
assign addr[61676]= -1951102334;
assign addr[61677]= -1934815911;
assign addr[61678]= -1917915825;
assign addr[61679]= -1900407434;
assign addr[61680]= -1882296293;
assign addr[61681]= -1863588145;
assign addr[61682]= -1844288924;
assign addr[61683]= -1824404752;
assign addr[61684]= -1803941934;
assign addr[61685]= -1782906961;
assign addr[61686]= -1761306505;
assign addr[61687]= -1739147417;
assign addr[61688]= -1716436725;
assign addr[61689]= -1693181631;
assign addr[61690]= -1669389513;
assign addr[61691]= -1645067915;
assign addr[61692]= -1620224553;
assign addr[61693]= -1594867305;
assign addr[61694]= -1569004214;
assign addr[61695]= -1542643483;
assign addr[61696]= -1515793473;
assign addr[61697]= -1488462700;
assign addr[61698]= -1460659832;
assign addr[61699]= -1432393688;
assign addr[61700]= -1403673233;
assign addr[61701]= -1374507575;
assign addr[61702]= -1344905966;
assign addr[61703]= -1314877795;
assign addr[61704]= -1284432584;
assign addr[61705]= -1253579991;
assign addr[61706]= -1222329801;
assign addr[61707]= -1190691925;
assign addr[61708]= -1158676398;
assign addr[61709]= -1126293375;
assign addr[61710]= -1093553126;
assign addr[61711]= -1060466036;
assign addr[61712]= -1027042599;
assign addr[61713]= -993293415;
assign addr[61714]= -959229189;
assign addr[61715]= -924860725;
assign addr[61716]= -890198924;
assign addr[61717]= -855254778;
assign addr[61718]= -820039373;
assign addr[61719]= -784563876;
assign addr[61720]= -748839539;
assign addr[61721]= -712877694;
assign addr[61722]= -676689746;
assign addr[61723]= -640287172;
assign addr[61724]= -603681519;
assign addr[61725]= -566884397;
assign addr[61726]= -529907477;
assign addr[61727]= -492762486;
assign addr[61728]= -455461206;
assign addr[61729]= -418015468;
assign addr[61730]= -380437148;
assign addr[61731]= -342738165;
assign addr[61732]= -304930476;
assign addr[61733]= -267026072;
assign addr[61734]= -229036977;
assign addr[61735]= -190975237;
assign addr[61736]= -152852926;
assign addr[61737]= -114682135;
assign addr[61738]= -76474970;
assign addr[61739]= -38243550;
assign addr[61740]= 0;
assign addr[61741]= 38243550;
assign addr[61742]= 76474970;
assign addr[61743]= 114682135;
assign addr[61744]= 152852926;
assign addr[61745]= 190975237;
assign addr[61746]= 229036977;
assign addr[61747]= 267026072;
assign addr[61748]= 304930476;
assign addr[61749]= 342738165;
assign addr[61750]= 380437148;
assign addr[61751]= 418015468;
assign addr[61752]= 455461206;
assign addr[61753]= 492762486;
assign addr[61754]= 529907477;
assign addr[61755]= 566884397;
assign addr[61756]= 603681519;
assign addr[61757]= 640287172;
assign addr[61758]= 676689746;
assign addr[61759]= 712877694;
assign addr[61760]= 748839539;
assign addr[61761]= 784563876;
assign addr[61762]= 820039373;
assign addr[61763]= 855254778;
assign addr[61764]= 890198924;
assign addr[61765]= 924860725;
assign addr[61766]= 959229189;
assign addr[61767]= 993293415;
assign addr[61768]= 1027042599;
assign addr[61769]= 1060466036;
assign addr[61770]= 1093553126;
assign addr[61771]= 1126293375;
assign addr[61772]= 1158676398;
assign addr[61773]= 1190691925;
assign addr[61774]= 1222329801;
assign addr[61775]= 1253579991;
assign addr[61776]= 1284432584;
assign addr[61777]= 1314877795;
assign addr[61778]= 1344905966;
assign addr[61779]= 1374507575;
assign addr[61780]= 1403673233;
assign addr[61781]= 1432393688;
assign addr[61782]= 1460659832;
assign addr[61783]= 1488462700;
assign addr[61784]= 1515793473;
assign addr[61785]= 1542643483;
assign addr[61786]= 1569004214;
assign addr[61787]= 1594867305;
assign addr[61788]= 1620224553;
assign addr[61789]= 1645067915;
assign addr[61790]= 1669389513;
assign addr[61791]= 1693181631;
assign addr[61792]= 1716436725;
assign addr[61793]= 1739147417;
assign addr[61794]= 1761306505;
assign addr[61795]= 1782906961;
assign addr[61796]= 1803941934;
assign addr[61797]= 1824404752;
assign addr[61798]= 1844288924;
assign addr[61799]= 1863588145;
assign addr[61800]= 1882296293;
assign addr[61801]= 1900407434;
assign addr[61802]= 1917915825;
assign addr[61803]= 1934815911;
assign addr[61804]= 1951102334;
assign addr[61805]= 1966769926;
assign addr[61806]= 1981813720;
assign addr[61807]= 1996228943;
assign addr[61808]= 2010011024;
assign addr[61809]= 2023155591;
assign addr[61810]= 2035658475;
assign addr[61811]= 2047515711;
assign addr[61812]= 2058723538;
assign addr[61813]= 2069278401;
assign addr[61814]= 2079176953;
assign addr[61815]= 2088416053;
assign addr[61816]= 2096992772;
assign addr[61817]= 2104904390;
assign addr[61818]= 2112148396;
assign addr[61819]= 2118722494;
assign addr[61820]= 2124624598;
assign addr[61821]= 2129852837;
assign addr[61822]= 2134405552;
assign addr[61823]= 2138281298;
assign addr[61824]= 2141478848;
assign addr[61825]= 2143997187;
assign addr[61826]= 2145835515;
assign addr[61827]= 2146993250;
assign addr[61828]= 2147470025;
assign addr[61829]= 2147265689;
assign addr[61830]= 2146380306;
assign addr[61831]= 2144814157;
assign addr[61832]= 2142567738;
assign addr[61833]= 2139641764;
assign addr[61834]= 2136037160;
assign addr[61835]= 2131755071;
assign addr[61836]= 2126796855;
assign addr[61837]= 2121164085;
assign addr[61838]= 2114858546;
assign addr[61839]= 2107882239;
assign addr[61840]= 2100237377;
assign addr[61841]= 2091926384;
assign addr[61842]= 2082951896;
assign addr[61843]= 2073316760;
assign addr[61844]= 2063024031;
assign addr[61845]= 2052076975;
assign addr[61846]= 2040479063;
assign addr[61847]= 2028233973;
assign addr[61848]= 2015345591;
assign addr[61849]= 2001818002;
assign addr[61850]= 1987655498;
assign addr[61851]= 1972862571;
assign addr[61852]= 1957443913;
assign addr[61853]= 1941404413;
assign addr[61854]= 1924749160;
assign addr[61855]= 1907483436;
assign addr[61856]= 1889612716;
assign addr[61857]= 1871142669;
assign addr[61858]= 1852079154;
assign addr[61859]= 1832428215;
assign addr[61860]= 1812196087;
assign addr[61861]= 1791389186;
assign addr[61862]= 1770014111;
assign addr[61863]= 1748077642;
assign addr[61864]= 1725586737;
assign addr[61865]= 1702548529;
assign addr[61866]= 1678970324;
assign addr[61867]= 1654859602;
assign addr[61868]= 1630224009;
assign addr[61869]= 1605071359;
assign addr[61870]= 1579409630;
assign addr[61871]= 1553246960;
assign addr[61872]= 1526591649;
assign addr[61873]= 1499452149;
assign addr[61874]= 1471837070;
assign addr[61875]= 1443755168;
assign addr[61876]= 1415215352;
assign addr[61877]= 1386226674;
assign addr[61878]= 1356798326;
assign addr[61879]= 1326939644;
assign addr[61880]= 1296660098;
assign addr[61881]= 1265969291;
assign addr[61882]= 1234876957;
assign addr[61883]= 1203392958;
assign addr[61884]= 1171527280;
assign addr[61885]= 1139290029;
assign addr[61886]= 1106691431;
assign addr[61887]= 1073741824;
assign addr[61888]= 1040451659;
assign addr[61889]= 1006831495;
assign addr[61890]= 972891995;
assign addr[61891]= 938643924;
assign addr[61892]= 904098143;
assign addr[61893]= 869265610;
assign addr[61894]= 834157373;
assign addr[61895]= 798784567;
assign addr[61896]= 763158411;
assign addr[61897]= 727290205;
assign addr[61898]= 691191324;
assign addr[61899]= 654873219;
assign addr[61900]= 618347408;
assign addr[61901]= 581625477;
assign addr[61902]= 544719071;
assign addr[61903]= 507639898;
assign addr[61904]= 470399716;
assign addr[61905]= 433010339;
assign addr[61906]= 395483624;
assign addr[61907]= 357831473;
assign addr[61908]= 320065829;
assign addr[61909]= 282198671;
assign addr[61910]= 244242007;
assign addr[61911]= 206207878;
assign addr[61912]= 168108346;
assign addr[61913]= 129955495;
assign addr[61914]= 91761426;
assign addr[61915]= 53538253;
assign addr[61916]= 15298099;
assign addr[61917]= -22946906;
assign addr[61918]= -61184634;
assign addr[61919]= -99402956;
assign addr[61920]= -137589750;
assign addr[61921]= -175732905;
assign addr[61922]= -213820322;
assign addr[61923]= -251839923;
assign addr[61924]= -289779648;
assign addr[61925]= -327627463;
assign addr[61926]= -365371365;
assign addr[61927]= -402999383;
assign addr[61928]= -440499581;
assign addr[61929]= -477860067;
assign addr[61930]= -515068990;
assign addr[61931]= -552114549;
assign addr[61932]= -588984994;
assign addr[61933]= -625668632;
assign addr[61934]= -662153826;
assign addr[61935]= -698429006;
assign addr[61936]= -734482665;
assign addr[61937]= -770303369;
assign addr[61938]= -805879757;
assign addr[61939]= -841200544;
assign addr[61940]= -876254528;
assign addr[61941]= -911030591;
assign addr[61942]= -945517704;
assign addr[61943]= -979704927;
assign addr[61944]= -1013581418;
assign addr[61945]= -1047136432;
assign addr[61946]= -1080359326;
assign addr[61947]= -1113239564;
assign addr[61948]= -1145766716;
assign addr[61949]= -1177930466;
assign addr[61950]= -1209720613;
assign addr[61951]= -1241127074;
assign addr[61952]= -1272139887;
assign addr[61953]= -1302749217;
assign addr[61954]= -1332945355;
assign addr[61955]= -1362718723;
assign addr[61956]= -1392059879;
assign addr[61957]= -1420959516;
assign addr[61958]= -1449408469;
assign addr[61959]= -1477397714;
assign addr[61960]= -1504918373;
assign addr[61961]= -1531961719;
assign addr[61962]= -1558519173;
assign addr[61963]= -1584582314;
assign addr[61964]= -1610142873;
assign addr[61965]= -1635192744;
assign addr[61966]= -1659723983;
assign addr[61967]= -1683728808;
assign addr[61968]= -1707199606;
assign addr[61969]= -1730128933;
assign addr[61970]= -1752509516;
assign addr[61971]= -1774334257;
assign addr[61972]= -1795596234;
assign addr[61973]= -1816288703;
assign addr[61974]= -1836405100;
assign addr[61975]= -1855939047;
assign addr[61976]= -1874884346;
assign addr[61977]= -1893234990;
assign addr[61978]= -1910985158;
assign addr[61979]= -1928129220;
assign addr[61980]= -1944661739;
assign addr[61981]= -1960577471;
assign addr[61982]= -1975871368;
assign addr[61983]= -1990538579;
assign addr[61984]= -2004574453;
assign addr[61985]= -2017974537;
assign addr[61986]= -2030734582;
assign addr[61987]= -2042850540;
assign addr[61988]= -2054318569;
assign addr[61989]= -2065135031;
assign addr[61990]= -2075296495;
assign addr[61991]= -2084799740;
assign addr[61992]= -2093641749;
assign addr[61993]= -2101819720;
assign addr[61994]= -2109331059;
assign addr[61995]= -2116173382;
assign addr[61996]= -2122344521;
assign addr[61997]= -2127842516;
assign addr[61998]= -2132665626;
assign addr[61999]= -2136812319;
assign addr[62000]= -2140281282;
assign addr[62001]= -2143071413;
assign addr[62002]= -2145181827;
assign addr[62003]= -2146611856;
assign addr[62004]= -2147361045;
assign addr[62005]= -2147429158;
assign addr[62006]= -2146816171;
assign addr[62007]= -2145522281;
assign addr[62008]= -2143547897;
assign addr[62009]= -2140893646;
assign addr[62010]= -2137560369;
assign addr[62011]= -2133549123;
assign addr[62012]= -2128861181;
assign addr[62013]= -2123498030;
assign addr[62014]= -2117461370;
assign addr[62015]= -2110753117;
assign addr[62016]= -2103375398;
assign addr[62017]= -2095330553;
assign addr[62018]= -2086621133;
assign addr[62019]= -2077249901;
assign addr[62020]= -2067219829;
assign addr[62021]= -2056534099;
assign addr[62022]= -2045196100;
assign addr[62023]= -2033209426;
assign addr[62024]= -2020577882;
assign addr[62025]= -2007305472;
assign addr[62026]= -1993396407;
assign addr[62027]= -1978855097;
assign addr[62028]= -1963686155;
assign addr[62029]= -1947894393;
assign addr[62030]= -1931484818;
assign addr[62031]= -1914462636;
assign addr[62032]= -1896833245;
assign addr[62033]= -1878602237;
assign addr[62034]= -1859775393;
assign addr[62035]= -1840358687;
assign addr[62036]= -1820358275;
assign addr[62037]= -1799780501;
assign addr[62038]= -1778631892;
assign addr[62039]= -1756919156;
assign addr[62040]= -1734649179;
assign addr[62041]= -1711829025;
assign addr[62042]= -1688465931;
assign addr[62043]= -1664567307;
assign addr[62044]= -1640140734;
assign addr[62045]= -1615193959;
assign addr[62046]= -1589734894;
assign addr[62047]= -1563771613;
assign addr[62048]= -1537312353;
assign addr[62049]= -1510365504;
assign addr[62050]= -1482939614;
assign addr[62051]= -1455043381;
assign addr[62052]= -1426685652;
assign addr[62053]= -1397875423;
assign addr[62054]= -1368621831;
assign addr[62055]= -1338934154;
assign addr[62056]= -1308821808;
assign addr[62057]= -1278294345;
assign addr[62058]= -1247361445;
assign addr[62059]= -1216032921;
assign addr[62060]= -1184318708;
assign addr[62061]= -1152228866;
assign addr[62062]= -1119773573;
assign addr[62063]= -1086963121;
assign addr[62064]= -1053807919;
assign addr[62065]= -1020318481;
assign addr[62066]= -986505429;
assign addr[62067]= -952379488;
assign addr[62068]= -917951481;
assign addr[62069]= -883232329;
assign addr[62070]= -848233042;
assign addr[62071]= -812964722;
assign addr[62072]= -777438554;
assign addr[62073]= -741665807;
assign addr[62074]= -705657826;
assign addr[62075]= -669426032;
assign addr[62076]= -632981917;
assign addr[62077]= -596337040;
assign addr[62078]= -559503022;
assign addr[62079]= -522491548;
assign addr[62080]= -485314355;
assign addr[62081]= -447983235;
assign addr[62082]= -410510029;
assign addr[62083]= -372906622;
assign addr[62084]= -335184940;
assign addr[62085]= -297356948;
assign addr[62086]= -259434643;
assign addr[62087]= -221430054;
assign addr[62088]= -183355234;
assign addr[62089]= -145222259;
assign addr[62090]= -107043224;
assign addr[62091]= -68830239;
assign addr[62092]= -30595422;
assign addr[62093]= 7649098;
assign addr[62094]= 45891193;
assign addr[62095]= 84118732;
assign addr[62096]= 122319591;
assign addr[62097]= 160481654;
assign addr[62098]= 198592817;
assign addr[62099]= 236640993;
assign addr[62100]= 274614114;
assign addr[62101]= 312500135;
assign addr[62102]= 350287041;
assign addr[62103]= 387962847;
assign addr[62104]= 425515602;
assign addr[62105]= 462933398;
assign addr[62106]= 500204365;
assign addr[62107]= 537316682;
assign addr[62108]= 574258580;
assign addr[62109]= 611018340;
assign addr[62110]= 647584304;
assign addr[62111]= 683944874;
assign addr[62112]= 720088517;
assign addr[62113]= 756003771;
assign addr[62114]= 791679244;
assign addr[62115]= 827103620;
assign addr[62116]= 862265664;
assign addr[62117]= 897154224;
assign addr[62118]= 931758235;
assign addr[62119]= 966066720;
assign addr[62120]= 1000068799;
assign addr[62121]= 1033753687;
assign addr[62122]= 1067110699;
assign addr[62123]= 1100129257;
assign addr[62124]= 1132798888;
assign addr[62125]= 1165109230;
assign addr[62126]= 1197050035;
assign addr[62127]= 1228611172;
assign addr[62128]= 1259782632;
assign addr[62129]= 1290554528;
assign addr[62130]= 1320917099;
assign addr[62131]= 1350860716;
assign addr[62132]= 1380375881;
assign addr[62133]= 1409453233;
assign addr[62134]= 1438083551;
assign addr[62135]= 1466257752;
assign addr[62136]= 1493966902;
assign addr[62137]= 1521202211;
assign addr[62138]= 1547955041;
assign addr[62139]= 1574216908;
assign addr[62140]= 1599979481;
assign addr[62141]= 1625234591;
assign addr[62142]= 1649974225;
assign addr[62143]= 1674190539;
assign addr[62144]= 1697875851;
assign addr[62145]= 1721022648;
assign addr[62146]= 1743623590;
assign addr[62147]= 1765671509;
assign addr[62148]= 1787159411;
assign addr[62149]= 1808080480;
assign addr[62150]= 1828428082;
assign addr[62151]= 1848195763;
assign addr[62152]= 1867377253;
assign addr[62153]= 1885966468;
assign addr[62154]= 1903957513;
assign addr[62155]= 1921344681;
assign addr[62156]= 1938122457;
assign addr[62157]= 1954285520;
assign addr[62158]= 1969828744;
assign addr[62159]= 1984747199;
assign addr[62160]= 1999036154;
assign addr[62161]= 2012691075;
assign addr[62162]= 2025707632;
assign addr[62163]= 2038081698;
assign addr[62164]= 2049809346;
assign addr[62165]= 2060886858;
assign addr[62166]= 2071310720;
assign addr[62167]= 2081077626;
assign addr[62168]= 2090184478;
assign addr[62169]= 2098628387;
assign addr[62170]= 2106406677;
assign addr[62171]= 2113516878;
assign addr[62172]= 2119956737;
assign addr[62173]= 2125724211;
assign addr[62174]= 2130817471;
assign addr[62175]= 2135234901;
assign addr[62176]= 2138975100;
assign addr[62177]= 2142036881;
assign addr[62178]= 2144419275;
assign addr[62179]= 2146121524;
assign addr[62180]= 2147143090;
assign addr[62181]= 2147483648;
assign addr[62182]= 2147143090;
assign addr[62183]= 2146121524;
assign addr[62184]= 2144419275;
assign addr[62185]= 2142036881;
assign addr[62186]= 2138975100;
assign addr[62187]= 2135234901;
assign addr[62188]= 2130817471;
assign addr[62189]= 2125724211;
assign addr[62190]= 2119956737;
assign addr[62191]= 2113516878;
assign addr[62192]= 2106406677;
assign addr[62193]= 2098628387;
assign addr[62194]= 2090184478;
assign addr[62195]= 2081077626;
assign addr[62196]= 2071310720;
assign addr[62197]= 2060886858;
assign addr[62198]= 2049809346;
assign addr[62199]= 2038081698;
assign addr[62200]= 2025707632;
assign addr[62201]= 2012691075;
assign addr[62202]= 1999036154;
assign addr[62203]= 1984747199;
assign addr[62204]= 1969828744;
assign addr[62205]= 1954285520;
assign addr[62206]= 1938122457;
assign addr[62207]= 1921344681;
assign addr[62208]= 1903957513;
assign addr[62209]= 1885966468;
assign addr[62210]= 1867377253;
assign addr[62211]= 1848195763;
assign addr[62212]= 1828428082;
assign addr[62213]= 1808080480;
assign addr[62214]= 1787159411;
assign addr[62215]= 1765671509;
assign addr[62216]= 1743623590;
assign addr[62217]= 1721022648;
assign addr[62218]= 1697875851;
assign addr[62219]= 1674190539;
assign addr[62220]= 1649974225;
assign addr[62221]= 1625234591;
assign addr[62222]= 1599979481;
assign addr[62223]= 1574216908;
assign addr[62224]= 1547955041;
assign addr[62225]= 1521202211;
assign addr[62226]= 1493966902;
assign addr[62227]= 1466257752;
assign addr[62228]= 1438083551;
assign addr[62229]= 1409453233;
assign addr[62230]= 1380375881;
assign addr[62231]= 1350860716;
assign addr[62232]= 1320917099;
assign addr[62233]= 1290554528;
assign addr[62234]= 1259782632;
assign addr[62235]= 1228611172;
assign addr[62236]= 1197050035;
assign addr[62237]= 1165109230;
assign addr[62238]= 1132798888;
assign addr[62239]= 1100129257;
assign addr[62240]= 1067110699;
assign addr[62241]= 1033753687;
assign addr[62242]= 1000068799;
assign addr[62243]= 966066720;
assign addr[62244]= 931758235;
assign addr[62245]= 897154224;
assign addr[62246]= 862265664;
assign addr[62247]= 827103620;
assign addr[62248]= 791679244;
assign addr[62249]= 756003771;
assign addr[62250]= 720088517;
assign addr[62251]= 683944874;
assign addr[62252]= 647584304;
assign addr[62253]= 611018340;
assign addr[62254]= 574258580;
assign addr[62255]= 537316682;
assign addr[62256]= 500204365;
assign addr[62257]= 462933398;
assign addr[62258]= 425515602;
assign addr[62259]= 387962847;
assign addr[62260]= 350287041;
assign addr[62261]= 312500135;
assign addr[62262]= 274614114;
assign addr[62263]= 236640993;
assign addr[62264]= 198592817;
assign addr[62265]= 160481654;
assign addr[62266]= 122319591;
assign addr[62267]= 84118732;
assign addr[62268]= 45891193;
assign addr[62269]= 7649098;
assign addr[62270]= -30595422;
assign addr[62271]= -68830239;
assign addr[62272]= -107043224;
assign addr[62273]= -145222259;
assign addr[62274]= -183355234;
assign addr[62275]= -221430054;
assign addr[62276]= -259434643;
assign addr[62277]= -297356948;
assign addr[62278]= -335184940;
assign addr[62279]= -372906622;
assign addr[62280]= -410510029;
assign addr[62281]= -447983235;
assign addr[62282]= -485314355;
assign addr[62283]= -522491548;
assign addr[62284]= -559503022;
assign addr[62285]= -596337040;
assign addr[62286]= -632981917;
assign addr[62287]= -669426032;
assign addr[62288]= -705657826;
assign addr[62289]= -741665807;
assign addr[62290]= -777438554;
assign addr[62291]= -812964722;
assign addr[62292]= -848233042;
assign addr[62293]= -883232329;
assign addr[62294]= -917951481;
assign addr[62295]= -952379488;
assign addr[62296]= -986505429;
assign addr[62297]= -1020318481;
assign addr[62298]= -1053807919;
assign addr[62299]= -1086963121;
assign addr[62300]= -1119773573;
assign addr[62301]= -1152228866;
assign addr[62302]= -1184318708;
assign addr[62303]= -1216032921;
assign addr[62304]= -1247361445;
assign addr[62305]= -1278294345;
assign addr[62306]= -1308821808;
assign addr[62307]= -1338934154;
assign addr[62308]= -1368621831;
assign addr[62309]= -1397875423;
assign addr[62310]= -1426685652;
assign addr[62311]= -1455043381;
assign addr[62312]= -1482939614;
assign addr[62313]= -1510365504;
assign addr[62314]= -1537312353;
assign addr[62315]= -1563771613;
assign addr[62316]= -1589734894;
assign addr[62317]= -1615193959;
assign addr[62318]= -1640140734;
assign addr[62319]= -1664567307;
assign addr[62320]= -1688465931;
assign addr[62321]= -1711829025;
assign addr[62322]= -1734649179;
assign addr[62323]= -1756919156;
assign addr[62324]= -1778631892;
assign addr[62325]= -1799780501;
assign addr[62326]= -1820358275;
assign addr[62327]= -1840358687;
assign addr[62328]= -1859775393;
assign addr[62329]= -1878602237;
assign addr[62330]= -1896833245;
assign addr[62331]= -1914462636;
assign addr[62332]= -1931484818;
assign addr[62333]= -1947894393;
assign addr[62334]= -1963686155;
assign addr[62335]= -1978855097;
assign addr[62336]= -1993396407;
assign addr[62337]= -2007305472;
assign addr[62338]= -2020577882;
assign addr[62339]= -2033209426;
assign addr[62340]= -2045196100;
assign addr[62341]= -2056534099;
assign addr[62342]= -2067219829;
assign addr[62343]= -2077249901;
assign addr[62344]= -2086621133;
assign addr[62345]= -2095330553;
assign addr[62346]= -2103375398;
assign addr[62347]= -2110753117;
assign addr[62348]= -2117461370;
assign addr[62349]= -2123498030;
assign addr[62350]= -2128861181;
assign addr[62351]= -2133549123;
assign addr[62352]= -2137560369;
assign addr[62353]= -2140893646;
assign addr[62354]= -2143547897;
assign addr[62355]= -2145522281;
assign addr[62356]= -2146816171;
assign addr[62357]= -2147429158;
assign addr[62358]= -2147361045;
assign addr[62359]= -2146611856;
assign addr[62360]= -2145181827;
assign addr[62361]= -2143071413;
assign addr[62362]= -2140281282;
assign addr[62363]= -2136812319;
assign addr[62364]= -2132665626;
assign addr[62365]= -2127842516;
assign addr[62366]= -2122344521;
assign addr[62367]= -2116173382;
assign addr[62368]= -2109331059;
assign addr[62369]= -2101819720;
assign addr[62370]= -2093641749;
assign addr[62371]= -2084799740;
assign addr[62372]= -2075296495;
assign addr[62373]= -2065135031;
assign addr[62374]= -2054318569;
assign addr[62375]= -2042850540;
assign addr[62376]= -2030734582;
assign addr[62377]= -2017974537;
assign addr[62378]= -2004574453;
assign addr[62379]= -1990538579;
assign addr[62380]= -1975871368;
assign addr[62381]= -1960577471;
assign addr[62382]= -1944661739;
assign addr[62383]= -1928129220;
assign addr[62384]= -1910985158;
assign addr[62385]= -1893234990;
assign addr[62386]= -1874884346;
assign addr[62387]= -1855939047;
assign addr[62388]= -1836405100;
assign addr[62389]= -1816288703;
assign addr[62390]= -1795596234;
assign addr[62391]= -1774334257;
assign addr[62392]= -1752509516;
assign addr[62393]= -1730128933;
assign addr[62394]= -1707199606;
assign addr[62395]= -1683728808;
assign addr[62396]= -1659723983;
assign addr[62397]= -1635192744;
assign addr[62398]= -1610142873;
assign addr[62399]= -1584582314;
assign addr[62400]= -1558519173;
assign addr[62401]= -1531961719;
assign addr[62402]= -1504918373;
assign addr[62403]= -1477397714;
assign addr[62404]= -1449408469;
assign addr[62405]= -1420959516;
assign addr[62406]= -1392059879;
assign addr[62407]= -1362718723;
assign addr[62408]= -1332945355;
assign addr[62409]= -1302749217;
assign addr[62410]= -1272139887;
assign addr[62411]= -1241127074;
assign addr[62412]= -1209720613;
assign addr[62413]= -1177930466;
assign addr[62414]= -1145766716;
assign addr[62415]= -1113239564;
assign addr[62416]= -1080359326;
assign addr[62417]= -1047136432;
assign addr[62418]= -1013581418;
assign addr[62419]= -979704927;
assign addr[62420]= -945517704;
assign addr[62421]= -911030591;
assign addr[62422]= -876254528;
assign addr[62423]= -841200544;
assign addr[62424]= -805879757;
assign addr[62425]= -770303369;
assign addr[62426]= -734482665;
assign addr[62427]= -698429006;
assign addr[62428]= -662153826;
assign addr[62429]= -625668632;
assign addr[62430]= -588984994;
assign addr[62431]= -552114549;
assign addr[62432]= -515068990;
assign addr[62433]= -477860067;
assign addr[62434]= -440499581;
assign addr[62435]= -402999383;
assign addr[62436]= -365371365;
assign addr[62437]= -327627463;
assign addr[62438]= -289779648;
assign addr[62439]= -251839923;
assign addr[62440]= -213820322;
assign addr[62441]= -175732905;
assign addr[62442]= -137589750;
assign addr[62443]= -99402956;
assign addr[62444]= -61184634;
assign addr[62445]= -22946906;
assign addr[62446]= 15298099;
assign addr[62447]= 53538253;
assign addr[62448]= 91761426;
assign addr[62449]= 129955495;
assign addr[62450]= 168108346;
assign addr[62451]= 206207878;
assign addr[62452]= 244242007;
assign addr[62453]= 282198671;
assign addr[62454]= 320065829;
assign addr[62455]= 357831473;
assign addr[62456]= 395483624;
assign addr[62457]= 433010339;
assign addr[62458]= 470399716;
assign addr[62459]= 507639898;
assign addr[62460]= 544719071;
assign addr[62461]= 581625477;
assign addr[62462]= 618347408;
assign addr[62463]= 654873219;
assign addr[62464]= 691191324;
assign addr[62465]= 727290205;
assign addr[62466]= 763158411;
assign addr[62467]= 798784567;
assign addr[62468]= 834157373;
assign addr[62469]= 869265610;
assign addr[62470]= 904098143;
assign addr[62471]= 938643924;
assign addr[62472]= 972891995;
assign addr[62473]= 1006831495;
assign addr[62474]= 1040451659;
assign addr[62475]= 1073741824;
assign addr[62476]= 1106691431;
assign addr[62477]= 1139290029;
assign addr[62478]= 1171527280;
assign addr[62479]= 1203392958;
assign addr[62480]= 1234876957;
assign addr[62481]= 1265969291;
assign addr[62482]= 1296660098;
assign addr[62483]= 1326939644;
assign addr[62484]= 1356798326;
assign addr[62485]= 1386226674;
assign addr[62486]= 1415215352;
assign addr[62487]= 1443755168;
assign addr[62488]= 1471837070;
assign addr[62489]= 1499452149;
assign addr[62490]= 1526591649;
assign addr[62491]= 1553246960;
assign addr[62492]= 1579409630;
assign addr[62493]= 1605071359;
assign addr[62494]= 1630224009;
assign addr[62495]= 1654859602;
assign addr[62496]= 1678970324;
assign addr[62497]= 1702548529;
assign addr[62498]= 1725586737;
assign addr[62499]= 1748077642;
assign addr[62500]= 1770014111;
assign addr[62501]= 1791389186;
assign addr[62502]= 1812196087;
assign addr[62503]= 1832428215;
assign addr[62504]= 1852079154;
assign addr[62505]= 1871142669;
assign addr[62506]= 1889612716;
assign addr[62507]= 1907483436;
assign addr[62508]= 1924749160;
assign addr[62509]= 1941404413;
assign addr[62510]= 1957443913;
assign addr[62511]= 1972862571;
assign addr[62512]= 1987655498;
assign addr[62513]= 2001818002;
assign addr[62514]= 2015345591;
assign addr[62515]= 2028233973;
assign addr[62516]= 2040479063;
assign addr[62517]= 2052076975;
assign addr[62518]= 2063024031;
assign addr[62519]= 2073316760;
assign addr[62520]= 2082951896;
assign addr[62521]= 2091926384;
assign addr[62522]= 2100237377;
assign addr[62523]= 2107882239;
assign addr[62524]= 2114858546;
assign addr[62525]= 2121164085;
assign addr[62526]= 2126796855;
assign addr[62527]= 2131755071;
assign addr[62528]= 2136037160;
assign addr[62529]= 2139641764;
assign addr[62530]= 2142567738;
assign addr[62531]= 2144814157;
assign addr[62532]= 2146380306;
assign addr[62533]= 2147265689;
assign addr[62534]= 2147470025;
assign addr[62535]= 2146993250;
assign addr[62536]= 2145835515;
assign addr[62537]= 2143997187;
assign addr[62538]= 2141478848;
assign addr[62539]= 2138281298;
assign addr[62540]= 2134405552;
assign addr[62541]= 2129852837;
assign addr[62542]= 2124624598;
assign addr[62543]= 2118722494;
assign addr[62544]= 2112148396;
assign addr[62545]= 2104904390;
assign addr[62546]= 2096992772;
assign addr[62547]= 2088416053;
assign addr[62548]= 2079176953;
assign addr[62549]= 2069278401;
assign addr[62550]= 2058723538;
assign addr[62551]= 2047515711;
assign addr[62552]= 2035658475;
assign addr[62553]= 2023155591;
assign addr[62554]= 2010011024;
assign addr[62555]= 1996228943;
assign addr[62556]= 1981813720;
assign addr[62557]= 1966769926;
assign addr[62558]= 1951102334;
assign addr[62559]= 1934815911;
assign addr[62560]= 1917915825;
assign addr[62561]= 1900407434;
assign addr[62562]= 1882296293;
assign addr[62563]= 1863588145;
assign addr[62564]= 1844288924;
assign addr[62565]= 1824404752;
assign addr[62566]= 1803941934;
assign addr[62567]= 1782906961;
assign addr[62568]= 1761306505;
assign addr[62569]= 1739147417;
assign addr[62570]= 1716436725;
assign addr[62571]= 1693181631;
assign addr[62572]= 1669389513;
assign addr[62573]= 1645067915;
assign addr[62574]= 1620224553;
assign addr[62575]= 1594867305;
assign addr[62576]= 1569004214;
assign addr[62577]= 1542643483;
assign addr[62578]= 1515793473;
assign addr[62579]= 1488462700;
assign addr[62580]= 1460659832;
assign addr[62581]= 1432393688;
assign addr[62582]= 1403673233;
assign addr[62583]= 1374507575;
assign addr[62584]= 1344905966;
assign addr[62585]= 1314877795;
assign addr[62586]= 1284432584;
assign addr[62587]= 1253579991;
assign addr[62588]= 1222329801;
assign addr[62589]= 1190691925;
assign addr[62590]= 1158676398;
assign addr[62591]= 1126293375;
assign addr[62592]= 1093553126;
assign addr[62593]= 1060466036;
assign addr[62594]= 1027042599;
assign addr[62595]= 993293415;
assign addr[62596]= 959229189;
assign addr[62597]= 924860725;
assign addr[62598]= 890198924;
assign addr[62599]= 855254778;
assign addr[62600]= 820039373;
assign addr[62601]= 784563876;
assign addr[62602]= 748839539;
assign addr[62603]= 712877694;
assign addr[62604]= 676689746;
assign addr[62605]= 640287172;
assign addr[62606]= 603681519;
assign addr[62607]= 566884397;
assign addr[62608]= 529907477;
assign addr[62609]= 492762486;
assign addr[62610]= 455461206;
assign addr[62611]= 418015468;
assign addr[62612]= 380437148;
assign addr[62613]= 342738165;
assign addr[62614]= 304930476;
assign addr[62615]= 267026072;
assign addr[62616]= 229036977;
assign addr[62617]= 190975237;
assign addr[62618]= 152852926;
assign addr[62619]= 114682135;
assign addr[62620]= 76474970;
assign addr[62621]= 38243550;
assign addr[62622]= 0;
assign addr[62623]= -38243550;
assign addr[62624]= -76474970;
assign addr[62625]= -114682135;
assign addr[62626]= -152852926;
assign addr[62627]= -190975237;
assign addr[62628]= -229036977;
assign addr[62629]= -267026072;
assign addr[62630]= -304930476;
assign addr[62631]= -342738165;
assign addr[62632]= -380437148;
assign addr[62633]= -418015468;
assign addr[62634]= -455461206;
assign addr[62635]= -492762486;
assign addr[62636]= -529907477;
assign addr[62637]= -566884397;
assign addr[62638]= -603681519;
assign addr[62639]= -640287172;
assign addr[62640]= -676689746;
assign addr[62641]= -712877694;
assign addr[62642]= -748839539;
assign addr[62643]= -784563876;
assign addr[62644]= -820039373;
assign addr[62645]= -855254778;
assign addr[62646]= -890198924;
assign addr[62647]= -924860725;
assign addr[62648]= -959229189;
assign addr[62649]= -993293415;
assign addr[62650]= -1027042599;
assign addr[62651]= -1060466036;
assign addr[62652]= -1093553126;
assign addr[62653]= -1126293375;
assign addr[62654]= -1158676398;
assign addr[62655]= -1190691925;
assign addr[62656]= -1222329801;
assign addr[62657]= -1253579991;
assign addr[62658]= -1284432584;
assign addr[62659]= -1314877795;
assign addr[62660]= -1344905966;
assign addr[62661]= -1374507575;
assign addr[62662]= -1403673233;
assign addr[62663]= -1432393688;
assign addr[62664]= -1460659832;
assign addr[62665]= -1488462700;
assign addr[62666]= -1515793473;
assign addr[62667]= -1542643483;
assign addr[62668]= -1569004214;
assign addr[62669]= -1594867305;
assign addr[62670]= -1620224553;
assign addr[62671]= -1645067915;
assign addr[62672]= -1669389513;
assign addr[62673]= -1693181631;
assign addr[62674]= -1716436725;
assign addr[62675]= -1739147417;
assign addr[62676]= -1761306505;
assign addr[62677]= -1782906961;
assign addr[62678]= -1803941934;
assign addr[62679]= -1824404752;
assign addr[62680]= -1844288924;
assign addr[62681]= -1863588145;
assign addr[62682]= -1882296293;
assign addr[62683]= -1900407434;
assign addr[62684]= -1917915825;
assign addr[62685]= -1934815911;
assign addr[62686]= -1951102334;
assign addr[62687]= -1966769926;
assign addr[62688]= -1981813720;
assign addr[62689]= -1996228943;
assign addr[62690]= -2010011024;
assign addr[62691]= -2023155591;
assign addr[62692]= -2035658475;
assign addr[62693]= -2047515711;
assign addr[62694]= -2058723538;
assign addr[62695]= -2069278401;
assign addr[62696]= -2079176953;
assign addr[62697]= -2088416053;
assign addr[62698]= -2096992772;
assign addr[62699]= -2104904390;
assign addr[62700]= -2112148396;
assign addr[62701]= -2118722494;
assign addr[62702]= -2124624598;
assign addr[62703]= -2129852837;
assign addr[62704]= -2134405552;
assign addr[62705]= -2138281298;
assign addr[62706]= -2141478848;
assign addr[62707]= -2143997187;
assign addr[62708]= -2145835515;
assign addr[62709]= -2146993250;
assign addr[62710]= -2147470025;
assign addr[62711]= -2147265689;
assign addr[62712]= -2146380306;
assign addr[62713]= -2144814157;
assign addr[62714]= -2142567738;
assign addr[62715]= -2139641764;
assign addr[62716]= -2136037160;
assign addr[62717]= -2131755071;
assign addr[62718]= -2126796855;
assign addr[62719]= -2121164085;
assign addr[62720]= -2114858546;
assign addr[62721]= -2107882239;
assign addr[62722]= -2100237377;
assign addr[62723]= -2091926384;
assign addr[62724]= -2082951896;
assign addr[62725]= -2073316760;
assign addr[62726]= -2063024031;
assign addr[62727]= -2052076975;
assign addr[62728]= -2040479063;
assign addr[62729]= -2028233973;
assign addr[62730]= -2015345591;
assign addr[62731]= -2001818002;
assign addr[62732]= -1987655498;
assign addr[62733]= -1972862571;
assign addr[62734]= -1957443913;
assign addr[62735]= -1941404413;
assign addr[62736]= -1924749160;
assign addr[62737]= -1907483436;
assign addr[62738]= -1889612716;
assign addr[62739]= -1871142669;
assign addr[62740]= -1852079154;
assign addr[62741]= -1832428215;
assign addr[62742]= -1812196087;
assign addr[62743]= -1791389186;
assign addr[62744]= -1770014111;
assign addr[62745]= -1748077642;
assign addr[62746]= -1725586737;
assign addr[62747]= -1702548529;
assign addr[62748]= -1678970324;
assign addr[62749]= -1654859602;
assign addr[62750]= -1630224009;
assign addr[62751]= -1605071359;
assign addr[62752]= -1579409630;
assign addr[62753]= -1553246960;
assign addr[62754]= -1526591649;
assign addr[62755]= -1499452149;
assign addr[62756]= -1471837070;
assign addr[62757]= -1443755168;
assign addr[62758]= -1415215352;
assign addr[62759]= -1386226674;
assign addr[62760]= -1356798326;
assign addr[62761]= -1326939644;
assign addr[62762]= -1296660098;
assign addr[62763]= -1265969291;
assign addr[62764]= -1234876957;
assign addr[62765]= -1203392958;
assign addr[62766]= -1171527280;
assign addr[62767]= -1139290029;
assign addr[62768]= -1106691431;
assign addr[62769]= -1073741824;
assign addr[62770]= -1040451659;
assign addr[62771]= -1006831495;
assign addr[62772]= -972891995;
assign addr[62773]= -938643924;
assign addr[62774]= -904098143;
assign addr[62775]= -869265610;
assign addr[62776]= -834157373;
assign addr[62777]= -798784567;
assign addr[62778]= -763158411;
assign addr[62779]= -727290205;
assign addr[62780]= -691191324;
assign addr[62781]= -654873219;
assign addr[62782]= -618347408;
assign addr[62783]= -581625477;
assign addr[62784]= -544719071;
assign addr[62785]= -507639898;
assign addr[62786]= -470399716;
assign addr[62787]= -433010339;
assign addr[62788]= -395483624;
assign addr[62789]= -357831473;
assign addr[62790]= -320065829;
assign addr[62791]= -282198671;
assign addr[62792]= -244242007;
assign addr[62793]= -206207878;
assign addr[62794]= -168108346;
assign addr[62795]= -129955495;
assign addr[62796]= -91761426;
assign addr[62797]= -53538253;
assign addr[62798]= -15298099;
assign addr[62799]= 22946906;
assign addr[62800]= 61184634;
assign addr[62801]= 99402956;
assign addr[62802]= 137589750;
assign addr[62803]= 175732905;
assign addr[62804]= 213820322;
assign addr[62805]= 251839923;
assign addr[62806]= 289779648;
assign addr[62807]= 327627463;
assign addr[62808]= 365371365;
assign addr[62809]= 402999383;
assign addr[62810]= 440499581;
assign addr[62811]= 477860067;
assign addr[62812]= 515068990;
assign addr[62813]= 552114549;
assign addr[62814]= 588984994;
assign addr[62815]= 625668632;
assign addr[62816]= 662153826;
assign addr[62817]= 698429006;
assign addr[62818]= 734482665;
assign addr[62819]= 770303369;
assign addr[62820]= 805879757;
assign addr[62821]= 841200544;
assign addr[62822]= 876254528;
assign addr[62823]= 911030591;
assign addr[62824]= 945517704;
assign addr[62825]= 979704927;
assign addr[62826]= 1013581418;
assign addr[62827]= 1047136432;
assign addr[62828]= 1080359326;
assign addr[62829]= 1113239564;
assign addr[62830]= 1145766716;
assign addr[62831]= 1177930466;
assign addr[62832]= 1209720613;
assign addr[62833]= 1241127074;
assign addr[62834]= 1272139887;
assign addr[62835]= 1302749217;
assign addr[62836]= 1332945355;
assign addr[62837]= 1362718723;
assign addr[62838]= 1392059879;
assign addr[62839]= 1420959516;
assign addr[62840]= 1449408469;
assign addr[62841]= 1477397714;
assign addr[62842]= 1504918373;
assign addr[62843]= 1531961719;
assign addr[62844]= 1558519173;
assign addr[62845]= 1584582314;
assign addr[62846]= 1610142873;
assign addr[62847]= 1635192744;
assign addr[62848]= 1659723983;
assign addr[62849]= 1683728808;
assign addr[62850]= 1707199606;
assign addr[62851]= 1730128933;
assign addr[62852]= 1752509516;
assign addr[62853]= 1774334257;
assign addr[62854]= 1795596234;
assign addr[62855]= 1816288703;
assign addr[62856]= 1836405100;
assign addr[62857]= 1855939047;
assign addr[62858]= 1874884346;
assign addr[62859]= 1893234990;
assign addr[62860]= 1910985158;
assign addr[62861]= 1928129220;
assign addr[62862]= 1944661739;
assign addr[62863]= 1960577471;
assign addr[62864]= 1975871368;
assign addr[62865]= 1990538579;
assign addr[62866]= 2004574453;
assign addr[62867]= 2017974537;
assign addr[62868]= 2030734582;
assign addr[62869]= 2042850540;
assign addr[62870]= 2054318569;
assign addr[62871]= 2065135031;
assign addr[62872]= 2075296495;
assign addr[62873]= 2084799740;
assign addr[62874]= 2093641749;
assign addr[62875]= 2101819720;
assign addr[62876]= 2109331059;
assign addr[62877]= 2116173382;
assign addr[62878]= 2122344521;
assign addr[62879]= 2127842516;
assign addr[62880]= 2132665626;
assign addr[62881]= 2136812319;
assign addr[62882]= 2140281282;
assign addr[62883]= 2143071413;
assign addr[62884]= 2145181827;
assign addr[62885]= 2146611856;
assign addr[62886]= 2147361045;
assign addr[62887]= 2147429158;
assign addr[62888]= 2146816171;
assign addr[62889]= 2145522281;
assign addr[62890]= 2143547897;
assign addr[62891]= 2140893646;
assign addr[62892]= 2137560369;
assign addr[62893]= 2133549123;
assign addr[62894]= 2128861181;
assign addr[62895]= 2123498030;
assign addr[62896]= 2117461370;
assign addr[62897]= 2110753117;
assign addr[62898]= 2103375398;
assign addr[62899]= 2095330553;
assign addr[62900]= 2086621133;
assign addr[62901]= 2077249901;
assign addr[62902]= 2067219829;
assign addr[62903]= 2056534099;
assign addr[62904]= 2045196100;
assign addr[62905]= 2033209426;
assign addr[62906]= 2020577882;
assign addr[62907]= 2007305472;
assign addr[62908]= 1993396407;
assign addr[62909]= 1978855097;
assign addr[62910]= 1963686155;
assign addr[62911]= 1947894393;
assign addr[62912]= 1931484818;
assign addr[62913]= 1914462636;
assign addr[62914]= 1896833245;
assign addr[62915]= 1878602237;
assign addr[62916]= 1859775393;
assign addr[62917]= 1840358687;
assign addr[62918]= 1820358275;
assign addr[62919]= 1799780501;
assign addr[62920]= 1778631892;
assign addr[62921]= 1756919156;
assign addr[62922]= 1734649179;
assign addr[62923]= 1711829025;
assign addr[62924]= 1688465931;
assign addr[62925]= 1664567307;
assign addr[62926]= 1640140734;
assign addr[62927]= 1615193959;
assign addr[62928]= 1589734894;
assign addr[62929]= 1563771613;
assign addr[62930]= 1537312353;
assign addr[62931]= 1510365504;
assign addr[62932]= 1482939614;
assign addr[62933]= 1455043381;
assign addr[62934]= 1426685652;
assign addr[62935]= 1397875423;
assign addr[62936]= 1368621831;
assign addr[62937]= 1338934154;
assign addr[62938]= 1308821808;
assign addr[62939]= 1278294345;
assign addr[62940]= 1247361445;
assign addr[62941]= 1216032921;
assign addr[62942]= 1184318708;
assign addr[62943]= 1152228866;
assign addr[62944]= 1119773573;
assign addr[62945]= 1086963121;
assign addr[62946]= 1053807919;
assign addr[62947]= 1020318481;
assign addr[62948]= 986505429;
assign addr[62949]= 952379488;
assign addr[62950]= 917951481;
assign addr[62951]= 883232329;
assign addr[62952]= 848233042;
assign addr[62953]= 812964722;
assign addr[62954]= 777438554;
assign addr[62955]= 741665807;
assign addr[62956]= 705657826;
assign addr[62957]= 669426032;
assign addr[62958]= 632981917;
assign addr[62959]= 596337040;
assign addr[62960]= 559503022;
assign addr[62961]= 522491548;
assign addr[62962]= 485314355;
assign addr[62963]= 447983235;
assign addr[62964]= 410510029;
assign addr[62965]= 372906622;
assign addr[62966]= 335184940;
assign addr[62967]= 297356948;
assign addr[62968]= 259434643;
assign addr[62969]= 221430054;
assign addr[62970]= 183355234;
assign addr[62971]= 145222259;
assign addr[62972]= 107043224;
assign addr[62973]= 68830239;
assign addr[62974]= 30595422;
assign addr[62975]= -7649098;
assign addr[62976]= -45891193;
assign addr[62977]= -84118732;
assign addr[62978]= -122319591;
assign addr[62979]= -160481654;
assign addr[62980]= -198592817;
assign addr[62981]= -236640993;
assign addr[62982]= -274614114;
assign addr[62983]= -312500135;
assign addr[62984]= -350287041;
assign addr[62985]= -387962847;
assign addr[62986]= -425515602;
assign addr[62987]= -462933398;
assign addr[62988]= -500204365;
assign addr[62989]= -537316682;
assign addr[62990]= -574258580;
assign addr[62991]= -611018340;
assign addr[62992]= -647584304;
assign addr[62993]= -683944874;
assign addr[62994]= -720088517;
assign addr[62995]= -756003771;
assign addr[62996]= -791679244;
assign addr[62997]= -827103620;
assign addr[62998]= -862265664;
assign addr[62999]= -897154224;
assign addr[63000]= -931758235;
assign addr[63001]= -966066720;
assign addr[63002]= -1000068799;
assign addr[63003]= -1033753687;
assign addr[63004]= -1067110699;
assign addr[63005]= -1100129257;
assign addr[63006]= -1132798888;
assign addr[63007]= -1165109230;
assign addr[63008]= -1197050035;
assign addr[63009]= -1228611172;
assign addr[63010]= -1259782632;
assign addr[63011]= -1290554528;
assign addr[63012]= -1320917099;
assign addr[63013]= -1350860716;
assign addr[63014]= -1380375881;
assign addr[63015]= -1409453233;
assign addr[63016]= -1438083551;
assign addr[63017]= -1466257752;
assign addr[63018]= -1493966902;
assign addr[63019]= -1521202211;
assign addr[63020]= -1547955041;
assign addr[63021]= -1574216908;
assign addr[63022]= -1599979481;
assign addr[63023]= -1625234591;
assign addr[63024]= -1649974225;
assign addr[63025]= -1674190539;
assign addr[63026]= -1697875851;
assign addr[63027]= -1721022648;
assign addr[63028]= -1743623590;
assign addr[63029]= -1765671509;
assign addr[63030]= -1787159411;
assign addr[63031]= -1808080480;
assign addr[63032]= -1828428082;
assign addr[63033]= -1848195763;
assign addr[63034]= -1867377253;
assign addr[63035]= -1885966468;
assign addr[63036]= -1903957513;
assign addr[63037]= -1921344681;
assign addr[63038]= -1938122457;
assign addr[63039]= -1954285520;
assign addr[63040]= -1969828744;
assign addr[63041]= -1984747199;
assign addr[63042]= -1999036154;
assign addr[63043]= -2012691075;
assign addr[63044]= -2025707632;
assign addr[63045]= -2038081698;
assign addr[63046]= -2049809346;
assign addr[63047]= -2060886858;
assign addr[63048]= -2071310720;
assign addr[63049]= -2081077626;
assign addr[63050]= -2090184478;
assign addr[63051]= -2098628387;
assign addr[63052]= -2106406677;
assign addr[63053]= -2113516878;
assign addr[63054]= -2119956737;
assign addr[63055]= -2125724211;
assign addr[63056]= -2130817471;
assign addr[63057]= -2135234901;
assign addr[63058]= -2138975100;
assign addr[63059]= -2142036881;
assign addr[63060]= -2144419275;
assign addr[63061]= -2146121524;
assign addr[63062]= -2147143090;
assign addr[63063]= -2147483648;
assign addr[63064]= -2147143090;
assign addr[63065]= -2146121524;
assign addr[63066]= -2144419275;
assign addr[63067]= -2142036881;
assign addr[63068]= -2138975100;
assign addr[63069]= -2135234901;
assign addr[63070]= -2130817471;
assign addr[63071]= -2125724211;
assign addr[63072]= -2119956737;
assign addr[63073]= -2113516878;
assign addr[63074]= -2106406677;
assign addr[63075]= -2098628387;
assign addr[63076]= -2090184478;
assign addr[63077]= -2081077626;
assign addr[63078]= -2071310720;
assign addr[63079]= -2060886858;
assign addr[63080]= -2049809346;
assign addr[63081]= -2038081698;
assign addr[63082]= -2025707632;
assign addr[63083]= -2012691075;
assign addr[63084]= -1999036154;
assign addr[63085]= -1984747199;
assign addr[63086]= -1969828744;
assign addr[63087]= -1954285520;
assign addr[63088]= -1938122457;
assign addr[63089]= -1921344681;
assign addr[63090]= -1903957513;
assign addr[63091]= -1885966468;
assign addr[63092]= -1867377253;
assign addr[63093]= -1848195763;
assign addr[63094]= -1828428082;
assign addr[63095]= -1808080480;
assign addr[63096]= -1787159411;
assign addr[63097]= -1765671509;
assign addr[63098]= -1743623590;
assign addr[63099]= -1721022648;
assign addr[63100]= -1697875851;
assign addr[63101]= -1674190539;
assign addr[63102]= -1649974225;
assign addr[63103]= -1625234591;
assign addr[63104]= -1599979481;
assign addr[63105]= -1574216908;
assign addr[63106]= -1547955041;
assign addr[63107]= -1521202211;
assign addr[63108]= -1493966902;
assign addr[63109]= -1466257752;
assign addr[63110]= -1438083551;
assign addr[63111]= -1409453233;
assign addr[63112]= -1380375881;
assign addr[63113]= -1350860716;
assign addr[63114]= -1320917099;
assign addr[63115]= -1290554528;
assign addr[63116]= -1259782632;
assign addr[63117]= -1228611172;
assign addr[63118]= -1197050035;
assign addr[63119]= -1165109230;
assign addr[63120]= -1132798888;
assign addr[63121]= -1100129257;
assign addr[63122]= -1067110699;
assign addr[63123]= -1033753687;
assign addr[63124]= -1000068799;
assign addr[63125]= -966066720;
assign addr[63126]= -931758235;
assign addr[63127]= -897154224;
assign addr[63128]= -862265664;
assign addr[63129]= -827103620;
assign addr[63130]= -791679244;
assign addr[63131]= -756003771;
assign addr[63132]= -720088517;
assign addr[63133]= -683944874;
assign addr[63134]= -647584304;
assign addr[63135]= -611018340;
assign addr[63136]= -574258580;
assign addr[63137]= -537316682;
assign addr[63138]= -500204365;
assign addr[63139]= -462933398;
assign addr[63140]= -425515602;
assign addr[63141]= -387962847;
assign addr[63142]= -350287041;
assign addr[63143]= -312500135;
assign addr[63144]= -274614114;
assign addr[63145]= -236640993;
assign addr[63146]= -198592817;
assign addr[63147]= -160481654;
assign addr[63148]= -122319591;
assign addr[63149]= -84118732;
assign addr[63150]= -45891193;
assign addr[63151]= -7649098;
assign addr[63152]= 30595422;
assign addr[63153]= 68830239;
assign addr[63154]= 107043224;
assign addr[63155]= 145222259;
assign addr[63156]= 183355234;
assign addr[63157]= 221430054;
assign addr[63158]= 259434643;
assign addr[63159]= 297356948;
assign addr[63160]= 335184940;
assign addr[63161]= 372906622;
assign addr[63162]= 410510029;
assign addr[63163]= 447983235;
assign addr[63164]= 485314355;
assign addr[63165]= 522491548;
assign addr[63166]= 559503022;
assign addr[63167]= 596337040;
assign addr[63168]= 632981917;
assign addr[63169]= 669426032;
assign addr[63170]= 705657826;
assign addr[63171]= 741665807;
assign addr[63172]= 777438554;
assign addr[63173]= 812964722;
assign addr[63174]= 848233042;
assign addr[63175]= 883232329;
assign addr[63176]= 917951481;
assign addr[63177]= 952379488;
assign addr[63178]= 986505429;
assign addr[63179]= 1020318481;
assign addr[63180]= 1053807919;
assign addr[63181]= 1086963121;
assign addr[63182]= 1119773573;
assign addr[63183]= 1152228866;
assign addr[63184]= 1184318708;
assign addr[63185]= 1216032921;
assign addr[63186]= 1247361445;
assign addr[63187]= 1278294345;
assign addr[63188]= 1308821808;
assign addr[63189]= 1338934154;
assign addr[63190]= 1368621831;
assign addr[63191]= 1397875423;
assign addr[63192]= 1426685652;
assign addr[63193]= 1455043381;
assign addr[63194]= 1482939614;
assign addr[63195]= 1510365504;
assign addr[63196]= 1537312353;
assign addr[63197]= 1563771613;
assign addr[63198]= 1589734894;
assign addr[63199]= 1615193959;
assign addr[63200]= 1640140734;
assign addr[63201]= 1664567307;
assign addr[63202]= 1688465931;
assign addr[63203]= 1711829025;
assign addr[63204]= 1734649179;
assign addr[63205]= 1756919156;
assign addr[63206]= 1778631892;
assign addr[63207]= 1799780501;
assign addr[63208]= 1820358275;
assign addr[63209]= 1840358687;
assign addr[63210]= 1859775393;
assign addr[63211]= 1878602237;
assign addr[63212]= 1896833245;
assign addr[63213]= 1914462636;
assign addr[63214]= 1931484818;
assign addr[63215]= 1947894393;
assign addr[63216]= 1963686155;
assign addr[63217]= 1978855097;
assign addr[63218]= 1993396407;
assign addr[63219]= 2007305472;
assign addr[63220]= 2020577882;
assign addr[63221]= 2033209426;
assign addr[63222]= 2045196100;
assign addr[63223]= 2056534099;
assign addr[63224]= 2067219829;
assign addr[63225]= 2077249901;
assign addr[63226]= 2086621133;
assign addr[63227]= 2095330553;
assign addr[63228]= 2103375398;
assign addr[63229]= 2110753117;
assign addr[63230]= 2117461370;
assign addr[63231]= 2123498030;
assign addr[63232]= 2128861181;
assign addr[63233]= 2133549123;
assign addr[63234]= 2137560369;
assign addr[63235]= 2140893646;
assign addr[63236]= 2143547897;
assign addr[63237]= 2145522281;
assign addr[63238]= 2146816171;
assign addr[63239]= 2147429158;
assign addr[63240]= 2147361045;
assign addr[63241]= 2146611856;
assign addr[63242]= 2145181827;
assign addr[63243]= 2143071413;
assign addr[63244]= 2140281282;
assign addr[63245]= 2136812319;
assign addr[63246]= 2132665626;
assign addr[63247]= 2127842516;
assign addr[63248]= 2122344521;
assign addr[63249]= 2116173382;
assign addr[63250]= 2109331059;
assign addr[63251]= 2101819720;
assign addr[63252]= 2093641749;
assign addr[63253]= 2084799740;
assign addr[63254]= 2075296495;
assign addr[63255]= 2065135031;
assign addr[63256]= 2054318569;
assign addr[63257]= 2042850540;
assign addr[63258]= 2030734582;
assign addr[63259]= 2017974537;
assign addr[63260]= 2004574453;
assign addr[63261]= 1990538579;
assign addr[63262]= 1975871368;
assign addr[63263]= 1960577471;
assign addr[63264]= 1944661739;
assign addr[63265]= 1928129220;
assign addr[63266]= 1910985158;
assign addr[63267]= 1893234990;
assign addr[63268]= 1874884346;
assign addr[63269]= 1855939047;
assign addr[63270]= 1836405100;
assign addr[63271]= 1816288703;
assign addr[63272]= 1795596234;
assign addr[63273]= 1774334257;
assign addr[63274]= 1752509516;
assign addr[63275]= 1730128933;
assign addr[63276]= 1707199606;
assign addr[63277]= 1683728808;
assign addr[63278]= 1659723983;
assign addr[63279]= 1635192744;
assign addr[63280]= 1610142873;
assign addr[63281]= 1584582314;
assign addr[63282]= 1558519173;
assign addr[63283]= 1531961719;
assign addr[63284]= 1504918373;
assign addr[63285]= 1477397714;
assign addr[63286]= 1449408469;
assign addr[63287]= 1420959516;
assign addr[63288]= 1392059879;
assign addr[63289]= 1362718723;
assign addr[63290]= 1332945355;
assign addr[63291]= 1302749217;
assign addr[63292]= 1272139887;
assign addr[63293]= 1241127074;
assign addr[63294]= 1209720613;
assign addr[63295]= 1177930466;
assign addr[63296]= 1145766716;
assign addr[63297]= 1113239564;
assign addr[63298]= 1080359326;
assign addr[63299]= 1047136432;
assign addr[63300]= 1013581418;
assign addr[63301]= 979704927;
assign addr[63302]= 945517704;
assign addr[63303]= 911030591;
assign addr[63304]= 876254528;
assign addr[63305]= 841200544;
assign addr[63306]= 805879757;
assign addr[63307]= 770303369;
assign addr[63308]= 734482665;
assign addr[63309]= 698429006;
assign addr[63310]= 662153826;
assign addr[63311]= 625668632;
assign addr[63312]= 588984994;
assign addr[63313]= 552114549;
assign addr[63314]= 515068990;
assign addr[63315]= 477860067;
assign addr[63316]= 440499581;
assign addr[63317]= 402999383;
assign addr[63318]= 365371365;
assign addr[63319]= 327627463;
assign addr[63320]= 289779648;
assign addr[63321]= 251839923;
assign addr[63322]= 213820322;
assign addr[63323]= 175732905;
assign addr[63324]= 137589750;
assign addr[63325]= 99402956;
assign addr[63326]= 61184634;
assign addr[63327]= 22946906;
assign addr[63328]= -15298099;
assign addr[63329]= -53538253;
assign addr[63330]= -91761426;
assign addr[63331]= -129955495;
assign addr[63332]= -168108346;
assign addr[63333]= -206207878;
assign addr[63334]= -244242007;
assign addr[63335]= -282198671;
assign addr[63336]= -320065829;
assign addr[63337]= -357831473;
assign addr[63338]= -395483624;
assign addr[63339]= -433010339;
assign addr[63340]= -470399716;
assign addr[63341]= -507639898;
assign addr[63342]= -544719071;
assign addr[63343]= -581625477;
assign addr[63344]= -618347408;
assign addr[63345]= -654873219;
assign addr[63346]= -691191324;
assign addr[63347]= -727290205;
assign addr[63348]= -763158411;
assign addr[63349]= -798784567;
assign addr[63350]= -834157373;
assign addr[63351]= -869265610;
assign addr[63352]= -904098143;
assign addr[63353]= -938643924;
assign addr[63354]= -972891995;
assign addr[63355]= -1006831495;
assign addr[63356]= -1040451659;
assign addr[63357]= -1073741824;
assign addr[63358]= -1106691431;
assign addr[63359]= -1139290029;
assign addr[63360]= -1171527280;
assign addr[63361]= -1203392958;
assign addr[63362]= -1234876957;
assign addr[63363]= -1265969291;
assign addr[63364]= -1296660098;
assign addr[63365]= -1326939644;
assign addr[63366]= -1356798326;
assign addr[63367]= -1386226674;
assign addr[63368]= -1415215352;
assign addr[63369]= -1443755168;
assign addr[63370]= -1471837070;
assign addr[63371]= -1499452149;
assign addr[63372]= -1526591649;
assign addr[63373]= -1553246960;
assign addr[63374]= -1579409630;
assign addr[63375]= -1605071359;
assign addr[63376]= -1630224009;
assign addr[63377]= -1654859602;
assign addr[63378]= -1678970324;
assign addr[63379]= -1702548529;
assign addr[63380]= -1725586737;
assign addr[63381]= -1748077642;
assign addr[63382]= -1770014111;
assign addr[63383]= -1791389186;
assign addr[63384]= -1812196087;
assign addr[63385]= -1832428215;
assign addr[63386]= -1852079154;
assign addr[63387]= -1871142669;
assign addr[63388]= -1889612716;
assign addr[63389]= -1907483436;
assign addr[63390]= -1924749160;
assign addr[63391]= -1941404413;
assign addr[63392]= -1957443913;
assign addr[63393]= -1972862571;
assign addr[63394]= -1987655498;
assign addr[63395]= -2001818002;
assign addr[63396]= -2015345591;
assign addr[63397]= -2028233973;
assign addr[63398]= -2040479063;
assign addr[63399]= -2052076975;
assign addr[63400]= -2063024031;
assign addr[63401]= -2073316760;
assign addr[63402]= -2082951896;
assign addr[63403]= -2091926384;
assign addr[63404]= -2100237377;
assign addr[63405]= -2107882239;
assign addr[63406]= -2114858546;
assign addr[63407]= -2121164085;
assign addr[63408]= -2126796855;
assign addr[63409]= -2131755071;
assign addr[63410]= -2136037160;
assign addr[63411]= -2139641764;
assign addr[63412]= -2142567738;
assign addr[63413]= -2144814157;
assign addr[63414]= -2146380306;
assign addr[63415]= -2147265689;
assign addr[63416]= -2147470025;
assign addr[63417]= -2146993250;
assign addr[63418]= -2145835515;
assign addr[63419]= -2143997187;
assign addr[63420]= -2141478848;
assign addr[63421]= -2138281298;
assign addr[63422]= -2134405552;
assign addr[63423]= -2129852837;
assign addr[63424]= -2124624598;
assign addr[63425]= -2118722494;
assign addr[63426]= -2112148396;
assign addr[63427]= -2104904390;
assign addr[63428]= -2096992772;
assign addr[63429]= -2088416053;
assign addr[63430]= -2079176953;
assign addr[63431]= -2069278401;
assign addr[63432]= -2058723538;
assign addr[63433]= -2047515711;
assign addr[63434]= -2035658475;
assign addr[63435]= -2023155591;
assign addr[63436]= -2010011024;
assign addr[63437]= -1996228943;
assign addr[63438]= -1981813720;
assign addr[63439]= -1966769926;
assign addr[63440]= -1951102334;
assign addr[63441]= -1934815911;
assign addr[63442]= -1917915825;
assign addr[63443]= -1900407434;
assign addr[63444]= -1882296293;
assign addr[63445]= -1863588145;
assign addr[63446]= -1844288924;
assign addr[63447]= -1824404752;
assign addr[63448]= -1803941934;
assign addr[63449]= -1782906961;
assign addr[63450]= -1761306505;
assign addr[63451]= -1739147417;
assign addr[63452]= -1716436725;
assign addr[63453]= -1693181631;
assign addr[63454]= -1669389513;
assign addr[63455]= -1645067915;
assign addr[63456]= -1620224553;
assign addr[63457]= -1594867305;
assign addr[63458]= -1569004214;
assign addr[63459]= -1542643483;
assign addr[63460]= -1515793473;
assign addr[63461]= -1488462700;
assign addr[63462]= -1460659832;
assign addr[63463]= -1432393688;
assign addr[63464]= -1403673233;
assign addr[63465]= -1374507575;
assign addr[63466]= -1344905966;
assign addr[63467]= -1314877795;
assign addr[63468]= -1284432584;
assign addr[63469]= -1253579991;
assign addr[63470]= -1222329801;
assign addr[63471]= -1190691925;
assign addr[63472]= -1158676398;
assign addr[63473]= -1126293375;
assign addr[63474]= -1093553126;
assign addr[63475]= -1060466036;
assign addr[63476]= -1027042599;
assign addr[63477]= -993293415;
assign addr[63478]= -959229189;
assign addr[63479]= -924860725;
assign addr[63480]= -890198924;
assign addr[63481]= -855254778;
assign addr[63482]= -820039373;
assign addr[63483]= -784563876;
assign addr[63484]= -748839539;
assign addr[63485]= -712877694;
assign addr[63486]= -676689746;
assign addr[63487]= -640287172;
assign addr[63488]= -603681519;
assign addr[63489]= -566884397;
assign addr[63490]= -529907477;
assign addr[63491]= -492762486;
assign addr[63492]= -455461206;
assign addr[63493]= -418015468;
assign addr[63494]= -380437148;
assign addr[63495]= -342738165;
assign addr[63496]= -304930476;
assign addr[63497]= -267026072;
assign addr[63498]= -229036977;
assign addr[63499]= -190975237;
assign addr[63500]= -152852926;
assign addr[63501]= -114682135;
assign addr[63502]= -76474970;
assign addr[63503]= -38243550;
assign addr[63504]= 0;
assign addr[63505]= 38243550;
assign addr[63506]= 76474970;
assign addr[63507]= 114682135;
assign addr[63508]= 152852926;
assign addr[63509]= 190975237;
assign addr[63510]= 229036977;
assign addr[63511]= 267026072;
assign addr[63512]= 304930476;
assign addr[63513]= 342738165;
assign addr[63514]= 380437148;
assign addr[63515]= 418015468;
assign addr[63516]= 455461206;
assign addr[63517]= 492762486;
assign addr[63518]= 529907477;
assign addr[63519]= 566884397;
assign addr[63520]= 603681519;
assign addr[63521]= 640287172;
assign addr[63522]= 676689746;
assign addr[63523]= 712877694;
assign addr[63524]= 748839539;
assign addr[63525]= 784563876;
assign addr[63526]= 820039373;
assign addr[63527]= 855254778;
assign addr[63528]= 890198924;
assign addr[63529]= 924860725;
assign addr[63530]= 959229189;
assign addr[63531]= 993293415;
assign addr[63532]= 1027042599;
assign addr[63533]= 1060466036;
assign addr[63534]= 1093553126;
assign addr[63535]= 1126293375;
assign addr[63536]= 1158676398;
assign addr[63537]= 1190691925;
assign addr[63538]= 1222329801;
assign addr[63539]= 1253579991;
assign addr[63540]= 1284432584;
assign addr[63541]= 1314877795;
assign addr[63542]= 1344905966;
assign addr[63543]= 1374507575;
assign addr[63544]= 1403673233;
assign addr[63545]= 1432393688;
assign addr[63546]= 1460659832;
assign addr[63547]= 1488462700;
assign addr[63548]= 1515793473;
assign addr[63549]= 1542643483;
assign addr[63550]= 1569004214;
assign addr[63551]= 1594867305;
assign addr[63552]= 1620224553;
assign addr[63553]= 1645067915;
assign addr[63554]= 1669389513;
assign addr[63555]= 1693181631;
assign addr[63556]= 1716436725;
assign addr[63557]= 1739147417;
assign addr[63558]= 1761306505;
assign addr[63559]= 1782906961;
assign addr[63560]= 1803941934;
assign addr[63561]= 1824404752;
assign addr[63562]= 1844288924;
assign addr[63563]= 1863588145;
assign addr[63564]= 1882296293;
assign addr[63565]= 1900407434;
assign addr[63566]= 1917915825;
assign addr[63567]= 1934815911;
assign addr[63568]= 1951102334;
assign addr[63569]= 1966769926;
assign addr[63570]= 1981813720;
assign addr[63571]= 1996228943;
assign addr[63572]= 2010011024;
assign addr[63573]= 2023155591;
assign addr[63574]= 2035658475;
assign addr[63575]= 2047515711;
assign addr[63576]= 2058723538;
assign addr[63577]= 2069278401;
assign addr[63578]= 2079176953;
assign addr[63579]= 2088416053;
assign addr[63580]= 2096992772;
assign addr[63581]= 2104904390;
assign addr[63582]= 2112148396;
assign addr[63583]= 2118722494;
assign addr[63584]= 2124624598;
assign addr[63585]= 2129852837;
assign addr[63586]= 2134405552;
assign addr[63587]= 2138281298;
assign addr[63588]= 2141478848;
assign addr[63589]= 2143997187;
assign addr[63590]= 2145835515;
assign addr[63591]= 2146993250;
assign addr[63592]= 2147470025;
assign addr[63593]= 2147265689;
assign addr[63594]= 2146380306;
assign addr[63595]= 2144814157;
assign addr[63596]= 2142567738;
assign addr[63597]= 2139641764;
assign addr[63598]= 2136037160;
assign addr[63599]= 2131755071;
assign addr[63600]= 2126796855;
assign addr[63601]= 2121164085;
assign addr[63602]= 2114858546;
assign addr[63603]= 2107882239;
assign addr[63604]= 2100237377;
assign addr[63605]= 2091926384;
assign addr[63606]= 2082951896;
assign addr[63607]= 2073316760;
assign addr[63608]= 2063024031;
assign addr[63609]= 2052076975;
assign addr[63610]= 2040479063;
assign addr[63611]= 2028233973;
assign addr[63612]= 2015345591;
assign addr[63613]= 2001818002;
assign addr[63614]= 1987655498;
assign addr[63615]= 1972862571;
assign addr[63616]= 1957443913;
assign addr[63617]= 1941404413;
assign addr[63618]= 1924749160;
assign addr[63619]= 1907483436;
assign addr[63620]= 1889612716;
assign addr[63621]= 1871142669;
assign addr[63622]= 1852079154;
assign addr[63623]= 1832428215;
assign addr[63624]= 1812196087;
assign addr[63625]= 1791389186;
assign addr[63626]= 1770014111;
assign addr[63627]= 1748077642;
assign addr[63628]= 1725586737;
assign addr[63629]= 1702548529;
assign addr[63630]= 1678970324;
assign addr[63631]= 1654859602;
assign addr[63632]= 1630224009;
assign addr[63633]= 1605071359;
assign addr[63634]= 1579409630;
assign addr[63635]= 1553246960;
assign addr[63636]= 1526591649;
assign addr[63637]= 1499452149;
assign addr[63638]= 1471837070;
assign addr[63639]= 1443755168;
assign addr[63640]= 1415215352;
assign addr[63641]= 1386226674;
assign addr[63642]= 1356798326;
assign addr[63643]= 1326939644;
assign addr[63644]= 1296660098;
assign addr[63645]= 1265969291;
assign addr[63646]= 1234876957;
assign addr[63647]= 1203392958;
assign addr[63648]= 1171527280;
assign addr[63649]= 1139290029;
assign addr[63650]= 1106691431;
assign addr[63651]= 1073741824;
assign addr[63652]= 1040451659;
assign addr[63653]= 1006831495;
assign addr[63654]= 972891995;
assign addr[63655]= 938643924;
assign addr[63656]= 904098143;
assign addr[63657]= 869265610;
assign addr[63658]= 834157373;
assign addr[63659]= 798784567;
assign addr[63660]= 763158411;
assign addr[63661]= 727290205;
assign addr[63662]= 691191324;
assign addr[63663]= 654873219;
assign addr[63664]= 618347408;
assign addr[63665]= 581625477;
assign addr[63666]= 544719071;
assign addr[63667]= 507639898;
assign addr[63668]= 470399716;
assign addr[63669]= 433010339;
assign addr[63670]= 395483624;
assign addr[63671]= 357831473;
assign addr[63672]= 320065829;
assign addr[63673]= 282198671;
assign addr[63674]= 244242007;
assign addr[63675]= 206207878;
assign addr[63676]= 168108346;
assign addr[63677]= 129955495;
assign addr[63678]= 91761426;
assign addr[63679]= 53538253;
assign addr[63680]= 15298099;
assign addr[63681]= -22946906;
assign addr[63682]= -61184634;
assign addr[63683]= -99402956;
assign addr[63684]= -137589750;
assign addr[63685]= -175732905;
assign addr[63686]= -213820322;
assign addr[63687]= -251839923;
assign addr[63688]= -289779648;
assign addr[63689]= -327627463;
assign addr[63690]= -365371365;
assign addr[63691]= -402999383;
assign addr[63692]= -440499581;
assign addr[63693]= -477860067;
assign addr[63694]= -515068990;
assign addr[63695]= -552114549;
assign addr[63696]= -588984994;
assign addr[63697]= -625668632;
assign addr[63698]= -662153826;
assign addr[63699]= -698429006;
assign addr[63700]= -734482665;
assign addr[63701]= -770303369;
assign addr[63702]= -805879757;
assign addr[63703]= -841200544;
assign addr[63704]= -876254528;
assign addr[63705]= -911030591;
assign addr[63706]= -945517704;
assign addr[63707]= -979704927;
assign addr[63708]= -1013581418;
assign addr[63709]= -1047136432;
assign addr[63710]= -1080359326;
assign addr[63711]= -1113239564;
assign addr[63712]= -1145766716;
assign addr[63713]= -1177930466;
assign addr[63714]= -1209720613;
assign addr[63715]= -1241127074;
assign addr[63716]= -1272139887;
assign addr[63717]= -1302749217;
assign addr[63718]= -1332945355;
assign addr[63719]= -1362718723;
assign addr[63720]= -1392059879;
assign addr[63721]= -1420959516;
assign addr[63722]= -1449408469;
assign addr[63723]= -1477397714;
assign addr[63724]= -1504918373;
assign addr[63725]= -1531961719;
assign addr[63726]= -1558519173;
assign addr[63727]= -1584582314;
assign addr[63728]= -1610142873;
assign addr[63729]= -1635192744;
assign addr[63730]= -1659723983;
assign addr[63731]= -1683728808;
assign addr[63732]= -1707199606;
assign addr[63733]= -1730128933;
assign addr[63734]= -1752509516;
assign addr[63735]= -1774334257;
assign addr[63736]= -1795596234;
assign addr[63737]= -1816288703;
assign addr[63738]= -1836405100;
assign addr[63739]= -1855939047;
assign addr[63740]= -1874884346;
assign addr[63741]= -1893234990;
assign addr[63742]= -1910985158;
assign addr[63743]= -1928129220;
assign addr[63744]= -1944661739;
assign addr[63745]= -1960577471;
assign addr[63746]= -1975871368;
assign addr[63747]= -1990538579;
assign addr[63748]= -2004574453;
assign addr[63749]= -2017974537;
assign addr[63750]= -2030734582;
assign addr[63751]= -2042850540;
assign addr[63752]= -2054318569;
assign addr[63753]= -2065135031;
assign addr[63754]= -2075296495;
assign addr[63755]= -2084799740;
assign addr[63756]= -2093641749;
assign addr[63757]= -2101819720;
assign addr[63758]= -2109331059;
assign addr[63759]= -2116173382;
assign addr[63760]= -2122344521;
assign addr[63761]= -2127842516;
assign addr[63762]= -2132665626;
assign addr[63763]= -2136812319;
assign addr[63764]= -2140281282;
assign addr[63765]= -2143071413;
assign addr[63766]= -2145181827;
assign addr[63767]= -2146611856;
assign addr[63768]= -2147361045;
assign addr[63769]= -2147429158;
assign addr[63770]= -2146816171;
assign addr[63771]= -2145522281;
assign addr[63772]= -2143547897;
assign addr[63773]= -2140893646;
assign addr[63774]= -2137560369;
assign addr[63775]= -2133549123;
assign addr[63776]= -2128861181;
assign addr[63777]= -2123498030;
assign addr[63778]= -2117461370;
assign addr[63779]= -2110753117;
assign addr[63780]= -2103375398;
assign addr[63781]= -2095330553;
assign addr[63782]= -2086621133;
assign addr[63783]= -2077249901;
assign addr[63784]= -2067219829;
assign addr[63785]= -2056534099;
assign addr[63786]= -2045196100;
assign addr[63787]= -2033209426;
assign addr[63788]= -2020577882;
assign addr[63789]= -2007305472;
assign addr[63790]= -1993396407;
assign addr[63791]= -1978855097;
assign addr[63792]= -1963686155;
assign addr[63793]= -1947894393;
assign addr[63794]= -1931484818;
assign addr[63795]= -1914462636;
assign addr[63796]= -1896833245;
assign addr[63797]= -1878602237;
assign addr[63798]= -1859775393;
assign addr[63799]= -1840358687;
assign addr[63800]= -1820358275;
assign addr[63801]= -1799780501;
assign addr[63802]= -1778631892;
assign addr[63803]= -1756919156;
assign addr[63804]= -1734649179;
assign addr[63805]= -1711829025;
assign addr[63806]= -1688465931;
assign addr[63807]= -1664567307;
assign addr[63808]= -1640140734;
assign addr[63809]= -1615193959;
assign addr[63810]= -1589734894;
assign addr[63811]= -1563771613;
assign addr[63812]= -1537312353;
assign addr[63813]= -1510365504;
assign addr[63814]= -1482939614;
assign addr[63815]= -1455043381;
assign addr[63816]= -1426685652;
assign addr[63817]= -1397875423;
assign addr[63818]= -1368621831;
assign addr[63819]= -1338934154;
assign addr[63820]= -1308821808;
assign addr[63821]= -1278294345;
assign addr[63822]= -1247361445;
assign addr[63823]= -1216032921;
assign addr[63824]= -1184318708;
assign addr[63825]= -1152228866;
assign addr[63826]= -1119773573;
assign addr[63827]= -1086963121;
assign addr[63828]= -1053807919;
assign addr[63829]= -1020318481;
assign addr[63830]= -986505429;
assign addr[63831]= -952379488;
assign addr[63832]= -917951481;
assign addr[63833]= -883232329;
assign addr[63834]= -848233042;
assign addr[63835]= -812964722;
assign addr[63836]= -777438554;
assign addr[63837]= -741665807;
assign addr[63838]= -705657826;
assign addr[63839]= -669426032;
assign addr[63840]= -632981917;
assign addr[63841]= -596337040;
assign addr[63842]= -559503022;
assign addr[63843]= -522491548;
assign addr[63844]= -485314355;
assign addr[63845]= -447983235;
assign addr[63846]= -410510029;
assign addr[63847]= -372906622;
assign addr[63848]= -335184940;
assign addr[63849]= -297356948;
assign addr[63850]= -259434643;
assign addr[63851]= -221430054;
assign addr[63852]= -183355234;
assign addr[63853]= -145222259;
assign addr[63854]= -107043224;
assign addr[63855]= -68830239;
assign addr[63856]= -30595422;
assign addr[63857]= 7649098;
assign addr[63858]= 45891193;
assign addr[63859]= 84118732;
assign addr[63860]= 122319591;
assign addr[63861]= 160481654;
assign addr[63862]= 198592817;
assign addr[63863]= 236640993;
assign addr[63864]= 274614114;
assign addr[63865]= 312500135;
assign addr[63866]= 350287041;
assign addr[63867]= 387962847;
assign addr[63868]= 425515602;
assign addr[63869]= 462933398;
assign addr[63870]= 500204365;
assign addr[63871]= 537316682;
assign addr[63872]= 574258580;
assign addr[63873]= 611018340;
assign addr[63874]= 647584304;
assign addr[63875]= 683944874;
assign addr[63876]= 720088517;
assign addr[63877]= 756003771;
assign addr[63878]= 791679244;
assign addr[63879]= 827103620;
assign addr[63880]= 862265664;
assign addr[63881]= 897154224;
assign addr[63882]= 931758235;
assign addr[63883]= 966066720;
assign addr[63884]= 1000068799;
assign addr[63885]= 1033753687;
assign addr[63886]= 1067110699;
assign addr[63887]= 1100129257;
assign addr[63888]= 1132798888;
assign addr[63889]= 1165109230;
assign addr[63890]= 1197050035;
assign addr[63891]= 1228611172;
assign addr[63892]= 1259782632;
assign addr[63893]= 1290554528;
assign addr[63894]= 1320917099;
assign addr[63895]= 1350860716;
assign addr[63896]= 1380375881;
assign addr[63897]= 1409453233;
assign addr[63898]= 1438083551;
assign addr[63899]= 1466257752;
assign addr[63900]= 1493966902;
assign addr[63901]= 1521202211;
assign addr[63902]= 1547955041;
assign addr[63903]= 1574216908;
assign addr[63904]= 1599979481;
assign addr[63905]= 1625234591;
assign addr[63906]= 1649974225;
assign addr[63907]= 1674190539;
assign addr[63908]= 1697875851;
assign addr[63909]= 1721022648;
assign addr[63910]= 1743623590;
assign addr[63911]= 1765671509;
assign addr[63912]= 1787159411;
assign addr[63913]= 1808080480;
assign addr[63914]= 1828428082;
assign addr[63915]= 1848195763;
assign addr[63916]= 1867377253;
assign addr[63917]= 1885966468;
assign addr[63918]= 1903957513;
assign addr[63919]= 1921344681;
assign addr[63920]= 1938122457;
assign addr[63921]= 1954285520;
assign addr[63922]= 1969828744;
assign addr[63923]= 1984747199;
assign addr[63924]= 1999036154;
assign addr[63925]= 2012691075;
assign addr[63926]= 2025707632;
assign addr[63927]= 2038081698;
assign addr[63928]= 2049809346;
assign addr[63929]= 2060886858;
assign addr[63930]= 2071310720;
assign addr[63931]= 2081077626;
assign addr[63932]= 2090184478;
assign addr[63933]= 2098628387;
assign addr[63934]= 2106406677;
assign addr[63935]= 2113516878;
assign addr[63936]= 2119956737;
assign addr[63937]= 2125724211;
assign addr[63938]= 2130817471;
assign addr[63939]= 2135234901;
assign addr[63940]= 2138975100;
assign addr[63941]= 2142036881;
assign addr[63942]= 2144419275;
assign addr[63943]= 2146121524;
assign addr[63944]= 2147143090;
assign addr[63945]= 2147483648;
assign addr[63946]= 2147143090;
assign addr[63947]= 2146121524;
assign addr[63948]= 2144419275;
assign addr[63949]= 2142036881;
assign addr[63950]= 2138975100;
assign addr[63951]= 2135234901;
assign addr[63952]= 2130817471;
assign addr[63953]= 2125724211;
assign addr[63954]= 2119956737;
assign addr[63955]= 2113516878;
assign addr[63956]= 2106406677;
assign addr[63957]= 2098628387;
assign addr[63958]= 2090184478;
assign addr[63959]= 2081077626;
assign addr[63960]= 2071310720;
assign addr[63961]= 2060886858;
assign addr[63962]= 2049809346;
assign addr[63963]= 2038081698;
assign addr[63964]= 2025707632;
assign addr[63965]= 2012691075;
assign addr[63966]= 1999036154;
assign addr[63967]= 1984747199;
assign addr[63968]= 1969828744;
assign addr[63969]= 1954285520;
assign addr[63970]= 1938122457;
assign addr[63971]= 1921344681;
assign addr[63972]= 1903957513;
assign addr[63973]= 1885966468;
assign addr[63974]= 1867377253;
assign addr[63975]= 1848195763;
assign addr[63976]= 1828428082;
assign addr[63977]= 1808080480;
assign addr[63978]= 1787159411;
assign addr[63979]= 1765671509;
assign addr[63980]= 1743623590;
assign addr[63981]= 1721022648;
assign addr[63982]= 1697875851;
assign addr[63983]= 1674190539;
assign addr[63984]= 1649974225;
assign addr[63985]= 1625234591;
assign addr[63986]= 1599979481;
assign addr[63987]= 1574216908;
assign addr[63988]= 1547955041;
assign addr[63989]= 1521202211;
assign addr[63990]= 1493966902;
assign addr[63991]= 1466257752;
assign addr[63992]= 1438083551;
assign addr[63993]= 1409453233;
assign addr[63994]= 1380375881;
assign addr[63995]= 1350860716;
assign addr[63996]= 1320917099;
assign addr[63997]= 1290554528;
assign addr[63998]= 1259782632;
assign addr[63999]= 1228611172;
assign addr[64000]= 1197050035;
assign addr[64001]= 1165109230;
assign addr[64002]= 1132798888;
assign addr[64003]= 1100129257;
assign addr[64004]= 1067110699;
assign addr[64005]= 1033753687;
assign addr[64006]= 1000068799;
assign addr[64007]= 966066720;
assign addr[64008]= 931758235;
assign addr[64009]= 897154224;
assign addr[64010]= 862265664;
assign addr[64011]= 827103620;
assign addr[64012]= 791679244;
assign addr[64013]= 756003771;
assign addr[64014]= 720088517;
assign addr[64015]= 683944874;
assign addr[64016]= 647584304;
assign addr[64017]= 611018340;
assign addr[64018]= 574258580;
assign addr[64019]= 537316682;
assign addr[64020]= 500204365;
assign addr[64021]= 462933398;
assign addr[64022]= 425515602;
assign addr[64023]= 387962847;
assign addr[64024]= 350287041;
assign addr[64025]= 312500135;
assign addr[64026]= 274614114;
assign addr[64027]= 236640993;
assign addr[64028]= 198592817;
assign addr[64029]= 160481654;
assign addr[64030]= 122319591;
assign addr[64031]= 84118732;
assign addr[64032]= 45891193;
assign addr[64033]= 7649098;
assign addr[64034]= -30595422;
assign addr[64035]= -68830239;
assign addr[64036]= -107043224;
assign addr[64037]= -145222259;
assign addr[64038]= -183355234;
assign addr[64039]= -221430054;
assign addr[64040]= -259434643;
assign addr[64041]= -297356948;
assign addr[64042]= -335184940;
assign addr[64043]= -372906622;
assign addr[64044]= -410510029;
assign addr[64045]= -447983235;
assign addr[64046]= -485314355;
assign addr[64047]= -522491548;
assign addr[64048]= -559503022;
assign addr[64049]= -596337040;
assign addr[64050]= -632981917;
assign addr[64051]= -669426032;
assign addr[64052]= -705657826;
assign addr[64053]= -741665807;
assign addr[64054]= -777438554;
assign addr[64055]= -812964722;
assign addr[64056]= -848233042;
assign addr[64057]= -883232329;
assign addr[64058]= -917951481;
assign addr[64059]= -952379488;
assign addr[64060]= -986505429;
assign addr[64061]= -1020318481;
assign addr[64062]= -1053807919;
assign addr[64063]= -1086963121;
assign addr[64064]= -1119773573;
assign addr[64065]= -1152228866;
assign addr[64066]= -1184318708;
assign addr[64067]= -1216032921;
assign addr[64068]= -1247361445;
assign addr[64069]= -1278294345;
assign addr[64070]= -1308821808;
assign addr[64071]= -1338934154;
assign addr[64072]= -1368621831;
assign addr[64073]= -1397875423;
assign addr[64074]= -1426685652;
assign addr[64075]= -1455043381;
assign addr[64076]= -1482939614;
assign addr[64077]= -1510365504;
assign addr[64078]= -1537312353;
assign addr[64079]= -1563771613;
assign addr[64080]= -1589734894;
assign addr[64081]= -1615193959;
assign addr[64082]= -1640140734;
assign addr[64083]= -1664567307;
assign addr[64084]= -1688465931;
assign addr[64085]= -1711829025;
assign addr[64086]= -1734649179;
assign addr[64087]= -1756919156;
assign addr[64088]= -1778631892;
assign addr[64089]= -1799780501;
assign addr[64090]= -1820358275;
assign addr[64091]= -1840358687;
assign addr[64092]= -1859775393;
assign addr[64093]= -1878602237;
assign addr[64094]= -1896833245;
assign addr[64095]= -1914462636;
assign addr[64096]= -1931484818;
assign addr[64097]= -1947894393;
assign addr[64098]= -1963686155;
assign addr[64099]= -1978855097;
assign addr[64100]= -1993396407;
assign addr[64101]= -2007305472;
assign addr[64102]= -2020577882;
assign addr[64103]= -2033209426;
assign addr[64104]= -2045196100;
assign addr[64105]= -2056534099;
assign addr[64106]= -2067219829;
assign addr[64107]= -2077249901;
assign addr[64108]= -2086621133;
assign addr[64109]= -2095330553;
assign addr[64110]= -2103375398;
assign addr[64111]= -2110753117;
assign addr[64112]= -2117461370;
assign addr[64113]= -2123498030;
assign addr[64114]= -2128861181;
assign addr[64115]= -2133549123;
assign addr[64116]= -2137560369;
assign addr[64117]= -2140893646;
assign addr[64118]= -2143547897;
assign addr[64119]= -2145522281;
assign addr[64120]= -2146816171;
assign addr[64121]= -2147429158;
assign addr[64122]= -2147361045;
assign addr[64123]= -2146611856;
assign addr[64124]= -2145181827;
assign addr[64125]= -2143071413;
assign addr[64126]= -2140281282;
assign addr[64127]= -2136812319;
assign addr[64128]= -2132665626;
assign addr[64129]= -2127842516;
assign addr[64130]= -2122344521;
assign addr[64131]= -2116173382;
assign addr[64132]= -2109331059;
assign addr[64133]= -2101819720;
assign addr[64134]= -2093641749;
assign addr[64135]= -2084799740;
assign addr[64136]= -2075296495;
assign addr[64137]= -2065135031;
assign addr[64138]= -2054318569;
assign addr[64139]= -2042850540;
assign addr[64140]= -2030734582;
assign addr[64141]= -2017974537;
assign addr[64142]= -2004574453;
assign addr[64143]= -1990538579;
assign addr[64144]= -1975871368;
assign addr[64145]= -1960577471;
assign addr[64146]= -1944661739;
assign addr[64147]= -1928129220;
assign addr[64148]= -1910985158;
assign addr[64149]= -1893234990;
assign addr[64150]= -1874884346;
assign addr[64151]= -1855939047;
assign addr[64152]= -1836405100;
assign addr[64153]= -1816288703;
assign addr[64154]= -1795596234;
assign addr[64155]= -1774334257;
assign addr[64156]= -1752509516;
assign addr[64157]= -1730128933;
assign addr[64158]= -1707199606;
assign addr[64159]= -1683728808;
assign addr[64160]= -1659723983;
assign addr[64161]= -1635192744;
assign addr[64162]= -1610142873;
assign addr[64163]= -1584582314;
assign addr[64164]= -1558519173;
assign addr[64165]= -1531961719;
assign addr[64166]= -1504918373;
assign addr[64167]= -1477397714;
assign addr[64168]= -1449408469;
assign addr[64169]= -1420959516;
assign addr[64170]= -1392059879;
assign addr[64171]= -1362718723;
assign addr[64172]= -1332945355;
assign addr[64173]= -1302749217;
assign addr[64174]= -1272139887;
assign addr[64175]= -1241127074;
assign addr[64176]= -1209720613;
assign addr[64177]= -1177930466;
assign addr[64178]= -1145766716;
assign addr[64179]= -1113239564;
assign addr[64180]= -1080359326;
assign addr[64181]= -1047136432;
assign addr[64182]= -1013581418;
assign addr[64183]= -979704927;
assign addr[64184]= -945517704;
assign addr[64185]= -911030591;
assign addr[64186]= -876254528;
assign addr[64187]= -841200544;
assign addr[64188]= -805879757;
assign addr[64189]= -770303369;
assign addr[64190]= -734482665;
assign addr[64191]= -698429006;
assign addr[64192]= -662153826;
assign addr[64193]= -625668632;
assign addr[64194]= -588984994;
assign addr[64195]= -552114549;
assign addr[64196]= -515068990;
assign addr[64197]= -477860067;
assign addr[64198]= -440499581;
assign addr[64199]= -402999383;
assign addr[64200]= -365371365;
assign addr[64201]= -327627463;
assign addr[64202]= -289779648;
assign addr[64203]= -251839923;
assign addr[64204]= -213820322;
assign addr[64205]= -175732905;
assign addr[64206]= -137589750;
assign addr[64207]= -99402956;
assign addr[64208]= -61184634;
assign addr[64209]= -22946906;
assign addr[64210]= 15298099;
assign addr[64211]= 53538253;
assign addr[64212]= 91761426;
assign addr[64213]= 129955495;
assign addr[64214]= 168108346;
assign addr[64215]= 206207878;
assign addr[64216]= 244242007;
assign addr[64217]= 282198671;
assign addr[64218]= 320065829;
assign addr[64219]= 357831473;
assign addr[64220]= 395483624;
assign addr[64221]= 433010339;
assign addr[64222]= 470399716;
assign addr[64223]= 507639898;
assign addr[64224]= 544719071;
assign addr[64225]= 581625477;
assign addr[64226]= 618347408;
assign addr[64227]= 654873219;
assign addr[64228]= 691191324;
assign addr[64229]= 727290205;
assign addr[64230]= 763158411;
assign addr[64231]= 798784567;
assign addr[64232]= 834157373;
assign addr[64233]= 869265610;
assign addr[64234]= 904098143;
assign addr[64235]= 938643924;
assign addr[64236]= 972891995;
assign addr[64237]= 1006831495;
assign addr[64238]= 1040451659;
assign addr[64239]= 1073741824;
assign addr[64240]= 1106691431;
assign addr[64241]= 1139290029;
assign addr[64242]= 1171527280;
assign addr[64243]= 1203392958;
assign addr[64244]= 1234876957;
assign addr[64245]= 1265969291;
assign addr[64246]= 1296660098;
assign addr[64247]= 1326939644;
assign addr[64248]= 1356798326;
assign addr[64249]= 1386226674;
assign addr[64250]= 1415215352;
assign addr[64251]= 1443755168;
assign addr[64252]= 1471837070;
assign addr[64253]= 1499452149;
assign addr[64254]= 1526591649;
assign addr[64255]= 1553246960;
assign addr[64256]= 1579409630;
assign addr[64257]= 1605071359;
assign addr[64258]= 1630224009;
assign addr[64259]= 1654859602;
assign addr[64260]= 1678970324;
assign addr[64261]= 1702548529;
assign addr[64262]= 1725586737;
assign addr[64263]= 1748077642;
assign addr[64264]= 1770014111;
assign addr[64265]= 1791389186;
assign addr[64266]= 1812196087;
assign addr[64267]= 1832428215;
assign addr[64268]= 1852079154;
assign addr[64269]= 1871142669;
assign addr[64270]= 1889612716;
assign addr[64271]= 1907483436;
assign addr[64272]= 1924749160;
assign addr[64273]= 1941404413;
assign addr[64274]= 1957443913;
assign addr[64275]= 1972862571;
assign addr[64276]= 1987655498;
assign addr[64277]= 2001818002;
assign addr[64278]= 2015345591;
assign addr[64279]= 2028233973;
assign addr[64280]= 2040479063;
assign addr[64281]= 2052076975;
assign addr[64282]= 2063024031;
assign addr[64283]= 2073316760;
assign addr[64284]= 2082951896;
assign addr[64285]= 2091926384;
assign addr[64286]= 2100237377;
assign addr[64287]= 2107882239;
assign addr[64288]= 2114858546;
assign addr[64289]= 2121164085;
assign addr[64290]= 2126796855;
assign addr[64291]= 2131755071;
assign addr[64292]= 2136037160;
assign addr[64293]= 2139641764;
assign addr[64294]= 2142567738;
assign addr[64295]= 2144814157;
assign addr[64296]= 2146380306;
assign addr[64297]= 2147265689;
assign addr[64298]= 2147470025;
assign addr[64299]= 2146993250;
assign addr[64300]= 2145835515;
assign addr[64301]= 2143997187;
assign addr[64302]= 2141478848;
assign addr[64303]= 2138281298;
assign addr[64304]= 2134405552;
assign addr[64305]= 2129852837;
assign addr[64306]= 2124624598;
assign addr[64307]= 2118722494;
assign addr[64308]= 2112148396;
assign addr[64309]= 2104904390;
assign addr[64310]= 2096992772;
assign addr[64311]= 2088416053;
assign addr[64312]= 2079176953;
assign addr[64313]= 2069278401;
assign addr[64314]= 2058723538;
assign addr[64315]= 2047515711;
assign addr[64316]= 2035658475;
assign addr[64317]= 2023155591;
assign addr[64318]= 2010011024;
assign addr[64319]= 1996228943;
assign addr[64320]= 1981813720;
assign addr[64321]= 1966769926;
assign addr[64322]= 1951102334;
assign addr[64323]= 1934815911;
assign addr[64324]= 1917915825;
assign addr[64325]= 1900407434;
assign addr[64326]= 1882296293;
assign addr[64327]= 1863588145;
assign addr[64328]= 1844288924;
assign addr[64329]= 1824404752;
assign addr[64330]= 1803941934;
assign addr[64331]= 1782906961;
assign addr[64332]= 1761306505;
assign addr[64333]= 1739147417;
assign addr[64334]= 1716436725;
assign addr[64335]= 1693181631;
assign addr[64336]= 1669389513;
assign addr[64337]= 1645067915;
assign addr[64338]= 1620224553;
assign addr[64339]= 1594867305;
assign addr[64340]= 1569004214;
assign addr[64341]= 1542643483;
assign addr[64342]= 1515793473;
assign addr[64343]= 1488462700;
assign addr[64344]= 1460659832;
assign addr[64345]= 1432393688;
assign addr[64346]= 1403673233;
assign addr[64347]= 1374507575;
assign addr[64348]= 1344905966;
assign addr[64349]= 1314877795;
assign addr[64350]= 1284432584;
assign addr[64351]= 1253579991;
assign addr[64352]= 1222329801;
assign addr[64353]= 1190691925;
assign addr[64354]= 1158676398;
assign addr[64355]= 1126293375;
assign addr[64356]= 1093553126;
assign addr[64357]= 1060466036;
assign addr[64358]= 1027042599;
assign addr[64359]= 993293415;
assign addr[64360]= 959229189;
assign addr[64361]= 924860725;
assign addr[64362]= 890198924;
assign addr[64363]= 855254778;
assign addr[64364]= 820039373;
assign addr[64365]= 784563876;
assign addr[64366]= 748839539;
assign addr[64367]= 712877694;
assign addr[64368]= 676689746;
assign addr[64369]= 640287172;
assign addr[64370]= 603681519;
assign addr[64371]= 566884397;
assign addr[64372]= 529907477;
assign addr[64373]= 492762486;
assign addr[64374]= 455461206;
assign addr[64375]= 418015468;
assign addr[64376]= 380437148;
assign addr[64377]= 342738165;
assign addr[64378]= 304930476;
assign addr[64379]= 267026072;
assign addr[64380]= 229036977;
assign addr[64381]= 190975237;
assign addr[64382]= 152852926;
assign addr[64383]= 114682135;
assign addr[64384]= 76474970;
assign addr[64385]= 38243550;
assign addr[64386]= 0;
assign addr[64387]= -38243550;
assign addr[64388]= -76474970;
assign addr[64389]= -114682135;
assign addr[64390]= -152852926;
assign addr[64391]= -190975237;
assign addr[64392]= -229036977;
assign addr[64393]= -267026072;
assign addr[64394]= -304930476;
assign addr[64395]= -342738165;
assign addr[64396]= -380437148;
assign addr[64397]= -418015468;
assign addr[64398]= -455461206;
assign addr[64399]= -492762486;
assign addr[64400]= -529907477;
assign addr[64401]= -566884397;
assign addr[64402]= -603681519;
assign addr[64403]= -640287172;
assign addr[64404]= -676689746;
assign addr[64405]= -712877694;
assign addr[64406]= -748839539;
assign addr[64407]= -784563876;
assign addr[64408]= -820039373;
assign addr[64409]= -855254778;
assign addr[64410]= -890198924;
assign addr[64411]= -924860725;
assign addr[64412]= -959229189;
assign addr[64413]= -993293415;
assign addr[64414]= -1027042599;
assign addr[64415]= -1060466036;
assign addr[64416]= -1093553126;
assign addr[64417]= -1126293375;
assign addr[64418]= -1158676398;
assign addr[64419]= -1190691925;
assign addr[64420]= -1222329801;
assign addr[64421]= -1253579991;
assign addr[64422]= -1284432584;
assign addr[64423]= -1314877795;
assign addr[64424]= -1344905966;
assign addr[64425]= -1374507575;
assign addr[64426]= -1403673233;
assign addr[64427]= -1432393688;
assign addr[64428]= -1460659832;
assign addr[64429]= -1488462700;
assign addr[64430]= -1515793473;
assign addr[64431]= -1542643483;
assign addr[64432]= -1569004214;
assign addr[64433]= -1594867305;
assign addr[64434]= -1620224553;
assign addr[64435]= -1645067915;
assign addr[64436]= -1669389513;
assign addr[64437]= -1693181631;
assign addr[64438]= -1716436725;
assign addr[64439]= -1739147417;
assign addr[64440]= -1761306505;
assign addr[64441]= -1782906961;
assign addr[64442]= -1803941934;
assign addr[64443]= -1824404752;
assign addr[64444]= -1844288924;
assign addr[64445]= -1863588145;
assign addr[64446]= -1882296293;
assign addr[64447]= -1900407434;
assign addr[64448]= -1917915825;
assign addr[64449]= -1934815911;
assign addr[64450]= -1951102334;
assign addr[64451]= -1966769926;
assign addr[64452]= -1981813720;
assign addr[64453]= -1996228943;
assign addr[64454]= -2010011024;
assign addr[64455]= -2023155591;
assign addr[64456]= -2035658475;
assign addr[64457]= -2047515711;
assign addr[64458]= -2058723538;
assign addr[64459]= -2069278401;
assign addr[64460]= -2079176953;
assign addr[64461]= -2088416053;
assign addr[64462]= -2096992772;
assign addr[64463]= -2104904390;
assign addr[64464]= -2112148396;
assign addr[64465]= -2118722494;
assign addr[64466]= -2124624598;
assign addr[64467]= -2129852837;
assign addr[64468]= -2134405552;
assign addr[64469]= -2138281298;
assign addr[64470]= -2141478848;
assign addr[64471]= -2143997187;
assign addr[64472]= -2145835515;
assign addr[64473]= -2146993250;
assign addr[64474]= -2147470025;
assign addr[64475]= -2147265689;
assign addr[64476]= -2146380306;
assign addr[64477]= -2144814157;
assign addr[64478]= -2142567738;
assign addr[64479]= -2139641764;
assign addr[64480]= -2136037160;
assign addr[64481]= -2131755071;
assign addr[64482]= -2126796855;
assign addr[64483]= -2121164085;
assign addr[64484]= -2114858546;
assign addr[64485]= -2107882239;
assign addr[64486]= -2100237377;
assign addr[64487]= -2091926384;
assign addr[64488]= -2082951896;
assign addr[64489]= -2073316760;
assign addr[64490]= -2063024031;
assign addr[64491]= -2052076975;
assign addr[64492]= -2040479063;
assign addr[64493]= -2028233973;
assign addr[64494]= -2015345591;
assign addr[64495]= -2001818002;
assign addr[64496]= -1987655498;
assign addr[64497]= -1972862571;
assign addr[64498]= -1957443913;
assign addr[64499]= -1941404413;
assign addr[64500]= -1924749160;
assign addr[64501]= -1907483436;
assign addr[64502]= -1889612716;
assign addr[64503]= -1871142669;
assign addr[64504]= -1852079154;
assign addr[64505]= -1832428215;
assign addr[64506]= -1812196087;
assign addr[64507]= -1791389186;
assign addr[64508]= -1770014111;
assign addr[64509]= -1748077642;
assign addr[64510]= -1725586737;
assign addr[64511]= -1702548529;
assign addr[64512]= -1678970324;
assign addr[64513]= -1654859602;
assign addr[64514]= -1630224009;
assign addr[64515]= -1605071359;
assign addr[64516]= -1579409630;
assign addr[64517]= -1553246960;
assign addr[64518]= -1526591649;
assign addr[64519]= -1499452149;
assign addr[64520]= -1471837070;
assign addr[64521]= -1443755168;
assign addr[64522]= -1415215352;
assign addr[64523]= -1386226674;
assign addr[64524]= -1356798326;
assign addr[64525]= -1326939644;
assign addr[64526]= -1296660098;
assign addr[64527]= -1265969291;
assign addr[64528]= -1234876957;
assign addr[64529]= -1203392958;
assign addr[64530]= -1171527280;
assign addr[64531]= -1139290029;
assign addr[64532]= -1106691431;
assign addr[64533]= -1073741824;
assign addr[64534]= -1040451659;
assign addr[64535]= -1006831495;
assign addr[64536]= -972891995;
assign addr[64537]= -938643924;
assign addr[64538]= -904098143;
assign addr[64539]= -869265610;
assign addr[64540]= -834157373;
assign addr[64541]= -798784567;
assign addr[64542]= -763158411;
assign addr[64543]= -727290205;
assign addr[64544]= -691191324;
assign addr[64545]= -654873219;
assign addr[64546]= -618347408;
assign addr[64547]= -581625477;
assign addr[64548]= -544719071;
assign addr[64549]= -507639898;
assign addr[64550]= -470399716;
assign addr[64551]= -433010339;
assign addr[64552]= -395483624;
assign addr[64553]= -357831473;
assign addr[64554]= -320065829;
assign addr[64555]= -282198671;
assign addr[64556]= -244242007;
assign addr[64557]= -206207878;
assign addr[64558]= -168108346;
assign addr[64559]= -129955495;
assign addr[64560]= -91761426;
assign addr[64561]= -53538253;
assign addr[64562]= -15298099;
assign addr[64563]= 22946906;
assign addr[64564]= 61184634;
assign addr[64565]= 99402956;
assign addr[64566]= 137589750;
assign addr[64567]= 175732905;
assign addr[64568]= 213820322;
assign addr[64569]= 251839923;
assign addr[64570]= 289779648;
assign addr[64571]= 327627463;
assign addr[64572]= 365371365;
assign addr[64573]= 402999383;
assign addr[64574]= 440499581;
assign addr[64575]= 477860067;
assign addr[64576]= 515068990;
assign addr[64577]= 552114549;
assign addr[64578]= 588984994;
assign addr[64579]= 625668632;
assign addr[64580]= 662153826;
assign addr[64581]= 698429006;
assign addr[64582]= 734482665;
assign addr[64583]= 770303369;
assign addr[64584]= 805879757;
assign addr[64585]= 841200544;
assign addr[64586]= 876254528;
assign addr[64587]= 911030591;
assign addr[64588]= 945517704;
assign addr[64589]= 979704927;
assign addr[64590]= 1013581418;
assign addr[64591]= 1047136432;
assign addr[64592]= 1080359326;
assign addr[64593]= 1113239564;
assign addr[64594]= 1145766716;
assign addr[64595]= 1177930466;
assign addr[64596]= 1209720613;
assign addr[64597]= 1241127074;
assign addr[64598]= 1272139887;
assign addr[64599]= 1302749217;
assign addr[64600]= 1332945355;
assign addr[64601]= 1362718723;
assign addr[64602]= 1392059879;
assign addr[64603]= 1420959516;
assign addr[64604]= 1449408469;
assign addr[64605]= 1477397714;
assign addr[64606]= 1504918373;
assign addr[64607]= 1531961719;
assign addr[64608]= 1558519173;
assign addr[64609]= 1584582314;
assign addr[64610]= 1610142873;
assign addr[64611]= 1635192744;
assign addr[64612]= 1659723983;
assign addr[64613]= 1683728808;
assign addr[64614]= 1707199606;
assign addr[64615]= 1730128933;
assign addr[64616]= 1752509516;
assign addr[64617]= 1774334257;
assign addr[64618]= 1795596234;
assign addr[64619]= 1816288703;
assign addr[64620]= 1836405100;
assign addr[64621]= 1855939047;
assign addr[64622]= 1874884346;
assign addr[64623]= 1893234990;
assign addr[64624]= 1910985158;
assign addr[64625]= 1928129220;
assign addr[64626]= 1944661739;
assign addr[64627]= 1960577471;
assign addr[64628]= 1975871368;
assign addr[64629]= 1990538579;
assign addr[64630]= 2004574453;
assign addr[64631]= 2017974537;
assign addr[64632]= 2030734582;
assign addr[64633]= 2042850540;
assign addr[64634]= 2054318569;
assign addr[64635]= 2065135031;
assign addr[64636]= 2075296495;
assign addr[64637]= 2084799740;
assign addr[64638]= 2093641749;
assign addr[64639]= 2101819720;
assign addr[64640]= 2109331059;
assign addr[64641]= 2116173382;
assign addr[64642]= 2122344521;
assign addr[64643]= 2127842516;
assign addr[64644]= 2132665626;
assign addr[64645]= 2136812319;
assign addr[64646]= 2140281282;
assign addr[64647]= 2143071413;
assign addr[64648]= 2145181827;
assign addr[64649]= 2146611856;
assign addr[64650]= 2147361045;
assign addr[64651]= 2147429158;
assign addr[64652]= 2146816171;
assign addr[64653]= 2145522281;
assign addr[64654]= 2143547897;
assign addr[64655]= 2140893646;
assign addr[64656]= 2137560369;
assign addr[64657]= 2133549123;
assign addr[64658]= 2128861181;
assign addr[64659]= 2123498030;
assign addr[64660]= 2117461370;
assign addr[64661]= 2110753117;
assign addr[64662]= 2103375398;
assign addr[64663]= 2095330553;
assign addr[64664]= 2086621133;
assign addr[64665]= 2077249901;
assign addr[64666]= 2067219829;
assign addr[64667]= 2056534099;
assign addr[64668]= 2045196100;
assign addr[64669]= 2033209426;
assign addr[64670]= 2020577882;
assign addr[64671]= 2007305472;
assign addr[64672]= 1993396407;
assign addr[64673]= 1978855097;
assign addr[64674]= 1963686155;
assign addr[64675]= 1947894393;
assign addr[64676]= 1931484818;
assign addr[64677]= 1914462636;
assign addr[64678]= 1896833245;
assign addr[64679]= 1878602237;
assign addr[64680]= 1859775393;
assign addr[64681]= 1840358687;
assign addr[64682]= 1820358275;
assign addr[64683]= 1799780501;
assign addr[64684]= 1778631892;
assign addr[64685]= 1756919156;
assign addr[64686]= 1734649179;
assign addr[64687]= 1711829025;
assign addr[64688]= 1688465931;
assign addr[64689]= 1664567307;
assign addr[64690]= 1640140734;
assign addr[64691]= 1615193959;
assign addr[64692]= 1589734894;
assign addr[64693]= 1563771613;
assign addr[64694]= 1537312353;
assign addr[64695]= 1510365504;
assign addr[64696]= 1482939614;
assign addr[64697]= 1455043381;
assign addr[64698]= 1426685652;
assign addr[64699]= 1397875423;
assign addr[64700]= 1368621831;
assign addr[64701]= 1338934154;
assign addr[64702]= 1308821808;
assign addr[64703]= 1278294345;
assign addr[64704]= 1247361445;
assign addr[64705]= 1216032921;
assign addr[64706]= 1184318708;
assign addr[64707]= 1152228866;
assign addr[64708]= 1119773573;
assign addr[64709]= 1086963121;
assign addr[64710]= 1053807919;
assign addr[64711]= 1020318481;
assign addr[64712]= 986505429;
assign addr[64713]= 952379488;
assign addr[64714]= 917951481;
assign addr[64715]= 883232329;
assign addr[64716]= 848233042;
assign addr[64717]= 812964722;
assign addr[64718]= 777438554;
assign addr[64719]= 741665807;
assign addr[64720]= 705657826;
assign addr[64721]= 669426032;
assign addr[64722]= 632981917;
assign addr[64723]= 596337040;
assign addr[64724]= 559503022;
assign addr[64725]= 522491548;
assign addr[64726]= 485314355;
assign addr[64727]= 447983235;
assign addr[64728]= 410510029;
assign addr[64729]= 372906622;
assign addr[64730]= 335184940;
assign addr[64731]= 297356948;
assign addr[64732]= 259434643;
assign addr[64733]= 221430054;
assign addr[64734]= 183355234;
assign addr[64735]= 145222259;
assign addr[64736]= 107043224;
assign addr[64737]= 68830239;
assign addr[64738]= 30595422;
assign addr[64739]= -7649098;
assign addr[64740]= -45891193;
assign addr[64741]= -84118732;
assign addr[64742]= -122319591;
assign addr[64743]= -160481654;
assign addr[64744]= -198592817;
assign addr[64745]= -236640993;
assign addr[64746]= -274614114;
assign addr[64747]= -312500135;
assign addr[64748]= -350287041;
assign addr[64749]= -387962847;
assign addr[64750]= -425515602;
assign addr[64751]= -462933398;
assign addr[64752]= -500204365;
assign addr[64753]= -537316682;
assign addr[64754]= -574258580;
assign addr[64755]= -611018340;
assign addr[64756]= -647584304;
assign addr[64757]= -683944874;
assign addr[64758]= -720088517;
assign addr[64759]= -756003771;
assign addr[64760]= -791679244;
assign addr[64761]= -827103620;
assign addr[64762]= -862265664;
assign addr[64763]= -897154224;
assign addr[64764]= -931758235;
assign addr[64765]= -966066720;
assign addr[64766]= -1000068799;
assign addr[64767]= -1033753687;
assign addr[64768]= -1067110699;
assign addr[64769]= -1100129257;
assign addr[64770]= -1132798888;
assign addr[64771]= -1165109230;
assign addr[64772]= -1197050035;
assign addr[64773]= -1228611172;
assign addr[64774]= -1259782632;
assign addr[64775]= -1290554528;
assign addr[64776]= -1320917099;
assign addr[64777]= -1350860716;
assign addr[64778]= -1380375881;
assign addr[64779]= -1409453233;
assign addr[64780]= -1438083551;
assign addr[64781]= -1466257752;
assign addr[64782]= -1493966902;
assign addr[64783]= -1521202211;
assign addr[64784]= -1547955041;
assign addr[64785]= -1574216908;
assign addr[64786]= -1599979481;
assign addr[64787]= -1625234591;
assign addr[64788]= -1649974225;
assign addr[64789]= -1674190539;
assign addr[64790]= -1697875851;
assign addr[64791]= -1721022648;
assign addr[64792]= -1743623590;
assign addr[64793]= -1765671509;
assign addr[64794]= -1787159411;
assign addr[64795]= -1808080480;
assign addr[64796]= -1828428082;
assign addr[64797]= -1848195763;
assign addr[64798]= -1867377253;
assign addr[64799]= -1885966468;
assign addr[64800]= -1903957513;
assign addr[64801]= -1921344681;
assign addr[64802]= -1938122457;
assign addr[64803]= -1954285520;
assign addr[64804]= -1969828744;
assign addr[64805]= -1984747199;
assign addr[64806]= -1999036154;
assign addr[64807]= -2012691075;
assign addr[64808]= -2025707632;
assign addr[64809]= -2038081698;
assign addr[64810]= -2049809346;
assign addr[64811]= -2060886858;
assign addr[64812]= -2071310720;
assign addr[64813]= -2081077626;
assign addr[64814]= -2090184478;
assign addr[64815]= -2098628387;
assign addr[64816]= -2106406677;
assign addr[64817]= -2113516878;
assign addr[64818]= -2119956737;
assign addr[64819]= -2125724211;
assign addr[64820]= -2130817471;
assign addr[64821]= -2135234901;
assign addr[64822]= -2138975100;
assign addr[64823]= -2142036881;
assign addr[64824]= -2144419275;
assign addr[64825]= -2146121524;
assign addr[64826]= -2147143090;
assign addr[64827]= -2147483648;
assign addr[64828]= -2147143090;
assign addr[64829]= -2146121524;
assign addr[64830]= -2144419275;
assign addr[64831]= -2142036881;
assign addr[64832]= -2138975100;
assign addr[64833]= -2135234901;
assign addr[64834]= -2130817471;
assign addr[64835]= -2125724211;
assign addr[64836]= -2119956737;
assign addr[64837]= -2113516878;
assign addr[64838]= -2106406677;
assign addr[64839]= -2098628387;
assign addr[64840]= -2090184478;
assign addr[64841]= -2081077626;
assign addr[64842]= -2071310720;
assign addr[64843]= -2060886858;
assign addr[64844]= -2049809346;
assign addr[64845]= -2038081698;
assign addr[64846]= -2025707632;
assign addr[64847]= -2012691075;
assign addr[64848]= -1999036154;
assign addr[64849]= -1984747199;
assign addr[64850]= -1969828744;
assign addr[64851]= -1954285520;
assign addr[64852]= -1938122457;
assign addr[64853]= -1921344681;
assign addr[64854]= -1903957513;
assign addr[64855]= -1885966468;
assign addr[64856]= -1867377253;
assign addr[64857]= -1848195763;
assign addr[64858]= -1828428082;
assign addr[64859]= -1808080480;
assign addr[64860]= -1787159411;
assign addr[64861]= -1765671509;
assign addr[64862]= -1743623590;
assign addr[64863]= -1721022648;
assign addr[64864]= -1697875851;
assign addr[64865]= -1674190539;
assign addr[64866]= -1649974225;
assign addr[64867]= -1625234591;
assign addr[64868]= -1599979481;
assign addr[64869]= -1574216908;
assign addr[64870]= -1547955041;
assign addr[64871]= -1521202211;
assign addr[64872]= -1493966902;
assign addr[64873]= -1466257752;
assign addr[64874]= -1438083551;
assign addr[64875]= -1409453233;
assign addr[64876]= -1380375881;
assign addr[64877]= -1350860716;
assign addr[64878]= -1320917099;
assign addr[64879]= -1290554528;
assign addr[64880]= -1259782632;
assign addr[64881]= -1228611172;
assign addr[64882]= -1197050035;
assign addr[64883]= -1165109230;
assign addr[64884]= -1132798888;
assign addr[64885]= -1100129257;
assign addr[64886]= -1067110699;
assign addr[64887]= -1033753687;
assign addr[64888]= -1000068799;
assign addr[64889]= -966066720;
assign addr[64890]= -931758235;
assign addr[64891]= -897154224;
assign addr[64892]= -862265664;
assign addr[64893]= -827103620;
assign addr[64894]= -791679244;
assign addr[64895]= -756003771;
assign addr[64896]= -720088517;
assign addr[64897]= -683944874;
assign addr[64898]= -647584304;
assign addr[64899]= -611018340;
assign addr[64900]= -574258580;
assign addr[64901]= -537316682;
assign addr[64902]= -500204365;
assign addr[64903]= -462933398;
assign addr[64904]= -425515602;
assign addr[64905]= -387962847;
assign addr[64906]= -350287041;
assign addr[64907]= -312500135;
assign addr[64908]= -274614114;
assign addr[64909]= -236640993;
assign addr[64910]= -198592817;
assign addr[64911]= -160481654;
assign addr[64912]= -122319591;
assign addr[64913]= -84118732;
assign addr[64914]= -45891193;
assign addr[64915]= -7649098;
assign addr[64916]= 30595422;
assign addr[64917]= 68830239;
assign addr[64918]= 107043224;
assign addr[64919]= 145222259;
assign addr[64920]= 183355234;
assign addr[64921]= 221430054;
assign addr[64922]= 259434643;
assign addr[64923]= 297356948;
assign addr[64924]= 335184940;
assign addr[64925]= 372906622;
assign addr[64926]= 410510029;
assign addr[64927]= 447983235;
assign addr[64928]= 485314355;
assign addr[64929]= 522491548;
assign addr[64930]= 559503022;
assign addr[64931]= 596337040;
assign addr[64932]= 632981917;
assign addr[64933]= 669426032;
assign addr[64934]= 705657826;
assign addr[64935]= 741665807;
assign addr[64936]= 777438554;
assign addr[64937]= 812964722;
assign addr[64938]= 848233042;
assign addr[64939]= 883232329;
assign addr[64940]= 917951481;
assign addr[64941]= 952379488;
assign addr[64942]= 986505429;
assign addr[64943]= 1020318481;
assign addr[64944]= 1053807919;
assign addr[64945]= 1086963121;
assign addr[64946]= 1119773573;
assign addr[64947]= 1152228866;
assign addr[64948]= 1184318708;
assign addr[64949]= 1216032921;
assign addr[64950]= 1247361445;
assign addr[64951]= 1278294345;
assign addr[64952]= 1308821808;
assign addr[64953]= 1338934154;
assign addr[64954]= 1368621831;
assign addr[64955]= 1397875423;
assign addr[64956]= 1426685652;
assign addr[64957]= 1455043381;
assign addr[64958]= 1482939614;
assign addr[64959]= 1510365504;
assign addr[64960]= 1537312353;
assign addr[64961]= 1563771613;
assign addr[64962]= 1589734894;
assign addr[64963]= 1615193959;
assign addr[64964]= 1640140734;
assign addr[64965]= 1664567307;
assign addr[64966]= 1688465931;
assign addr[64967]= 1711829025;
assign addr[64968]= 1734649179;
assign addr[64969]= 1756919156;
assign addr[64970]= 1778631892;
assign addr[64971]= 1799780501;
assign addr[64972]= 1820358275;
assign addr[64973]= 1840358687;
assign addr[64974]= 1859775393;
assign addr[64975]= 1878602237;
assign addr[64976]= 1896833245;
assign addr[64977]= 1914462636;
assign addr[64978]= 1931484818;
assign addr[64979]= 1947894393;
assign addr[64980]= 1963686155;
assign addr[64981]= 1978855097;
assign addr[64982]= 1993396407;
assign addr[64983]= 2007305472;
assign addr[64984]= 2020577882;
assign addr[64985]= 2033209426;
assign addr[64986]= 2045196100;
assign addr[64987]= 2056534099;
assign addr[64988]= 2067219829;
assign addr[64989]= 2077249901;
assign addr[64990]= 2086621133;
assign addr[64991]= 2095330553;
assign addr[64992]= 2103375398;
assign addr[64993]= 2110753117;
assign addr[64994]= 2117461370;
assign addr[64995]= 2123498030;
assign addr[64996]= 2128861181;
assign addr[64997]= 2133549123;
assign addr[64998]= 2137560369;
assign addr[64999]= 2140893646;
assign addr[65000]= 2143547897;
assign addr[65001]= 2145522281;
assign addr[65002]= 2146816171;
assign addr[65003]= 2147429158;
assign addr[65004]= 2147361045;
assign addr[65005]= 2146611856;
assign addr[65006]= 2145181827;
assign addr[65007]= 2143071413;
assign addr[65008]= 2140281282;
assign addr[65009]= 2136812319;
assign addr[65010]= 2132665626;
assign addr[65011]= 2127842516;
assign addr[65012]= 2122344521;
assign addr[65013]= 2116173382;
assign addr[65014]= 2109331059;
assign addr[65015]= 2101819720;
assign addr[65016]= 2093641749;
assign addr[65017]= 2084799740;
assign addr[65018]= 2075296495;
assign addr[65019]= 2065135031;
assign addr[65020]= 2054318569;
assign addr[65021]= 2042850540;
assign addr[65022]= 2030734582;
assign addr[65023]= 2017974537;
assign addr[65024]= 2004574453;
assign addr[65025]= 1990538579;
assign addr[65026]= 1975871368;
assign addr[65027]= 1960577471;
assign addr[65028]= 1944661739;
assign addr[65029]= 1928129220;
assign addr[65030]= 1910985158;
assign addr[65031]= 1893234990;
assign addr[65032]= 1874884346;
assign addr[65033]= 1855939047;
assign addr[65034]= 1836405100;
assign addr[65035]= 1816288703;
assign addr[65036]= 1795596234;
assign addr[65037]= 1774334257;
assign addr[65038]= 1752509516;
assign addr[65039]= 1730128933;
assign addr[65040]= 1707199606;
assign addr[65041]= 1683728808;
assign addr[65042]= 1659723983;
assign addr[65043]= 1635192744;
assign addr[65044]= 1610142873;
assign addr[65045]= 1584582314;
assign addr[65046]= 1558519173;
assign addr[65047]= 1531961719;
assign addr[65048]= 1504918373;
assign addr[65049]= 1477397714;
assign addr[65050]= 1449408469;
assign addr[65051]= 1420959516;
assign addr[65052]= 1392059879;
assign addr[65053]= 1362718723;
assign addr[65054]= 1332945355;
assign addr[65055]= 1302749217;
assign addr[65056]= 1272139887;
assign addr[65057]= 1241127074;
assign addr[65058]= 1209720613;
assign addr[65059]= 1177930466;
assign addr[65060]= 1145766716;
assign addr[65061]= 1113239564;
assign addr[65062]= 1080359326;
assign addr[65063]= 1047136432;
assign addr[65064]= 1013581418;
assign addr[65065]= 979704927;
assign addr[65066]= 945517704;
assign addr[65067]= 911030591;
assign addr[65068]= 876254528;
assign addr[65069]= 841200544;
assign addr[65070]= 805879757;
assign addr[65071]= 770303369;
assign addr[65072]= 734482665;
assign addr[65073]= 698429006;
assign addr[65074]= 662153826;
assign addr[65075]= 625668632;
assign addr[65076]= 588984994;
assign addr[65077]= 552114549;
assign addr[65078]= 515068990;
assign addr[65079]= 477860067;
assign addr[65080]= 440499581;
assign addr[65081]= 402999383;
assign addr[65082]= 365371365;
assign addr[65083]= 327627463;
assign addr[65084]= 289779648;
assign addr[65085]= 251839923;
assign addr[65086]= 213820322;
assign addr[65087]= 175732905;
assign addr[65088]= 137589750;
assign addr[65089]= 99402956;
assign addr[65090]= 61184634;
assign addr[65091]= 22946906;
assign addr[65092]= -15298099;
assign addr[65093]= -53538253;
assign addr[65094]= -91761426;
assign addr[65095]= -129955495;
assign addr[65096]= -168108346;
assign addr[65097]= -206207878;
assign addr[65098]= -244242007;
assign addr[65099]= -282198671;
assign addr[65100]= -320065829;
assign addr[65101]= -357831473;
assign addr[65102]= -395483624;
assign addr[65103]= -433010339;
assign addr[65104]= -470399716;
assign addr[65105]= -507639898;
assign addr[65106]= -544719071;
assign addr[65107]= -581625477;
assign addr[65108]= -618347408;
assign addr[65109]= -654873219;
assign addr[65110]= -691191324;
assign addr[65111]= -727290205;
assign addr[65112]= -763158411;
assign addr[65113]= -798784567;
assign addr[65114]= -834157373;
assign addr[65115]= -869265610;
assign addr[65116]= -904098143;
assign addr[65117]= -938643924;
assign addr[65118]= -972891995;
assign addr[65119]= -1006831495;
assign addr[65120]= -1040451659;
assign addr[65121]= -1073741824;
assign addr[65122]= -1106691431;
assign addr[65123]= -1139290029;
assign addr[65124]= -1171527280;
assign addr[65125]= -1203392958;
assign addr[65126]= -1234876957;
assign addr[65127]= -1265969291;
assign addr[65128]= -1296660098;
assign addr[65129]= -1326939644;
assign addr[65130]= -1356798326;
assign addr[65131]= -1386226674;
assign addr[65132]= -1415215352;
assign addr[65133]= -1443755168;
assign addr[65134]= -1471837070;
assign addr[65135]= -1499452149;
assign addr[65136]= -1526591649;
assign addr[65137]= -1553246960;
assign addr[65138]= -1579409630;
assign addr[65139]= -1605071359;
assign addr[65140]= -1630224009;
assign addr[65141]= -1654859602;
assign addr[65142]= -1678970324;
assign addr[65143]= -1702548529;
assign addr[65144]= -1725586737;
assign addr[65145]= -1748077642;
assign addr[65146]= -1770014111;
assign addr[65147]= -1791389186;
assign addr[65148]= -1812196087;
assign addr[65149]= -1832428215;
assign addr[65150]= -1852079154;
assign addr[65151]= -1871142669;
assign addr[65152]= -1889612716;
assign addr[65153]= -1907483436;
assign addr[65154]= -1924749160;
assign addr[65155]= -1941404413;
assign addr[65156]= -1957443913;
assign addr[65157]= -1972862571;
assign addr[65158]= -1987655498;
assign addr[65159]= -2001818002;
assign addr[65160]= -2015345591;
assign addr[65161]= -2028233973;
assign addr[65162]= -2040479063;
assign addr[65163]= -2052076975;
assign addr[65164]= -2063024031;
assign addr[65165]= -2073316760;
assign addr[65166]= -2082951896;
assign addr[65167]= -2091926384;
assign addr[65168]= -2100237377;
assign addr[65169]= -2107882239;
assign addr[65170]= -2114858546;
assign addr[65171]= -2121164085;
assign addr[65172]= -2126796855;
assign addr[65173]= -2131755071;
assign addr[65174]= -2136037160;
assign addr[65175]= -2139641764;
assign addr[65176]= -2142567738;
assign addr[65177]= -2144814157;
assign addr[65178]= -2146380306;
assign addr[65179]= -2147265689;
assign addr[65180]= -2147470025;
assign addr[65181]= -2146993250;
assign addr[65182]= -2145835515;
assign addr[65183]= -2143997187;
assign addr[65184]= -2141478848;
assign addr[65185]= -2138281298;
assign addr[65186]= -2134405552;
assign addr[65187]= -2129852837;
assign addr[65188]= -2124624598;
assign addr[65189]= -2118722494;
assign addr[65190]= -2112148396;
assign addr[65191]= -2104904390;
assign addr[65192]= -2096992772;
assign addr[65193]= -2088416053;
assign addr[65194]= -2079176953;
assign addr[65195]= -2069278401;
assign addr[65196]= -2058723538;
assign addr[65197]= -2047515711;
assign addr[65198]= -2035658475;
assign addr[65199]= -2023155591;
assign addr[65200]= -2010011024;
assign addr[65201]= -1996228943;
assign addr[65202]= -1981813720;
assign addr[65203]= -1966769926;
assign addr[65204]= -1951102334;
assign addr[65205]= -1934815911;
assign addr[65206]= -1917915825;
assign addr[65207]= -1900407434;
assign addr[65208]= -1882296293;
assign addr[65209]= -1863588145;
assign addr[65210]= -1844288924;
assign addr[65211]= -1824404752;
assign addr[65212]= -1803941934;
assign addr[65213]= -1782906961;
assign addr[65214]= -1761306505;
assign addr[65215]= -1739147417;
assign addr[65216]= -1716436725;
assign addr[65217]= -1693181631;
assign addr[65218]= -1669389513;
assign addr[65219]= -1645067915;
assign addr[65220]= -1620224553;
assign addr[65221]= -1594867305;
assign addr[65222]= -1569004214;
assign addr[65223]= -1542643483;
assign addr[65224]= -1515793473;
assign addr[65225]= -1488462700;
assign addr[65226]= -1460659832;
assign addr[65227]= -1432393688;
assign addr[65228]= -1403673233;
assign addr[65229]= -1374507575;
assign addr[65230]= -1344905966;
assign addr[65231]= -1314877795;
assign addr[65232]= -1284432584;
assign addr[65233]= -1253579991;
assign addr[65234]= -1222329801;
assign addr[65235]= -1190691925;
assign addr[65236]= -1158676398;
assign addr[65237]= -1126293375;
assign addr[65238]= -1093553126;
assign addr[65239]= -1060466036;
assign addr[65240]= -1027042599;
assign addr[65241]= -993293415;
assign addr[65242]= -959229189;
assign addr[65243]= -924860725;
assign addr[65244]= -890198924;
assign addr[65245]= -855254778;
assign addr[65246]= -820039373;
assign addr[65247]= -784563876;
assign addr[65248]= -748839539;
assign addr[65249]= -712877694;
assign addr[65250]= -676689746;
assign addr[65251]= -640287172;
assign addr[65252]= -603681519;
assign addr[65253]= -566884397;
assign addr[65254]= -529907477;
assign addr[65255]= -492762486;
assign addr[65256]= -455461206;
assign addr[65257]= -418015468;
assign addr[65258]= -380437148;
assign addr[65259]= -342738165;
assign addr[65260]= -304930476;
assign addr[65261]= -267026072;
assign addr[65262]= -229036977;
assign addr[65263]= -190975237;
assign addr[65264]= -152852926;
assign addr[65265]= -114682135;
assign addr[65266]= -76474970;
assign addr[65267]= -38243550;
assign addr[65268]= 0;
assign addr[65269]= 38243550;
assign addr[65270]= 76474970;
assign addr[65271]= 114682135;
assign addr[65272]= 152852926;
assign addr[65273]= 190975237;
assign addr[65274]= 229036977;
assign addr[65275]= 267026072;
assign addr[65276]= 304930476;
assign addr[65277]= 342738165;
assign addr[65278]= 380437148;
assign addr[65279]= 418015468;
assign addr[65280]= 455461206;
assign addr[65281]= 492762486;
assign addr[65282]= 529907477;
assign addr[65283]= 566884397;
assign addr[65284]= 603681519;
assign addr[65285]= 640287172;
assign addr[65286]= 676689746;
assign addr[65287]= 712877694;
assign addr[65288]= 748839539;
assign addr[65289]= 784563876;
assign addr[65290]= 820039373;
assign addr[65291]= 855254778;
assign addr[65292]= 890198924;
assign addr[65293]= 924860725;
assign addr[65294]= 959229189;
assign addr[65295]= 993293415;
assign addr[65296]= 1027042599;
assign addr[65297]= 1060466036;
assign addr[65298]= 1093553126;
assign addr[65299]= 1126293375;
assign addr[65300]= 1158676398;
assign addr[65301]= 1190691925;
assign addr[65302]= 1222329801;
assign addr[65303]= 1253579991;
assign addr[65304]= 1284432584;
assign addr[65305]= 1314877795;
assign addr[65306]= 1344905966;
assign addr[65307]= 1374507575;
assign addr[65308]= 1403673233;
assign addr[65309]= 1432393688;
assign addr[65310]= 1460659832;
assign addr[65311]= 1488462700;
assign addr[65312]= 1515793473;
assign addr[65313]= 1542643483;
assign addr[65314]= 1569004214;
assign addr[65315]= 1594867305;
assign addr[65316]= 1620224553;
assign addr[65317]= 1645067915;
assign addr[65318]= 1669389513;
assign addr[65319]= 1693181631;
assign addr[65320]= 1716436725;
assign addr[65321]= 1739147417;
assign addr[65322]= 1761306505;
assign addr[65323]= 1782906961;
assign addr[65324]= 1803941934;
assign addr[65325]= 1824404752;
assign addr[65326]= 1844288924;
assign addr[65327]= 1863588145;
assign addr[65328]= 1882296293;
assign addr[65329]= 1900407434;
assign addr[65330]= 1917915825;
assign addr[65331]= 1934815911;
assign addr[65332]= 1951102334;
assign addr[65333]= 1966769926;
assign addr[65334]= 1981813720;
assign addr[65335]= 1996228943;
assign addr[65336]= 2010011024;
assign addr[65337]= 2023155591;
assign addr[65338]= 2035658475;
assign addr[65339]= 2047515711;
assign addr[65340]= 2058723538;
assign addr[65341]= 2069278401;
assign addr[65342]= 2079176953;
assign addr[65343]= 2088416053;
assign addr[65344]= 2096992772;
assign addr[65345]= 2104904390;
assign addr[65346]= 2112148396;
assign addr[65347]= 2118722494;
assign addr[65348]= 2124624598;
assign addr[65349]= 2129852837;
assign addr[65350]= 2134405552;
assign addr[65351]= 2138281298;
assign addr[65352]= 2141478848;
assign addr[65353]= 2143997187;
assign addr[65354]= 2145835515;
assign addr[65355]= 2146993250;
assign addr[65356]= 2147470025;
assign addr[65357]= 2147265689;
assign addr[65358]= 2146380306;
assign addr[65359]= 2144814157;
assign addr[65360]= 2142567738;
assign addr[65361]= 2139641764;
assign addr[65362]= 2136037160;
assign addr[65363]= 2131755071;
assign addr[65364]= 2126796855;
assign addr[65365]= 2121164085;
assign addr[65366]= 2114858546;
assign addr[65367]= 2107882239;
assign addr[65368]= 2100237377;
assign addr[65369]= 2091926384;
assign addr[65370]= 2082951896;
assign addr[65371]= 2073316760;
assign addr[65372]= 2063024031;
assign addr[65373]= 2052076975;
assign addr[65374]= 2040479063;
assign addr[65375]= 2028233973;
assign addr[65376]= 2015345591;
assign addr[65377]= 2001818002;
assign addr[65378]= 1987655498;
assign addr[65379]= 1972862571;
assign addr[65380]= 1957443913;
assign addr[65381]= 1941404413;
assign addr[65382]= 1924749160;
assign addr[65383]= 1907483436;
assign addr[65384]= 1889612716;
assign addr[65385]= 1871142669;
assign addr[65386]= 1852079154;
assign addr[65387]= 1832428215;
assign addr[65388]= 1812196087;
assign addr[65389]= 1791389186;
assign addr[65390]= 1770014111;
assign addr[65391]= 1748077642;
assign addr[65392]= 1725586737;
assign addr[65393]= 1702548529;
assign addr[65394]= 1678970324;
assign addr[65395]= 1654859602;
assign addr[65396]= 1630224009;
assign addr[65397]= 1605071359;
assign addr[65398]= 1579409630;
assign addr[65399]= 1553246960;
assign addr[65400]= 1526591649;
assign addr[65401]= 1499452149;
assign addr[65402]= 1471837070;
assign addr[65403]= 1443755168;
assign addr[65404]= 1415215352;
assign addr[65405]= 1386226674;
assign addr[65406]= 1356798326;
assign addr[65407]= 1326939644;
assign addr[65408]= 1296660098;
assign addr[65409]= 1265969291;
assign addr[65410]= 1234876957;
assign addr[65411]= 1203392958;
assign addr[65412]= 1171527280;
assign addr[65413]= 1139290029;
assign addr[65414]= 1106691431;
assign addr[65415]= 1073741824;
assign addr[65416]= 1040451659;
assign addr[65417]= 1006831495;
assign addr[65418]= 972891995;
assign addr[65419]= 938643924;
assign addr[65420]= 904098143;
assign addr[65421]= 869265610;
assign addr[65422]= 834157373;
assign addr[65423]= 798784567;
assign addr[65424]= 763158411;
assign addr[65425]= 727290205;
assign addr[65426]= 691191324;
assign addr[65427]= 654873219;
assign addr[65428]= 618347408;
assign addr[65429]= 581625477;
assign addr[65430]= 544719071;
assign addr[65431]= 507639898;
assign addr[65432]= 470399716;
assign addr[65433]= 433010339;
assign addr[65434]= 395483624;
assign addr[65435]= 357831473;
assign addr[65436]= 320065829;
assign addr[65437]= 282198671;
assign addr[65438]= 244242007;
assign addr[65439]= 206207878;
assign addr[65440]= 168108346;
assign addr[65441]= 129955495;
assign addr[65442]= 91761426;
assign addr[65443]= 53538253;
assign addr[65444]= 15298099;
assign addr[65445]= -22946906;
assign addr[65446]= -61184634;
assign addr[65447]= -99402956;
assign addr[65448]= -137589750;
assign addr[65449]= -175732905;
assign addr[65450]= -213820322;
assign addr[65451]= -251839923;
assign addr[65452]= -289779648;
assign addr[65453]= -327627463;
assign addr[65454]= -365371365;
assign addr[65455]= -402999383;
assign addr[65456]= -440499581;
assign addr[65457]= -477860067;
assign addr[65458]= -515068990;
assign addr[65459]= -552114549;
assign addr[65460]= -588984994;
assign addr[65461]= -625668632;
assign addr[65462]= -662153826;
assign addr[65463]= -698429006;
assign addr[65464]= -734482665;
assign addr[65465]= -770303369;
assign addr[65466]= -805879757;
assign addr[65467]= -841200544;
assign addr[65468]= -876254528;
assign addr[65469]= -911030591;
assign addr[65470]= -945517704;
assign addr[65471]= -979704927;
assign addr[65472]= -1013581418;
assign addr[65473]= -1047136432;
assign addr[65474]= -1080359326;
assign addr[65475]= -1113239564;
assign addr[65476]= -1145766716;
assign addr[65477]= -1177930466;
assign addr[65478]= -1209720613;
assign addr[65479]= -1241127074;
assign addr[65480]= -1272139887;
assign addr[65481]= -1302749217;
assign addr[65482]= -1332945355;
assign addr[65483]= -1362718723;
assign addr[65484]= -1392059879;
assign addr[65485]= -1420959516;
assign addr[65486]= -1449408469;
assign addr[65487]= -1477397714;
assign addr[65488]= -1504918373;
assign addr[65489]= -1531961719;
assign addr[65490]= -1558519173;
assign addr[65491]= -1584582314;
assign addr[65492]= -1610142873;
assign addr[65493]= -1635192744;
assign addr[65494]= -1659723983;
assign addr[65495]= -1683728808;
assign addr[65496]= -1707199606;
assign addr[65497]= -1730128933;
assign addr[65498]= -1752509516;
assign addr[65499]= -1774334257;
assign addr[65500]= -1795596234;
assign addr[65501]= -1816288703;
assign addr[65502]= -1836405100;
assign addr[65503]= -1855939047;
assign addr[65504]= -1874884346;
assign addr[65505]= -1893234990;
assign addr[65506]= -1910985158;
assign addr[65507]= -1928129220;
assign addr[65508]= -1944661739;
assign addr[65509]= -1960577471;
assign addr[65510]= -1975871368;
assign addr[65511]= -1990538579;
assign addr[65512]= -2004574453;
assign addr[65513]= -2017974537;
assign addr[65514]= -2030734582;
assign addr[65515]= -2042850540;
assign addr[65516]= -2054318569;
assign addr[65517]= -2065135031;
assign addr[65518]= -2075296495;
assign addr[65519]= -2084799740;
assign addr[65520]= -2093641749;
assign addr[65521]= -2101819720;
assign addr[65522]= -2109331059;
assign addr[65523]= -2116173382;
assign addr[65524]= -2122344521;
assign addr[65525]= -2127842516;
assign addr[65526]= -2132665626;
assign addr[65527]= -2136812319;
assign addr[65528]= -2140281282;
assign addr[65529]= -2143071413;
assign addr[65530]= -2145181827;
assign addr[65531]= -2146611856;
assign addr[65532]= -2147361045;
assign addr[65533]= -2147429158;
assign addr[65534]= -2146816171;
assign addr[65535]= -2145522281;
endmodule