module rompcm705_v3(
	input clk,//49m
	input reset_n,
	output signed [31:0]addrout
);

wire signed [31:0]addr[0:65535];
reg [5:0]k;
wire lrck;
always @(posedge clk or negedge reset_n)begin
	if(reset_n ==0) 
	k = 0;
	
	else
	k <= k+1;

end
assign lrck = k[5];
reg [15:0]i;
always @(posedge lrck or negedge reset_n)begin
	if(reset_n ==0)begin
		i <= 0;
	//	addrout <= 32'd0;
		end
	
	else begin
		i <= i+1;
	//	addrout <= addr[i];
		end
end
assign addrout = addr[i];
assign addr[0] = 0;
assign addr[1] = -16039;
assign addr[2] = -153364;
assign addr[3] = -640904;
assign addr[4] = -1430647;
assign addr[5] = -1301779;
assign addr[6] = 2355806;
assign addr[7] = 11917167;
assign addr[8] = 27381545;
assign addr[9] = 46372366;
assign addr[10] = 66278007;
assign addr[11] = 85876139;
assign addr[12] = 105117235;
assign addr[13] = 124228708;
assign addr[14] = 143314291;
assign addr[15] = 162388511;
assign addr[16] = 181449854;
assign addr[17] = 200496809;
assign addr[18] = 219527866;
assign addr[19] = 238541516;
assign addr[20] = 257536251;
assign addr[21] = 276510565;
assign addr[22] = 295462954;
assign addr[23] = 314391913;
assign addr[24] = 333295944;
assign addr[25] = 352173546;
assign addr[26] = 371023223;
assign addr[27] = 389843480;
assign addr[28] = 408632825;
assign addr[29] = 427389768;
assign addr[30] = 446112822;
assign addr[31] = 464800501;
assign addr[32] = 483451325;
assign addr[33] = 502063814;
assign addr[34] = 520636492;
assign addr[35] = 539167887;
assign addr[36] = 557656529;
assign addr[37] = 576100953;
assign addr[38] = 594499695;
assign addr[39] = 612851297;
assign addr[40] = 631154304;
assign addr[41] = 649407264;
assign addr[42] = 667608730;
assign addr[43] = 685757258;
assign addr[44] = 703851410;
assign addr[45] = 721889752;
assign addr[46] = 739870851;
assign addr[47] = 757793284;
assign addr[48] = 775655628;
assign addr[49] = 793456467;
assign addr[50] = 811194391;
assign addr[51] = 828867991;
assign addr[52] = 846475867;
assign addr[53] = 864016623;
assign addr[54] = 881488868;
assign addr[55] = 898891215;
assign addr[56] = 916222287;
assign addr[57] = 933480707;
assign addr[58] = 950665109;
assign addr[59] = 967774128;
assign addr[60] = 984806408;
assign addr[61] = 1001760600;
assign addr[62] = 1018635358;
assign addr[63] = 1035429345;
assign addr[64] = 1052141228;
assign addr[65] = 1068769683;
assign addr[66] = 1085313391;
assign addr[67] = 1101771040;
assign addr[68] = 1118141326;
assign addr[69] = 1134422949;
assign addr[70] = 1150614620;
assign addr[71] = 1166715055;
assign addr[72] = 1182722976;
assign addr[73] = 1198637114;
assign addr[74] = 1214456207;
assign addr[75] = 1230179002;
assign addr[76] = 1245804251;
assign addr[77] = 1261330715;
assign addr[78] = 1276757164;
assign addr[79] = 1292082373;
assign addr[80] = 1307305128;
assign addr[81] = 1322424222;
assign addr[82] = 1337438456;
assign addr[83] = 1352346639;
assign addr[84] = 1367147589;
assign addr[85] = 1381840133;
assign addr[86] = 1396423105;
assign addr[87] = 1410895350;
assign addr[88] = 1425255719;
assign addr[89] = 1439503074;
assign addr[90] = 1453636285;
assign addr[91] = 1467654232;
assign addr[92] = 1481555802;
assign addr[93] = 1495339895;
assign addr[94] = 1509005416;
assign addr[95] = 1522551282;
assign addr[96] = 1535976419;
assign addr[97] = 1549279763;
assign addr[98] = 1562460258;
assign addr[99] = 1575516860;
assign addr[100] = 1588448533;
assign addr[101] = 1601254251;
assign addr[102] = 1613933000;
assign addr[103] = 1626483774;
assign addr[104] = 1638905577;
assign addr[105] = 1651197426;
assign addr[106] = 1663358344;
assign addr[107] = 1675387369;
assign addr[108] = 1687283545;
assign addr[109] = 1699045930;
assign addr[110] = 1710673591;
assign addr[111] = 1722165606;
assign addr[112] = 1733521064;
assign addr[113] = 1744739065;
assign addr[114] = 1755818718;
assign addr[115] = 1766759146;
assign addr[116] = 1777559480;
assign addr[117] = 1788218865;
assign addr[118] = 1798736454;
assign addr[119] = 1809111415;
assign addr[120] = 1819342925;
assign addr[121] = 1829430172;
assign addr[122] = 1839372356;
assign addr[123] = 1849168689;
assign addr[124] = 1858818395;
assign addr[125] = 1868320707;
assign addr[126] = 1877674873;
assign addr[127] = 1886880151;
assign addr[128] = 1895935811;
assign addr[129] = 1904841135;
assign addr[130] = 1913595416;
assign addr[131] = 1922197961;
assign addr[132] = 1930648088;
assign addr[133] = 1938945125;
assign addr[134] = 1947088417;
assign addr[135] = 1955077316;
assign addr[136] = 1962911189;
assign addr[137] = 1970589416;
assign addr[138] = 1978111387;
assign addr[139] = 1985476506;
assign addr[140] = 1992684188;
assign addr[141] = 1999733863;
assign addr[142] = 2006624971;
assign addr[143] = 2013356967;
assign addr[144] = 2019929315;
assign addr[145] = 2026341495;
assign addr[146] = 2032592999;
assign addr[147] = 2038683330;
assign addr[148] = 2044612007;
assign addr[149] = 2050378558;
assign addr[150] = 2055982526;
assign addr[151] = 2061423468;
assign addr[152] = 2066700952;
assign addr[153] = 2071814558;
assign addr[154] = 2076763883;
assign addr[155] = 2081548533;
assign addr[156] = 2086168128;
assign addr[157] = 2090622304;
assign addr[158] = 2094910706;
assign addr[159] = 2099032994;
assign addr[160] = 2102988841;
assign addr[161] = 2106777935;
assign addr[162] = 2110399974;
assign addr[163] = 2113854671;
assign addr[164] = 2117141752;
assign addr[165] = 2120260957;
assign addr[166] = 2123212038;
assign addr[167] = 2125994762;
assign addr[168] = 2128608907;
assign addr[169] = 2131054266;
assign addr[170] = 2133330646;
assign addr[171] = 2135437865;
assign addr[172] = 2137375758;
assign addr[173] = 2139144169;
assign addr[174] = 2140742960;
assign addr[175] = 2142172003;
assign addr[176] = 2143431184;
assign addr[177] = 2144520405;
assign addr[178] = 2145439578;
assign addr[179] = 2146188631;
assign addr[180] = 2146767505;
assign addr[181] = 2147176152;
assign addr[182] = 2147414542;
assign addr[183] = 2147482655;
assign addr[184] = 2147380486;
assign addr[185] = 2147108043;
assign addr[186] = 2146665347;
assign addr[187] = 2146052433;
assign addr[188] = 2145269351;
assign addr[189] = 2144316162;
assign addr[190] = 2143192942;
assign addr[191] = 2141899780;
assign addr[192] = 2140436778;
assign addr[193] = 2138804053;
assign addr[194] = 2137001733;
assign addr[195] = 2135029962;
assign addr[196] = 2132888897;
assign addr[197] = 2130578706;
assign addr[198] = 2128099574;
assign addr[199] = 2125451696;
assign addr[200] = 2122635283;
assign addr[201] = 2119650558;
assign addr[202] = 2116497758;
assign addr[203] = 2113177132;
assign addr[204] = 2109688944;
assign addr[205] = 2106033471;
assign addr[206] = 2102211002;
assign addr[207] = 2098221841;
assign addr[208] = 2094066304;
assign addr[209] = 2089744719;
assign addr[210] = 2085257431;
assign addr[211] = 2080604795;
assign addr[212] = 2075787180;
assign addr[213] = 2070804967;
assign addr[214] = 2065658552;
assign addr[215] = 2060348343;
assign addr[216] = 2054874761;
assign addr[217] = 2049238240;
assign addr[218] = 2043439226;
assign addr[219] = 2037478181;
assign addr[220] = 2031355576;
assign addr[221] = 2025071897;
assign addr[222] = 2018627642;
assign addr[223] = 2012023322;
assign addr[224] = 2005259462;
assign addr[225] = 1998336596;
assign addr[226] = 1991255274;
assign addr[227] = 1984016058;
assign addr[228] = 1976619522;
assign addr[229] = 1969066252;
assign addr[230] = 1961356847;
assign addr[231] = 1953491918;
assign addr[232] = 1945472089;
assign addr[233] = 1937297997;
assign addr[234] = 1928970288;
assign addr[235] = 1920489624;
assign addr[236] = 1911856677;
assign addr[237] = 1903072131;
assign addr[238] = 1894136683;
assign addr[239] = 1885051042;
assign addr[240] = 1875815927;
assign addr[241] = 1866432072;
assign addr[242] = 1856900221;
assign addr[243] = 1847221128;
assign addr[244] = 1837395562;
assign addr[245] = 1827424302;
assign addr[246] = 1817308138;
assign addr[247] = 1807047873;
assign addr[248] = 1796644320;
assign addr[249] = 1786098304;
assign addr[250] = 1775410662;
assign addr[251] = 1764582240;
assign addr[252] = 1753613897;
assign addr[253] = 1742506504;
assign addr[254] = 1731260941;
assign addr[255] = 1719878099;
assign addr[256] = 1708358881;
assign addr[257] = 1696704201;
assign addr[258] = 1684914983;
assign addr[259] = 1672992161;
assign addr[260] = 1660936681;
assign addr[261] = 1648749499;
assign addr[262] = 1636431582;
assign addr[263] = 1623983905;
assign addr[264] = 1611407456;
assign addr[265] = 1598703233;
assign addr[266] = 1585872242;
assign addr[267] = 1572915501;
assign addr[268] = 1559834037;
assign addr[269] = 1546628888;
assign addr[270] = 1533301101;
assign addr[271] = 1519851733;
assign addr[272] = 1506281850;
assign addr[273] = 1492592527;
assign addr[274] = 1478784851;
assign addr[275] = 1464859917;
assign addr[276] = 1450818828;
assign addr[277] = 1436662698;
assign addr[278] = 1422392650;
assign addr[279] = 1408009814;
assign addr[280] = 1393515332;
assign addr[281] = 1378910353;
assign addr[282] = 1364196034;
assign addr[283] = 1349373543;
assign addr[284] = 1334444055;
assign addr[285] = 1319408754;
assign addr[286] = 1304268832;
assign addr[287] = 1289025489;
assign addr[288] = 1273679934;
assign addr[289] = 1258233384;
assign addr[290] = 1242687064;
assign addr[291] = 1227042207;
assign addr[292] = 1211300053;
assign addr[293] = 1195461849;
assign addr[294] = 1179528853;
assign addr[295] = 1163502328;
assign addr[296] = 1147383544;
assign addr[297] = 1131173780;
assign addr[298] = 1114874320;
assign addr[299] = 1098486458;
assign addr[300] = 1082011492;
assign addr[301] = 1065450729;
assign addr[302] = 1048805483;
assign addr[303] = 1032077073;
assign addr[304] = 1015266825;
assign addr[305] = 998376073;
assign addr[306] = 981406156;
assign addr[307] = 964358420;
assign addr[308] = 947234215;
assign addr[309] = 930034901;
assign addr[310] = 912761841;
assign addr[311] = 895416404;
assign addr[312] = 877999966;
assign addr[313] = 860513908;
assign addr[314] = 842959617;
assign addr[315] = 825338484;
assign addr[316] = 807651907;
assign addr[317] = 789901288;
assign addr[318] = 772088034;
assign addr[319] = 754213559;
assign addr[320] = 736279279;
assign addr[321] = 718286617;
assign addr[322] = 700236999;
assign addr[323] = 682131857;
assign addr[324] = 663972625;
assign addr[325] = 645760745;
assign addr[326] = 627497660;
assign addr[327] = 609184818;
assign addr[328] = 590823671;
assign addr[329] = 572415676;
assign addr[330] = 553962291;
assign addr[331] = 535464981;
assign addr[332] = 516925212;
assign addr[333] = 498344454;
assign addr[334] = 479724180;
assign addr[335] = 461065866;
assign addr[336] = 442370993;
assign addr[337] = 423641043;
assign addr[338] = 404877501;
assign addr[339] = 386081854;
assign addr[340] = 367255594;
assign addr[341] = 348400212;
assign addr[342] = 329517204;
assign addr[343] = 310608068;
assign addr[344] = 291674302;
assign addr[345] = 272717408;
assign addr[346] = 253738890;
assign addr[347] = 234740251;
assign addr[348] = 215722999;
assign addr[349] = 196688642;
assign addr[350] = 177638688;
assign addr[351] = 158574649;
assign addr[352] = 139498035;
assign addr[353] = 120410361;
assign addr[354] = 101313138;
assign addr[355] = 82207882;
assign addr[356] = 63096108;
assign addr[357] = 43979330;
assign addr[358] = 24859065;
assign addr[359] = 5736829;
assign addr[360] = -13385863;
assign addr[361] = -32507492;
assign addr[362] = -51626544;
assign addr[363] = -70741503;
assign addr[364] = -89850852;
assign addr[365] = -108953076;
assign addr[366] = -128046661;
assign addr[367] = -147130093;
assign addr[368] = -166201858;
assign addr[369] = -185260444;
assign addr[370] = -204304341;
assign addr[371] = -223332037;
assign addr[372] = -242342025;
assign addr[373] = -261332796;
assign addr[374] = -280302845;
assign addr[375] = -299250668;
assign addr[376] = -318174762;
assign addr[377] = -337073627;
assign addr[378] = -355945764;
assign addr[379] = -374789676;
assign addr[380] = -393603870;
assign addr[381] = -412386854;
assign addr[382] = -431137138;
assign addr[383] = -449853235;
assign addr[384] = -468533662;
assign addr[385] = -487176937;
assign addr[386] = -505781581;
assign addr[387] = -524346121;
assign addr[388] = -542869083;
assign addr[389] = -561348998;
assign addr[390] = -579784402;
assign addr[391] = -598173833;
assign addr[392] = -616515832;
assign addr[393] = -634808946;
assign addr[394] = -653051723;
assign addr[395] = -671242716;
assign addr[396] = -689380485;
assign addr[397] = -707463589;
assign addr[398] = -725490597;
assign addr[399] = -743460077;
assign addr[400] = -761370605;
assign addr[401] = -779220762;
assign addr[402] = -797009130;
assign addr[403] = -814734301;
assign addr[404] = -832394869;
assign addr[405] = -849989433;
assign addr[406] = -867516597;
assign addr[407] = -884974973;
assign addr[408] = -902363176;
assign addr[409] = -919679827;
assign addr[410] = -936923553;
assign addr[411] = -954092986;
assign addr[412] = -971186766;
assign addr[413] = -988203537;
assign addr[414] = -1005141949;
assign addr[415] = -1022000660;
assign addr[416] = -1038778332;
assign addr[417] = -1055473635;
assign addr[418] = -1072085246;
assign addr[419] = -1088611847;
assign addr[420] = -1105052128;
assign addr[421] = -1121404785;
assign addr[422] = -1137668521;
assign addr[423] = -1153842047;
assign addr[424] = -1169924081;
assign addr[425] = -1185913346;
assign addr[426] = -1201808576;
assign addr[427] = -1217608510;
assign addr[428] = -1233311895;
assign addr[429] = -1248917486;
assign addr[430] = -1264424045;
assign addr[431] = -1279830344;
assign addr[432] = -1295135159;
assign addr[433] = -1310337279;
assign addr[434] = -1325435496;
assign addr[435] = -1340428615;
assign addr[436] = -1355315445;
assign addr[437] = -1370094808;
assign addr[438] = -1384765530;
assign addr[439] = -1399326449;
assign addr[440] = -1413776410;
assign addr[441] = -1428114267;
assign addr[442] = -1442338884;
assign addr[443] = -1456449131;
assign addr[444] = -1470443891;
assign addr[445] = -1484322054;
assign addr[446] = -1498082520;
assign addr[447] = -1511724196;
assign addr[448] = -1525246002;
assign addr[449] = -1538646865;
assign addr[450] = -1551925723;
assign addr[451] = -1565081523;
assign addr[452] = -1578113222;
assign addr[453] = -1591019785;
assign addr[454] = -1603800191;
assign addr[455] = -1616453425;
assign addr[456] = -1628978484;
assign addr[457] = -1641374375;
assign addr[458] = -1653640115;
assign addr[459] = -1665774731;
assign addr[460] = -1677777262;
assign addr[461] = -1689646755;
assign addr[462] = -1701382270;
assign addr[463] = -1712982875;
assign addr[464] = -1724447652;
assign addr[465] = -1735775690;
assign addr[466] = -1746966091;
assign addr[467] = -1758017969;
assign addr[468] = -1768930447;
assign addr[469] = -1779702660;
assign addr[470] = -1790333753;
assign addr[471] = -1800822883;
assign addr[472] = -1811169220;
assign addr[473] = -1821371941;
assign addr[474] = -1831430239;
assign addr[475] = -1841343316;
assign addr[476] = -1851110385;
assign addr[477] = -1860730673;
assign addr[478] = -1870203416;
assign addr[479] = -1879527863;
assign addr[480] = -1888703276;
assign addr[481] = -1897728925;
assign addr[482] = -1906604097;
assign addr[483] = -1915328086;
assign addr[484] = -1923900201;
assign addr[485] = -1932319763;
assign addr[486] = -1940586104;
assign addr[487] = -1948698568;
assign addr[488] = -1956656513;
assign addr[489] = -1964459306;
assign addr[490] = -1972106330;
assign addr[491] = -1979596978;
assign addr[492] = -1986930656;
assign addr[493] = -1994106782;
assign addr[494] = -2001124788;
assign addr[495] = -2007984117;
assign addr[496] = -2014684225;
assign addr[497] = -2021224581;
assign addr[498] = -2027604666;
assign addr[499] = -2033823974;
assign addr[500] = -2039882013;
assign addr[501] = -2045778302;
assign addr[502] = -2051512372;
assign addr[503] = -2057083771;
assign addr[504] = -2062492055;
assign addr[505] = -2067736796;
assign addr[506] = -2072817579;
assign addr[507] = -2077733999;
assign addr[508] = -2082485668;
assign addr[509] = -2087072209;
assign addr[510] = -2091493257;
assign addr[511] = -2095748463;
assign addr[512] = -2099837489;
assign addr[513] = -2103760010;
assign addr[514] = -2107515716;
assign addr[515] = -2111104309;
assign addr[516] = -2114525505;
assign addr[517] = -2117779031;
assign addr[518] = -2120864631;
assign addr[519] = -2123782059;
assign addr[520] = -2126531084;
assign addr[521] = -2129111488;
assign addr[522] = -2131523066;
assign addr[523] = -2133765628;
assign addr[524] = -2135838995;
assign addr[525] = -2137743003;
assign addr[526] = -2139477502;
assign addr[527] = -2141042352;
assign addr[528] = -2142437431;
assign addr[529] = -2143662628;
assign addr[530] = -2144717846;
assign addr[531] = -2145603001;
assign addr[532] = -2146318022;
assign addr[533] = -2146862854;
assign addr[534] = -2147237452;
assign addr[535] = -2147441787;
assign addr[536] = -2147475844;
assign addr[537] = -2147339619;
assign addr[538] = -2147033123;
assign addr[539] = -2146556380;
assign addr[540] = -2145909429;
assign addr[541] = -2145092320;
assign addr[542] = -2144105118;
assign addr[543] = -2142947902;
assign addr[544] = -2141620763;
assign addr[545] = -2140123807;
assign addr[546] = -2138457152;
assign addr[547] = -2136620930;
assign addr[548] = -2134615288;
assign addr[549] = -2132440383;
assign addr[550] = -2130096389;
assign addr[551] = -2127583492;
assign addr[552] = -2124901890;
assign addr[553] = -2122051796;
assign addr[554] = -2119033436;
assign addr[555] = -2115847050;
assign addr[556] = -2112492891;
assign addr[557] = -2108971223;
assign addr[558] = -2105282327;
assign addr[559] = -2101426496;
assign addr[560] = -2097404033;
assign addr[561] = -2093215260;
assign addr[562] = -2088860507;
assign addr[563] = -2084340120;
assign addr[564] = -2079654458;
assign addr[565] = -2074803892;
assign addr[566] = -2069788807;
assign addr[567] = -2064609600;
assign addr[568] = -2059266683;
assign addr[569] = -2053760478;
assign addr[570] = -2048091422;
assign addr[571] = -2042259965;
assign addr[572] = -2036266570;
assign addr[573] = -2030111710;
assign addr[574] = -2023795876;
assign addr[575] = -2017319567;
assign addr[576] = -2010683297;
assign addr[577] = -2003887591;
assign addr[578] = -1996932990;
assign addr[579] = -1989820044;
assign addr[580] = -1982549318;
assign addr[581] = -1975121388;
assign addr[582] = -1967536842;
assign addr[583] = -1959796283;
assign addr[584] = -1951900324;
assign addr[585] = -1943849591;
assign addr[586] = -1935644723;
assign addr[587] = -1927286370;
assign addr[588] = -1918775195;
assign addr[589] = -1910111873;
assign addr[590] = -1901297091;
assign addr[591] = -1892331547;
assign addr[592] = -1883215953;
assign addr[593] = -1873951032;
assign addr[594] = -1864537518;
assign addr[595] = -1854976157;
assign addr[596] = -1845267708;
assign addr[597] = -1835412941;
assign addr[598] = -1825412636;
assign addr[599] = -1815267588;
assign addr[600] = -1804978599;
assign addr[601] = -1794546487;
assign addr[602] = -1783972079;
assign addr[603] = -1773256212;
assign addr[604] = -1762399737;
assign addr[605] = -1751403515;
assign addr[606] = -1740268417;
assign addr[607] = -1728995326;
assign addr[608] = -1717585136;
assign addr[609] = -1706038753;
assign addr[610] = -1694357091;
assign addr[611] = -1682541077;
assign addr[612] = -1670591647;
assign addr[613] = -1658509750;
assign addr[614] = -1646296344;
assign addr[615] = -1633952396;
assign addr[616] = -1621478885;
assign addr[617] = -1608876801;
assign addr[618] = -1596147143;
assign addr[619] = -1583290921;
assign addr[620] = -1570309153;
assign addr[621] = -1557202869;
assign addr[622] = -1543973108;
assign addr[623] = -1530620920;
assign addr[624] = -1517147363;
assign addr[625] = -1503553506;
assign addr[626] = -1489840425;
assign addr[627] = -1476009210;
assign addr[628] = -1462060956;
assign addr[629] = -1447996770;
assign addr[630] = -1433817766;
assign addr[631] = -1419525069;
assign addr[632] = -1405119813;
assign addr[633] = -1390603139;
assign addr[634] = -1375976199;
assign addr[635] = -1361240152;
assign addr[636] = -1346396168;
assign addr[637] = -1331445422;
assign addr[638] = -1316389101;
assign addr[639] = -1301228398;
assign addr[640] = -1285964516;
assign addr[641] = -1270598665;
assign addr[642] = -1255132063;
assign addr[643] = -1239565936;
assign addr[644] = -1223901520;
assign addr[645] = -1208140056;
assign addr[646] = -1192282793;
assign addr[647] = -1176330990;
assign addr[648] = -1160285911;
assign addr[649] = -1144148829;
assign addr[650] = -1127921022;
assign addr[651] = -1111603778;
assign addr[652] = -1095198391;
assign addr[653] = -1078706161;
assign addr[654] = -1062128397;
assign addr[655] = -1045466412;
assign addr[656] = -1028721528;
assign addr[657] = -1011895073;
assign addr[658] = -994988380;
assign addr[659] = -978002791;
assign addr[660] = -960939653;
assign addr[661] = -943800318;
assign addr[662] = -926586145;
assign addr[663] = -909298500;
assign addr[664] = -891938752;
assign addr[665] = -874508280;
assign addr[666] = -857008464;
assign addr[667] = -839440693;
assign addr[668] = -821806359;
assign addr[669] = -804106861;
assign addr[670] = -786343603;
assign addr[671] = -768517992;
assign addr[672] = -750631442;
assign addr[673] = -732685372;
assign addr[674] = -714681204;
assign addr[675] = -696620367;
assign addr[676] = -678504291;
assign addr[677] = -660334415;
assign addr[678] = -642112178;
assign addr[679] = -623839025;
assign addr[680] = -605516406;
assign addr[681] = -587145773;
assign addr[682] = -568728583;
assign addr[683] = -550266296;
assign addr[684] = -531760377;
assign addr[685] = -513212292;
assign addr[686] = -494623513;
assign addr[687] = -475995513;
assign addr[688] = -457329769;
assign addr[689] = -438627762;
assign addr[690] = -419890975;
assign addr[691] = -401120892;
assign addr[692] = -382319004;
assign addr[693] = -363486799;
assign addr[694] = -344625773;
assign addr[695] = -325737419;
assign addr[696] = -306823237;
assign addr[697] = -287884725;
assign addr[698] = -268923386;
assign addr[699] = -249940723;
assign addr[700] = -230938242;
assign addr[701] = -211917448;
assign addr[702] = -192879850;
assign addr[703] = -173826959;
assign addr[704] = -154760284;
assign addr[705] = -135681337;
assign addr[706] = -116591632;
assign addr[707] = -97492681;
assign addr[708] = -78386000;
assign addr[709] = -59273104;
assign addr[710] = -40155507;
assign addr[711] = -21034727;
assign addr[712] = -1912278;
assign addr[713] = 17210322;
assign addr[714] = 36331557;
assign addr[715] = 55449912;
assign addr[716] = 74563870;
assign addr[717] = 93671915;
assign addr[718] = 112772533;
assign addr[719] = 131864208;
assign addr[720] = 150945428;
assign addr[721] = 170014678;
assign addr[722] = 189070447;
assign addr[723] = 208111224;
assign addr[724] = 227135500;
assign addr[725] = 246141764;
assign addr[726] = 265128512;
assign addr[727] = 284094236;
assign addr[728] = 303037433;
assign addr[729] = 321956601;
assign addr[730] = 340850240;
assign addr[731] = 359716852;
assign addr[732] = 378554940;
assign addr[733] = 397363011;
assign addr[734] = 416139574;
assign addr[735] = 434883140;
assign addr[736] = 453592221;
assign addr[737] = 472265336;
assign addr[738] = 490901003;
assign addr[739] = 509497745;
assign addr[740] = 528054086;
assign addr[741] = 546568556;
assign addr[742] = 565039687;
assign addr[743] = 583466013;
assign addr[744] = 601846074;
assign addr[745] = 620178412;
assign addr[746] = 638461574;
assign addr[747] = 656694110;
assign addr[748] = 674874574;
assign addr[749] = 693001525;
assign addr[750] = 711073524;
assign addr[751] = 729089140;
assign addr[752] = 747046944;
assign addr[753] = 764945512;
assign addr[754] = 782783424;
assign addr[755] = 800559266;
assign addr[756] = 818271628;
assign addr[757] = 835919107;
assign addr[758] = 853500302;
assign addr[759] = 871013820;
assign addr[760] = 888458272;
assign addr[761] = 905832274;
assign addr[762] = 923134450;
assign addr[763] = 940363427;
assign addr[764] = 957517838;
assign addr[765] = 974596324;
assign addr[766] = 991597531;
assign addr[767] = 1008520110;
assign addr[768] = 1025362720;
assign addr[769] = 1042124025;
assign addr[770] = 1058802695;
assign addr[771] = 1075397409;
assign addr[772] = 1091906851;
assign addr[773] = 1108329711;
assign addr[774] = 1124664687;
assign addr[775] = 1140910484;
assign addr[776] = 1157065814;
assign addr[777] = 1173129396;
assign addr[778] = 1189099956;
assign addr[779] = 1204976227;
assign addr[780] = 1220756951;
assign addr[781] = 1236440877;
assign addr[782] = 1252026760;
assign addr[783] = 1267513365;
assign addr[784] = 1282899464;
assign addr[785] = 1298183838;
assign addr[786] = 1313365273;
assign addr[787] = 1328442566;
assign addr[788] = 1343414522;
assign addr[789] = 1358279953;
assign addr[790] = 1373037681;
assign addr[791] = 1387686535;
assign addr[792] = 1402225355;
assign addr[793] = 1416652986;
assign addr[794] = 1430968286;
assign addr[795] = 1445170118;
assign addr[796] = 1459257358;
assign addr[797] = 1473228887;
assign addr[798] = 1487083598;
assign addr[799] = 1500820393;
assign addr[800] = 1514438181;
assign addr[801] = 1527935884;
assign addr[802] = 1541312431;
assign addr[803] = 1554566762;
assign addr[804] = 1567697824;
assign addr[805] = 1580704578;
assign addr[806] = 1593585992;
assign addr[807] = 1606341043;
assign addr[808] = 1618968722;
assign addr[809] = 1631468027;
assign addr[810] = 1643837966;
assign addr[811] = 1656077559;
assign addr[812] = 1668185835;
assign addr[813] = 1680161834;
assign addr[814] = 1692004606;
assign addr[815] = 1703713213;
assign addr[816] = 1715286726;
assign addr[817] = 1726724227;
assign addr[818] = 1738024810;
assign addr[819] = 1749187577;
assign addr[820] = 1760211645;
assign addr[821] = 1771096139;
assign addr[822] = 1781840195;
assign addr[823] = 1792442963;
assign addr[824] = 1802903601;
assign addr[825] = 1813221279;
assign addr[826] = 1823395180;
assign addr[827] = 1833424497;
assign addr[828] = 1843308435;
assign addr[829] = 1853046210;
assign addr[830] = 1862637049;
assign addr[831] = 1872080193;
assign addr[832] = 1881374892;
assign addr[833] = 1890520410;
assign addr[834] = 1899516021;
assign addr[835] = 1908361011;
assign addr[836] = 1917054681;
assign addr[837] = 1925596340;
assign addr[838] = 1933985310;
assign addr[839] = 1942220928;
assign addr[840] = 1950302539;
assign addr[841] = 1958229503;
assign addr[842] = 1966001192;
assign addr[843] = 1973616989;
assign addr[844] = 1981076290;
assign addr[845] = 1988378503;
assign addr[846] = 1995523051;
assign addr[847] = 2002509365;
assign addr[848] = 2009336893;
assign addr[849] = 2016005093;
assign addr[850] = 2022513436;
assign addr[851] = 2028861406;
assign addr[852] = 2035048499;
assign addr[853] = 2041074226;
assign addr[854] = 2046938108;
assign addr[855] = 2052639680;
assign addr[856] = 2058178491;
assign addr[857] = 2063554100;
assign addr[858] = 2068766083;
assign addr[859] = 2073814024;
assign addr[860] = 2078697525;
assign addr[861] = 2083416198;
assign addr[862] = 2087969669;
assign addr[863] = 2092357577;
assign addr[864] = 2096579573;
assign addr[865] = 2100635323;
assign addr[866] = 2104524506;
assign addr[867] = 2108246813;
assign addr[868] = 2111801949;
assign addr[869] = 2115189632;
assign addr[870] = 2118409593;
assign addr[871] = 2121461578;
assign addr[872] = 2124345343;
assign addr[873] = 2127060661;
assign addr[874] = 2129607316;
assign addr[875] = 2131985106;
assign addr[876] = 2134193842;
assign addr[877] = 2136233350;
assign addr[878] = 2138103468;
assign addr[879] = 2139804048;
assign addr[880] = 2141334954;
assign addr[881] = 2142696065;
assign addr[882] = 2143887273;
assign addr[883] = 2144908484;
assign addr[884] = 2145759618;
assign addr[885] = 2146440605;
assign addr[886] = 2146951393;
assign addr[887] = 2147291941;
assign addr[888] = 2147462221;
assign addr[889] = 2147462221;
assign addr[890] = 2147291941;
assign addr[891] = 2146951393;
assign addr[892] = 2146440605;
assign addr[893] = 2145759618;
assign addr[894] = 2144908484;
assign addr[895] = 2143887273;
assign addr[896] = 2142696065;
assign addr[897] = 2141334954;
assign addr[898] = 2139804048;
assign addr[899] = 2138103468;
assign addr[900] = 2136233350;
assign addr[901] = 2134193842;
assign addr[902] = 2131985106;
assign addr[903] = 2129607316;
assign addr[904] = 2127060661;
assign addr[905] = 2124345343;
assign addr[906] = 2121461578;
assign addr[907] = 2118409593;
assign addr[908] = 2115189632;
assign addr[909] = 2111801949;
assign addr[910] = 2108246813;
assign addr[911] = 2104524506;
assign addr[912] = 2100635323;
assign addr[913] = 2096579573;
assign addr[914] = 2092357577;
assign addr[915] = 2087969669;
assign addr[916] = 2083416198;
assign addr[917] = 2078697525;
assign addr[918] = 2073814024;
assign addr[919] = 2068766083;
assign addr[920] = 2063554100;
assign addr[921] = 2058178491;
assign addr[922] = 2052639680;
assign addr[923] = 2046938108;
assign addr[924] = 2041074226;
assign addr[925] = 2035048499;
assign addr[926] = 2028861406;
assign addr[927] = 2022513436;
assign addr[928] = 2016005093;
assign addr[929] = 2009336893;
assign addr[930] = 2002509365;
assign addr[931] = 1995523051;
assign addr[932] = 1988378503;
assign addr[933] = 1981076290;
assign addr[934] = 1973616989;
assign addr[935] = 1966001192;
assign addr[936] = 1958229503;
assign addr[937] = 1950302539;
assign addr[938] = 1942220928;
assign addr[939] = 1933985310;
assign addr[940] = 1925596340;
assign addr[941] = 1917054681;
assign addr[942] = 1908361011;
assign addr[943] = 1899516021;
assign addr[944] = 1890520410;
assign addr[945] = 1881374892;
assign addr[946] = 1872080193;
assign addr[947] = 1862637049;
assign addr[948] = 1853046210;
assign addr[949] = 1843308435;
assign addr[950] = 1833424497;
assign addr[951] = 1823395180;
assign addr[952] = 1813221279;
assign addr[953] = 1802903601;
assign addr[954] = 1792442963;
assign addr[955] = 1781840195;
assign addr[956] = 1771096139;
assign addr[957] = 1760211645;
assign addr[958] = 1749187577;
assign addr[959] = 1738024810;
assign addr[960] = 1726724227;
assign addr[961] = 1715286726;
assign addr[962] = 1703713213;
assign addr[963] = 1692004606;
assign addr[964] = 1680161834;
assign addr[965] = 1668185835;
assign addr[966] = 1656077559;
assign addr[967] = 1643837966;
assign addr[968] = 1631468027;
assign addr[969] = 1618968722;
assign addr[970] = 1606341043;
assign addr[971] = 1593585992;
assign addr[972] = 1580704578;
assign addr[973] = 1567697824;
assign addr[974] = 1554566762;
assign addr[975] = 1541312431;
assign addr[976] = 1527935884;
assign addr[977] = 1514438181;
assign addr[978] = 1500820393;
assign addr[979] = 1487083598;
assign addr[980] = 1473228887;
assign addr[981] = 1459257358;
assign addr[982] = 1445170118;
assign addr[983] = 1430968286;
assign addr[984] = 1416652986;
assign addr[985] = 1402225355;
assign addr[986] = 1387686535;
assign addr[987] = 1373037681;
assign addr[988] = 1358279953;
assign addr[989] = 1343414522;
assign addr[990] = 1328442566;
assign addr[991] = 1313365273;
assign addr[992] = 1298183838;
assign addr[993] = 1282899464;
assign addr[994] = 1267513365;
assign addr[995] = 1252026760;
assign addr[996] = 1236440877;
assign addr[997] = 1220756951;
assign addr[998] = 1204976227;
assign addr[999] = 1189099956;
assign addr[1000] = 1173129396;
assign addr[1001] = 1157065814;
assign addr[1002] = 1140910484;
assign addr[1003] = 1124664687;
assign addr[1004] = 1108329711;
assign addr[1005] = 1091906851;
assign addr[1006] = 1075397409;
assign addr[1007] = 1058802695;
assign addr[1008] = 1042124025;
assign addr[1009] = 1025362720;
assign addr[1010] = 1008520110;
assign addr[1011] = 991597531;
assign addr[1012] = 974596324;
assign addr[1013] = 957517838;
assign addr[1014] = 940363427;
assign addr[1015] = 923134450;
assign addr[1016] = 905832274;
assign addr[1017] = 888458272;
assign addr[1018] = 871013820;
assign addr[1019] = 853500302;
assign addr[1020] = 835919107;
assign addr[1021] = 818271628;
assign addr[1022] = 800559266;
assign addr[1023] = 782783424;
assign addr[1024] = 764945512;
assign addr[1025] = 747046944;
assign addr[1026] = 729089140;
assign addr[1027] = 711073524;
assign addr[1028] = 693001525;
assign addr[1029] = 674874574;
assign addr[1030] = 656694110;
assign addr[1031] = 638461574;
assign addr[1032] = 620178412;
assign addr[1033] = 601846074;
assign addr[1034] = 583466013;
assign addr[1035] = 565039687;
assign addr[1036] = 546568556;
assign addr[1037] = 528054086;
assign addr[1038] = 509497745;
assign addr[1039] = 490901003;
assign addr[1040] = 472265336;
assign addr[1041] = 453592221;
assign addr[1042] = 434883140;
assign addr[1043] = 416139574;
assign addr[1044] = 397363011;
assign addr[1045] = 378554940;
assign addr[1046] = 359716852;
assign addr[1047] = 340850240;
assign addr[1048] = 321956601;
assign addr[1049] = 303037433;
assign addr[1050] = 284094236;
assign addr[1051] = 265128512;
assign addr[1052] = 246141764;
assign addr[1053] = 227135500;
assign addr[1054] = 208111224;
assign addr[1055] = 189070447;
assign addr[1056] = 170014678;
assign addr[1057] = 150945428;
assign addr[1058] = 131864208;
assign addr[1059] = 112772533;
assign addr[1060] = 93671915;
assign addr[1061] = 74563870;
assign addr[1062] = 55449912;
assign addr[1063] = 36331557;
assign addr[1064] = 17210322;
assign addr[1065] = -1912278;
assign addr[1066] = -21034727;
assign addr[1067] = -40155507;
assign addr[1068] = -59273104;
assign addr[1069] = -78386000;
assign addr[1070] = -97492681;
assign addr[1071] = -116591632;
assign addr[1072] = -135681337;
assign addr[1073] = -154760284;
assign addr[1074] = -173826959;
assign addr[1075] = -192879850;
assign addr[1076] = -211917448;
assign addr[1077] = -230938242;
assign addr[1078] = -249940723;
assign addr[1079] = -268923386;
assign addr[1080] = -287884725;
assign addr[1081] = -306823237;
assign addr[1082] = -325737419;
assign addr[1083] = -344625773;
assign addr[1084] = -363486799;
assign addr[1085] = -382319004;
assign addr[1086] = -401120892;
assign addr[1087] = -419890975;
assign addr[1088] = -438627762;
assign addr[1089] = -457329769;
assign addr[1090] = -475995513;
assign addr[1091] = -494623513;
assign addr[1092] = -513212292;
assign addr[1093] = -531760377;
assign addr[1094] = -550266296;
assign addr[1095] = -568728583;
assign addr[1096] = -587145773;
assign addr[1097] = -605516406;
assign addr[1098] = -623839025;
assign addr[1099] = -642112178;
assign addr[1100] = -660334415;
assign addr[1101] = -678504291;
assign addr[1102] = -696620367;
assign addr[1103] = -714681204;
assign addr[1104] = -732685372;
assign addr[1105] = -750631442;
assign addr[1106] = -768517992;
assign addr[1107] = -786343603;
assign addr[1108] = -804106861;
assign addr[1109] = -821806359;
assign addr[1110] = -839440693;
assign addr[1111] = -857008464;
assign addr[1112] = -874508280;
assign addr[1113] = -891938752;
assign addr[1114] = -909298500;
assign addr[1115] = -926586145;
assign addr[1116] = -943800318;
assign addr[1117] = -960939653;
assign addr[1118] = -978002791;
assign addr[1119] = -994988380;
assign addr[1120] = -1011895073;
assign addr[1121] = -1028721528;
assign addr[1122] = -1045466412;
assign addr[1123] = -1062128397;
assign addr[1124] = -1078706161;
assign addr[1125] = -1095198391;
assign addr[1126] = -1111603778;
assign addr[1127] = -1127921022;
assign addr[1128] = -1144148829;
assign addr[1129] = -1160285911;
assign addr[1130] = -1176330990;
assign addr[1131] = -1192282793;
assign addr[1132] = -1208140056;
assign addr[1133] = -1223901520;
assign addr[1134] = -1239565936;
assign addr[1135] = -1255132063;
assign addr[1136] = -1270598665;
assign addr[1137] = -1285964516;
assign addr[1138] = -1301228398;
assign addr[1139] = -1316389101;
assign addr[1140] = -1331445422;
assign addr[1141] = -1346396168;
assign addr[1142] = -1361240152;
assign addr[1143] = -1375976199;
assign addr[1144] = -1390603139;
assign addr[1145] = -1405119813;
assign addr[1146] = -1419525069;
assign addr[1147] = -1433817766;
assign addr[1148] = -1447996770;
assign addr[1149] = -1462060956;
assign addr[1150] = -1476009210;
assign addr[1151] = -1489840425;
assign addr[1152] = -1503553506;
assign addr[1153] = -1517147363;
assign addr[1154] = -1530620920;
assign addr[1155] = -1543973108;
assign addr[1156] = -1557202869;
assign addr[1157] = -1570309153;
assign addr[1158] = -1583290921;
assign addr[1159] = -1596147143;
assign addr[1160] = -1608876801;
assign addr[1161] = -1621478885;
assign addr[1162] = -1633952396;
assign addr[1163] = -1646296344;
assign addr[1164] = -1658509750;
assign addr[1165] = -1670591647;
assign addr[1166] = -1682541077;
assign addr[1167] = -1694357091;
assign addr[1168] = -1706038753;
assign addr[1169] = -1717585136;
assign addr[1170] = -1728995326;
assign addr[1171] = -1740268417;
assign addr[1172] = -1751403515;
assign addr[1173] = -1762399737;
assign addr[1174] = -1773256212;
assign addr[1175] = -1783972079;
assign addr[1176] = -1794546487;
assign addr[1177] = -1804978599;
assign addr[1178] = -1815267588;
assign addr[1179] = -1825412636;
assign addr[1180] = -1835412941;
assign addr[1181] = -1845267708;
assign addr[1182] = -1854976157;
assign addr[1183] = -1864537518;
assign addr[1184] = -1873951032;
assign addr[1185] = -1883215953;
assign addr[1186] = -1892331547;
assign addr[1187] = -1901297091;
assign addr[1188] = -1910111873;
assign addr[1189] = -1918775195;
assign addr[1190] = -1927286370;
assign addr[1191] = -1935644723;
assign addr[1192] = -1943849591;
assign addr[1193] = -1951900324;
assign addr[1194] = -1959796283;
assign addr[1195] = -1967536842;
assign addr[1196] = -1975121388;
assign addr[1197] = -1982549318;
assign addr[1198] = -1989820044;
assign addr[1199] = -1996932990;
assign addr[1200] = -2003887591;
assign addr[1201] = -2010683297;
assign addr[1202] = -2017319567;
assign addr[1203] = -2023795876;
assign addr[1204] = -2030111710;
assign addr[1205] = -2036266570;
assign addr[1206] = -2042259965;
assign addr[1207] = -2048091422;
assign addr[1208] = -2053760478;
assign addr[1209] = -2059266683;
assign addr[1210] = -2064609600;
assign addr[1211] = -2069788807;
assign addr[1212] = -2074803892;
assign addr[1213] = -2079654458;
assign addr[1214] = -2084340120;
assign addr[1215] = -2088860507;
assign addr[1216] = -2093215260;
assign addr[1217] = -2097404033;
assign addr[1218] = -2101426496;
assign addr[1219] = -2105282327;
assign addr[1220] = -2108971223;
assign addr[1221] = -2112492891;
assign addr[1222] = -2115847050;
assign addr[1223] = -2119033436;
assign addr[1224] = -2122051796;
assign addr[1225] = -2124901890;
assign addr[1226] = -2127583492;
assign addr[1227] = -2130096389;
assign addr[1228] = -2132440383;
assign addr[1229] = -2134615288;
assign addr[1230] = -2136620930;
assign addr[1231] = -2138457152;
assign addr[1232] = -2140123807;
assign addr[1233] = -2141620763;
assign addr[1234] = -2142947902;
assign addr[1235] = -2144105118;
assign addr[1236] = -2145092320;
assign addr[1237] = -2145909429;
assign addr[1238] = -2146556380;
assign addr[1239] = -2147033123;
assign addr[1240] = -2147339619;
assign addr[1241] = -2147475844;
assign addr[1242] = -2147441787;
assign addr[1243] = -2147237452;
assign addr[1244] = -2146862854;
assign addr[1245] = -2146318022;
assign addr[1246] = -2145603001;
assign addr[1247] = -2144717846;
assign addr[1248] = -2143662628;
assign addr[1249] = -2142437431;
assign addr[1250] = -2141042352;
assign addr[1251] = -2139477502;
assign addr[1252] = -2137743003;
assign addr[1253] = -2135838995;
assign addr[1254] = -2133765628;
assign addr[1255] = -2131523066;
assign addr[1256] = -2129111488;
assign addr[1257] = -2126531084;
assign addr[1258] = -2123782059;
assign addr[1259] = -2120864631;
assign addr[1260] = -2117779031;
assign addr[1261] = -2114525505;
assign addr[1262] = -2111104309;
assign addr[1263] = -2107515716;
assign addr[1264] = -2103760010;
assign addr[1265] = -2099837489;
assign addr[1266] = -2095748463;
assign addr[1267] = -2091493257;
assign addr[1268] = -2087072209;
assign addr[1269] = -2082485668;
assign addr[1270] = -2077733999;
assign addr[1271] = -2072817579;
assign addr[1272] = -2067736796;
assign addr[1273] = -2062492055;
assign addr[1274] = -2057083771;
assign addr[1275] = -2051512372;
assign addr[1276] = -2045778302;
assign addr[1277] = -2039882013;
assign addr[1278] = -2033823974;
assign addr[1279] = -2027604666;
assign addr[1280] = -2021224581;
assign addr[1281] = -2014684225;
assign addr[1282] = -2007984117;
assign addr[1283] = -2001124788;
assign addr[1284] = -1994106782;
assign addr[1285] = -1986930656;
assign addr[1286] = -1979596978;
assign addr[1287] = -1972106330;
assign addr[1288] = -1964459306;
assign addr[1289] = -1956656513;
assign addr[1290] = -1948698568;
assign addr[1291] = -1940586104;
assign addr[1292] = -1932319763;
assign addr[1293] = -1923900201;
assign addr[1294] = -1915328086;
assign addr[1295] = -1906604097;
assign addr[1296] = -1897728925;
assign addr[1297] = -1888703276;
assign addr[1298] = -1879527863;
assign addr[1299] = -1870203416;
assign addr[1300] = -1860730673;
assign addr[1301] = -1851110385;
assign addr[1302] = -1841343316;
assign addr[1303] = -1831430239;
assign addr[1304] = -1821371941;
assign addr[1305] = -1811169220;
assign addr[1306] = -1800822883;
assign addr[1307] = -1790333753;
assign addr[1308] = -1779702660;
assign addr[1309] = -1768930447;
assign addr[1310] = -1758017969;
assign addr[1311] = -1746966091;
assign addr[1312] = -1735775690;
assign addr[1313] = -1724447652;
assign addr[1314] = -1712982875;
assign addr[1315] = -1701382270;
assign addr[1316] = -1689646755;
assign addr[1317] = -1677777262;
assign addr[1318] = -1665774731;
assign addr[1319] = -1653640115;
assign addr[1320] = -1641374375;
assign addr[1321] = -1628978484;
assign addr[1322] = -1616453425;
assign addr[1323] = -1603800191;
assign addr[1324] = -1591019785;
assign addr[1325] = -1578113222;
assign addr[1326] = -1565081523;
assign addr[1327] = -1551925723;
assign addr[1328] = -1538646865;
assign addr[1329] = -1525246002;
assign addr[1330] = -1511724196;
assign addr[1331] = -1498082520;
assign addr[1332] = -1484322054;
assign addr[1333] = -1470443891;
assign addr[1334] = -1456449131;
assign addr[1335] = -1442338884;
assign addr[1336] = -1428114267;
assign addr[1337] = -1413776410;
assign addr[1338] = -1399326449;
assign addr[1339] = -1384765530;
assign addr[1340] = -1370094808;
assign addr[1341] = -1355315445;
assign addr[1342] = -1340428615;
assign addr[1343] = -1325435496;
assign addr[1344] = -1310337279;
assign addr[1345] = -1295135159;
assign addr[1346] = -1279830344;
assign addr[1347] = -1264424045;
assign addr[1348] = -1248917486;
assign addr[1349] = -1233311895;
assign addr[1350] = -1217608510;
assign addr[1351] = -1201808576;
assign addr[1352] = -1185913346;
assign addr[1353] = -1169924081;
assign addr[1354] = -1153842047;
assign addr[1355] = -1137668521;
assign addr[1356] = -1121404785;
assign addr[1357] = -1105052128;
assign addr[1358] = -1088611847;
assign addr[1359] = -1072085246;
assign addr[1360] = -1055473635;
assign addr[1361] = -1038778332;
assign addr[1362] = -1022000660;
assign addr[1363] = -1005141949;
assign addr[1364] = -988203537;
assign addr[1365] = -971186766;
assign addr[1366] = -954092986;
assign addr[1367] = -936923553;
assign addr[1368] = -919679827;
assign addr[1369] = -902363176;
assign addr[1370] = -884974973;
assign addr[1371] = -867516597;
assign addr[1372] = -849989433;
assign addr[1373] = -832394869;
assign addr[1374] = -814734301;
assign addr[1375] = -797009130;
assign addr[1376] = -779220762;
assign addr[1377] = -761370605;
assign addr[1378] = -743460077;
assign addr[1379] = -725490597;
assign addr[1380] = -707463589;
assign addr[1381] = -689380485;
assign addr[1382] = -671242716;
assign addr[1383] = -653051723;
assign addr[1384] = -634808946;
assign addr[1385] = -616515832;
assign addr[1386] = -598173833;
assign addr[1387] = -579784402;
assign addr[1388] = -561348998;
assign addr[1389] = -542869083;
assign addr[1390] = -524346121;
assign addr[1391] = -505781581;
assign addr[1392] = -487176937;
assign addr[1393] = -468533662;
assign addr[1394] = -449853235;
assign addr[1395] = -431137138;
assign addr[1396] = -412386854;
assign addr[1397] = -393603870;
assign addr[1398] = -374789676;
assign addr[1399] = -355945764;
assign addr[1400] = -337073627;
assign addr[1401] = -318174762;
assign addr[1402] = -299250668;
assign addr[1403] = -280302845;
assign addr[1404] = -261332796;
assign addr[1405] = -242342025;
assign addr[1406] = -223332037;
assign addr[1407] = -204304341;
assign addr[1408] = -185260444;
assign addr[1409] = -166201858;
assign addr[1410] = -147130093;
assign addr[1411] = -128046661;
assign addr[1412] = -108953076;
assign addr[1413] = -89850852;
assign addr[1414] = -70741503;
assign addr[1415] = -51626544;
assign addr[1416] = -32507492;
assign addr[1417] = -13385863;
assign addr[1418] = 5736829;
assign addr[1419] = 24859065;
assign addr[1420] = 43979330;
assign addr[1421] = 63096108;
assign addr[1422] = 82207882;
assign addr[1423] = 101313138;
assign addr[1424] = 120410361;
assign addr[1425] = 139498035;
assign addr[1426] = 158574649;
assign addr[1427] = 177638688;
assign addr[1428] = 196688642;
assign addr[1429] = 215722999;
assign addr[1430] = 234740251;
assign addr[1431] = 253738890;
assign addr[1432] = 272717408;
assign addr[1433] = 291674302;
assign addr[1434] = 310608068;
assign addr[1435] = 329517204;
assign addr[1436] = 348400212;
assign addr[1437] = 367255594;
assign addr[1438] = 386081854;
assign addr[1439] = 404877501;
assign addr[1440] = 423641043;
assign addr[1441] = 442370993;
assign addr[1442] = 461065866;
assign addr[1443] = 479724180;
assign addr[1444] = 498344454;
assign addr[1445] = 516925212;
assign addr[1446] = 535464981;
assign addr[1447] = 553962291;
assign addr[1448] = 572415676;
assign addr[1449] = 590823671;
assign addr[1450] = 609184818;
assign addr[1451] = 627497660;
assign addr[1452] = 645760745;
assign addr[1453] = 663972625;
assign addr[1454] = 682131857;
assign addr[1455] = 700236999;
assign addr[1456] = 718286617;
assign addr[1457] = 736279279;
assign addr[1458] = 754213559;
assign addr[1459] = 772088034;
assign addr[1460] = 789901288;
assign addr[1461] = 807651907;
assign addr[1462] = 825338484;
assign addr[1463] = 842959617;
assign addr[1464] = 860513908;
assign addr[1465] = 877999966;
assign addr[1466] = 895416404;
assign addr[1467] = 912761841;
assign addr[1468] = 930034901;
assign addr[1469] = 947234215;
assign addr[1470] = 964358420;
assign addr[1471] = 981406156;
assign addr[1472] = 998376073;
assign addr[1473] = 1015266825;
assign addr[1474] = 1032077073;
assign addr[1475] = 1048805483;
assign addr[1476] = 1065450729;
assign addr[1477] = 1082011492;
assign addr[1478] = 1098486458;
assign addr[1479] = 1114874320;
assign addr[1480] = 1131173780;
assign addr[1481] = 1147383544;
assign addr[1482] = 1163502328;
assign addr[1483] = 1179528853;
assign addr[1484] = 1195461849;
assign addr[1485] = 1211300053;
assign addr[1486] = 1227042207;
assign addr[1487] = 1242687064;
assign addr[1488] = 1258233384;
assign addr[1489] = 1273679934;
assign addr[1490] = 1289025489;
assign addr[1491] = 1304268832;
assign addr[1492] = 1319408754;
assign addr[1493] = 1334444055;
assign addr[1494] = 1349373543;
assign addr[1495] = 1364196034;
assign addr[1496] = 1378910353;
assign addr[1497] = 1393515332;
assign addr[1498] = 1408009814;
assign addr[1499] = 1422392650;
assign addr[1500] = 1436662698;
assign addr[1501] = 1450818828;
assign addr[1502] = 1464859917;
assign addr[1503] = 1478784851;
assign addr[1504] = 1492592527;
assign addr[1505] = 1506281850;
assign addr[1506] = 1519851733;
assign addr[1507] = 1533301101;
assign addr[1508] = 1546628888;
assign addr[1509] = 1559834037;
assign addr[1510] = 1572915501;
assign addr[1511] = 1585872242;
assign addr[1512] = 1598703233;
assign addr[1513] = 1611407456;
assign addr[1514] = 1623983905;
assign addr[1515] = 1636431582;
assign addr[1516] = 1648749499;
assign addr[1517] = 1660936681;
assign addr[1518] = 1672992161;
assign addr[1519] = 1684914983;
assign addr[1520] = 1696704201;
assign addr[1521] = 1708358881;
assign addr[1522] = 1719878099;
assign addr[1523] = 1731260941;
assign addr[1524] = 1742506504;
assign addr[1525] = 1753613897;
assign addr[1526] = 1764582240;
assign addr[1527] = 1775410662;
assign addr[1528] = 1786098304;
assign addr[1529] = 1796644320;
assign addr[1530] = 1807047873;
assign addr[1531] = 1817308138;
assign addr[1532] = 1827424302;
assign addr[1533] = 1837395562;
assign addr[1534] = 1847221128;
assign addr[1535] = 1856900221;
assign addr[1536] = 1866432072;
assign addr[1537] = 1875815927;
assign addr[1538] = 1885051042;
assign addr[1539] = 1894136683;
assign addr[1540] = 1903072131;
assign addr[1541] = 1911856677;
assign addr[1542] = 1920489624;
assign addr[1543] = 1928970288;
assign addr[1544] = 1937297997;
assign addr[1545] = 1945472089;
assign addr[1546] = 1953491918;
assign addr[1547] = 1961356847;
assign addr[1548] = 1969066252;
assign addr[1549] = 1976619522;
assign addr[1550] = 1984016058;
assign addr[1551] = 1991255274;
assign addr[1552] = 1998336596;
assign addr[1553] = 2005259462;
assign addr[1554] = 2012023322;
assign addr[1555] = 2018627642;
assign addr[1556] = 2025071897;
assign addr[1557] = 2031355576;
assign addr[1558] = 2037478181;
assign addr[1559] = 2043439226;
assign addr[1560] = 2049238240;
assign addr[1561] = 2054874761;
assign addr[1562] = 2060348343;
assign addr[1563] = 2065658552;
assign addr[1564] = 2070804967;
assign addr[1565] = 2075787180;
assign addr[1566] = 2080604795;
assign addr[1567] = 2085257431;
assign addr[1568] = 2089744719;
assign addr[1569] = 2094066304;
assign addr[1570] = 2098221841;
assign addr[1571] = 2102211002;
assign addr[1572] = 2106033471;
assign addr[1573] = 2109688944;
assign addr[1574] = 2113177132;
assign addr[1575] = 2116497758;
assign addr[1576] = 2119650558;
assign addr[1577] = 2122635283;
assign addr[1578] = 2125451696;
assign addr[1579] = 2128099574;
assign addr[1580] = 2130578706;
assign addr[1581] = 2132888897;
assign addr[1582] = 2135029962;
assign addr[1583] = 2137001733;
assign addr[1584] = 2138804053;
assign addr[1585] = 2140436778;
assign addr[1586] = 2141899780;
assign addr[1587] = 2143192942;
assign addr[1588] = 2144316162;
assign addr[1589] = 2145269351;
assign addr[1590] = 2146052433;
assign addr[1591] = 2146665347;
assign addr[1592] = 2147108043;
assign addr[1593] = 2147380486;
assign addr[1594] = 2147482655;
assign addr[1595] = 2147414542;
assign addr[1596] = 2147176152;
assign addr[1597] = 2146767505;
assign addr[1598] = 2146188631;
assign addr[1599] = 2145439578;
assign addr[1600] = 2144520405;
assign addr[1601] = 2143431184;
assign addr[1602] = 2142172003;
assign addr[1603] = 2140742960;
assign addr[1604] = 2139144169;
assign addr[1605] = 2137375758;
assign addr[1606] = 2135437865;
assign addr[1607] = 2133330646;
assign addr[1608] = 2131054266;
assign addr[1609] = 2128608907;
assign addr[1610] = 2125994762;
assign addr[1611] = 2123212038;
assign addr[1612] = 2120260957;
assign addr[1613] = 2117141752;
assign addr[1614] = 2113854671;
assign addr[1615] = 2110399974;
assign addr[1616] = 2106777935;
assign addr[1617] = 2102988841;
assign addr[1618] = 2099032994;
assign addr[1619] = 2094910706;
assign addr[1620] = 2090622304;
assign addr[1621] = 2086168128;
assign addr[1622] = 2081548533;
assign addr[1623] = 2076763883;
assign addr[1624] = 2071814558;
assign addr[1625] = 2066700952;
assign addr[1626] = 2061423468;
assign addr[1627] = 2055982526;
assign addr[1628] = 2050378558;
assign addr[1629] = 2044612007;
assign addr[1630] = 2038683330;
assign addr[1631] = 2032592999;
assign addr[1632] = 2026341495;
assign addr[1633] = 2019929315;
assign addr[1634] = 2013356967;
assign addr[1635] = 2006624971;
assign addr[1636] = 1999733863;
assign addr[1637] = 1992684188;
assign addr[1638] = 1985476506;
assign addr[1639] = 1978111387;
assign addr[1640] = 1970589416;
assign addr[1641] = 1962911189;
assign addr[1642] = 1955077316;
assign addr[1643] = 1947088417;
assign addr[1644] = 1938945125;
assign addr[1645] = 1930648088;
assign addr[1646] = 1922197961;
assign addr[1647] = 1913595416;
assign addr[1648] = 1904841135;
assign addr[1649] = 1895935811;
assign addr[1650] = 1886880151;
assign addr[1651] = 1877674873;
assign addr[1652] = 1868320707;
assign addr[1653] = 1858818395;
assign addr[1654] = 1849168689;
assign addr[1655] = 1839372356;
assign addr[1656] = 1829430172;
assign addr[1657] = 1819342925;
assign addr[1658] = 1809111415;
assign addr[1659] = 1798736454;
assign addr[1660] = 1788218865;
assign addr[1661] = 1777559480;
assign addr[1662] = 1766759146;
assign addr[1663] = 1755818718;
assign addr[1664] = 1744739065;
assign addr[1665] = 1733521064;
assign addr[1666] = 1722165606;
assign addr[1667] = 1710673591;
assign addr[1668] = 1699045930;
assign addr[1669] = 1687283545;
assign addr[1670] = 1675387369;
assign addr[1671] = 1663358344;
assign addr[1672] = 1651197426;
assign addr[1673] = 1638905577;
assign addr[1674] = 1626483774;
assign addr[1675] = 1613933000;
assign addr[1676] = 1601254251;
assign addr[1677] = 1588448533;
assign addr[1678] = 1575516860;
assign addr[1679] = 1562460258;
assign addr[1680] = 1549279763;
assign addr[1681] = 1535976419;
assign addr[1682] = 1522551282;
assign addr[1683] = 1509005416;
assign addr[1684] = 1495339895;
assign addr[1685] = 1481555802;
assign addr[1686] = 1467654232;
assign addr[1687] = 1453636285;
assign addr[1688] = 1439503074;
assign addr[1689] = 1425255719;
assign addr[1690] = 1410895350;
assign addr[1691] = 1396423105;
assign addr[1692] = 1381840133;
assign addr[1693] = 1367147589;
assign addr[1694] = 1352346639;
assign addr[1695] = 1337438456;
assign addr[1696] = 1322424222;
assign addr[1697] = 1307305128;
assign addr[1698] = 1292082373;
assign addr[1699] = 1276757164;
assign addr[1700] = 1261330715;
assign addr[1701] = 1245804251;
assign addr[1702] = 1230179002;
assign addr[1703] = 1214456207;
assign addr[1704] = 1198637114;
assign addr[1705] = 1182722976;
assign addr[1706] = 1166715055;
assign addr[1707] = 1150614620;
assign addr[1708] = 1134422949;
assign addr[1709] = 1118141326;
assign addr[1710] = 1101771040;
assign addr[1711] = 1085313391;
assign addr[1712] = 1068769683;
assign addr[1713] = 1052141228;
assign addr[1714] = 1035429345;
assign addr[1715] = 1018635358;
assign addr[1716] = 1001760600;
assign addr[1717] = 984806408;
assign addr[1718] = 967774128;
assign addr[1719] = 950665109;
assign addr[1720] = 933480707;
assign addr[1721] = 916222287;
assign addr[1722] = 898891215;
assign addr[1723] = 881488868;
assign addr[1724] = 864016623;
assign addr[1725] = 846475867;
assign addr[1726] = 828867991;
assign addr[1727] = 811194391;
assign addr[1728] = 793456467;
assign addr[1729] = 775655628;
assign addr[1730] = 757793284;
assign addr[1731] = 739870851;
assign addr[1732] = 721889752;
assign addr[1733] = 703851410;
assign addr[1734] = 685757258;
assign addr[1735] = 667608730;
assign addr[1736] = 649407264;
assign addr[1737] = 631154304;
assign addr[1738] = 612851297;
assign addr[1739] = 594499695;
assign addr[1740] = 576100953;
assign addr[1741] = 557656529;
assign addr[1742] = 539167887;
assign addr[1743] = 520636492;
assign addr[1744] = 502063814;
assign addr[1745] = 483451325;
assign addr[1746] = 464800501;
assign addr[1747] = 446112822;
assign addr[1748] = 427389768;
assign addr[1749] = 408632825;
assign addr[1750] = 389843480;
assign addr[1751] = 371023223;
assign addr[1752] = 352173546;
assign addr[1753] = 333295944;
assign addr[1754] = 314391913;
assign addr[1755] = 295462954;
assign addr[1756] = 276510565;
assign addr[1757] = 257536251;
assign addr[1758] = 238541516;
assign addr[1759] = 219527866;
assign addr[1760] = 200496809;
assign addr[1761] = 181449854;
assign addr[1762] = 162388511;
assign addr[1763] = 143314291;
assign addr[1764] = 124228708;
assign addr[1765] = 105133274;
assign addr[1766] = 86029503;
assign addr[1767] = 66918911;
assign addr[1768] = 47803013;
assign addr[1769] = 28683324;
assign addr[1770] = 9561361;
assign addr[1771] = -9561361;
assign addr[1772] = -28683324;
assign addr[1773] = -47803013;
assign addr[1774] = -66918911;
assign addr[1775] = -86029503;
assign addr[1776] = -105133274;
assign addr[1777] = -124228708;
assign addr[1778] = -143314291;
assign addr[1779] = -162388511;
assign addr[1780] = -181449854;
assign addr[1781] = -200496809;
assign addr[1782] = -219527866;
assign addr[1783] = -238541516;
assign addr[1784] = -257536251;
assign addr[1785] = -276510565;
assign addr[1786] = -295462954;
assign addr[1787] = -314391913;
assign addr[1788] = -333295944;
assign addr[1789] = -352173546;
assign addr[1790] = -371023223;
assign addr[1791] = -389843480;
assign addr[1792] = -408632825;
assign addr[1793] = -427389768;
assign addr[1794] = -446112822;
assign addr[1795] = -464800501;
assign addr[1796] = -483451325;
assign addr[1797] = -502063814;
assign addr[1798] = -520636492;
assign addr[1799] = -539167887;
assign addr[1800] = -557656529;
assign addr[1801] = -576100953;
assign addr[1802] = -594499695;
assign addr[1803] = -612851297;
assign addr[1804] = -631154304;
assign addr[1805] = -649407264;
assign addr[1806] = -667608730;
assign addr[1807] = -685757258;
assign addr[1808] = -703851410;
assign addr[1809] = -721889752;
assign addr[1810] = -739870851;
assign addr[1811] = -757793284;
assign addr[1812] = -775655628;
assign addr[1813] = -793456467;
assign addr[1814] = -811194391;
assign addr[1815] = -828867991;
assign addr[1816] = -846475867;
assign addr[1817] = -864016623;
assign addr[1818] = -881488868;
assign addr[1819] = -898891215;
assign addr[1820] = -916222287;
assign addr[1821] = -933480707;
assign addr[1822] = -950665109;
assign addr[1823] = -967774128;
assign addr[1824] = -984806408;
assign addr[1825] = -1001760600;
assign addr[1826] = -1018635358;
assign addr[1827] = -1035429345;
assign addr[1828] = -1052141228;
assign addr[1829] = -1068769683;
assign addr[1830] = -1085313391;
assign addr[1831] = -1101771040;
assign addr[1832] = -1118141326;
assign addr[1833] = -1134422949;
assign addr[1834] = -1150614620;
assign addr[1835] = -1166715055;
assign addr[1836] = -1182722976;
assign addr[1837] = -1198637114;
assign addr[1838] = -1214456207;
assign addr[1839] = -1230179002;
assign addr[1840] = -1245804251;
assign addr[1841] = -1261330715;
assign addr[1842] = -1276757164;
assign addr[1843] = -1292082373;
assign addr[1844] = -1307305128;
assign addr[1845] = -1322424222;
assign addr[1846] = -1337438456;
assign addr[1847] = -1352346639;
assign addr[1848] = -1367147589;
assign addr[1849] = -1381840133;
assign addr[1850] = -1396423105;
assign addr[1851] = -1410895350;
assign addr[1852] = -1425255719;
assign addr[1853] = -1439503074;
assign addr[1854] = -1453636285;
assign addr[1855] = -1467654232;
assign addr[1856] = -1481555802;
assign addr[1857] = -1495339895;
assign addr[1858] = -1509005416;
assign addr[1859] = -1522551282;
assign addr[1860] = -1535976419;
assign addr[1861] = -1549279763;
assign addr[1862] = -1562460258;
assign addr[1863] = -1575516860;
assign addr[1864] = -1588448533;
assign addr[1865] = -1601254251;
assign addr[1866] = -1613933000;
assign addr[1867] = -1626483774;
assign addr[1868] = -1638905577;
assign addr[1869] = -1651197426;
assign addr[1870] = -1663358344;
assign addr[1871] = -1675387369;
assign addr[1872] = -1687283545;
assign addr[1873] = -1699045930;
assign addr[1874] = -1710673591;
assign addr[1875] = -1722165606;
assign addr[1876] = -1733521064;
assign addr[1877] = -1744739065;
assign addr[1878] = -1755818718;
assign addr[1879] = -1766759146;
assign addr[1880] = -1777559480;
assign addr[1881] = -1788218865;
assign addr[1882] = -1798736454;
assign addr[1883] = -1809111415;
assign addr[1884] = -1819342925;
assign addr[1885] = -1829430172;
assign addr[1886] = -1839372356;
assign addr[1887] = -1849168689;
assign addr[1888] = -1858818395;
assign addr[1889] = -1868320707;
assign addr[1890] = -1877674873;
assign addr[1891] = -1886880151;
assign addr[1892] = -1895935811;
assign addr[1893] = -1904841135;
assign addr[1894] = -1913595416;
assign addr[1895] = -1922197961;
assign addr[1896] = -1930648088;
assign addr[1897] = -1938945125;
assign addr[1898] = -1947088417;
assign addr[1899] = -1955077316;
assign addr[1900] = -1962911189;
assign addr[1901] = -1970589416;
assign addr[1902] = -1978111387;
assign addr[1903] = -1985476506;
assign addr[1904] = -1992684188;
assign addr[1905] = -1999733863;
assign addr[1906] = -2006624971;
assign addr[1907] = -2013356967;
assign addr[1908] = -2019929315;
assign addr[1909] = -2026341495;
assign addr[1910] = -2032592999;
assign addr[1911] = -2038683330;
assign addr[1912] = -2044612007;
assign addr[1913] = -2050378558;
assign addr[1914] = -2055982526;
assign addr[1915] = -2061423468;
assign addr[1916] = -2066700952;
assign addr[1917] = -2071814558;
assign addr[1918] = -2076763883;
assign addr[1919] = -2081548533;
assign addr[1920] = -2086168128;
assign addr[1921] = -2090622304;
assign addr[1922] = -2094910706;
assign addr[1923] = -2099032994;
assign addr[1924] = -2102988841;
assign addr[1925] = -2106777935;
assign addr[1926] = -2110399974;
assign addr[1927] = -2113854671;
assign addr[1928] = -2117141752;
assign addr[1929] = -2120260957;
assign addr[1930] = -2123212038;
assign addr[1931] = -2125994762;
assign addr[1932] = -2128608907;
assign addr[1933] = -2131054266;
assign addr[1934] = -2133330646;
assign addr[1935] = -2135437865;
assign addr[1936] = -2137375758;
assign addr[1937] = -2139144169;
assign addr[1938] = -2140742960;
assign addr[1939] = -2142172003;
assign addr[1940] = -2143431184;
assign addr[1941] = -2144520405;
assign addr[1942] = -2145439578;
assign addr[1943] = -2146188631;
assign addr[1944] = -2146767505;
assign addr[1945] = -2147176152;
assign addr[1946] = -2147414542;
assign addr[1947] = -2147482655;
assign addr[1948] = -2147380486;
assign addr[1949] = -2147108043;
assign addr[1950] = -2146665347;
assign addr[1951] = -2146052433;
assign addr[1952] = -2145269351;
assign addr[1953] = -2144316162;
assign addr[1954] = -2143192942;
assign addr[1955] = -2141899780;
assign addr[1956] = -2140436778;
assign addr[1957] = -2138804053;
assign addr[1958] = -2137001733;
assign addr[1959] = -2135029962;
assign addr[1960] = -2132888897;
assign addr[1961] = -2130578706;
assign addr[1962] = -2128099574;
assign addr[1963] = -2125451696;
assign addr[1964] = -2122635283;
assign addr[1965] = -2119650558;
assign addr[1966] = -2116497758;
assign addr[1967] = -2113177132;
assign addr[1968] = -2109688944;
assign addr[1969] = -2106033471;
assign addr[1970] = -2102211002;
assign addr[1971] = -2098221841;
assign addr[1972] = -2094066304;
assign addr[1973] = -2089744719;
assign addr[1974] = -2085257431;
assign addr[1975] = -2080604795;
assign addr[1976] = -2075787180;
assign addr[1977] = -2070804967;
assign addr[1978] = -2065658552;
assign addr[1979] = -2060348343;
assign addr[1980] = -2054874761;
assign addr[1981] = -2049238240;
assign addr[1982] = -2043439226;
assign addr[1983] = -2037478181;
assign addr[1984] = -2031355576;
assign addr[1985] = -2025071897;
assign addr[1986] = -2018627642;
assign addr[1987] = -2012023322;
assign addr[1988] = -2005259462;
assign addr[1989] = -1998336596;
assign addr[1990] = -1991255274;
assign addr[1991] = -1984016058;
assign addr[1992] = -1976619522;
assign addr[1993] = -1969066252;
assign addr[1994] = -1961356847;
assign addr[1995] = -1953491918;
assign addr[1996] = -1945472089;
assign addr[1997] = -1937297997;
assign addr[1998] = -1928970288;
assign addr[1999] = -1920489624;
assign addr[2000] = -1911856677;
assign addr[2001] = -1903072131;
assign addr[2002] = -1894136683;
assign addr[2003] = -1885051042;
assign addr[2004] = -1875815927;
assign addr[2005] = -1866432072;
assign addr[2006] = -1856900221;
assign addr[2007] = -1847221128;
assign addr[2008] = -1837395562;
assign addr[2009] = -1827424302;
assign addr[2010] = -1817308138;
assign addr[2011] = -1807047873;
assign addr[2012] = -1796644320;
assign addr[2013] = -1786098304;
assign addr[2014] = -1775410662;
assign addr[2015] = -1764582240;
assign addr[2016] = -1753613897;
assign addr[2017] = -1742506504;
assign addr[2018] = -1731260941;
assign addr[2019] = -1719878099;
assign addr[2020] = -1708358881;
assign addr[2021] = -1696704201;
assign addr[2022] = -1684914983;
assign addr[2023] = -1672992161;
assign addr[2024] = -1660936681;
assign addr[2025] = -1648749499;
assign addr[2026] = -1636431582;
assign addr[2027] = -1623983905;
assign addr[2028] = -1611407456;
assign addr[2029] = -1598703233;
assign addr[2030] = -1585872242;
assign addr[2031] = -1572915501;
assign addr[2032] = -1559834037;
assign addr[2033] = -1546628888;
assign addr[2034] = -1533301101;
assign addr[2035] = -1519851733;
assign addr[2036] = -1506281850;
assign addr[2037] = -1492592527;
assign addr[2038] = -1478784851;
assign addr[2039] = -1464859917;
assign addr[2040] = -1450818828;
assign addr[2041] = -1436662698;
assign addr[2042] = -1422392650;
assign addr[2043] = -1408009814;
assign addr[2044] = -1393515332;
assign addr[2045] = -1378910353;
assign addr[2046] = -1364196034;
assign addr[2047] = -1349373543;
assign addr[2048] = -1334444055;
assign addr[2049] = -1319408754;
assign addr[2050] = -1304268832;
assign addr[2051] = -1289025489;
assign addr[2052] = -1273679934;
assign addr[2053] = -1258233384;
assign addr[2054] = -1242687064;
assign addr[2055] = -1227042207;
assign addr[2056] = -1211300053;
assign addr[2057] = -1195461849;
assign addr[2058] = -1179528853;
assign addr[2059] = -1163502328;
assign addr[2060] = -1147383544;
assign addr[2061] = -1131173780;
assign addr[2062] = -1114874320;
assign addr[2063] = -1098486458;
assign addr[2064] = -1082011492;
assign addr[2065] = -1065450729;
assign addr[2066] = -1048805483;
assign addr[2067] = -1032077073;
assign addr[2068] = -1015266825;
assign addr[2069] = -998376073;
assign addr[2070] = -981406156;
assign addr[2071] = -964358420;
assign addr[2072] = -947234215;
assign addr[2073] = -930034901;
assign addr[2074] = -912761841;
assign addr[2075] = -895416404;
assign addr[2076] = -877999966;
assign addr[2077] = -860513908;
assign addr[2078] = -842959617;
assign addr[2079] = -825338484;
assign addr[2080] = -807651907;
assign addr[2081] = -789901288;
assign addr[2082] = -772088034;
assign addr[2083] = -754213559;
assign addr[2084] = -736279279;
assign addr[2085] = -718286617;
assign addr[2086] = -700236999;
assign addr[2087] = -682131857;
assign addr[2088] = -663972625;
assign addr[2089] = -645760745;
assign addr[2090] = -627497660;
assign addr[2091] = -609184818;
assign addr[2092] = -590823671;
assign addr[2093] = -572415676;
assign addr[2094] = -553962291;
assign addr[2095] = -535464981;
assign addr[2096] = -516925212;
assign addr[2097] = -498344454;
assign addr[2098] = -479724180;
assign addr[2099] = -461065866;
assign addr[2100] = -442370993;
assign addr[2101] = -423641043;
assign addr[2102] = -404877501;
assign addr[2103] = -386081854;
assign addr[2104] = -367255594;
assign addr[2105] = -348400212;
assign addr[2106] = -329517204;
assign addr[2107] = -310608068;
assign addr[2108] = -291674302;
assign addr[2109] = -272717408;
assign addr[2110] = -253738890;
assign addr[2111] = -234740251;
assign addr[2112] = -215722999;
assign addr[2113] = -196688642;
assign addr[2114] = -177638688;
assign addr[2115] = -158574649;
assign addr[2116] = -139498035;
assign addr[2117] = -120410361;
assign addr[2118] = -101313138;
assign addr[2119] = -82207882;
assign addr[2120] = -63096108;
assign addr[2121] = -43979330;
assign addr[2122] = -24859065;
assign addr[2123] = -5736829;
assign addr[2124] = 13385863;
assign addr[2125] = 32507492;
assign addr[2126] = 51626544;
assign addr[2127] = 70741503;
assign addr[2128] = 89850852;
assign addr[2129] = 108953076;
assign addr[2130] = 128046661;
assign addr[2131] = 147130093;
assign addr[2132] = 166201858;
assign addr[2133] = 185260444;
assign addr[2134] = 204304341;
assign addr[2135] = 223332037;
assign addr[2136] = 242342025;
assign addr[2137] = 261332796;
assign addr[2138] = 280302845;
assign addr[2139] = 299250668;
assign addr[2140] = 318174762;
assign addr[2141] = 337073627;
assign addr[2142] = 355945764;
assign addr[2143] = 374789676;
assign addr[2144] = 393603870;
assign addr[2145] = 412386854;
assign addr[2146] = 431137138;
assign addr[2147] = 449853235;
assign addr[2148] = 468533662;
assign addr[2149] = 487176937;
assign addr[2150] = 505781581;
assign addr[2151] = 524346121;
assign addr[2152] = 542869083;
assign addr[2153] = 561348998;
assign addr[2154] = 579784402;
assign addr[2155] = 598173833;
assign addr[2156] = 616515832;
assign addr[2157] = 634808946;
assign addr[2158] = 653051723;
assign addr[2159] = 671242716;
assign addr[2160] = 689380485;
assign addr[2161] = 707463589;
assign addr[2162] = 725490597;
assign addr[2163] = 743460077;
assign addr[2164] = 761370605;
assign addr[2165] = 779220762;
assign addr[2166] = 797009130;
assign addr[2167] = 814734301;
assign addr[2168] = 832394869;
assign addr[2169] = 849989433;
assign addr[2170] = 867516597;
assign addr[2171] = 884974973;
assign addr[2172] = 902363176;
assign addr[2173] = 919679827;
assign addr[2174] = 936923553;
assign addr[2175] = 954092986;
assign addr[2176] = 971186766;
assign addr[2177] = 988203537;
assign addr[2178] = 1005141949;
assign addr[2179] = 1022000660;
assign addr[2180] = 1038778332;
assign addr[2181] = 1055473635;
assign addr[2182] = 1072085246;
assign addr[2183] = 1088611847;
assign addr[2184] = 1105052128;
assign addr[2185] = 1121404785;
assign addr[2186] = 1137668521;
assign addr[2187] = 1153842047;
assign addr[2188] = 1169924081;
assign addr[2189] = 1185913346;
assign addr[2190] = 1201808576;
assign addr[2191] = 1217608510;
assign addr[2192] = 1233311895;
assign addr[2193] = 1248917486;
assign addr[2194] = 1264424045;
assign addr[2195] = 1279830344;
assign addr[2196] = 1295135159;
assign addr[2197] = 1310337279;
assign addr[2198] = 1325435496;
assign addr[2199] = 1340428615;
assign addr[2200] = 1355315445;
assign addr[2201] = 1370094808;
assign addr[2202] = 1384765530;
assign addr[2203] = 1399326449;
assign addr[2204] = 1413776410;
assign addr[2205] = 1428114267;
assign addr[2206] = 1442338884;
assign addr[2207] = 1456449131;
assign addr[2208] = 1470443891;
assign addr[2209] = 1484322054;
assign addr[2210] = 1498082520;
assign addr[2211] = 1511724196;
assign addr[2212] = 1525246002;
assign addr[2213] = 1538646865;
assign addr[2214] = 1551925723;
assign addr[2215] = 1565081523;
assign addr[2216] = 1578113222;
assign addr[2217] = 1591019785;
assign addr[2218] = 1603800191;
assign addr[2219] = 1616453425;
assign addr[2220] = 1628978484;
assign addr[2221] = 1641374375;
assign addr[2222] = 1653640115;
assign addr[2223] = 1665774731;
assign addr[2224] = 1677777262;
assign addr[2225] = 1689646755;
assign addr[2226] = 1701382270;
assign addr[2227] = 1712982875;
assign addr[2228] = 1724447652;
assign addr[2229] = 1735775690;
assign addr[2230] = 1746966091;
assign addr[2231] = 1758017969;
assign addr[2232] = 1768930447;
assign addr[2233] = 1779702660;
assign addr[2234] = 1790333753;
assign addr[2235] = 1800822883;
assign addr[2236] = 1811169220;
assign addr[2237] = 1821371941;
assign addr[2238] = 1831430239;
assign addr[2239] = 1841343316;
assign addr[2240] = 1851110385;
assign addr[2241] = 1860730673;
assign addr[2242] = 1870203416;
assign addr[2243] = 1879527863;
assign addr[2244] = 1888703276;
assign addr[2245] = 1897728925;
assign addr[2246] = 1906604097;
assign addr[2247] = 1915328086;
assign addr[2248] = 1923900201;
assign addr[2249] = 1932319763;
assign addr[2250] = 1940586104;
assign addr[2251] = 1948698568;
assign addr[2252] = 1956656513;
assign addr[2253] = 1964459306;
assign addr[2254] = 1972106330;
assign addr[2255] = 1979596978;
assign addr[2256] = 1986930656;
assign addr[2257] = 1994106782;
assign addr[2258] = 2001124788;
assign addr[2259] = 2007984117;
assign addr[2260] = 2014684225;
assign addr[2261] = 2021224581;
assign addr[2262] = 2027604666;
assign addr[2263] = 2033823974;
assign addr[2264] = 2039882013;
assign addr[2265] = 2045778302;
assign addr[2266] = 2051512372;
assign addr[2267] = 2057083771;
assign addr[2268] = 2062492055;
assign addr[2269] = 2067736796;
assign addr[2270] = 2072817579;
assign addr[2271] = 2077733999;
assign addr[2272] = 2082485668;
assign addr[2273] = 2087072209;
assign addr[2274] = 2091493257;
assign addr[2275] = 2095748463;
assign addr[2276] = 2099837489;
assign addr[2277] = 2103760010;
assign addr[2278] = 2107515716;
assign addr[2279] = 2111104309;
assign addr[2280] = 2114525505;
assign addr[2281] = 2117779031;
assign addr[2282] = 2120864631;
assign addr[2283] = 2123782059;
assign addr[2284] = 2126531084;
assign addr[2285] = 2129111488;
assign addr[2286] = 2131523066;
assign addr[2287] = 2133765628;
assign addr[2288] = 2135838995;
assign addr[2289] = 2137743003;
assign addr[2290] = 2139477502;
assign addr[2291] = 2141042352;
assign addr[2292] = 2142437431;
assign addr[2293] = 2143662628;
assign addr[2294] = 2144717846;
assign addr[2295] = 2145603001;
assign addr[2296] = 2146318022;
assign addr[2297] = 2146862854;
assign addr[2298] = 2147237452;
assign addr[2299] = 2147441787;
assign addr[2300] = 2147475844;
assign addr[2301] = 2147339619;
assign addr[2302] = 2147033123;
assign addr[2303] = 2146556380;
assign addr[2304] = 2145909429;
assign addr[2305] = 2145092320;
assign addr[2306] = 2144105118;
assign addr[2307] = 2142947902;
assign addr[2308] = 2141620763;
assign addr[2309] = 2140123807;
assign addr[2310] = 2138457152;
assign addr[2311] = 2136620930;
assign addr[2312] = 2134615288;
assign addr[2313] = 2132440383;
assign addr[2314] = 2130096389;
assign addr[2315] = 2127583492;
assign addr[2316] = 2124901890;
assign addr[2317] = 2122051796;
assign addr[2318] = 2119033436;
assign addr[2319] = 2115847050;
assign addr[2320] = 2112492891;
assign addr[2321] = 2108971223;
assign addr[2322] = 2105282327;
assign addr[2323] = 2101426496;
assign addr[2324] = 2097404033;
assign addr[2325] = 2093215260;
assign addr[2326] = 2088860507;
assign addr[2327] = 2084340120;
assign addr[2328] = 2079654458;
assign addr[2329] = 2074803892;
assign addr[2330] = 2069788807;
assign addr[2331] = 2064609600;
assign addr[2332] = 2059266683;
assign addr[2333] = 2053760478;
assign addr[2334] = 2048091422;
assign addr[2335] = 2042259965;
assign addr[2336] = 2036266570;
assign addr[2337] = 2030111710;
assign addr[2338] = 2023795876;
assign addr[2339] = 2017319567;
assign addr[2340] = 2010683297;
assign addr[2341] = 2003887591;
assign addr[2342] = 1996932990;
assign addr[2343] = 1989820044;
assign addr[2344] = 1982549318;
assign addr[2345] = 1975121388;
assign addr[2346] = 1967536842;
assign addr[2347] = 1959796283;
assign addr[2348] = 1951900324;
assign addr[2349] = 1943849591;
assign addr[2350] = 1935644723;
assign addr[2351] = 1927286370;
assign addr[2352] = 1918775195;
assign addr[2353] = 1910111873;
assign addr[2354] = 1901297091;
assign addr[2355] = 1892331547;
assign addr[2356] = 1883215953;
assign addr[2357] = 1873951032;
assign addr[2358] = 1864537518;
assign addr[2359] = 1854976157;
assign addr[2360] = 1845267708;
assign addr[2361] = 1835412941;
assign addr[2362] = 1825412636;
assign addr[2363] = 1815267588;
assign addr[2364] = 1804978599;
assign addr[2365] = 1794546487;
assign addr[2366] = 1783972079;
assign addr[2367] = 1773256212;
assign addr[2368] = 1762399737;
assign addr[2369] = 1751403515;
assign addr[2370] = 1740268417;
assign addr[2371] = 1728995326;
assign addr[2372] = 1717585136;
assign addr[2373] = 1706038753;
assign addr[2374] = 1694357091;
assign addr[2375] = 1682541077;
assign addr[2376] = 1670591647;
assign addr[2377] = 1658509750;
assign addr[2378] = 1646296344;
assign addr[2379] = 1633952396;
assign addr[2380] = 1621478885;
assign addr[2381] = 1608876801;
assign addr[2382] = 1596147143;
assign addr[2383] = 1583290921;
assign addr[2384] = 1570309153;
assign addr[2385] = 1557202869;
assign addr[2386] = 1543973108;
assign addr[2387] = 1530620920;
assign addr[2388] = 1517147363;
assign addr[2389] = 1503553506;
assign addr[2390] = 1489840425;
assign addr[2391] = 1476009210;
assign addr[2392] = 1462060956;
assign addr[2393] = 1447996770;
assign addr[2394] = 1433817766;
assign addr[2395] = 1419525069;
assign addr[2396] = 1405119813;
assign addr[2397] = 1390603139;
assign addr[2398] = 1375976199;
assign addr[2399] = 1361240152;
assign addr[2400] = 1346396168;
assign addr[2401] = 1331445422;
assign addr[2402] = 1316389101;
assign addr[2403] = 1301228398;
assign addr[2404] = 1285964516;
assign addr[2405] = 1270598665;
assign addr[2406] = 1255132063;
assign addr[2407] = 1239565936;
assign addr[2408] = 1223901520;
assign addr[2409] = 1208140056;
assign addr[2410] = 1192282793;
assign addr[2411] = 1176330990;
assign addr[2412] = 1160285911;
assign addr[2413] = 1144148829;
assign addr[2414] = 1127921022;
assign addr[2415] = 1111603778;
assign addr[2416] = 1095198391;
assign addr[2417] = 1078706161;
assign addr[2418] = 1062128397;
assign addr[2419] = 1045466412;
assign addr[2420] = 1028721528;
assign addr[2421] = 1011895073;
assign addr[2422] = 994988380;
assign addr[2423] = 978002791;
assign addr[2424] = 960939653;
assign addr[2425] = 943800318;
assign addr[2426] = 926586145;
assign addr[2427] = 909298500;
assign addr[2428] = 891938752;
assign addr[2429] = 874508280;
assign addr[2430] = 857008464;
assign addr[2431] = 839440693;
assign addr[2432] = 821806359;
assign addr[2433] = 804106861;
assign addr[2434] = 786343603;
assign addr[2435] = 768517992;
assign addr[2436] = 750631442;
assign addr[2437] = 732685372;
assign addr[2438] = 714681204;
assign addr[2439] = 696620367;
assign addr[2440] = 678504291;
assign addr[2441] = 660334415;
assign addr[2442] = 642112178;
assign addr[2443] = 623839025;
assign addr[2444] = 605516406;
assign addr[2445] = 587145773;
assign addr[2446] = 568728583;
assign addr[2447] = 550266296;
assign addr[2448] = 531760377;
assign addr[2449] = 513212292;
assign addr[2450] = 494623513;
assign addr[2451] = 475995513;
assign addr[2452] = 457329769;
assign addr[2453] = 438627762;
assign addr[2454] = 419890975;
assign addr[2455] = 401120892;
assign addr[2456] = 382319004;
assign addr[2457] = 363486799;
assign addr[2458] = 344625773;
assign addr[2459] = 325737419;
assign addr[2460] = 306823237;
assign addr[2461] = 287884725;
assign addr[2462] = 268923386;
assign addr[2463] = 249940723;
assign addr[2464] = 230938242;
assign addr[2465] = 211917448;
assign addr[2466] = 192879850;
assign addr[2467] = 173826959;
assign addr[2468] = 154760284;
assign addr[2469] = 135681337;
assign addr[2470] = 116591632;
assign addr[2471] = 97492681;
assign addr[2472] = 78386000;
assign addr[2473] = 59273104;
assign addr[2474] = 40155507;
assign addr[2475] = 21034727;
assign addr[2476] = 1912278;
assign addr[2477] = -17210322;
assign addr[2478] = -36331557;
assign addr[2479] = -55449912;
assign addr[2480] = -74563870;
assign addr[2481] = -93671915;
assign addr[2482] = -112772533;
assign addr[2483] = -131864208;
assign addr[2484] = -150945428;
assign addr[2485] = -170014678;
assign addr[2486] = -189070447;
assign addr[2487] = -208111224;
assign addr[2488] = -227135500;
assign addr[2489] = -246141764;
assign addr[2490] = -265128512;
assign addr[2491] = -284094236;
assign addr[2492] = -303037433;
assign addr[2493] = -321956601;
assign addr[2494] = -340850240;
assign addr[2495] = -359716852;
assign addr[2496] = -378554940;
assign addr[2497] = -397363011;
assign addr[2498] = -416139574;
assign addr[2499] = -434883140;
assign addr[2500] = -453592221;
assign addr[2501] = -472265336;
assign addr[2502] = -490901003;
assign addr[2503] = -509497745;
assign addr[2504] = -528054086;
assign addr[2505] = -546568556;
assign addr[2506] = -565039687;
assign addr[2507] = -583466013;
assign addr[2508] = -601846074;
assign addr[2509] = -620178412;
assign addr[2510] = -638461574;
assign addr[2511] = -656694110;
assign addr[2512] = -674874574;
assign addr[2513] = -693001525;
assign addr[2514] = -711073524;
assign addr[2515] = -729089140;
assign addr[2516] = -747046944;
assign addr[2517] = -764945512;
assign addr[2518] = -782783424;
assign addr[2519] = -800559266;
assign addr[2520] = -818271628;
assign addr[2521] = -835919107;
assign addr[2522] = -853500302;
assign addr[2523] = -871013820;
assign addr[2524] = -888458272;
assign addr[2525] = -905832274;
assign addr[2526] = -923134450;
assign addr[2527] = -940363427;
assign addr[2528] = -957517838;
assign addr[2529] = -974596324;
assign addr[2530] = -991597531;
assign addr[2531] = -1008520110;
assign addr[2532] = -1025362720;
assign addr[2533] = -1042124025;
assign addr[2534] = -1058802695;
assign addr[2535] = -1075397409;
assign addr[2536] = -1091906851;
assign addr[2537] = -1108329711;
assign addr[2538] = -1124664687;
assign addr[2539] = -1140910484;
assign addr[2540] = -1157065814;
assign addr[2541] = -1173129396;
assign addr[2542] = -1189099956;
assign addr[2543] = -1204976227;
assign addr[2544] = -1220756951;
assign addr[2545] = -1236440877;
assign addr[2546] = -1252026760;
assign addr[2547] = -1267513365;
assign addr[2548] = -1282899464;
assign addr[2549] = -1298183838;
assign addr[2550] = -1313365273;
assign addr[2551] = -1328442566;
assign addr[2552] = -1343414522;
assign addr[2553] = -1358279953;
assign addr[2554] = -1373037681;
assign addr[2555] = -1387686535;
assign addr[2556] = -1402225355;
assign addr[2557] = -1416652986;
assign addr[2558] = -1430968286;
assign addr[2559] = -1445170118;
assign addr[2560] = -1459257358;
assign addr[2561] = -1473228887;
assign addr[2562] = -1487083598;
assign addr[2563] = -1500820393;
assign addr[2564] = -1514438181;
assign addr[2565] = -1527935884;
assign addr[2566] = -1541312431;
assign addr[2567] = -1554566762;
assign addr[2568] = -1567697824;
assign addr[2569] = -1580704578;
assign addr[2570] = -1593585992;
assign addr[2571] = -1606341043;
assign addr[2572] = -1618968722;
assign addr[2573] = -1631468027;
assign addr[2574] = -1643837966;
assign addr[2575] = -1656077559;
assign addr[2576] = -1668185835;
assign addr[2577] = -1680161834;
assign addr[2578] = -1692004606;
assign addr[2579] = -1703713213;
assign addr[2580] = -1715286726;
assign addr[2581] = -1726724227;
assign addr[2582] = -1738024810;
assign addr[2583] = -1749187577;
assign addr[2584] = -1760211645;
assign addr[2585] = -1771096139;
assign addr[2586] = -1781840195;
assign addr[2587] = -1792442963;
assign addr[2588] = -1802903601;
assign addr[2589] = -1813221279;
assign addr[2590] = -1823395180;
assign addr[2591] = -1833424497;
assign addr[2592] = -1843308435;
assign addr[2593] = -1853046210;
assign addr[2594] = -1862637049;
assign addr[2595] = -1872080193;
assign addr[2596] = -1881374892;
assign addr[2597] = -1890520410;
assign addr[2598] = -1899516021;
assign addr[2599] = -1908361011;
assign addr[2600] = -1917054681;
assign addr[2601] = -1925596340;
assign addr[2602] = -1933985310;
assign addr[2603] = -1942220928;
assign addr[2604] = -1950302539;
assign addr[2605] = -1958229503;
assign addr[2606] = -1966001192;
assign addr[2607] = -1973616989;
assign addr[2608] = -1981076290;
assign addr[2609] = -1988378503;
assign addr[2610] = -1995523051;
assign addr[2611] = -2002509365;
assign addr[2612] = -2009336893;
assign addr[2613] = -2016005093;
assign addr[2614] = -2022513436;
assign addr[2615] = -2028861406;
assign addr[2616] = -2035048499;
assign addr[2617] = -2041074226;
assign addr[2618] = -2046938108;
assign addr[2619] = -2052639680;
assign addr[2620] = -2058178491;
assign addr[2621] = -2063554100;
assign addr[2622] = -2068766083;
assign addr[2623] = -2073814024;
assign addr[2624] = -2078697525;
assign addr[2625] = -2083416198;
assign addr[2626] = -2087969669;
assign addr[2627] = -2092357577;
assign addr[2628] = -2096579573;
assign addr[2629] = -2100635323;
assign addr[2630] = -2104524506;
assign addr[2631] = -2108246813;
assign addr[2632] = -2111801949;
assign addr[2633] = -2115189632;
assign addr[2634] = -2118409593;
assign addr[2635] = -2121461578;
assign addr[2636] = -2124345343;
assign addr[2637] = -2127060661;
assign addr[2638] = -2129607316;
assign addr[2639] = -2131985106;
assign addr[2640] = -2134193842;
assign addr[2641] = -2136233350;
assign addr[2642] = -2138103468;
assign addr[2643] = -2139804048;
assign addr[2644] = -2141334954;
assign addr[2645] = -2142696065;
assign addr[2646] = -2143887273;
assign addr[2647] = -2144908484;
assign addr[2648] = -2145759618;
assign addr[2649] = -2146440605;
assign addr[2650] = -2146951393;
assign addr[2651] = -2147291941;
assign addr[2652] = -2147462221;
assign addr[2653] = -2147462221;
assign addr[2654] = -2147291941;
assign addr[2655] = -2146951393;
assign addr[2656] = -2146440605;
assign addr[2657] = -2145759618;
assign addr[2658] = -2144908484;
assign addr[2659] = -2143887273;
assign addr[2660] = -2142696065;
assign addr[2661] = -2141334954;
assign addr[2662] = -2139804048;
assign addr[2663] = -2138103468;
assign addr[2664] = -2136233350;
assign addr[2665] = -2134193842;
assign addr[2666] = -2131985106;
assign addr[2667] = -2129607316;
assign addr[2668] = -2127060661;
assign addr[2669] = -2124345343;
assign addr[2670] = -2121461578;
assign addr[2671] = -2118409593;
assign addr[2672] = -2115189632;
assign addr[2673] = -2111801949;
assign addr[2674] = -2108246813;
assign addr[2675] = -2104524506;
assign addr[2676] = -2100635323;
assign addr[2677] = -2096579573;
assign addr[2678] = -2092357577;
assign addr[2679] = -2087969669;
assign addr[2680] = -2083416198;
assign addr[2681] = -2078697525;
assign addr[2682] = -2073814024;
assign addr[2683] = -2068766083;
assign addr[2684] = -2063554100;
assign addr[2685] = -2058178491;
assign addr[2686] = -2052639680;
assign addr[2687] = -2046938108;
assign addr[2688] = -2041074226;
assign addr[2689] = -2035048499;
assign addr[2690] = -2028861406;
assign addr[2691] = -2022513436;
assign addr[2692] = -2016005093;
assign addr[2693] = -2009336893;
assign addr[2694] = -2002509365;
assign addr[2695] = -1995523051;
assign addr[2696] = -1988378503;
assign addr[2697] = -1981076290;
assign addr[2698] = -1973616989;
assign addr[2699] = -1966001192;
assign addr[2700] = -1958229503;
assign addr[2701] = -1950302539;
assign addr[2702] = -1942220928;
assign addr[2703] = -1933985310;
assign addr[2704] = -1925596340;
assign addr[2705] = -1917054681;
assign addr[2706] = -1908361011;
assign addr[2707] = -1899516021;
assign addr[2708] = -1890520410;
assign addr[2709] = -1881374892;
assign addr[2710] = -1872080193;
assign addr[2711] = -1862637049;
assign addr[2712] = -1853046210;
assign addr[2713] = -1843308435;
assign addr[2714] = -1833424497;
assign addr[2715] = -1823395180;
assign addr[2716] = -1813221279;
assign addr[2717] = -1802903601;
assign addr[2718] = -1792442963;
assign addr[2719] = -1781840195;
assign addr[2720] = -1771096139;
assign addr[2721] = -1760211645;
assign addr[2722] = -1749187577;
assign addr[2723] = -1738024810;
assign addr[2724] = -1726724227;
assign addr[2725] = -1715286726;
assign addr[2726] = -1703713213;
assign addr[2727] = -1692004606;
assign addr[2728] = -1680161834;
assign addr[2729] = -1668185835;
assign addr[2730] = -1656077559;
assign addr[2731] = -1643837966;
assign addr[2732] = -1631468027;
assign addr[2733] = -1618968722;
assign addr[2734] = -1606341043;
assign addr[2735] = -1593585992;
assign addr[2736] = -1580704578;
assign addr[2737] = -1567697824;
assign addr[2738] = -1554566762;
assign addr[2739] = -1541312431;
assign addr[2740] = -1527935884;
assign addr[2741] = -1514438181;
assign addr[2742] = -1500820393;
assign addr[2743] = -1487083598;
assign addr[2744] = -1473228887;
assign addr[2745] = -1459257358;
assign addr[2746] = -1445170118;
assign addr[2747] = -1430968286;
assign addr[2748] = -1416652986;
assign addr[2749] = -1402225355;
assign addr[2750] = -1387686535;
assign addr[2751] = -1373037681;
assign addr[2752] = -1358279953;
assign addr[2753] = -1343414522;
assign addr[2754] = -1328442566;
assign addr[2755] = -1313365273;
assign addr[2756] = -1298183838;
assign addr[2757] = -1282899464;
assign addr[2758] = -1267513365;
assign addr[2759] = -1252026760;
assign addr[2760] = -1236440877;
assign addr[2761] = -1220756951;
assign addr[2762] = -1204976227;
assign addr[2763] = -1189099956;
assign addr[2764] = -1173129396;
assign addr[2765] = -1157065814;
assign addr[2766] = -1140910484;
assign addr[2767] = -1124664687;
assign addr[2768] = -1108329711;
assign addr[2769] = -1091906851;
assign addr[2770] = -1075397409;
assign addr[2771] = -1058802695;
assign addr[2772] = -1042124025;
assign addr[2773] = -1025362720;
assign addr[2774] = -1008520110;
assign addr[2775] = -991597531;
assign addr[2776] = -974596324;
assign addr[2777] = -957517838;
assign addr[2778] = -940363427;
assign addr[2779] = -923134450;
assign addr[2780] = -905832274;
assign addr[2781] = -888458272;
assign addr[2782] = -871013820;
assign addr[2783] = -853500302;
assign addr[2784] = -835919107;
assign addr[2785] = -818271628;
assign addr[2786] = -800559266;
assign addr[2787] = -782783424;
assign addr[2788] = -764945512;
assign addr[2789] = -747046944;
assign addr[2790] = -729089140;
assign addr[2791] = -711073524;
assign addr[2792] = -693001525;
assign addr[2793] = -674874574;
assign addr[2794] = -656694110;
assign addr[2795] = -638461574;
assign addr[2796] = -620178412;
assign addr[2797] = -601846074;
assign addr[2798] = -583466013;
assign addr[2799] = -565039687;
assign addr[2800] = -546568556;
assign addr[2801] = -528054086;
assign addr[2802] = -509497745;
assign addr[2803] = -490901003;
assign addr[2804] = -472265336;
assign addr[2805] = -453592221;
assign addr[2806] = -434883140;
assign addr[2807] = -416139574;
assign addr[2808] = -397363011;
assign addr[2809] = -378554940;
assign addr[2810] = -359716852;
assign addr[2811] = -340850240;
assign addr[2812] = -321956601;
assign addr[2813] = -303037433;
assign addr[2814] = -284094236;
assign addr[2815] = -265128512;
assign addr[2816] = -246141764;
assign addr[2817] = -227135500;
assign addr[2818] = -208111224;
assign addr[2819] = -189070447;
assign addr[2820] = -170014678;
assign addr[2821] = -150945428;
assign addr[2822] = -131864208;
assign addr[2823] = -112772533;
assign addr[2824] = -93671915;
assign addr[2825] = -74563870;
assign addr[2826] = -55449912;
assign addr[2827] = -36331557;
assign addr[2828] = -17210322;
assign addr[2829] = 1912278;
assign addr[2830] = 21034727;
assign addr[2831] = 40155507;
assign addr[2832] = 59273104;
assign addr[2833] = 78386000;
assign addr[2834] = 97492681;
assign addr[2835] = 116591632;
assign addr[2836] = 135681337;
assign addr[2837] = 154760284;
assign addr[2838] = 173826959;
assign addr[2839] = 192879850;
assign addr[2840] = 211917448;
assign addr[2841] = 230938242;
assign addr[2842] = 249940723;
assign addr[2843] = 268923386;
assign addr[2844] = 287884725;
assign addr[2845] = 306823237;
assign addr[2846] = 325737419;
assign addr[2847] = 344625773;
assign addr[2848] = 363486799;
assign addr[2849] = 382319004;
assign addr[2850] = 401120892;
assign addr[2851] = 419890975;
assign addr[2852] = 438627762;
assign addr[2853] = 457329769;
assign addr[2854] = 475995513;
assign addr[2855] = 494623513;
assign addr[2856] = 513212292;
assign addr[2857] = 531760377;
assign addr[2858] = 550266296;
assign addr[2859] = 568728583;
assign addr[2860] = 587145773;
assign addr[2861] = 605516406;
assign addr[2862] = 623839025;
assign addr[2863] = 642112178;
assign addr[2864] = 660334415;
assign addr[2865] = 678504291;
assign addr[2866] = 696620367;
assign addr[2867] = 714681204;
assign addr[2868] = 732685372;
assign addr[2869] = 750631442;
assign addr[2870] = 768517992;
assign addr[2871] = 786343603;
assign addr[2872] = 804106861;
assign addr[2873] = 821806359;
assign addr[2874] = 839440693;
assign addr[2875] = 857008464;
assign addr[2876] = 874508280;
assign addr[2877] = 891938752;
assign addr[2878] = 909298500;
assign addr[2879] = 926586145;
assign addr[2880] = 943800318;
assign addr[2881] = 960939653;
assign addr[2882] = 978002791;
assign addr[2883] = 994988380;
assign addr[2884] = 1011895073;
assign addr[2885] = 1028721528;
assign addr[2886] = 1045466412;
assign addr[2887] = 1062128397;
assign addr[2888] = 1078706161;
assign addr[2889] = 1095198391;
assign addr[2890] = 1111603778;
assign addr[2891] = 1127921022;
assign addr[2892] = 1144148829;
assign addr[2893] = 1160285911;
assign addr[2894] = 1176330990;
assign addr[2895] = 1192282793;
assign addr[2896] = 1208140056;
assign addr[2897] = 1223901520;
assign addr[2898] = 1239565936;
assign addr[2899] = 1255132063;
assign addr[2900] = 1270598665;
assign addr[2901] = 1285964516;
assign addr[2902] = 1301228398;
assign addr[2903] = 1316389101;
assign addr[2904] = 1331445422;
assign addr[2905] = 1346396168;
assign addr[2906] = 1361240152;
assign addr[2907] = 1375976199;
assign addr[2908] = 1390603139;
assign addr[2909] = 1405119813;
assign addr[2910] = 1419525069;
assign addr[2911] = 1433817766;
assign addr[2912] = 1447996770;
assign addr[2913] = 1462060956;
assign addr[2914] = 1476009210;
assign addr[2915] = 1489840425;
assign addr[2916] = 1503553506;
assign addr[2917] = 1517147363;
assign addr[2918] = 1530620920;
assign addr[2919] = 1543973108;
assign addr[2920] = 1557202869;
assign addr[2921] = 1570309153;
assign addr[2922] = 1583290921;
assign addr[2923] = 1596147143;
assign addr[2924] = 1608876801;
assign addr[2925] = 1621478885;
assign addr[2926] = 1633952396;
assign addr[2927] = 1646296344;
assign addr[2928] = 1658509750;
assign addr[2929] = 1670591647;
assign addr[2930] = 1682541077;
assign addr[2931] = 1694357091;
assign addr[2932] = 1706038753;
assign addr[2933] = 1717585136;
assign addr[2934] = 1728995326;
assign addr[2935] = 1740268417;
assign addr[2936] = 1751403515;
assign addr[2937] = 1762399737;
assign addr[2938] = 1773256212;
assign addr[2939] = 1783972079;
assign addr[2940] = 1794546487;
assign addr[2941] = 1804978599;
assign addr[2942] = 1815267588;
assign addr[2943] = 1825412636;
assign addr[2944] = 1835412941;
assign addr[2945] = 1845267708;
assign addr[2946] = 1854976157;
assign addr[2947] = 1864537518;
assign addr[2948] = 1873951032;
assign addr[2949] = 1883215953;
assign addr[2950] = 1892331547;
assign addr[2951] = 1901297091;
assign addr[2952] = 1910111873;
assign addr[2953] = 1918775195;
assign addr[2954] = 1927286370;
assign addr[2955] = 1935644723;
assign addr[2956] = 1943849591;
assign addr[2957] = 1951900324;
assign addr[2958] = 1959796283;
assign addr[2959] = 1967536842;
assign addr[2960] = 1975121388;
assign addr[2961] = 1982549318;
assign addr[2962] = 1989820044;
assign addr[2963] = 1996932990;
assign addr[2964] = 2003887591;
assign addr[2965] = 2010683297;
assign addr[2966] = 2017319567;
assign addr[2967] = 2023795876;
assign addr[2968] = 2030111710;
assign addr[2969] = 2036266570;
assign addr[2970] = 2042259965;
assign addr[2971] = 2048091422;
assign addr[2972] = 2053760478;
assign addr[2973] = 2059266683;
assign addr[2974] = 2064609600;
assign addr[2975] = 2069788807;
assign addr[2976] = 2074803892;
assign addr[2977] = 2079654458;
assign addr[2978] = 2084340120;
assign addr[2979] = 2088860507;
assign addr[2980] = 2093215260;
assign addr[2981] = 2097404033;
assign addr[2982] = 2101426496;
assign addr[2983] = 2105282327;
assign addr[2984] = 2108971223;
assign addr[2985] = 2112492891;
assign addr[2986] = 2115847050;
assign addr[2987] = 2119033436;
assign addr[2988] = 2122051796;
assign addr[2989] = 2124901890;
assign addr[2990] = 2127583492;
assign addr[2991] = 2130096389;
assign addr[2992] = 2132440383;
assign addr[2993] = 2134615288;
assign addr[2994] = 2136620930;
assign addr[2995] = 2138457152;
assign addr[2996] = 2140123807;
assign addr[2997] = 2141620763;
assign addr[2998] = 2142947902;
assign addr[2999] = 2144105118;
assign addr[3000] = 2145092320;
assign addr[3001] = 2145909429;
assign addr[3002] = 2146556380;
assign addr[3003] = 2147033123;
assign addr[3004] = 2147339619;
assign addr[3005] = 2147475844;
assign addr[3006] = 2147441787;
assign addr[3007] = 2147237452;
assign addr[3008] = 2146862854;
assign addr[3009] = 2146318022;
assign addr[3010] = 2145603001;
assign addr[3011] = 2144717846;
assign addr[3012] = 2143662628;
assign addr[3013] = 2142437431;
assign addr[3014] = 2141042352;
assign addr[3015] = 2139477502;
assign addr[3016] = 2137743003;
assign addr[3017] = 2135838995;
assign addr[3018] = 2133765628;
assign addr[3019] = 2131523066;
assign addr[3020] = 2129111488;
assign addr[3021] = 2126531084;
assign addr[3022] = 2123782059;
assign addr[3023] = 2120864631;
assign addr[3024] = 2117779031;
assign addr[3025] = 2114525505;
assign addr[3026] = 2111104309;
assign addr[3027] = 2107515716;
assign addr[3028] = 2103760010;
assign addr[3029] = 2099837489;
assign addr[3030] = 2095748463;
assign addr[3031] = 2091493257;
assign addr[3032] = 2087072209;
assign addr[3033] = 2082485668;
assign addr[3034] = 2077733999;
assign addr[3035] = 2072817579;
assign addr[3036] = 2067736796;
assign addr[3037] = 2062492055;
assign addr[3038] = 2057083771;
assign addr[3039] = 2051512372;
assign addr[3040] = 2045778302;
assign addr[3041] = 2039882013;
assign addr[3042] = 2033823974;
assign addr[3043] = 2027604666;
assign addr[3044] = 2021224581;
assign addr[3045] = 2014684225;
assign addr[3046] = 2007984117;
assign addr[3047] = 2001124788;
assign addr[3048] = 1994106782;
assign addr[3049] = 1986930656;
assign addr[3050] = 1979596978;
assign addr[3051] = 1972106330;
assign addr[3052] = 1964459306;
assign addr[3053] = 1956656513;
assign addr[3054] = 1948698568;
assign addr[3055] = 1940586104;
assign addr[3056] = 1932319763;
assign addr[3057] = 1923900201;
assign addr[3058] = 1915328086;
assign addr[3059] = 1906604097;
assign addr[3060] = 1897728925;
assign addr[3061] = 1888703276;
assign addr[3062] = 1879527863;
assign addr[3063] = 1870203416;
assign addr[3064] = 1860730673;
assign addr[3065] = 1851110385;
assign addr[3066] = 1841343316;
assign addr[3067] = 1831430239;
assign addr[3068] = 1821371941;
assign addr[3069] = 1811169220;
assign addr[3070] = 1800822883;
assign addr[3071] = 1790333753;
assign addr[3072] = 1779702660;
assign addr[3073] = 1768930447;
assign addr[3074] = 1758017969;
assign addr[3075] = 1746966091;
assign addr[3076] = 1735775690;
assign addr[3077] = 1724447652;
assign addr[3078] = 1712982875;
assign addr[3079] = 1701382270;
assign addr[3080] = 1689646755;
assign addr[3081] = 1677777262;
assign addr[3082] = 1665774731;
assign addr[3083] = 1653640115;
assign addr[3084] = 1641374375;
assign addr[3085] = 1628978484;
assign addr[3086] = 1616453425;
assign addr[3087] = 1603800191;
assign addr[3088] = 1591019785;
assign addr[3089] = 1578113222;
assign addr[3090] = 1565081523;
assign addr[3091] = 1551925723;
assign addr[3092] = 1538646865;
assign addr[3093] = 1525246002;
assign addr[3094] = 1511724196;
assign addr[3095] = 1498082520;
assign addr[3096] = 1484322054;
assign addr[3097] = 1470443891;
assign addr[3098] = 1456449131;
assign addr[3099] = 1442338884;
assign addr[3100] = 1428114267;
assign addr[3101] = 1413776410;
assign addr[3102] = 1399326449;
assign addr[3103] = 1384765530;
assign addr[3104] = 1370094808;
assign addr[3105] = 1355315445;
assign addr[3106] = 1340428615;
assign addr[3107] = 1325435496;
assign addr[3108] = 1310337279;
assign addr[3109] = 1295135159;
assign addr[3110] = 1279830344;
assign addr[3111] = 1264424045;
assign addr[3112] = 1248917486;
assign addr[3113] = 1233311895;
assign addr[3114] = 1217608510;
assign addr[3115] = 1201808576;
assign addr[3116] = 1185913346;
assign addr[3117] = 1169924081;
assign addr[3118] = 1153842047;
assign addr[3119] = 1137668521;
assign addr[3120] = 1121404785;
assign addr[3121] = 1105052128;
assign addr[3122] = 1088611847;
assign addr[3123] = 1072085246;
assign addr[3124] = 1055473635;
assign addr[3125] = 1038778332;
assign addr[3126] = 1022000660;
assign addr[3127] = 1005141949;
assign addr[3128] = 988203537;
assign addr[3129] = 971186766;
assign addr[3130] = 954092986;
assign addr[3131] = 936923553;
assign addr[3132] = 919679827;
assign addr[3133] = 902363176;
assign addr[3134] = 884974973;
assign addr[3135] = 867516597;
assign addr[3136] = 849989433;
assign addr[3137] = 832394869;
assign addr[3138] = 814734301;
assign addr[3139] = 797009130;
assign addr[3140] = 779220762;
assign addr[3141] = 761370605;
assign addr[3142] = 743460077;
assign addr[3143] = 725490597;
assign addr[3144] = 707463589;
assign addr[3145] = 689380485;
assign addr[3146] = 671242716;
assign addr[3147] = 653051723;
assign addr[3148] = 634808946;
assign addr[3149] = 616515832;
assign addr[3150] = 598173833;
assign addr[3151] = 579784402;
assign addr[3152] = 561348998;
assign addr[3153] = 542869083;
assign addr[3154] = 524346121;
assign addr[3155] = 505781581;
assign addr[3156] = 487176937;
assign addr[3157] = 468533662;
assign addr[3158] = 449853235;
assign addr[3159] = 431137138;
assign addr[3160] = 412386854;
assign addr[3161] = 393603870;
assign addr[3162] = 374789676;
assign addr[3163] = 355945764;
assign addr[3164] = 337073627;
assign addr[3165] = 318174762;
assign addr[3166] = 299250668;
assign addr[3167] = 280302845;
assign addr[3168] = 261332796;
assign addr[3169] = 242342025;
assign addr[3170] = 223332037;
assign addr[3171] = 204304341;
assign addr[3172] = 185260444;
assign addr[3173] = 166201858;
assign addr[3174] = 147130093;
assign addr[3175] = 128046661;
assign addr[3176] = 108953076;
assign addr[3177] = 89850852;
assign addr[3178] = 70741503;
assign addr[3179] = 51626544;
assign addr[3180] = 32507492;
assign addr[3181] = 13385863;
assign addr[3182] = -5736829;
assign addr[3183] = -24859065;
assign addr[3184] = -43979330;
assign addr[3185] = -63096108;
assign addr[3186] = -82207882;
assign addr[3187] = -101313138;
assign addr[3188] = -120410361;
assign addr[3189] = -139498035;
assign addr[3190] = -158574649;
assign addr[3191] = -177638688;
assign addr[3192] = -196688642;
assign addr[3193] = -215722999;
assign addr[3194] = -234740251;
assign addr[3195] = -253738890;
assign addr[3196] = -272717408;
assign addr[3197] = -291674302;
assign addr[3198] = -310608068;
assign addr[3199] = -329517204;
assign addr[3200] = -348400212;
assign addr[3201] = -367255594;
assign addr[3202] = -386081854;
assign addr[3203] = -404877501;
assign addr[3204] = -423641043;
assign addr[3205] = -442370993;
assign addr[3206] = -461065866;
assign addr[3207] = -479724180;
assign addr[3208] = -498344454;
assign addr[3209] = -516925212;
assign addr[3210] = -535464981;
assign addr[3211] = -553962291;
assign addr[3212] = -572415676;
assign addr[3213] = -590823671;
assign addr[3214] = -609184818;
assign addr[3215] = -627497660;
assign addr[3216] = -645760745;
assign addr[3217] = -663972625;
assign addr[3218] = -682131857;
assign addr[3219] = -700236999;
assign addr[3220] = -718286617;
assign addr[3221] = -736279279;
assign addr[3222] = -754213559;
assign addr[3223] = -772088034;
assign addr[3224] = -789901288;
assign addr[3225] = -807651907;
assign addr[3226] = -825338484;
assign addr[3227] = -842959617;
assign addr[3228] = -860513908;
assign addr[3229] = -877999966;
assign addr[3230] = -895416404;
assign addr[3231] = -912761841;
assign addr[3232] = -930034901;
assign addr[3233] = -947234215;
assign addr[3234] = -964358420;
assign addr[3235] = -981406156;
assign addr[3236] = -998376073;
assign addr[3237] = -1015266825;
assign addr[3238] = -1032077073;
assign addr[3239] = -1048805483;
assign addr[3240] = -1065450729;
assign addr[3241] = -1082011492;
assign addr[3242] = -1098486458;
assign addr[3243] = -1114874320;
assign addr[3244] = -1131173780;
assign addr[3245] = -1147383544;
assign addr[3246] = -1163502328;
assign addr[3247] = -1179528853;
assign addr[3248] = -1195461849;
assign addr[3249] = -1211300053;
assign addr[3250] = -1227042207;
assign addr[3251] = -1242687064;
assign addr[3252] = -1258233384;
assign addr[3253] = -1273679934;
assign addr[3254] = -1289025489;
assign addr[3255] = -1304268832;
assign addr[3256] = -1319408754;
assign addr[3257] = -1334444055;
assign addr[3258] = -1349373543;
assign addr[3259] = -1364196034;
assign addr[3260] = -1378910353;
assign addr[3261] = -1393515332;
assign addr[3262] = -1408009814;
assign addr[3263] = -1422392650;
assign addr[3264] = -1436662698;
assign addr[3265] = -1450818828;
assign addr[3266] = -1464859917;
assign addr[3267] = -1478784851;
assign addr[3268] = -1492592527;
assign addr[3269] = -1506281850;
assign addr[3270] = -1519851733;
assign addr[3271] = -1533301101;
assign addr[3272] = -1546628888;
assign addr[3273] = -1559834037;
assign addr[3274] = -1572915501;
assign addr[3275] = -1585872242;
assign addr[3276] = -1598703233;
assign addr[3277] = -1611407456;
assign addr[3278] = -1623983905;
assign addr[3279] = -1636431582;
assign addr[3280] = -1648749499;
assign addr[3281] = -1660936681;
assign addr[3282] = -1672992161;
assign addr[3283] = -1684914983;
assign addr[3284] = -1696704201;
assign addr[3285] = -1708358881;
assign addr[3286] = -1719878099;
assign addr[3287] = -1731260941;
assign addr[3288] = -1742506504;
assign addr[3289] = -1753613897;
assign addr[3290] = -1764582240;
assign addr[3291] = -1775410662;
assign addr[3292] = -1786098304;
assign addr[3293] = -1796644320;
assign addr[3294] = -1807047873;
assign addr[3295] = -1817308138;
assign addr[3296] = -1827424302;
assign addr[3297] = -1837395562;
assign addr[3298] = -1847221128;
assign addr[3299] = -1856900221;
assign addr[3300] = -1866432072;
assign addr[3301] = -1875815927;
assign addr[3302] = -1885051042;
assign addr[3303] = -1894136683;
assign addr[3304] = -1903072131;
assign addr[3305] = -1911856677;
assign addr[3306] = -1920489624;
assign addr[3307] = -1928970288;
assign addr[3308] = -1937297997;
assign addr[3309] = -1945472089;
assign addr[3310] = -1953491918;
assign addr[3311] = -1961356847;
assign addr[3312] = -1969066252;
assign addr[3313] = -1976619522;
assign addr[3314] = -1984016058;
assign addr[3315] = -1991255274;
assign addr[3316] = -1998336596;
assign addr[3317] = -2005259462;
assign addr[3318] = -2012023322;
assign addr[3319] = -2018627642;
assign addr[3320] = -2025071897;
assign addr[3321] = -2031355576;
assign addr[3322] = -2037478181;
assign addr[3323] = -2043439226;
assign addr[3324] = -2049238240;
assign addr[3325] = -2054874761;
assign addr[3326] = -2060348343;
assign addr[3327] = -2065658552;
assign addr[3328] = -2070804967;
assign addr[3329] = -2075787180;
assign addr[3330] = -2080604795;
assign addr[3331] = -2085257431;
assign addr[3332] = -2089744719;
assign addr[3333] = -2094066304;
assign addr[3334] = -2098221841;
assign addr[3335] = -2102211002;
assign addr[3336] = -2106033471;
assign addr[3337] = -2109688944;
assign addr[3338] = -2113177132;
assign addr[3339] = -2116497758;
assign addr[3340] = -2119650558;
assign addr[3341] = -2122635283;
assign addr[3342] = -2125451696;
assign addr[3343] = -2128099574;
assign addr[3344] = -2130578706;
assign addr[3345] = -2132888897;
assign addr[3346] = -2135029962;
assign addr[3347] = -2137001733;
assign addr[3348] = -2138804053;
assign addr[3349] = -2140436778;
assign addr[3350] = -2141899780;
assign addr[3351] = -2143192942;
assign addr[3352] = -2144316162;
assign addr[3353] = -2145269351;
assign addr[3354] = -2146052433;
assign addr[3355] = -2146665347;
assign addr[3356] = -2147108043;
assign addr[3357] = -2147380486;
assign addr[3358] = -2147482655;
assign addr[3359] = -2147414542;
assign addr[3360] = -2147176152;
assign addr[3361] = -2146767505;
assign addr[3362] = -2146188631;
assign addr[3363] = -2145439578;
assign addr[3364] = -2144520405;
assign addr[3365] = -2143431184;
assign addr[3366] = -2142172003;
assign addr[3367] = -2140742960;
assign addr[3368] = -2139144169;
assign addr[3369] = -2137375758;
assign addr[3370] = -2135437865;
assign addr[3371] = -2133330646;
assign addr[3372] = -2131054266;
assign addr[3373] = -2128608907;
assign addr[3374] = -2125994762;
assign addr[3375] = -2123212038;
assign addr[3376] = -2120260957;
assign addr[3377] = -2117141752;
assign addr[3378] = -2113854671;
assign addr[3379] = -2110399974;
assign addr[3380] = -2106777935;
assign addr[3381] = -2102988841;
assign addr[3382] = -2099032994;
assign addr[3383] = -2094910706;
assign addr[3384] = -2090622304;
assign addr[3385] = -2086168128;
assign addr[3386] = -2081548533;
assign addr[3387] = -2076763883;
assign addr[3388] = -2071814558;
assign addr[3389] = -2066700952;
assign addr[3390] = -2061423468;
assign addr[3391] = -2055982526;
assign addr[3392] = -2050378558;
assign addr[3393] = -2044612007;
assign addr[3394] = -2038683330;
assign addr[3395] = -2032592999;
assign addr[3396] = -2026341495;
assign addr[3397] = -2019929315;
assign addr[3398] = -2013356967;
assign addr[3399] = -2006624971;
assign addr[3400] = -1999733863;
assign addr[3401] = -1992684188;
assign addr[3402] = -1985476506;
assign addr[3403] = -1978111387;
assign addr[3404] = -1970589416;
assign addr[3405] = -1962911189;
assign addr[3406] = -1955077316;
assign addr[3407] = -1947088417;
assign addr[3408] = -1938945125;
assign addr[3409] = -1930648088;
assign addr[3410] = -1922197961;
assign addr[3411] = -1913595416;
assign addr[3412] = -1904841135;
assign addr[3413] = -1895935811;
assign addr[3414] = -1886880151;
assign addr[3415] = -1877674873;
assign addr[3416] = -1868320707;
assign addr[3417] = -1858818395;
assign addr[3418] = -1849168689;
assign addr[3419] = -1839372356;
assign addr[3420] = -1829430172;
assign addr[3421] = -1819342925;
assign addr[3422] = -1809111415;
assign addr[3423] = -1798736454;
assign addr[3424] = -1788218865;
assign addr[3425] = -1777559480;
assign addr[3426] = -1766759146;
assign addr[3427] = -1755818718;
assign addr[3428] = -1744739065;
assign addr[3429] = -1733521064;
assign addr[3430] = -1722165606;
assign addr[3431] = -1710673591;
assign addr[3432] = -1699045930;
assign addr[3433] = -1687283545;
assign addr[3434] = -1675387369;
assign addr[3435] = -1663358344;
assign addr[3436] = -1651197426;
assign addr[3437] = -1638905577;
assign addr[3438] = -1626483774;
assign addr[3439] = -1613933000;
assign addr[3440] = -1601254251;
assign addr[3441] = -1588448533;
assign addr[3442] = -1575516860;
assign addr[3443] = -1562460258;
assign addr[3444] = -1549279763;
assign addr[3445] = -1535976419;
assign addr[3446] = -1522551282;
assign addr[3447] = -1509005416;
assign addr[3448] = -1495339895;
assign addr[3449] = -1481555802;
assign addr[3450] = -1467654232;
assign addr[3451] = -1453636285;
assign addr[3452] = -1439503074;
assign addr[3453] = -1425255719;
assign addr[3454] = -1410895350;
assign addr[3455] = -1396423105;
assign addr[3456] = -1381840133;
assign addr[3457] = -1367147589;
assign addr[3458] = -1352346639;
assign addr[3459] = -1337438456;
assign addr[3460] = -1322424222;
assign addr[3461] = -1307305128;
assign addr[3462] = -1292082373;
assign addr[3463] = -1276757164;
assign addr[3464] = -1261330715;
assign addr[3465] = -1245804251;
assign addr[3466] = -1230179002;
assign addr[3467] = -1214456207;
assign addr[3468] = -1198637114;
assign addr[3469] = -1182722976;
assign addr[3470] = -1166715055;
assign addr[3471] = -1150614620;
assign addr[3472] = -1134422949;
assign addr[3473] = -1118141326;
assign addr[3474] = -1101771040;
assign addr[3475] = -1085313391;
assign addr[3476] = -1068769683;
assign addr[3477] = -1052141228;
assign addr[3478] = -1035429345;
assign addr[3479] = -1018635358;
assign addr[3480] = -1001760600;
assign addr[3481] = -984806408;
assign addr[3482] = -967774128;
assign addr[3483] = -950665109;
assign addr[3484] = -933480707;
assign addr[3485] = -916222287;
assign addr[3486] = -898891215;
assign addr[3487] = -881488868;
assign addr[3488] = -864016623;
assign addr[3489] = -846475867;
assign addr[3490] = -828867991;
assign addr[3491] = -811194391;
assign addr[3492] = -793456467;
assign addr[3493] = -775655628;
assign addr[3494] = -757793284;
assign addr[3495] = -739870851;
assign addr[3496] = -721889752;
assign addr[3497] = -703851410;
assign addr[3498] = -685757258;
assign addr[3499] = -667608730;
assign addr[3500] = -649407264;
assign addr[3501] = -631154304;
assign addr[3502] = -612851297;
assign addr[3503] = -594499695;
assign addr[3504] = -576100953;
assign addr[3505] = -557656529;
assign addr[3506] = -539167887;
assign addr[3507] = -520636492;
assign addr[3508] = -502063814;
assign addr[3509] = -483451325;
assign addr[3510] = -464800501;
assign addr[3511] = -446112822;
assign addr[3512] = -427389768;
assign addr[3513] = -408632825;
assign addr[3514] = -389843480;
assign addr[3515] = -371023223;
assign addr[3516] = -352173546;
assign addr[3517] = -333295944;
assign addr[3518] = -314391913;
assign addr[3519] = -295462954;
assign addr[3520] = -276510565;
assign addr[3521] = -257536251;
assign addr[3522] = -238541516;
assign addr[3523] = -219527866;
assign addr[3524] = -200496809;
assign addr[3525] = -181449854;
assign addr[3526] = -162388511;
assign addr[3527] = -143314291;
assign addr[3528] = -124228708;
assign addr[3529] = -105133274;
assign addr[3530] = -86029503;
assign addr[3531] = -66918911;
assign addr[3532] = -47803013;
assign addr[3533] = -28683324;
assign addr[3534] = -9561361;
assign addr[3535] = 9561361;
assign addr[3536] = 28683324;
assign addr[3537] = 47803013;
assign addr[3538] = 66918911;
assign addr[3539] = 86029503;
assign addr[3540] = 105133274;
assign addr[3541] = 124228708;
assign addr[3542] = 143314291;
assign addr[3543] = 162388511;
assign addr[3544] = 181449854;
assign addr[3545] = 200496809;
assign addr[3546] = 219527866;
assign addr[3547] = 238541516;
assign addr[3548] = 257536251;
assign addr[3549] = 276510565;
assign addr[3550] = 295462954;
assign addr[3551] = 314391913;
assign addr[3552] = 333295944;
assign addr[3553] = 352173546;
assign addr[3554] = 371023223;
assign addr[3555] = 389843480;
assign addr[3556] = 408632825;
assign addr[3557] = 427389768;
assign addr[3558] = 446112822;
assign addr[3559] = 464800501;
assign addr[3560] = 483451325;
assign addr[3561] = 502063814;
assign addr[3562] = 520636492;
assign addr[3563] = 539167887;
assign addr[3564] = 557656529;
assign addr[3565] = 576100953;
assign addr[3566] = 594499695;
assign addr[3567] = 612851297;
assign addr[3568] = 631154304;
assign addr[3569] = 649407264;
assign addr[3570] = 667608730;
assign addr[3571] = 685757258;
assign addr[3572] = 703851410;
assign addr[3573] = 721889752;
assign addr[3574] = 739870851;
assign addr[3575] = 757793284;
assign addr[3576] = 775655628;
assign addr[3577] = 793456467;
assign addr[3578] = 811194391;
assign addr[3579] = 828867991;
assign addr[3580] = 846475867;
assign addr[3581] = 864016623;
assign addr[3582] = 881488868;
assign addr[3583] = 898891215;
assign addr[3584] = 916222287;
assign addr[3585] = 933480707;
assign addr[3586] = 950665109;
assign addr[3587] = 967774128;
assign addr[3588] = 984806408;
assign addr[3589] = 1001760600;
assign addr[3590] = 1018635358;
assign addr[3591] = 1035429345;
assign addr[3592] = 1052141228;
assign addr[3593] = 1068769683;
assign addr[3594] = 1085313391;
assign addr[3595] = 1101771040;
assign addr[3596] = 1118141326;
assign addr[3597] = 1134422949;
assign addr[3598] = 1150614620;
assign addr[3599] = 1166715055;
assign addr[3600] = 1182722976;
assign addr[3601] = 1198637114;
assign addr[3602] = 1214456207;
assign addr[3603] = 1230179002;
assign addr[3604] = 1245804251;
assign addr[3605] = 1261330715;
assign addr[3606] = 1276757164;
assign addr[3607] = 1292082373;
assign addr[3608] = 1307305128;
assign addr[3609] = 1322424222;
assign addr[3610] = 1337438456;
assign addr[3611] = 1352346639;
assign addr[3612] = 1367147589;
assign addr[3613] = 1381840133;
assign addr[3614] = 1396423105;
assign addr[3615] = 1410895350;
assign addr[3616] = 1425255719;
assign addr[3617] = 1439503074;
assign addr[3618] = 1453636285;
assign addr[3619] = 1467654232;
assign addr[3620] = 1481555802;
assign addr[3621] = 1495339895;
assign addr[3622] = 1509005416;
assign addr[3623] = 1522551282;
assign addr[3624] = 1535976419;
assign addr[3625] = 1549279763;
assign addr[3626] = 1562460258;
assign addr[3627] = 1575516860;
assign addr[3628] = 1588448533;
assign addr[3629] = 1601254251;
assign addr[3630] = 1613933000;
assign addr[3631] = 1626483774;
assign addr[3632] = 1638905577;
assign addr[3633] = 1651197426;
assign addr[3634] = 1663358344;
assign addr[3635] = 1675387369;
assign addr[3636] = 1687283545;
assign addr[3637] = 1699045930;
assign addr[3638] = 1710673591;
assign addr[3639] = 1722165606;
assign addr[3640] = 1733521064;
assign addr[3641] = 1744739065;
assign addr[3642] = 1755818718;
assign addr[3643] = 1766759146;
assign addr[3644] = 1777559480;
assign addr[3645] = 1788218865;
assign addr[3646] = 1798736454;
assign addr[3647] = 1809111415;
assign addr[3648] = 1819342925;
assign addr[3649] = 1829430172;
assign addr[3650] = 1839372356;
assign addr[3651] = 1849168689;
assign addr[3652] = 1858818395;
assign addr[3653] = 1868320707;
assign addr[3654] = 1877674873;
assign addr[3655] = 1886880151;
assign addr[3656] = 1895935811;
assign addr[3657] = 1904841135;
assign addr[3658] = 1913595416;
assign addr[3659] = 1922197961;
assign addr[3660] = 1930648088;
assign addr[3661] = 1938945125;
assign addr[3662] = 1947088417;
assign addr[3663] = 1955077316;
assign addr[3664] = 1962911189;
assign addr[3665] = 1970589416;
assign addr[3666] = 1978111387;
assign addr[3667] = 1985476506;
assign addr[3668] = 1992684188;
assign addr[3669] = 1999733863;
assign addr[3670] = 2006624971;
assign addr[3671] = 2013356967;
assign addr[3672] = 2019929315;
assign addr[3673] = 2026341495;
assign addr[3674] = 2032592999;
assign addr[3675] = 2038683330;
assign addr[3676] = 2044612007;
assign addr[3677] = 2050378558;
assign addr[3678] = 2055982526;
assign addr[3679] = 2061423468;
assign addr[3680] = 2066700952;
assign addr[3681] = 2071814558;
assign addr[3682] = 2076763883;
assign addr[3683] = 2081548533;
assign addr[3684] = 2086168128;
assign addr[3685] = 2090622304;
assign addr[3686] = 2094910706;
assign addr[3687] = 2099032994;
assign addr[3688] = 2102988841;
assign addr[3689] = 2106777935;
assign addr[3690] = 2110399974;
assign addr[3691] = 2113854671;
assign addr[3692] = 2117141752;
assign addr[3693] = 2120260957;
assign addr[3694] = 2123212038;
assign addr[3695] = 2125994762;
assign addr[3696] = 2128608907;
assign addr[3697] = 2131054266;
assign addr[3698] = 2133330646;
assign addr[3699] = 2135437865;
assign addr[3700] = 2137375758;
assign addr[3701] = 2139144169;
assign addr[3702] = 2140742960;
assign addr[3703] = 2142172003;
assign addr[3704] = 2143431184;
assign addr[3705] = 2144520405;
assign addr[3706] = 2145439578;
assign addr[3707] = 2146188631;
assign addr[3708] = 2146767505;
assign addr[3709] = 2147176152;
assign addr[3710] = 2147414542;
assign addr[3711] = 2147482655;
assign addr[3712] = 2147380486;
assign addr[3713] = 2147108043;
assign addr[3714] = 2146665347;
assign addr[3715] = 2146052433;
assign addr[3716] = 2145269351;
assign addr[3717] = 2144316162;
assign addr[3718] = 2143192942;
assign addr[3719] = 2141899780;
assign addr[3720] = 2140436778;
assign addr[3721] = 2138804053;
assign addr[3722] = 2137001733;
assign addr[3723] = 2135029962;
assign addr[3724] = 2132888897;
assign addr[3725] = 2130578706;
assign addr[3726] = 2128099574;
assign addr[3727] = 2125451696;
assign addr[3728] = 2122635283;
assign addr[3729] = 2119650558;
assign addr[3730] = 2116497758;
assign addr[3731] = 2113177132;
assign addr[3732] = 2109688944;
assign addr[3733] = 2106033471;
assign addr[3734] = 2102211002;
assign addr[3735] = 2098221841;
assign addr[3736] = 2094066304;
assign addr[3737] = 2089744719;
assign addr[3738] = 2085257431;
assign addr[3739] = 2080604795;
assign addr[3740] = 2075787180;
assign addr[3741] = 2070804967;
assign addr[3742] = 2065658552;
assign addr[3743] = 2060348343;
assign addr[3744] = 2054874761;
assign addr[3745] = 2049238240;
assign addr[3746] = 2043439226;
assign addr[3747] = 2037478181;
assign addr[3748] = 2031355576;
assign addr[3749] = 2025071897;
assign addr[3750] = 2018627642;
assign addr[3751] = 2012023322;
assign addr[3752] = 2005259462;
assign addr[3753] = 1998336596;
assign addr[3754] = 1991255274;
assign addr[3755] = 1984016058;
assign addr[3756] = 1976619522;
assign addr[3757] = 1969066252;
assign addr[3758] = 1961356847;
assign addr[3759] = 1953491918;
assign addr[3760] = 1945472089;
assign addr[3761] = 1937297997;
assign addr[3762] = 1928970288;
assign addr[3763] = 1920489624;
assign addr[3764] = 1911856677;
assign addr[3765] = 1903072131;
assign addr[3766] = 1894136683;
assign addr[3767] = 1885051042;
assign addr[3768] = 1875815927;
assign addr[3769] = 1866432072;
assign addr[3770] = 1856900221;
assign addr[3771] = 1847221128;
assign addr[3772] = 1837395562;
assign addr[3773] = 1827424302;
assign addr[3774] = 1817308138;
assign addr[3775] = 1807047873;
assign addr[3776] = 1796644320;
assign addr[3777] = 1786098304;
assign addr[3778] = 1775410662;
assign addr[3779] = 1764582240;
assign addr[3780] = 1753613897;
assign addr[3781] = 1742506504;
assign addr[3782] = 1731260941;
assign addr[3783] = 1719878099;
assign addr[3784] = 1708358881;
assign addr[3785] = 1696704201;
assign addr[3786] = 1684914983;
assign addr[3787] = 1672992161;
assign addr[3788] = 1660936681;
assign addr[3789] = 1648749499;
assign addr[3790] = 1636431582;
assign addr[3791] = 1623983905;
assign addr[3792] = 1611407456;
assign addr[3793] = 1598703233;
assign addr[3794] = 1585872242;
assign addr[3795] = 1572915501;
assign addr[3796] = 1559834037;
assign addr[3797] = 1546628888;
assign addr[3798] = 1533301101;
assign addr[3799] = 1519851733;
assign addr[3800] = 1506281850;
assign addr[3801] = 1492592527;
assign addr[3802] = 1478784851;
assign addr[3803] = 1464859917;
assign addr[3804] = 1450818828;
assign addr[3805] = 1436662698;
assign addr[3806] = 1422392650;
assign addr[3807] = 1408009814;
assign addr[3808] = 1393515332;
assign addr[3809] = 1378910353;
assign addr[3810] = 1364196034;
assign addr[3811] = 1349373543;
assign addr[3812] = 1334444055;
assign addr[3813] = 1319408754;
assign addr[3814] = 1304268832;
assign addr[3815] = 1289025489;
assign addr[3816] = 1273679934;
assign addr[3817] = 1258233384;
assign addr[3818] = 1242687064;
assign addr[3819] = 1227042207;
assign addr[3820] = 1211300053;
assign addr[3821] = 1195461849;
assign addr[3822] = 1179528853;
assign addr[3823] = 1163502328;
assign addr[3824] = 1147383544;
assign addr[3825] = 1131173780;
assign addr[3826] = 1114874320;
assign addr[3827] = 1098486458;
assign addr[3828] = 1082011492;
assign addr[3829] = 1065450729;
assign addr[3830] = 1048805483;
assign addr[3831] = 1032077073;
assign addr[3832] = 1015266825;
assign addr[3833] = 998376073;
assign addr[3834] = 981406156;
assign addr[3835] = 964358420;
assign addr[3836] = 947234215;
assign addr[3837] = 930034901;
assign addr[3838] = 912761841;
assign addr[3839] = 895416404;
assign addr[3840] = 877999966;
assign addr[3841] = 860513908;
assign addr[3842] = 842959617;
assign addr[3843] = 825338484;
assign addr[3844] = 807651907;
assign addr[3845] = 789901288;
assign addr[3846] = 772088034;
assign addr[3847] = 754213559;
assign addr[3848] = 736279279;
assign addr[3849] = 718286617;
assign addr[3850] = 700236999;
assign addr[3851] = 682131857;
assign addr[3852] = 663972625;
assign addr[3853] = 645760745;
assign addr[3854] = 627497660;
assign addr[3855] = 609184818;
assign addr[3856] = 590823671;
assign addr[3857] = 572415676;
assign addr[3858] = 553962291;
assign addr[3859] = 535464981;
assign addr[3860] = 516925212;
assign addr[3861] = 498344454;
assign addr[3862] = 479724180;
assign addr[3863] = 461065866;
assign addr[3864] = 442370993;
assign addr[3865] = 423641043;
assign addr[3866] = 404877501;
assign addr[3867] = 386081854;
assign addr[3868] = 367255594;
assign addr[3869] = 348400212;
assign addr[3870] = 329517204;
assign addr[3871] = 310608068;
assign addr[3872] = 291674302;
assign addr[3873] = 272717408;
assign addr[3874] = 253738890;
assign addr[3875] = 234740251;
assign addr[3876] = 215722999;
assign addr[3877] = 196688642;
assign addr[3878] = 177638688;
assign addr[3879] = 158574649;
assign addr[3880] = 139498035;
assign addr[3881] = 120410361;
assign addr[3882] = 101313138;
assign addr[3883] = 82207882;
assign addr[3884] = 63096108;
assign addr[3885] = 43979330;
assign addr[3886] = 24859065;
assign addr[3887] = 5736829;
assign addr[3888] = -13385863;
assign addr[3889] = -32507492;
assign addr[3890] = -51626544;
assign addr[3891] = -70741503;
assign addr[3892] = -89850852;
assign addr[3893] = -108953076;
assign addr[3894] = -128046661;
assign addr[3895] = -147130093;
assign addr[3896] = -166201858;
assign addr[3897] = -185260444;
assign addr[3898] = -204304341;
assign addr[3899] = -223332037;
assign addr[3900] = -242342025;
assign addr[3901] = -261332796;
assign addr[3902] = -280302845;
assign addr[3903] = -299250668;
assign addr[3904] = -318174762;
assign addr[3905] = -337073627;
assign addr[3906] = -355945764;
assign addr[3907] = -374789676;
assign addr[3908] = -393603870;
assign addr[3909] = -412386854;
assign addr[3910] = -431137138;
assign addr[3911] = -449853235;
assign addr[3912] = -468533662;
assign addr[3913] = -487176937;
assign addr[3914] = -505781581;
assign addr[3915] = -524346121;
assign addr[3916] = -542869083;
assign addr[3917] = -561348998;
assign addr[3918] = -579784402;
assign addr[3919] = -598173833;
assign addr[3920] = -616515832;
assign addr[3921] = -634808946;
assign addr[3922] = -653051723;
assign addr[3923] = -671242716;
assign addr[3924] = -689380485;
assign addr[3925] = -707463589;
assign addr[3926] = -725490597;
assign addr[3927] = -743460077;
assign addr[3928] = -761370605;
assign addr[3929] = -779220762;
assign addr[3930] = -797009130;
assign addr[3931] = -814734301;
assign addr[3932] = -832394869;
assign addr[3933] = -849989433;
assign addr[3934] = -867516597;
assign addr[3935] = -884974973;
assign addr[3936] = -902363176;
assign addr[3937] = -919679827;
assign addr[3938] = -936923553;
assign addr[3939] = -954092986;
assign addr[3940] = -971186766;
assign addr[3941] = -988203537;
assign addr[3942] = -1005141949;
assign addr[3943] = -1022000660;
assign addr[3944] = -1038778332;
assign addr[3945] = -1055473635;
assign addr[3946] = -1072085246;
assign addr[3947] = -1088611847;
assign addr[3948] = -1105052128;
assign addr[3949] = -1121404785;
assign addr[3950] = -1137668521;
assign addr[3951] = -1153842047;
assign addr[3952] = -1169924081;
assign addr[3953] = -1185913346;
assign addr[3954] = -1201808576;
assign addr[3955] = -1217608510;
assign addr[3956] = -1233311895;
assign addr[3957] = -1248917486;
assign addr[3958] = -1264424045;
assign addr[3959] = -1279830344;
assign addr[3960] = -1295135159;
assign addr[3961] = -1310337279;
assign addr[3962] = -1325435496;
assign addr[3963] = -1340428615;
assign addr[3964] = -1355315445;
assign addr[3965] = -1370094808;
assign addr[3966] = -1384765530;
assign addr[3967] = -1399326449;
assign addr[3968] = -1413776410;
assign addr[3969] = -1428114267;
assign addr[3970] = -1442338884;
assign addr[3971] = -1456449131;
assign addr[3972] = -1470443891;
assign addr[3973] = -1484322054;
assign addr[3974] = -1498082520;
assign addr[3975] = -1511724196;
assign addr[3976] = -1525246002;
assign addr[3977] = -1538646865;
assign addr[3978] = -1551925723;
assign addr[3979] = -1565081523;
assign addr[3980] = -1578113222;
assign addr[3981] = -1591019785;
assign addr[3982] = -1603800191;
assign addr[3983] = -1616453425;
assign addr[3984] = -1628978484;
assign addr[3985] = -1641374375;
assign addr[3986] = -1653640115;
assign addr[3987] = -1665774731;
assign addr[3988] = -1677777262;
assign addr[3989] = -1689646755;
assign addr[3990] = -1701382270;
assign addr[3991] = -1712982875;
assign addr[3992] = -1724447652;
assign addr[3993] = -1735775690;
assign addr[3994] = -1746966091;
assign addr[3995] = -1758017969;
assign addr[3996] = -1768930447;
assign addr[3997] = -1779702660;
assign addr[3998] = -1790333753;
assign addr[3999] = -1800822883;
assign addr[4000] = -1811169220;
assign addr[4001] = -1821371941;
assign addr[4002] = -1831430239;
assign addr[4003] = -1841343316;
assign addr[4004] = -1851110385;
assign addr[4005] = -1860730673;
assign addr[4006] = -1870203416;
assign addr[4007] = -1879527863;
assign addr[4008] = -1888703276;
assign addr[4009] = -1897728925;
assign addr[4010] = -1906604097;
assign addr[4011] = -1915328086;
assign addr[4012] = -1923900201;
assign addr[4013] = -1932319763;
assign addr[4014] = -1940586104;
assign addr[4015] = -1948698568;
assign addr[4016] = -1956656513;
assign addr[4017] = -1964459306;
assign addr[4018] = -1972106330;
assign addr[4019] = -1979596978;
assign addr[4020] = -1986930656;
assign addr[4021] = -1994106782;
assign addr[4022] = -2001124788;
assign addr[4023] = -2007984117;
assign addr[4024] = -2014684225;
assign addr[4025] = -2021224581;
assign addr[4026] = -2027604666;
assign addr[4027] = -2033823974;
assign addr[4028] = -2039882013;
assign addr[4029] = -2045778302;
assign addr[4030] = -2051512372;
assign addr[4031] = -2057083771;
assign addr[4032] = -2062492055;
assign addr[4033] = -2067736796;
assign addr[4034] = -2072817579;
assign addr[4035] = -2077733999;
assign addr[4036] = -2082485668;
assign addr[4037] = -2087072209;
assign addr[4038] = -2091493257;
assign addr[4039] = -2095748463;
assign addr[4040] = -2099837489;
assign addr[4041] = -2103760010;
assign addr[4042] = -2107515716;
assign addr[4043] = -2111104309;
assign addr[4044] = -2114525505;
assign addr[4045] = -2117779031;
assign addr[4046] = -2120864631;
assign addr[4047] = -2123782059;
assign addr[4048] = -2126531084;
assign addr[4049] = -2129111488;
assign addr[4050] = -2131523066;
assign addr[4051] = -2133765628;
assign addr[4052] = -2135838995;
assign addr[4053] = -2137743003;
assign addr[4054] = -2139477502;
assign addr[4055] = -2141042352;
assign addr[4056] = -2142437431;
assign addr[4057] = -2143662628;
assign addr[4058] = -2144717846;
assign addr[4059] = -2145603001;
assign addr[4060] = -2146318022;
assign addr[4061] = -2146862854;
assign addr[4062] = -2147237452;
assign addr[4063] = -2147441787;
assign addr[4064] = -2147475844;
assign addr[4065] = -2147339619;
assign addr[4066] = -2147033123;
assign addr[4067] = -2146556380;
assign addr[4068] = -2145909429;
assign addr[4069] = -2145092320;
assign addr[4070] = -2144105118;
assign addr[4071] = -2142947902;
assign addr[4072] = -2141620763;
assign addr[4073] = -2140123807;
assign addr[4074] = -2138457152;
assign addr[4075] = -2136620930;
assign addr[4076] = -2134615288;
assign addr[4077] = -2132440383;
assign addr[4078] = -2130096389;
assign addr[4079] = -2127583492;
assign addr[4080] = -2124901890;
assign addr[4081] = -2122051796;
assign addr[4082] = -2119033436;
assign addr[4083] = -2115847050;
assign addr[4084] = -2112492891;
assign addr[4085] = -2108971223;
assign addr[4086] = -2105282327;
assign addr[4087] = -2101426496;
assign addr[4088] = -2097404033;
assign addr[4089] = -2093215260;
assign addr[4090] = -2088860507;
assign addr[4091] = -2084340120;
assign addr[4092] = -2079654458;
assign addr[4093] = -2074803892;
assign addr[4094] = -2069788807;
assign addr[4095] = -2064609600;
assign addr[4096] = -2059266683;
assign addr[4097] = -2053760478;
assign addr[4098] = -2048091422;
assign addr[4099] = -2042259965;
assign addr[4100] = -2036266570;
assign addr[4101] = -2030111710;
assign addr[4102] = -2023795876;
assign addr[4103] = -2017319567;
assign addr[4104] = -2010683297;
assign addr[4105] = -2003887591;
assign addr[4106] = -1996932990;
assign addr[4107] = -1989820044;
assign addr[4108] = -1982549318;
assign addr[4109] = -1975121388;
assign addr[4110] = -1967536842;
assign addr[4111] = -1959796283;
assign addr[4112] = -1951900324;
assign addr[4113] = -1943849591;
assign addr[4114] = -1935644723;
assign addr[4115] = -1927286370;
assign addr[4116] = -1918775195;
assign addr[4117] = -1910111873;
assign addr[4118] = -1901297091;
assign addr[4119] = -1892331547;
assign addr[4120] = -1883215953;
assign addr[4121] = -1873951032;
assign addr[4122] = -1864537518;
assign addr[4123] = -1854976157;
assign addr[4124] = -1845267708;
assign addr[4125] = -1835412941;
assign addr[4126] = -1825412636;
assign addr[4127] = -1815267588;
assign addr[4128] = -1804978599;
assign addr[4129] = -1794546487;
assign addr[4130] = -1783972079;
assign addr[4131] = -1773256212;
assign addr[4132] = -1762399737;
assign addr[4133] = -1751403515;
assign addr[4134] = -1740268417;
assign addr[4135] = -1728995326;
assign addr[4136] = -1717585136;
assign addr[4137] = -1706038753;
assign addr[4138] = -1694357091;
assign addr[4139] = -1682541077;
assign addr[4140] = -1670591647;
assign addr[4141] = -1658509750;
assign addr[4142] = -1646296344;
assign addr[4143] = -1633952396;
assign addr[4144] = -1621478885;
assign addr[4145] = -1608876801;
assign addr[4146] = -1596147143;
assign addr[4147] = -1583290921;
assign addr[4148] = -1570309153;
assign addr[4149] = -1557202869;
assign addr[4150] = -1543973108;
assign addr[4151] = -1530620920;
assign addr[4152] = -1517147363;
assign addr[4153] = -1503553506;
assign addr[4154] = -1489840425;
assign addr[4155] = -1476009210;
assign addr[4156] = -1462060956;
assign addr[4157] = -1447996770;
assign addr[4158] = -1433817766;
assign addr[4159] = -1419525069;
assign addr[4160] = -1405119813;
assign addr[4161] = -1390603139;
assign addr[4162] = -1375976199;
assign addr[4163] = -1361240152;
assign addr[4164] = -1346396168;
assign addr[4165] = -1331445422;
assign addr[4166] = -1316389101;
assign addr[4167] = -1301228398;
assign addr[4168] = -1285964516;
assign addr[4169] = -1270598665;
assign addr[4170] = -1255132063;
assign addr[4171] = -1239565936;
assign addr[4172] = -1223901520;
assign addr[4173] = -1208140056;
assign addr[4174] = -1192282793;
assign addr[4175] = -1176330990;
assign addr[4176] = -1160285911;
assign addr[4177] = -1144148829;
assign addr[4178] = -1127921022;
assign addr[4179] = -1111603778;
assign addr[4180] = -1095198391;
assign addr[4181] = -1078706161;
assign addr[4182] = -1062128397;
assign addr[4183] = -1045466412;
assign addr[4184] = -1028721528;
assign addr[4185] = -1011895073;
assign addr[4186] = -994988380;
assign addr[4187] = -978002791;
assign addr[4188] = -960939653;
assign addr[4189] = -943800318;
assign addr[4190] = -926586145;
assign addr[4191] = -909298500;
assign addr[4192] = -891938752;
assign addr[4193] = -874508280;
assign addr[4194] = -857008464;
assign addr[4195] = -839440693;
assign addr[4196] = -821806359;
assign addr[4197] = -804106861;
assign addr[4198] = -786343603;
assign addr[4199] = -768517992;
assign addr[4200] = -750631442;
assign addr[4201] = -732685372;
assign addr[4202] = -714681204;
assign addr[4203] = -696620367;
assign addr[4204] = -678504291;
assign addr[4205] = -660334415;
assign addr[4206] = -642112178;
assign addr[4207] = -623839025;
assign addr[4208] = -605516406;
assign addr[4209] = -587145773;
assign addr[4210] = -568728583;
assign addr[4211] = -550266296;
assign addr[4212] = -531760377;
assign addr[4213] = -513212292;
assign addr[4214] = -494623513;
assign addr[4215] = -475995513;
assign addr[4216] = -457329769;
assign addr[4217] = -438627762;
assign addr[4218] = -419890975;
assign addr[4219] = -401120892;
assign addr[4220] = -382319004;
assign addr[4221] = -363486799;
assign addr[4222] = -344625773;
assign addr[4223] = -325737419;
assign addr[4224] = -306823237;
assign addr[4225] = -287884725;
assign addr[4226] = -268923386;
assign addr[4227] = -249940723;
assign addr[4228] = -230938242;
assign addr[4229] = -211917448;
assign addr[4230] = -192879850;
assign addr[4231] = -173826959;
assign addr[4232] = -154760284;
assign addr[4233] = -135681337;
assign addr[4234] = -116591632;
assign addr[4235] = -97492681;
assign addr[4236] = -78386000;
assign addr[4237] = -59273104;
assign addr[4238] = -40155507;
assign addr[4239] = -21034727;
assign addr[4240] = -1912278;
assign addr[4241] = 17210322;
assign addr[4242] = 36331557;
assign addr[4243] = 55449912;
assign addr[4244] = 74563870;
assign addr[4245] = 93671915;
assign addr[4246] = 112772533;
assign addr[4247] = 131864208;
assign addr[4248] = 150945428;
assign addr[4249] = 170014678;
assign addr[4250] = 189070447;
assign addr[4251] = 208111224;
assign addr[4252] = 227135500;
assign addr[4253] = 246141764;
assign addr[4254] = 265128512;
assign addr[4255] = 284094236;
assign addr[4256] = 303037433;
assign addr[4257] = 321956601;
assign addr[4258] = 340850240;
assign addr[4259] = 359716852;
assign addr[4260] = 378554940;
assign addr[4261] = 397363011;
assign addr[4262] = 416139574;
assign addr[4263] = 434883140;
assign addr[4264] = 453592221;
assign addr[4265] = 472265336;
assign addr[4266] = 490901003;
assign addr[4267] = 509497745;
assign addr[4268] = 528054086;
assign addr[4269] = 546568556;
assign addr[4270] = 565039687;
assign addr[4271] = 583466013;
assign addr[4272] = 601846074;
assign addr[4273] = 620178412;
assign addr[4274] = 638461574;
assign addr[4275] = 656694110;
assign addr[4276] = 674874574;
assign addr[4277] = 693001525;
assign addr[4278] = 711073524;
assign addr[4279] = 729089140;
assign addr[4280] = 747046944;
assign addr[4281] = 764945512;
assign addr[4282] = 782783424;
assign addr[4283] = 800559266;
assign addr[4284] = 818271628;
assign addr[4285] = 835919107;
assign addr[4286] = 853500302;
assign addr[4287] = 871013820;
assign addr[4288] = 888458272;
assign addr[4289] = 905832274;
assign addr[4290] = 923134450;
assign addr[4291] = 940363427;
assign addr[4292] = 957517838;
assign addr[4293] = 974596324;
assign addr[4294] = 991597531;
assign addr[4295] = 1008520110;
assign addr[4296] = 1025362720;
assign addr[4297] = 1042124025;
assign addr[4298] = 1058802695;
assign addr[4299] = 1075397409;
assign addr[4300] = 1091906851;
assign addr[4301] = 1108329711;
assign addr[4302] = 1124664687;
assign addr[4303] = 1140910484;
assign addr[4304] = 1157065814;
assign addr[4305] = 1173129396;
assign addr[4306] = 1189099956;
assign addr[4307] = 1204976227;
assign addr[4308] = 1220756951;
assign addr[4309] = 1236440877;
assign addr[4310] = 1252026760;
assign addr[4311] = 1267513365;
assign addr[4312] = 1282899464;
assign addr[4313] = 1298183838;
assign addr[4314] = 1313365273;
assign addr[4315] = 1328442566;
assign addr[4316] = 1343414522;
assign addr[4317] = 1358279953;
assign addr[4318] = 1373037681;
assign addr[4319] = 1387686535;
assign addr[4320] = 1402225355;
assign addr[4321] = 1416652986;
assign addr[4322] = 1430968286;
assign addr[4323] = 1445170118;
assign addr[4324] = 1459257358;
assign addr[4325] = 1473228887;
assign addr[4326] = 1487083598;
assign addr[4327] = 1500820393;
assign addr[4328] = 1514438181;
assign addr[4329] = 1527935884;
assign addr[4330] = 1541312431;
assign addr[4331] = 1554566762;
assign addr[4332] = 1567697824;
assign addr[4333] = 1580704578;
assign addr[4334] = 1593585992;
assign addr[4335] = 1606341043;
assign addr[4336] = 1618968722;
assign addr[4337] = 1631468027;
assign addr[4338] = 1643837966;
assign addr[4339] = 1656077559;
assign addr[4340] = 1668185835;
assign addr[4341] = 1680161834;
assign addr[4342] = 1692004606;
assign addr[4343] = 1703713213;
assign addr[4344] = 1715286726;
assign addr[4345] = 1726724227;
assign addr[4346] = 1738024810;
assign addr[4347] = 1749187577;
assign addr[4348] = 1760211645;
assign addr[4349] = 1771096139;
assign addr[4350] = 1781840195;
assign addr[4351] = 1792442963;
assign addr[4352] = 1802903601;
assign addr[4353] = 1813221279;
assign addr[4354] = 1823395180;
assign addr[4355] = 1833424497;
assign addr[4356] = 1843308435;
assign addr[4357] = 1853046210;
assign addr[4358] = 1862637049;
assign addr[4359] = 1872080193;
assign addr[4360] = 1881374892;
assign addr[4361] = 1890520410;
assign addr[4362] = 1899516021;
assign addr[4363] = 1908361011;
assign addr[4364] = 1917054681;
assign addr[4365] = 1925596340;
assign addr[4366] = 1933985310;
assign addr[4367] = 1942220928;
assign addr[4368] = 1950302539;
assign addr[4369] = 1958229503;
assign addr[4370] = 1966001192;
assign addr[4371] = 1973616989;
assign addr[4372] = 1981076290;
assign addr[4373] = 1988378503;
assign addr[4374] = 1995523051;
assign addr[4375] = 2002509365;
assign addr[4376] = 2009336893;
assign addr[4377] = 2016005093;
assign addr[4378] = 2022513436;
assign addr[4379] = 2028861406;
assign addr[4380] = 2035048499;
assign addr[4381] = 2041074226;
assign addr[4382] = 2046938108;
assign addr[4383] = 2052639680;
assign addr[4384] = 2058178491;
assign addr[4385] = 2063554100;
assign addr[4386] = 2068766083;
assign addr[4387] = 2073814024;
assign addr[4388] = 2078697525;
assign addr[4389] = 2083416198;
assign addr[4390] = 2087969669;
assign addr[4391] = 2092357577;
assign addr[4392] = 2096579573;
assign addr[4393] = 2100635323;
assign addr[4394] = 2104524506;
assign addr[4395] = 2108246813;
assign addr[4396] = 2111801949;
assign addr[4397] = 2115189632;
assign addr[4398] = 2118409593;
assign addr[4399] = 2121461578;
assign addr[4400] = 2124345343;
assign addr[4401] = 2127060661;
assign addr[4402] = 2129607316;
assign addr[4403] = 2131985106;
assign addr[4404] = 2134193842;
assign addr[4405] = 2136233350;
assign addr[4406] = 2138103468;
assign addr[4407] = 2139804048;
assign addr[4408] = 2141334954;
assign addr[4409] = 2142696065;
assign addr[4410] = 2143887273;
assign addr[4411] = 2144908484;
assign addr[4412] = 2145759618;
assign addr[4413] = 2146440605;
assign addr[4414] = 2146951393;
assign addr[4415] = 2147291941;
assign addr[4416] = 2147462221;
assign addr[4417] = 2147462221;
assign addr[4418] = 2147291941;
assign addr[4419] = 2146951393;
assign addr[4420] = 2146440605;
assign addr[4421] = 2145759618;
assign addr[4422] = 2144908484;
assign addr[4423] = 2143887273;
assign addr[4424] = 2142696065;
assign addr[4425] = 2141334954;
assign addr[4426] = 2139804048;
assign addr[4427] = 2138103468;
assign addr[4428] = 2136233350;
assign addr[4429] = 2134193842;
assign addr[4430] = 2131985106;
assign addr[4431] = 2129607316;
assign addr[4432] = 2127060661;
assign addr[4433] = 2124345343;
assign addr[4434] = 2121461578;
assign addr[4435] = 2118409593;
assign addr[4436] = 2115189632;
assign addr[4437] = 2111801949;
assign addr[4438] = 2108246813;
assign addr[4439] = 2104524506;
assign addr[4440] = 2100635323;
assign addr[4441] = 2096579573;
assign addr[4442] = 2092357577;
assign addr[4443] = 2087969669;
assign addr[4444] = 2083416198;
assign addr[4445] = 2078697525;
assign addr[4446] = 2073814024;
assign addr[4447] = 2068766083;
assign addr[4448] = 2063554100;
assign addr[4449] = 2058178491;
assign addr[4450] = 2052639680;
assign addr[4451] = 2046938108;
assign addr[4452] = 2041074226;
assign addr[4453] = 2035048499;
assign addr[4454] = 2028861406;
assign addr[4455] = 2022513436;
assign addr[4456] = 2016005093;
assign addr[4457] = 2009336893;
assign addr[4458] = 2002509365;
assign addr[4459] = 1995523051;
assign addr[4460] = 1988378503;
assign addr[4461] = 1981076290;
assign addr[4462] = 1973616989;
assign addr[4463] = 1966001192;
assign addr[4464] = 1958229503;
assign addr[4465] = 1950302539;
assign addr[4466] = 1942220928;
assign addr[4467] = 1933985310;
assign addr[4468] = 1925596340;
assign addr[4469] = 1917054681;
assign addr[4470] = 1908361011;
assign addr[4471] = 1899516021;
assign addr[4472] = 1890520410;
assign addr[4473] = 1881374892;
assign addr[4474] = 1872080193;
assign addr[4475] = 1862637049;
assign addr[4476] = 1853046210;
assign addr[4477] = 1843308435;
assign addr[4478] = 1833424497;
assign addr[4479] = 1823395180;
assign addr[4480] = 1813221279;
assign addr[4481] = 1802903601;
assign addr[4482] = 1792442963;
assign addr[4483] = 1781840195;
assign addr[4484] = 1771096139;
assign addr[4485] = 1760211645;
assign addr[4486] = 1749187577;
assign addr[4487] = 1738024810;
assign addr[4488] = 1726724227;
assign addr[4489] = 1715286726;
assign addr[4490] = 1703713213;
assign addr[4491] = 1692004606;
assign addr[4492] = 1680161834;
assign addr[4493] = 1668185835;
assign addr[4494] = 1656077559;
assign addr[4495] = 1643837966;
assign addr[4496] = 1631468027;
assign addr[4497] = 1618968722;
assign addr[4498] = 1606341043;
assign addr[4499] = 1593585992;
assign addr[4500] = 1580704578;
assign addr[4501] = 1567697824;
assign addr[4502] = 1554566762;
assign addr[4503] = 1541312431;
assign addr[4504] = 1527935884;
assign addr[4505] = 1514438181;
assign addr[4506] = 1500820393;
assign addr[4507] = 1487083598;
assign addr[4508] = 1473228887;
assign addr[4509] = 1459257358;
assign addr[4510] = 1445170118;
assign addr[4511] = 1430968286;
assign addr[4512] = 1416652986;
assign addr[4513] = 1402225355;
assign addr[4514] = 1387686535;
assign addr[4515] = 1373037681;
assign addr[4516] = 1358279953;
assign addr[4517] = 1343414522;
assign addr[4518] = 1328442566;
assign addr[4519] = 1313365273;
assign addr[4520] = 1298183838;
assign addr[4521] = 1282899464;
assign addr[4522] = 1267513365;
assign addr[4523] = 1252026760;
assign addr[4524] = 1236440877;
assign addr[4525] = 1220756951;
assign addr[4526] = 1204976227;
assign addr[4527] = 1189099956;
assign addr[4528] = 1173129396;
assign addr[4529] = 1157065814;
assign addr[4530] = 1140910484;
assign addr[4531] = 1124664687;
assign addr[4532] = 1108329711;
assign addr[4533] = 1091906851;
assign addr[4534] = 1075397409;
assign addr[4535] = 1058802695;
assign addr[4536] = 1042124025;
assign addr[4537] = 1025362720;
assign addr[4538] = 1008520110;
assign addr[4539] = 991597531;
assign addr[4540] = 974596324;
assign addr[4541] = 957517838;
assign addr[4542] = 940363427;
assign addr[4543] = 923134450;
assign addr[4544] = 905832274;
assign addr[4545] = 888458272;
assign addr[4546] = 871013820;
assign addr[4547] = 853500302;
assign addr[4548] = 835919107;
assign addr[4549] = 818271628;
assign addr[4550] = 800559266;
assign addr[4551] = 782783424;
assign addr[4552] = 764945512;
assign addr[4553] = 747046944;
assign addr[4554] = 729089140;
assign addr[4555] = 711073524;
assign addr[4556] = 693001525;
assign addr[4557] = 674874574;
assign addr[4558] = 656694110;
assign addr[4559] = 638461574;
assign addr[4560] = 620178412;
assign addr[4561] = 601846074;
assign addr[4562] = 583466013;
assign addr[4563] = 565039687;
assign addr[4564] = 546568556;
assign addr[4565] = 528054086;
assign addr[4566] = 509497745;
assign addr[4567] = 490901003;
assign addr[4568] = 472265336;
assign addr[4569] = 453592221;
assign addr[4570] = 434883140;
assign addr[4571] = 416139574;
assign addr[4572] = 397363011;
assign addr[4573] = 378554940;
assign addr[4574] = 359716852;
assign addr[4575] = 340850240;
assign addr[4576] = 321956601;
assign addr[4577] = 303037433;
assign addr[4578] = 284094236;
assign addr[4579] = 265128512;
assign addr[4580] = 246141764;
assign addr[4581] = 227135500;
assign addr[4582] = 208111224;
assign addr[4583] = 189070447;
assign addr[4584] = 170014678;
assign addr[4585] = 150945428;
assign addr[4586] = 131864208;
assign addr[4587] = 112772533;
assign addr[4588] = 93671915;
assign addr[4589] = 74563870;
assign addr[4590] = 55449912;
assign addr[4591] = 36331557;
assign addr[4592] = 17210322;
assign addr[4593] = -1912278;
assign addr[4594] = -21034727;
assign addr[4595] = -40155507;
assign addr[4596] = -59273104;
assign addr[4597] = -78386000;
assign addr[4598] = -97492681;
assign addr[4599] = -116591632;
assign addr[4600] = -135681337;
assign addr[4601] = -154760284;
assign addr[4602] = -173826959;
assign addr[4603] = -192879850;
assign addr[4604] = -211917448;
assign addr[4605] = -230938242;
assign addr[4606] = -249940723;
assign addr[4607] = -268923386;
assign addr[4608] = -287884725;
assign addr[4609] = -306823237;
assign addr[4610] = -325737419;
assign addr[4611] = -344625773;
assign addr[4612] = -363486799;
assign addr[4613] = -382319004;
assign addr[4614] = -401120892;
assign addr[4615] = -419890975;
assign addr[4616] = -438627762;
assign addr[4617] = -457329769;
assign addr[4618] = -475995513;
assign addr[4619] = -494623513;
assign addr[4620] = -513212292;
assign addr[4621] = -531760377;
assign addr[4622] = -550266296;
assign addr[4623] = -568728583;
assign addr[4624] = -587145773;
assign addr[4625] = -605516406;
assign addr[4626] = -623839025;
assign addr[4627] = -642112178;
assign addr[4628] = -660334415;
assign addr[4629] = -678504291;
assign addr[4630] = -696620367;
assign addr[4631] = -714681204;
assign addr[4632] = -732685372;
assign addr[4633] = -750631442;
assign addr[4634] = -768517992;
assign addr[4635] = -786343603;
assign addr[4636] = -804106861;
assign addr[4637] = -821806359;
assign addr[4638] = -839440693;
assign addr[4639] = -857008464;
assign addr[4640] = -874508280;
assign addr[4641] = -891938752;
assign addr[4642] = -909298500;
assign addr[4643] = -926586145;
assign addr[4644] = -943800318;
assign addr[4645] = -960939653;
assign addr[4646] = -978002791;
assign addr[4647] = -994988380;
assign addr[4648] = -1011895073;
assign addr[4649] = -1028721528;
assign addr[4650] = -1045466412;
assign addr[4651] = -1062128397;
assign addr[4652] = -1078706161;
assign addr[4653] = -1095198391;
assign addr[4654] = -1111603778;
assign addr[4655] = -1127921022;
assign addr[4656] = -1144148829;
assign addr[4657] = -1160285911;
assign addr[4658] = -1176330990;
assign addr[4659] = -1192282793;
assign addr[4660] = -1208140056;
assign addr[4661] = -1223901520;
assign addr[4662] = -1239565936;
assign addr[4663] = -1255132063;
assign addr[4664] = -1270598665;
assign addr[4665] = -1285964516;
assign addr[4666] = -1301228398;
assign addr[4667] = -1316389101;
assign addr[4668] = -1331445422;
assign addr[4669] = -1346396168;
assign addr[4670] = -1361240152;
assign addr[4671] = -1375976199;
assign addr[4672] = -1390603139;
assign addr[4673] = -1405119813;
assign addr[4674] = -1419525069;
assign addr[4675] = -1433817766;
assign addr[4676] = -1447996770;
assign addr[4677] = -1462060956;
assign addr[4678] = -1476009210;
assign addr[4679] = -1489840425;
assign addr[4680] = -1503553506;
assign addr[4681] = -1517147363;
assign addr[4682] = -1530620920;
assign addr[4683] = -1543973108;
assign addr[4684] = -1557202869;
assign addr[4685] = -1570309153;
assign addr[4686] = -1583290921;
assign addr[4687] = -1596147143;
assign addr[4688] = -1608876801;
assign addr[4689] = -1621478885;
assign addr[4690] = -1633952396;
assign addr[4691] = -1646296344;
assign addr[4692] = -1658509750;
assign addr[4693] = -1670591647;
assign addr[4694] = -1682541077;
assign addr[4695] = -1694357091;
assign addr[4696] = -1706038753;
assign addr[4697] = -1717585136;
assign addr[4698] = -1728995326;
assign addr[4699] = -1740268417;
assign addr[4700] = -1751403515;
assign addr[4701] = -1762399737;
assign addr[4702] = -1773256212;
assign addr[4703] = -1783972079;
assign addr[4704] = -1794546487;
assign addr[4705] = -1804978599;
assign addr[4706] = -1815267588;
assign addr[4707] = -1825412636;
assign addr[4708] = -1835412941;
assign addr[4709] = -1845267708;
assign addr[4710] = -1854976157;
assign addr[4711] = -1864537518;
assign addr[4712] = -1873951032;
assign addr[4713] = -1883215953;
assign addr[4714] = -1892331547;
assign addr[4715] = -1901297091;
assign addr[4716] = -1910111873;
assign addr[4717] = -1918775195;
assign addr[4718] = -1927286370;
assign addr[4719] = -1935644723;
assign addr[4720] = -1943849591;
assign addr[4721] = -1951900324;
assign addr[4722] = -1959796283;
assign addr[4723] = -1967536842;
assign addr[4724] = -1975121388;
assign addr[4725] = -1982549318;
assign addr[4726] = -1989820044;
assign addr[4727] = -1996932990;
assign addr[4728] = -2003887591;
assign addr[4729] = -2010683297;
assign addr[4730] = -2017319567;
assign addr[4731] = -2023795876;
assign addr[4732] = -2030111710;
assign addr[4733] = -2036266570;
assign addr[4734] = -2042259965;
assign addr[4735] = -2048091422;
assign addr[4736] = -2053760478;
assign addr[4737] = -2059266683;
assign addr[4738] = -2064609600;
assign addr[4739] = -2069788807;
assign addr[4740] = -2074803892;
assign addr[4741] = -2079654458;
assign addr[4742] = -2084340120;
assign addr[4743] = -2088860507;
assign addr[4744] = -2093215260;
assign addr[4745] = -2097404033;
assign addr[4746] = -2101426496;
assign addr[4747] = -2105282327;
assign addr[4748] = -2108971223;
assign addr[4749] = -2112492891;
assign addr[4750] = -2115847050;
assign addr[4751] = -2119033436;
assign addr[4752] = -2122051796;
assign addr[4753] = -2124901890;
assign addr[4754] = -2127583492;
assign addr[4755] = -2130096389;
assign addr[4756] = -2132440383;
assign addr[4757] = -2134615288;
assign addr[4758] = -2136620930;
assign addr[4759] = -2138457152;
assign addr[4760] = -2140123807;
assign addr[4761] = -2141620763;
assign addr[4762] = -2142947902;
assign addr[4763] = -2144105118;
assign addr[4764] = -2145092320;
assign addr[4765] = -2145909429;
assign addr[4766] = -2146556380;
assign addr[4767] = -2147033123;
assign addr[4768] = -2147339619;
assign addr[4769] = -2147475844;
assign addr[4770] = -2147441787;
assign addr[4771] = -2147237452;
assign addr[4772] = -2146862854;
assign addr[4773] = -2146318022;
assign addr[4774] = -2145603001;
assign addr[4775] = -2144717846;
assign addr[4776] = -2143662628;
assign addr[4777] = -2142437431;
assign addr[4778] = -2141042352;
assign addr[4779] = -2139477502;
assign addr[4780] = -2137743003;
assign addr[4781] = -2135838995;
assign addr[4782] = -2133765628;
assign addr[4783] = -2131523066;
assign addr[4784] = -2129111488;
assign addr[4785] = -2126531084;
assign addr[4786] = -2123782059;
assign addr[4787] = -2120864631;
assign addr[4788] = -2117779031;
assign addr[4789] = -2114525505;
assign addr[4790] = -2111104309;
assign addr[4791] = -2107515716;
assign addr[4792] = -2103760010;
assign addr[4793] = -2099837489;
assign addr[4794] = -2095748463;
assign addr[4795] = -2091493257;
assign addr[4796] = -2087072209;
assign addr[4797] = -2082485668;
assign addr[4798] = -2077733999;
assign addr[4799] = -2072817579;
assign addr[4800] = -2067736796;
assign addr[4801] = -2062492055;
assign addr[4802] = -2057083771;
assign addr[4803] = -2051512372;
assign addr[4804] = -2045778302;
assign addr[4805] = -2039882013;
assign addr[4806] = -2033823974;
assign addr[4807] = -2027604666;
assign addr[4808] = -2021224581;
assign addr[4809] = -2014684225;
assign addr[4810] = -2007984117;
assign addr[4811] = -2001124788;
assign addr[4812] = -1994106782;
assign addr[4813] = -1986930656;
assign addr[4814] = -1979596978;
assign addr[4815] = -1972106330;
assign addr[4816] = -1964459306;
assign addr[4817] = -1956656513;
assign addr[4818] = -1948698568;
assign addr[4819] = -1940586104;
assign addr[4820] = -1932319763;
assign addr[4821] = -1923900201;
assign addr[4822] = -1915328086;
assign addr[4823] = -1906604097;
assign addr[4824] = -1897728925;
assign addr[4825] = -1888703276;
assign addr[4826] = -1879527863;
assign addr[4827] = -1870203416;
assign addr[4828] = -1860730673;
assign addr[4829] = -1851110385;
assign addr[4830] = -1841343316;
assign addr[4831] = -1831430239;
assign addr[4832] = -1821371941;
assign addr[4833] = -1811169220;
assign addr[4834] = -1800822883;
assign addr[4835] = -1790333753;
assign addr[4836] = -1779702660;
assign addr[4837] = -1768930447;
assign addr[4838] = -1758017969;
assign addr[4839] = -1746966091;
assign addr[4840] = -1735775690;
assign addr[4841] = -1724447652;
assign addr[4842] = -1712982875;
assign addr[4843] = -1701382270;
assign addr[4844] = -1689646755;
assign addr[4845] = -1677777262;
assign addr[4846] = -1665774731;
assign addr[4847] = -1653640115;
assign addr[4848] = -1641374375;
assign addr[4849] = -1628978484;
assign addr[4850] = -1616453425;
assign addr[4851] = -1603800191;
assign addr[4852] = -1591019785;
assign addr[4853] = -1578113222;
assign addr[4854] = -1565081523;
assign addr[4855] = -1551925723;
assign addr[4856] = -1538646865;
assign addr[4857] = -1525246002;
assign addr[4858] = -1511724196;
assign addr[4859] = -1498082520;
assign addr[4860] = -1484322054;
assign addr[4861] = -1470443891;
assign addr[4862] = -1456449131;
assign addr[4863] = -1442338884;
assign addr[4864] = -1428114267;
assign addr[4865] = -1413776410;
assign addr[4866] = -1399326449;
assign addr[4867] = -1384765530;
assign addr[4868] = -1370094808;
assign addr[4869] = -1355315445;
assign addr[4870] = -1340428615;
assign addr[4871] = -1325435496;
assign addr[4872] = -1310337279;
assign addr[4873] = -1295135159;
assign addr[4874] = -1279830344;
assign addr[4875] = -1264424045;
assign addr[4876] = -1248917486;
assign addr[4877] = -1233311895;
assign addr[4878] = -1217608510;
assign addr[4879] = -1201808576;
assign addr[4880] = -1185913346;
assign addr[4881] = -1169924081;
assign addr[4882] = -1153842047;
assign addr[4883] = -1137668521;
assign addr[4884] = -1121404785;
assign addr[4885] = -1105052128;
assign addr[4886] = -1088611847;
assign addr[4887] = -1072085246;
assign addr[4888] = -1055473635;
assign addr[4889] = -1038778332;
assign addr[4890] = -1022000660;
assign addr[4891] = -1005141949;
assign addr[4892] = -988203537;
assign addr[4893] = -971186766;
assign addr[4894] = -954092986;
assign addr[4895] = -936923553;
assign addr[4896] = -919679827;
assign addr[4897] = -902363176;
assign addr[4898] = -884974973;
assign addr[4899] = -867516597;
assign addr[4900] = -849989433;
assign addr[4901] = -832394869;
assign addr[4902] = -814734301;
assign addr[4903] = -797009130;
assign addr[4904] = -779220762;
assign addr[4905] = -761370605;
assign addr[4906] = -743460077;
assign addr[4907] = -725490597;
assign addr[4908] = -707463589;
assign addr[4909] = -689380485;
assign addr[4910] = -671242716;
assign addr[4911] = -653051723;
assign addr[4912] = -634808946;
assign addr[4913] = -616515832;
assign addr[4914] = -598173833;
assign addr[4915] = -579784402;
assign addr[4916] = -561348998;
assign addr[4917] = -542869083;
assign addr[4918] = -524346121;
assign addr[4919] = -505781581;
assign addr[4920] = -487176937;
assign addr[4921] = -468533662;
assign addr[4922] = -449853235;
assign addr[4923] = -431137138;
assign addr[4924] = -412386854;
assign addr[4925] = -393603870;
assign addr[4926] = -374789676;
assign addr[4927] = -355945764;
assign addr[4928] = -337073627;
assign addr[4929] = -318174762;
assign addr[4930] = -299250668;
assign addr[4931] = -280302845;
assign addr[4932] = -261332796;
assign addr[4933] = -242342025;
assign addr[4934] = -223332037;
assign addr[4935] = -204304341;
assign addr[4936] = -185260444;
assign addr[4937] = -166201858;
assign addr[4938] = -147130093;
assign addr[4939] = -128046661;
assign addr[4940] = -108953076;
assign addr[4941] = -89850852;
assign addr[4942] = -70741503;
assign addr[4943] = -51626544;
assign addr[4944] = -32507492;
assign addr[4945] = -13385863;
assign addr[4946] = 5736829;
assign addr[4947] = 24859065;
assign addr[4948] = 43979330;
assign addr[4949] = 63096108;
assign addr[4950] = 82207882;
assign addr[4951] = 101313138;
assign addr[4952] = 120410361;
assign addr[4953] = 139498035;
assign addr[4954] = 158574649;
assign addr[4955] = 177638688;
assign addr[4956] = 196688642;
assign addr[4957] = 215722999;
assign addr[4958] = 234740251;
assign addr[4959] = 253738890;
assign addr[4960] = 272717408;
assign addr[4961] = 291674302;
assign addr[4962] = 310608068;
assign addr[4963] = 329517204;
assign addr[4964] = 348400212;
assign addr[4965] = 367255594;
assign addr[4966] = 386081854;
assign addr[4967] = 404877501;
assign addr[4968] = 423641043;
assign addr[4969] = 442370993;
assign addr[4970] = 461065866;
assign addr[4971] = 479724180;
assign addr[4972] = 498344454;
assign addr[4973] = 516925212;
assign addr[4974] = 535464981;
assign addr[4975] = 553962291;
assign addr[4976] = 572415676;
assign addr[4977] = 590823671;
assign addr[4978] = 609184818;
assign addr[4979] = 627497660;
assign addr[4980] = 645760745;
assign addr[4981] = 663972625;
assign addr[4982] = 682131857;
assign addr[4983] = 700236999;
assign addr[4984] = 718286617;
assign addr[4985] = 736279279;
assign addr[4986] = 754213559;
assign addr[4987] = 772088034;
assign addr[4988] = 789901288;
assign addr[4989] = 807651907;
assign addr[4990] = 825338484;
assign addr[4991] = 842959617;
assign addr[4992] = 860513908;
assign addr[4993] = 877999966;
assign addr[4994] = 895416404;
assign addr[4995] = 912761841;
assign addr[4996] = 930034901;
assign addr[4997] = 947234215;
assign addr[4998] = 964358420;
assign addr[4999] = 981406156;
assign addr[5000] = 998376073;
assign addr[5001] = 1015266825;
assign addr[5002] = 1032077073;
assign addr[5003] = 1048805483;
assign addr[5004] = 1065450729;
assign addr[5005] = 1082011492;
assign addr[5006] = 1098486458;
assign addr[5007] = 1114874320;
assign addr[5008] = 1131173780;
assign addr[5009] = 1147383544;
assign addr[5010] = 1163502328;
assign addr[5011] = 1179528853;
assign addr[5012] = 1195461849;
assign addr[5013] = 1211300053;
assign addr[5014] = 1227042207;
assign addr[5015] = 1242687064;
assign addr[5016] = 1258233384;
assign addr[5017] = 1273679934;
assign addr[5018] = 1289025489;
assign addr[5019] = 1304268832;
assign addr[5020] = 1319408754;
assign addr[5021] = 1334444055;
assign addr[5022] = 1349373543;
assign addr[5023] = 1364196034;
assign addr[5024] = 1378910353;
assign addr[5025] = 1393515332;
assign addr[5026] = 1408009814;
assign addr[5027] = 1422392650;
assign addr[5028] = 1436662698;
assign addr[5029] = 1450818828;
assign addr[5030] = 1464859917;
assign addr[5031] = 1478784851;
assign addr[5032] = 1492592527;
assign addr[5033] = 1506281850;
assign addr[5034] = 1519851733;
assign addr[5035] = 1533301101;
assign addr[5036] = 1546628888;
assign addr[5037] = 1559834037;
assign addr[5038] = 1572915501;
assign addr[5039] = 1585872242;
assign addr[5040] = 1598703233;
assign addr[5041] = 1611407456;
assign addr[5042] = 1623983905;
assign addr[5043] = 1636431582;
assign addr[5044] = 1648749499;
assign addr[5045] = 1660936681;
assign addr[5046] = 1672992161;
assign addr[5047] = 1684914983;
assign addr[5048] = 1696704201;
assign addr[5049] = 1708358881;
assign addr[5050] = 1719878099;
assign addr[5051] = 1731260941;
assign addr[5052] = 1742506504;
assign addr[5053] = 1753613897;
assign addr[5054] = 1764582240;
assign addr[5055] = 1775410662;
assign addr[5056] = 1786098304;
assign addr[5057] = 1796644320;
assign addr[5058] = 1807047873;
assign addr[5059] = 1817308138;
assign addr[5060] = 1827424302;
assign addr[5061] = 1837395562;
assign addr[5062] = 1847221128;
assign addr[5063] = 1856900221;
assign addr[5064] = 1866432072;
assign addr[5065] = 1875815927;
assign addr[5066] = 1885051042;
assign addr[5067] = 1894136683;
assign addr[5068] = 1903072131;
assign addr[5069] = 1911856677;
assign addr[5070] = 1920489624;
assign addr[5071] = 1928970288;
assign addr[5072] = 1937297997;
assign addr[5073] = 1945472089;
assign addr[5074] = 1953491918;
assign addr[5075] = 1961356847;
assign addr[5076] = 1969066252;
assign addr[5077] = 1976619522;
assign addr[5078] = 1984016058;
assign addr[5079] = 1991255274;
assign addr[5080] = 1998336596;
assign addr[5081] = 2005259462;
assign addr[5082] = 2012023322;
assign addr[5083] = 2018627642;
assign addr[5084] = 2025071897;
assign addr[5085] = 2031355576;
assign addr[5086] = 2037478181;
assign addr[5087] = 2043439226;
assign addr[5088] = 2049238240;
assign addr[5089] = 2054874761;
assign addr[5090] = 2060348343;
assign addr[5091] = 2065658552;
assign addr[5092] = 2070804967;
assign addr[5093] = 2075787180;
assign addr[5094] = 2080604795;
assign addr[5095] = 2085257431;
assign addr[5096] = 2089744719;
assign addr[5097] = 2094066304;
assign addr[5098] = 2098221841;
assign addr[5099] = 2102211002;
assign addr[5100] = 2106033471;
assign addr[5101] = 2109688944;
assign addr[5102] = 2113177132;
assign addr[5103] = 2116497758;
assign addr[5104] = 2119650558;
assign addr[5105] = 2122635283;
assign addr[5106] = 2125451696;
assign addr[5107] = 2128099574;
assign addr[5108] = 2130578706;
assign addr[5109] = 2132888897;
assign addr[5110] = 2135029962;
assign addr[5111] = 2137001733;
assign addr[5112] = 2138804053;
assign addr[5113] = 2140436778;
assign addr[5114] = 2141899780;
assign addr[5115] = 2143192942;
assign addr[5116] = 2144316162;
assign addr[5117] = 2145269351;
assign addr[5118] = 2146052433;
assign addr[5119] = 2146665347;
assign addr[5120] = 2147108043;
assign addr[5121] = 2147380486;
assign addr[5122] = 2147482655;
assign addr[5123] = 2147414542;
assign addr[5124] = 2147176152;
assign addr[5125] = 2146767505;
assign addr[5126] = 2146188631;
assign addr[5127] = 2145439578;
assign addr[5128] = 2144520405;
assign addr[5129] = 2143431184;
assign addr[5130] = 2142172003;
assign addr[5131] = 2140742960;
assign addr[5132] = 2139144169;
assign addr[5133] = 2137375758;
assign addr[5134] = 2135437865;
assign addr[5135] = 2133330646;
assign addr[5136] = 2131054266;
assign addr[5137] = 2128608907;
assign addr[5138] = 2125994762;
assign addr[5139] = 2123212038;
assign addr[5140] = 2120260957;
assign addr[5141] = 2117141752;
assign addr[5142] = 2113854671;
assign addr[5143] = 2110399974;
assign addr[5144] = 2106777935;
assign addr[5145] = 2102988841;
assign addr[5146] = 2099032994;
assign addr[5147] = 2094910706;
assign addr[5148] = 2090622304;
assign addr[5149] = 2086168128;
assign addr[5150] = 2081548533;
assign addr[5151] = 2076763883;
assign addr[5152] = 2071814558;
assign addr[5153] = 2066700952;
assign addr[5154] = 2061423468;
assign addr[5155] = 2055982526;
assign addr[5156] = 2050378558;
assign addr[5157] = 2044612007;
assign addr[5158] = 2038683330;
assign addr[5159] = 2032592999;
assign addr[5160] = 2026341495;
assign addr[5161] = 2019929315;
assign addr[5162] = 2013356967;
assign addr[5163] = 2006624971;
assign addr[5164] = 1999733863;
assign addr[5165] = 1992684188;
assign addr[5166] = 1985476506;
assign addr[5167] = 1978111387;
assign addr[5168] = 1970589416;
assign addr[5169] = 1962911189;
assign addr[5170] = 1955077316;
assign addr[5171] = 1947088417;
assign addr[5172] = 1938945125;
assign addr[5173] = 1930648088;
assign addr[5174] = 1922197961;
assign addr[5175] = 1913595416;
assign addr[5176] = 1904841135;
assign addr[5177] = 1895935811;
assign addr[5178] = 1886880151;
assign addr[5179] = 1877674873;
assign addr[5180] = 1868320707;
assign addr[5181] = 1858818395;
assign addr[5182] = 1849168689;
assign addr[5183] = 1839372356;
assign addr[5184] = 1829430172;
assign addr[5185] = 1819342925;
assign addr[5186] = 1809111415;
assign addr[5187] = 1798736454;
assign addr[5188] = 1788218865;
assign addr[5189] = 1777559480;
assign addr[5190] = 1766759146;
assign addr[5191] = 1755818718;
assign addr[5192] = 1744739065;
assign addr[5193] = 1733521064;
assign addr[5194] = 1722165606;
assign addr[5195] = 1710673591;
assign addr[5196] = 1699045930;
assign addr[5197] = 1687283545;
assign addr[5198] = 1675387369;
assign addr[5199] = 1663358344;
assign addr[5200] = 1651197426;
assign addr[5201] = 1638905577;
assign addr[5202] = 1626483774;
assign addr[5203] = 1613933000;
assign addr[5204] = 1601254251;
assign addr[5205] = 1588448533;
assign addr[5206] = 1575516860;
assign addr[5207] = 1562460258;
assign addr[5208] = 1549279763;
assign addr[5209] = 1535976419;
assign addr[5210] = 1522551282;
assign addr[5211] = 1509005416;
assign addr[5212] = 1495339895;
assign addr[5213] = 1481555802;
assign addr[5214] = 1467654232;
assign addr[5215] = 1453636285;
assign addr[5216] = 1439503074;
assign addr[5217] = 1425255719;
assign addr[5218] = 1410895350;
assign addr[5219] = 1396423105;
assign addr[5220] = 1381840133;
assign addr[5221] = 1367147589;
assign addr[5222] = 1352346639;
assign addr[5223] = 1337438456;
assign addr[5224] = 1322424222;
assign addr[5225] = 1307305128;
assign addr[5226] = 1292082373;
assign addr[5227] = 1276757164;
assign addr[5228] = 1261330715;
assign addr[5229] = 1245804251;
assign addr[5230] = 1230179002;
assign addr[5231] = 1214456207;
assign addr[5232] = 1198637114;
assign addr[5233] = 1182722976;
assign addr[5234] = 1166715055;
assign addr[5235] = 1150614620;
assign addr[5236] = 1134422949;
assign addr[5237] = 1118141326;
assign addr[5238] = 1101771040;
assign addr[5239] = 1085313391;
assign addr[5240] = 1068769683;
assign addr[5241] = 1052141228;
assign addr[5242] = 1035429345;
assign addr[5243] = 1018635358;
assign addr[5244] = 1001760600;
assign addr[5245] = 984806408;
assign addr[5246] = 967774128;
assign addr[5247] = 950665109;
assign addr[5248] = 933480707;
assign addr[5249] = 916222287;
assign addr[5250] = 898891215;
assign addr[5251] = 881488868;
assign addr[5252] = 864016623;
assign addr[5253] = 846475867;
assign addr[5254] = 828867991;
assign addr[5255] = 811194391;
assign addr[5256] = 793456467;
assign addr[5257] = 775655628;
assign addr[5258] = 757793284;
assign addr[5259] = 739870851;
assign addr[5260] = 721889752;
assign addr[5261] = 703851410;
assign addr[5262] = 685757258;
assign addr[5263] = 667608730;
assign addr[5264] = 649407264;
assign addr[5265] = 631154304;
assign addr[5266] = 612851297;
assign addr[5267] = 594499695;
assign addr[5268] = 576100953;
assign addr[5269] = 557656529;
assign addr[5270] = 539167887;
assign addr[5271] = 520636492;
assign addr[5272] = 502063814;
assign addr[5273] = 483451325;
assign addr[5274] = 464800501;
assign addr[5275] = 446112822;
assign addr[5276] = 427389768;
assign addr[5277] = 408632825;
assign addr[5278] = 389843480;
assign addr[5279] = 371023223;
assign addr[5280] = 352173546;
assign addr[5281] = 333295944;
assign addr[5282] = 314391913;
assign addr[5283] = 295462954;
assign addr[5284] = 276510565;
assign addr[5285] = 257536251;
assign addr[5286] = 238541516;
assign addr[5287] = 219527866;
assign addr[5288] = 200496809;
assign addr[5289] = 181449854;
assign addr[5290] = 162388511;
assign addr[5291] = 143314291;
assign addr[5292] = 124228708;
assign addr[5293] = 105133274;
assign addr[5294] = 86029503;
assign addr[5295] = 66918911;
assign addr[5296] = 47803013;
assign addr[5297] = 28683324;
assign addr[5298] = 9561361;
assign addr[5299] = -9561361;
assign addr[5300] = -28683324;
assign addr[5301] = -47803013;
assign addr[5302] = -66918911;
assign addr[5303] = -86029503;
assign addr[5304] = -105133274;
assign addr[5305] = -124228708;
assign addr[5306] = -143314291;
assign addr[5307] = -162388511;
assign addr[5308] = -181449854;
assign addr[5309] = -200496809;
assign addr[5310] = -219527866;
assign addr[5311] = -238541516;
assign addr[5312] = -257536251;
assign addr[5313] = -276510565;
assign addr[5314] = -295462954;
assign addr[5315] = -314391913;
assign addr[5316] = -333295944;
assign addr[5317] = -352173546;
assign addr[5318] = -371023223;
assign addr[5319] = -389843480;
assign addr[5320] = -408632825;
assign addr[5321] = -427389768;
assign addr[5322] = -446112822;
assign addr[5323] = -464800501;
assign addr[5324] = -483451325;
assign addr[5325] = -502063814;
assign addr[5326] = -520636492;
assign addr[5327] = -539167887;
assign addr[5328] = -557656529;
assign addr[5329] = -576100953;
assign addr[5330] = -594499695;
assign addr[5331] = -612851297;
assign addr[5332] = -631154304;
assign addr[5333] = -649407264;
assign addr[5334] = -667608730;
assign addr[5335] = -685757258;
assign addr[5336] = -703851410;
assign addr[5337] = -721889752;
assign addr[5338] = -739870851;
assign addr[5339] = -757793284;
assign addr[5340] = -775655628;
assign addr[5341] = -793456467;
assign addr[5342] = -811194391;
assign addr[5343] = -828867991;
assign addr[5344] = -846475867;
assign addr[5345] = -864016623;
assign addr[5346] = -881488868;
assign addr[5347] = -898891215;
assign addr[5348] = -916222287;
assign addr[5349] = -933480707;
assign addr[5350] = -950665109;
assign addr[5351] = -967774128;
assign addr[5352] = -984806408;
assign addr[5353] = -1001760600;
assign addr[5354] = -1018635358;
assign addr[5355] = -1035429345;
assign addr[5356] = -1052141228;
assign addr[5357] = -1068769683;
assign addr[5358] = -1085313391;
assign addr[5359] = -1101771040;
assign addr[5360] = -1118141326;
assign addr[5361] = -1134422949;
assign addr[5362] = -1150614620;
assign addr[5363] = -1166715055;
assign addr[5364] = -1182722976;
assign addr[5365] = -1198637114;
assign addr[5366] = -1214456207;
assign addr[5367] = -1230179002;
assign addr[5368] = -1245804251;
assign addr[5369] = -1261330715;
assign addr[5370] = -1276757164;
assign addr[5371] = -1292082373;
assign addr[5372] = -1307305128;
assign addr[5373] = -1322424222;
assign addr[5374] = -1337438456;
assign addr[5375] = -1352346639;
assign addr[5376] = -1367147589;
assign addr[5377] = -1381840133;
assign addr[5378] = -1396423105;
assign addr[5379] = -1410895350;
assign addr[5380] = -1425255719;
assign addr[5381] = -1439503074;
assign addr[5382] = -1453636285;
assign addr[5383] = -1467654232;
assign addr[5384] = -1481555802;
assign addr[5385] = -1495339895;
assign addr[5386] = -1509005416;
assign addr[5387] = -1522551282;
assign addr[5388] = -1535976419;
assign addr[5389] = -1549279763;
assign addr[5390] = -1562460258;
assign addr[5391] = -1575516860;
assign addr[5392] = -1588448533;
assign addr[5393] = -1601254251;
assign addr[5394] = -1613933000;
assign addr[5395] = -1626483774;
assign addr[5396] = -1638905577;
assign addr[5397] = -1651197426;
assign addr[5398] = -1663358344;
assign addr[5399] = -1675387369;
assign addr[5400] = -1687283545;
assign addr[5401] = -1699045930;
assign addr[5402] = -1710673591;
assign addr[5403] = -1722165606;
assign addr[5404] = -1733521064;
assign addr[5405] = -1744739065;
assign addr[5406] = -1755818718;
assign addr[5407] = -1766759146;
assign addr[5408] = -1777559480;
assign addr[5409] = -1788218865;
assign addr[5410] = -1798736454;
assign addr[5411] = -1809111415;
assign addr[5412] = -1819342925;
assign addr[5413] = -1829430172;
assign addr[5414] = -1839372356;
assign addr[5415] = -1849168689;
assign addr[5416] = -1858818395;
assign addr[5417] = -1868320707;
assign addr[5418] = -1877674873;
assign addr[5419] = -1886880151;
assign addr[5420] = -1895935811;
assign addr[5421] = -1904841135;
assign addr[5422] = -1913595416;
assign addr[5423] = -1922197961;
assign addr[5424] = -1930648088;
assign addr[5425] = -1938945125;
assign addr[5426] = -1947088417;
assign addr[5427] = -1955077316;
assign addr[5428] = -1962911189;
assign addr[5429] = -1970589416;
assign addr[5430] = -1978111387;
assign addr[5431] = -1985476506;
assign addr[5432] = -1992684188;
assign addr[5433] = -1999733863;
assign addr[5434] = -2006624971;
assign addr[5435] = -2013356967;
assign addr[5436] = -2019929315;
assign addr[5437] = -2026341495;
assign addr[5438] = -2032592999;
assign addr[5439] = -2038683330;
assign addr[5440] = -2044612007;
assign addr[5441] = -2050378558;
assign addr[5442] = -2055982526;
assign addr[5443] = -2061423468;
assign addr[5444] = -2066700952;
assign addr[5445] = -2071814558;
assign addr[5446] = -2076763883;
assign addr[5447] = -2081548533;
assign addr[5448] = -2086168128;
assign addr[5449] = -2090622304;
assign addr[5450] = -2094910706;
assign addr[5451] = -2099032994;
assign addr[5452] = -2102988841;
assign addr[5453] = -2106777935;
assign addr[5454] = -2110399974;
assign addr[5455] = -2113854671;
assign addr[5456] = -2117141752;
assign addr[5457] = -2120260957;
assign addr[5458] = -2123212038;
assign addr[5459] = -2125994762;
assign addr[5460] = -2128608907;
assign addr[5461] = -2131054266;
assign addr[5462] = -2133330646;
assign addr[5463] = -2135437865;
assign addr[5464] = -2137375758;
assign addr[5465] = -2139144169;
assign addr[5466] = -2140742960;
assign addr[5467] = -2142172003;
assign addr[5468] = -2143431184;
assign addr[5469] = -2144520405;
assign addr[5470] = -2145439578;
assign addr[5471] = -2146188631;
assign addr[5472] = -2146767505;
assign addr[5473] = -2147176152;
assign addr[5474] = -2147414542;
assign addr[5475] = -2147482655;
assign addr[5476] = -2147380486;
assign addr[5477] = -2147108043;
assign addr[5478] = -2146665347;
assign addr[5479] = -2146052433;
assign addr[5480] = -2145269351;
assign addr[5481] = -2144316162;
assign addr[5482] = -2143192942;
assign addr[5483] = -2141899780;
assign addr[5484] = -2140436778;
assign addr[5485] = -2138804053;
assign addr[5486] = -2137001733;
assign addr[5487] = -2135029962;
assign addr[5488] = -2132888897;
assign addr[5489] = -2130578706;
assign addr[5490] = -2128099574;
assign addr[5491] = -2125451696;
assign addr[5492] = -2122635283;
assign addr[5493] = -2119650558;
assign addr[5494] = -2116497758;
assign addr[5495] = -2113177132;
assign addr[5496] = -2109688944;
assign addr[5497] = -2106033471;
assign addr[5498] = -2102211002;
assign addr[5499] = -2098221841;
assign addr[5500] = -2094066304;
assign addr[5501] = -2089744719;
assign addr[5502] = -2085257431;
assign addr[5503] = -2080604795;
assign addr[5504] = -2075787180;
assign addr[5505] = -2070804967;
assign addr[5506] = -2065658552;
assign addr[5507] = -2060348343;
assign addr[5508] = -2054874761;
assign addr[5509] = -2049238240;
assign addr[5510] = -2043439226;
assign addr[5511] = -2037478181;
assign addr[5512] = -2031355576;
assign addr[5513] = -2025071897;
assign addr[5514] = -2018627642;
assign addr[5515] = -2012023322;
assign addr[5516] = -2005259462;
assign addr[5517] = -1998336596;
assign addr[5518] = -1991255274;
assign addr[5519] = -1984016058;
assign addr[5520] = -1976619522;
assign addr[5521] = -1969066252;
assign addr[5522] = -1961356847;
assign addr[5523] = -1953491918;
assign addr[5524] = -1945472089;
assign addr[5525] = -1937297997;
assign addr[5526] = -1928970288;
assign addr[5527] = -1920489624;
assign addr[5528] = -1911856677;
assign addr[5529] = -1903072131;
assign addr[5530] = -1894136683;
assign addr[5531] = -1885051042;
assign addr[5532] = -1875815927;
assign addr[5533] = -1866432072;
assign addr[5534] = -1856900221;
assign addr[5535] = -1847221128;
assign addr[5536] = -1837395562;
assign addr[5537] = -1827424302;
assign addr[5538] = -1817308138;
assign addr[5539] = -1807047873;
assign addr[5540] = -1796644320;
assign addr[5541] = -1786098304;
assign addr[5542] = -1775410662;
assign addr[5543] = -1764582240;
assign addr[5544] = -1753613897;
assign addr[5545] = -1742506504;
assign addr[5546] = -1731260941;
assign addr[5547] = -1719878099;
assign addr[5548] = -1708358881;
assign addr[5549] = -1696704201;
assign addr[5550] = -1684914983;
assign addr[5551] = -1672992161;
assign addr[5552] = -1660936681;
assign addr[5553] = -1648749499;
assign addr[5554] = -1636431582;
assign addr[5555] = -1623983905;
assign addr[5556] = -1611407456;
assign addr[5557] = -1598703233;
assign addr[5558] = -1585872242;
assign addr[5559] = -1572915501;
assign addr[5560] = -1559834037;
assign addr[5561] = -1546628888;
assign addr[5562] = -1533301101;
assign addr[5563] = -1519851733;
assign addr[5564] = -1506281850;
assign addr[5565] = -1492592527;
assign addr[5566] = -1478784851;
assign addr[5567] = -1464859917;
assign addr[5568] = -1450818828;
assign addr[5569] = -1436662698;
assign addr[5570] = -1422392650;
assign addr[5571] = -1408009814;
assign addr[5572] = -1393515332;
assign addr[5573] = -1378910353;
assign addr[5574] = -1364196034;
assign addr[5575] = -1349373543;
assign addr[5576] = -1334444055;
assign addr[5577] = -1319408754;
assign addr[5578] = -1304268832;
assign addr[5579] = -1289025489;
assign addr[5580] = -1273679934;
assign addr[5581] = -1258233384;
assign addr[5582] = -1242687064;
assign addr[5583] = -1227042207;
assign addr[5584] = -1211300053;
assign addr[5585] = -1195461849;
assign addr[5586] = -1179528853;
assign addr[5587] = -1163502328;
assign addr[5588] = -1147383544;
assign addr[5589] = -1131173780;
assign addr[5590] = -1114874320;
assign addr[5591] = -1098486458;
assign addr[5592] = -1082011492;
assign addr[5593] = -1065450729;
assign addr[5594] = -1048805483;
assign addr[5595] = -1032077073;
assign addr[5596] = -1015266825;
assign addr[5597] = -998376073;
assign addr[5598] = -981406156;
assign addr[5599] = -964358420;
assign addr[5600] = -947234215;
assign addr[5601] = -930034901;
assign addr[5602] = -912761841;
assign addr[5603] = -895416404;
assign addr[5604] = -877999966;
assign addr[5605] = -860513908;
assign addr[5606] = -842959617;
assign addr[5607] = -825338484;
assign addr[5608] = -807651907;
assign addr[5609] = -789901288;
assign addr[5610] = -772088034;
assign addr[5611] = -754213559;
assign addr[5612] = -736279279;
assign addr[5613] = -718286617;
assign addr[5614] = -700236999;
assign addr[5615] = -682131857;
assign addr[5616] = -663972625;
assign addr[5617] = -645760745;
assign addr[5618] = -627497660;
assign addr[5619] = -609184818;
assign addr[5620] = -590823671;
assign addr[5621] = -572415676;
assign addr[5622] = -553962291;
assign addr[5623] = -535464981;
assign addr[5624] = -516925212;
assign addr[5625] = -498344454;
assign addr[5626] = -479724180;
assign addr[5627] = -461065866;
assign addr[5628] = -442370993;
assign addr[5629] = -423641043;
assign addr[5630] = -404877501;
assign addr[5631] = -386081854;
assign addr[5632] = -367255594;
assign addr[5633] = -348400212;
assign addr[5634] = -329517204;
assign addr[5635] = -310608068;
assign addr[5636] = -291674302;
assign addr[5637] = -272717408;
assign addr[5638] = -253738890;
assign addr[5639] = -234740251;
assign addr[5640] = -215722999;
assign addr[5641] = -196688642;
assign addr[5642] = -177638688;
assign addr[5643] = -158574649;
assign addr[5644] = -139498035;
assign addr[5645] = -120410361;
assign addr[5646] = -101313138;
assign addr[5647] = -82207882;
assign addr[5648] = -63096108;
assign addr[5649] = -43979330;
assign addr[5650] = -24859065;
assign addr[5651] = -5736829;
assign addr[5652] = 13385863;
assign addr[5653] = 32507492;
assign addr[5654] = 51626544;
assign addr[5655] = 70741503;
assign addr[5656] = 89850852;
assign addr[5657] = 108953076;
assign addr[5658] = 128046661;
assign addr[5659] = 147130093;
assign addr[5660] = 166201858;
assign addr[5661] = 185260444;
assign addr[5662] = 204304341;
assign addr[5663] = 223332037;
assign addr[5664] = 242342025;
assign addr[5665] = 261332796;
assign addr[5666] = 280302845;
assign addr[5667] = 299250668;
assign addr[5668] = 318174762;
assign addr[5669] = 337073627;
assign addr[5670] = 355945764;
assign addr[5671] = 374789676;
assign addr[5672] = 393603870;
assign addr[5673] = 412386854;
assign addr[5674] = 431137138;
assign addr[5675] = 449853235;
assign addr[5676] = 468533662;
assign addr[5677] = 487176937;
assign addr[5678] = 505781581;
assign addr[5679] = 524346121;
assign addr[5680] = 542869083;
assign addr[5681] = 561348998;
assign addr[5682] = 579784402;
assign addr[5683] = 598173833;
assign addr[5684] = 616515832;
assign addr[5685] = 634808946;
assign addr[5686] = 653051723;
assign addr[5687] = 671242716;
assign addr[5688] = 689380485;
assign addr[5689] = 707463589;
assign addr[5690] = 725490597;
assign addr[5691] = 743460077;
assign addr[5692] = 761370605;
assign addr[5693] = 779220762;
assign addr[5694] = 797009130;
assign addr[5695] = 814734301;
assign addr[5696] = 832394869;
assign addr[5697] = 849989433;
assign addr[5698] = 867516597;
assign addr[5699] = 884974973;
assign addr[5700] = 902363176;
assign addr[5701] = 919679827;
assign addr[5702] = 936923553;
assign addr[5703] = 954092986;
assign addr[5704] = 971186766;
assign addr[5705] = 988203537;
assign addr[5706] = 1005141949;
assign addr[5707] = 1022000660;
assign addr[5708] = 1038778332;
assign addr[5709] = 1055473635;
assign addr[5710] = 1072085246;
assign addr[5711] = 1088611847;
assign addr[5712] = 1105052128;
assign addr[5713] = 1121404785;
assign addr[5714] = 1137668521;
assign addr[5715] = 1153842047;
assign addr[5716] = 1169924081;
assign addr[5717] = 1185913346;
assign addr[5718] = 1201808576;
assign addr[5719] = 1217608510;
assign addr[5720] = 1233311895;
assign addr[5721] = 1248917486;
assign addr[5722] = 1264424045;
assign addr[5723] = 1279830344;
assign addr[5724] = 1295135159;
assign addr[5725] = 1310337279;
assign addr[5726] = 1325435496;
assign addr[5727] = 1340428615;
assign addr[5728] = 1355315445;
assign addr[5729] = 1370094808;
assign addr[5730] = 1384765530;
assign addr[5731] = 1399326449;
assign addr[5732] = 1413776410;
assign addr[5733] = 1428114267;
assign addr[5734] = 1442338884;
assign addr[5735] = 1456449131;
assign addr[5736] = 1470443891;
assign addr[5737] = 1484322054;
assign addr[5738] = 1498082520;
assign addr[5739] = 1511724196;
assign addr[5740] = 1525246002;
assign addr[5741] = 1538646865;
assign addr[5742] = 1551925723;
assign addr[5743] = 1565081523;
assign addr[5744] = 1578113222;
assign addr[5745] = 1591019785;
assign addr[5746] = 1603800191;
assign addr[5747] = 1616453425;
assign addr[5748] = 1628978484;
assign addr[5749] = 1641374375;
assign addr[5750] = 1653640115;
assign addr[5751] = 1665774731;
assign addr[5752] = 1677777262;
assign addr[5753] = 1689646755;
assign addr[5754] = 1701382270;
assign addr[5755] = 1712982875;
assign addr[5756] = 1724447652;
assign addr[5757] = 1735775690;
assign addr[5758] = 1746966091;
assign addr[5759] = 1758017969;
assign addr[5760] = 1768930447;
assign addr[5761] = 1779702660;
assign addr[5762] = 1790333753;
assign addr[5763] = 1800822883;
assign addr[5764] = 1811169220;
assign addr[5765] = 1821371941;
assign addr[5766] = 1831430239;
assign addr[5767] = 1841343316;
assign addr[5768] = 1851110385;
assign addr[5769] = 1860730673;
assign addr[5770] = 1870203416;
assign addr[5771] = 1879527863;
assign addr[5772] = 1888703276;
assign addr[5773] = 1897728925;
assign addr[5774] = 1906604097;
assign addr[5775] = 1915328086;
assign addr[5776] = 1923900201;
assign addr[5777] = 1932319763;
assign addr[5778] = 1940586104;
assign addr[5779] = 1948698568;
assign addr[5780] = 1956656513;
assign addr[5781] = 1964459306;
assign addr[5782] = 1972106330;
assign addr[5783] = 1979596978;
assign addr[5784] = 1986930656;
assign addr[5785] = 1994106782;
assign addr[5786] = 2001124788;
assign addr[5787] = 2007984117;
assign addr[5788] = 2014684225;
assign addr[5789] = 2021224581;
assign addr[5790] = 2027604666;
assign addr[5791] = 2033823974;
assign addr[5792] = 2039882013;
assign addr[5793] = 2045778302;
assign addr[5794] = 2051512372;
assign addr[5795] = 2057083771;
assign addr[5796] = 2062492055;
assign addr[5797] = 2067736796;
assign addr[5798] = 2072817579;
assign addr[5799] = 2077733999;
assign addr[5800] = 2082485668;
assign addr[5801] = 2087072209;
assign addr[5802] = 2091493257;
assign addr[5803] = 2095748463;
assign addr[5804] = 2099837489;
assign addr[5805] = 2103760010;
assign addr[5806] = 2107515716;
assign addr[5807] = 2111104309;
assign addr[5808] = 2114525505;
assign addr[5809] = 2117779031;
assign addr[5810] = 2120864631;
assign addr[5811] = 2123782059;
assign addr[5812] = 2126531084;
assign addr[5813] = 2129111488;
assign addr[5814] = 2131523066;
assign addr[5815] = 2133765628;
assign addr[5816] = 2135838995;
assign addr[5817] = 2137743003;
assign addr[5818] = 2139477502;
assign addr[5819] = 2141042352;
assign addr[5820] = 2142437431;
assign addr[5821] = 2143662628;
assign addr[5822] = 2144717846;
assign addr[5823] = 2145603001;
assign addr[5824] = 2146318022;
assign addr[5825] = 2146862854;
assign addr[5826] = 2147237452;
assign addr[5827] = 2147441787;
assign addr[5828] = 2147475844;
assign addr[5829] = 2147339619;
assign addr[5830] = 2147033123;
assign addr[5831] = 2146556380;
assign addr[5832] = 2145909429;
assign addr[5833] = 2145092320;
assign addr[5834] = 2144105118;
assign addr[5835] = 2142947902;
assign addr[5836] = 2141620763;
assign addr[5837] = 2140123807;
assign addr[5838] = 2138457152;
assign addr[5839] = 2136620930;
assign addr[5840] = 2134615288;
assign addr[5841] = 2132440383;
assign addr[5842] = 2130096389;
assign addr[5843] = 2127583492;
assign addr[5844] = 2124901890;
assign addr[5845] = 2122051796;
assign addr[5846] = 2119033436;
assign addr[5847] = 2115847050;
assign addr[5848] = 2112492891;
assign addr[5849] = 2108971223;
assign addr[5850] = 2105282327;
assign addr[5851] = 2101426496;
assign addr[5852] = 2097404033;
assign addr[5853] = 2093215260;
assign addr[5854] = 2088860507;
assign addr[5855] = 2084340120;
assign addr[5856] = 2079654458;
assign addr[5857] = 2074803892;
assign addr[5858] = 2069788807;
assign addr[5859] = 2064609600;
assign addr[5860] = 2059266683;
assign addr[5861] = 2053760478;
assign addr[5862] = 2048091422;
assign addr[5863] = 2042259965;
assign addr[5864] = 2036266570;
assign addr[5865] = 2030111710;
assign addr[5866] = 2023795876;
assign addr[5867] = 2017319567;
assign addr[5868] = 2010683297;
assign addr[5869] = 2003887591;
assign addr[5870] = 1996932990;
assign addr[5871] = 1989820044;
assign addr[5872] = 1982549318;
assign addr[5873] = 1975121388;
assign addr[5874] = 1967536842;
assign addr[5875] = 1959796283;
assign addr[5876] = 1951900324;
assign addr[5877] = 1943849591;
assign addr[5878] = 1935644723;
assign addr[5879] = 1927286370;
assign addr[5880] = 1918775195;
assign addr[5881] = 1910111873;
assign addr[5882] = 1901297091;
assign addr[5883] = 1892331547;
assign addr[5884] = 1883215953;
assign addr[5885] = 1873951032;
assign addr[5886] = 1864537518;
assign addr[5887] = 1854976157;
assign addr[5888] = 1845267708;
assign addr[5889] = 1835412941;
assign addr[5890] = 1825412636;
assign addr[5891] = 1815267588;
assign addr[5892] = 1804978599;
assign addr[5893] = 1794546487;
assign addr[5894] = 1783972079;
assign addr[5895] = 1773256212;
assign addr[5896] = 1762399737;
assign addr[5897] = 1751403515;
assign addr[5898] = 1740268417;
assign addr[5899] = 1728995326;
assign addr[5900] = 1717585136;
assign addr[5901] = 1706038753;
assign addr[5902] = 1694357091;
assign addr[5903] = 1682541077;
assign addr[5904] = 1670591647;
assign addr[5905] = 1658509750;
assign addr[5906] = 1646296344;
assign addr[5907] = 1633952396;
assign addr[5908] = 1621478885;
assign addr[5909] = 1608876801;
assign addr[5910] = 1596147143;
assign addr[5911] = 1583290921;
assign addr[5912] = 1570309153;
assign addr[5913] = 1557202869;
assign addr[5914] = 1543973108;
assign addr[5915] = 1530620920;
assign addr[5916] = 1517147363;
assign addr[5917] = 1503553506;
assign addr[5918] = 1489840425;
assign addr[5919] = 1476009210;
assign addr[5920] = 1462060956;
assign addr[5921] = 1447996770;
assign addr[5922] = 1433817766;
assign addr[5923] = 1419525069;
assign addr[5924] = 1405119813;
assign addr[5925] = 1390603139;
assign addr[5926] = 1375976199;
assign addr[5927] = 1361240152;
assign addr[5928] = 1346396168;
assign addr[5929] = 1331445422;
assign addr[5930] = 1316389101;
assign addr[5931] = 1301228398;
assign addr[5932] = 1285964516;
assign addr[5933] = 1270598665;
assign addr[5934] = 1255132063;
assign addr[5935] = 1239565936;
assign addr[5936] = 1223901520;
assign addr[5937] = 1208140056;
assign addr[5938] = 1192282793;
assign addr[5939] = 1176330990;
assign addr[5940] = 1160285911;
assign addr[5941] = 1144148829;
assign addr[5942] = 1127921022;
assign addr[5943] = 1111603778;
assign addr[5944] = 1095198391;
assign addr[5945] = 1078706161;
assign addr[5946] = 1062128397;
assign addr[5947] = 1045466412;
assign addr[5948] = 1028721528;
assign addr[5949] = 1011895073;
assign addr[5950] = 994988380;
assign addr[5951] = 978002791;
assign addr[5952] = 960939653;
assign addr[5953] = 943800318;
assign addr[5954] = 926586145;
assign addr[5955] = 909298500;
assign addr[5956] = 891938752;
assign addr[5957] = 874508280;
assign addr[5958] = 857008464;
assign addr[5959] = 839440693;
assign addr[5960] = 821806359;
assign addr[5961] = 804106861;
assign addr[5962] = 786343603;
assign addr[5963] = 768517992;
assign addr[5964] = 750631442;
assign addr[5965] = 732685372;
assign addr[5966] = 714681204;
assign addr[5967] = 696620367;
assign addr[5968] = 678504291;
assign addr[5969] = 660334415;
assign addr[5970] = 642112178;
assign addr[5971] = 623839025;
assign addr[5972] = 605516406;
assign addr[5973] = 587145773;
assign addr[5974] = 568728583;
assign addr[5975] = 550266296;
assign addr[5976] = 531760377;
assign addr[5977] = 513212292;
assign addr[5978] = 494623513;
assign addr[5979] = 475995513;
assign addr[5980] = 457329769;
assign addr[5981] = 438627762;
assign addr[5982] = 419890975;
assign addr[5983] = 401120892;
assign addr[5984] = 382319004;
assign addr[5985] = 363486799;
assign addr[5986] = 344625773;
assign addr[5987] = 325737419;
assign addr[5988] = 306823237;
assign addr[5989] = 287884725;
assign addr[5990] = 268923386;
assign addr[5991] = 249940723;
assign addr[5992] = 230938242;
assign addr[5993] = 211917448;
assign addr[5994] = 192879850;
assign addr[5995] = 173826959;
assign addr[5996] = 154760284;
assign addr[5997] = 135681337;
assign addr[5998] = 116591632;
assign addr[5999] = 97492681;
assign addr[6000] = 78386000;
assign addr[6001] = 59273104;
assign addr[6002] = 40155507;
assign addr[6003] = 21034727;
assign addr[6004] = 1912278;
assign addr[6005] = -17210322;
assign addr[6006] = -36331557;
assign addr[6007] = -55449912;
assign addr[6008] = -74563870;
assign addr[6009] = -93671915;
assign addr[6010] = -112772533;
assign addr[6011] = -131864208;
assign addr[6012] = -150945428;
assign addr[6013] = -170014678;
assign addr[6014] = -189070447;
assign addr[6015] = -208111224;
assign addr[6016] = -227135500;
assign addr[6017] = -246141764;
assign addr[6018] = -265128512;
assign addr[6019] = -284094236;
assign addr[6020] = -303037433;
assign addr[6021] = -321956601;
assign addr[6022] = -340850240;
assign addr[6023] = -359716852;
assign addr[6024] = -378554940;
assign addr[6025] = -397363011;
assign addr[6026] = -416139574;
assign addr[6027] = -434883140;
assign addr[6028] = -453592221;
assign addr[6029] = -472265336;
assign addr[6030] = -490901003;
assign addr[6031] = -509497745;
assign addr[6032] = -528054086;
assign addr[6033] = -546568556;
assign addr[6034] = -565039687;
assign addr[6035] = -583466013;
assign addr[6036] = -601846074;
assign addr[6037] = -620178412;
assign addr[6038] = -638461574;
assign addr[6039] = -656694110;
assign addr[6040] = -674874574;
assign addr[6041] = -693001525;
assign addr[6042] = -711073524;
assign addr[6043] = -729089140;
assign addr[6044] = -747046944;
assign addr[6045] = -764945512;
assign addr[6046] = -782783424;
assign addr[6047] = -800559266;
assign addr[6048] = -818271628;
assign addr[6049] = -835919107;
assign addr[6050] = -853500302;
assign addr[6051] = -871013820;
assign addr[6052] = -888458272;
assign addr[6053] = -905832274;
assign addr[6054] = -923134450;
assign addr[6055] = -940363427;
assign addr[6056] = -957517838;
assign addr[6057] = -974596324;
assign addr[6058] = -991597531;
assign addr[6059] = -1008520110;
assign addr[6060] = -1025362720;
assign addr[6061] = -1042124025;
assign addr[6062] = -1058802695;
assign addr[6063] = -1075397409;
assign addr[6064] = -1091906851;
assign addr[6065] = -1108329711;
assign addr[6066] = -1124664687;
assign addr[6067] = -1140910484;
assign addr[6068] = -1157065814;
assign addr[6069] = -1173129396;
assign addr[6070] = -1189099956;
assign addr[6071] = -1204976227;
assign addr[6072] = -1220756951;
assign addr[6073] = -1236440877;
assign addr[6074] = -1252026760;
assign addr[6075] = -1267513365;
assign addr[6076] = -1282899464;
assign addr[6077] = -1298183838;
assign addr[6078] = -1313365273;
assign addr[6079] = -1328442566;
assign addr[6080] = -1343414522;
assign addr[6081] = -1358279953;
assign addr[6082] = -1373037681;
assign addr[6083] = -1387686535;
assign addr[6084] = -1402225355;
assign addr[6085] = -1416652986;
assign addr[6086] = -1430968286;
assign addr[6087] = -1445170118;
assign addr[6088] = -1459257358;
assign addr[6089] = -1473228887;
assign addr[6090] = -1487083598;
assign addr[6091] = -1500820393;
assign addr[6092] = -1514438181;
assign addr[6093] = -1527935884;
assign addr[6094] = -1541312431;
assign addr[6095] = -1554566762;
assign addr[6096] = -1567697824;
assign addr[6097] = -1580704578;
assign addr[6098] = -1593585992;
assign addr[6099] = -1606341043;
assign addr[6100] = -1618968722;
assign addr[6101] = -1631468027;
assign addr[6102] = -1643837966;
assign addr[6103] = -1656077559;
assign addr[6104] = -1668185835;
assign addr[6105] = -1680161834;
assign addr[6106] = -1692004606;
assign addr[6107] = -1703713213;
assign addr[6108] = -1715286726;
assign addr[6109] = -1726724227;
assign addr[6110] = -1738024810;
assign addr[6111] = -1749187577;
assign addr[6112] = -1760211645;
assign addr[6113] = -1771096139;
assign addr[6114] = -1781840195;
assign addr[6115] = -1792442963;
assign addr[6116] = -1802903601;
assign addr[6117] = -1813221279;
assign addr[6118] = -1823395180;
assign addr[6119] = -1833424497;
assign addr[6120] = -1843308435;
assign addr[6121] = -1853046210;
assign addr[6122] = -1862637049;
assign addr[6123] = -1872080193;
assign addr[6124] = -1881374892;
assign addr[6125] = -1890520410;
assign addr[6126] = -1899516021;
assign addr[6127] = -1908361011;
assign addr[6128] = -1917054681;
assign addr[6129] = -1925596340;
assign addr[6130] = -1933985310;
assign addr[6131] = -1942220928;
assign addr[6132] = -1950302539;
assign addr[6133] = -1958229503;
assign addr[6134] = -1966001192;
assign addr[6135] = -1973616989;
assign addr[6136] = -1981076290;
assign addr[6137] = -1988378503;
assign addr[6138] = -1995523051;
assign addr[6139] = -2002509365;
assign addr[6140] = -2009336893;
assign addr[6141] = -2016005093;
assign addr[6142] = -2022513436;
assign addr[6143] = -2028861406;
assign addr[6144] = -2035048499;
assign addr[6145] = -2041074226;
assign addr[6146] = -2046938108;
assign addr[6147] = -2052639680;
assign addr[6148] = -2058178491;
assign addr[6149] = -2063554100;
assign addr[6150] = -2068766083;
assign addr[6151] = -2073814024;
assign addr[6152] = -2078697525;
assign addr[6153] = -2083416198;
assign addr[6154] = -2087969669;
assign addr[6155] = -2092357577;
assign addr[6156] = -2096579573;
assign addr[6157] = -2100635323;
assign addr[6158] = -2104524506;
assign addr[6159] = -2108246813;
assign addr[6160] = -2111801949;
assign addr[6161] = -2115189632;
assign addr[6162] = -2118409593;
assign addr[6163] = -2121461578;
assign addr[6164] = -2124345343;
assign addr[6165] = -2127060661;
assign addr[6166] = -2129607316;
assign addr[6167] = -2131985106;
assign addr[6168] = -2134193842;
assign addr[6169] = -2136233350;
assign addr[6170] = -2138103468;
assign addr[6171] = -2139804048;
assign addr[6172] = -2141334954;
assign addr[6173] = -2142696065;
assign addr[6174] = -2143887273;
assign addr[6175] = -2144908484;
assign addr[6176] = -2145759618;
assign addr[6177] = -2146440605;
assign addr[6178] = -2146951393;
assign addr[6179] = -2147291941;
assign addr[6180] = -2147462221;
assign addr[6181] = -2147462221;
assign addr[6182] = -2147291941;
assign addr[6183] = -2146951393;
assign addr[6184] = -2146440605;
assign addr[6185] = -2145759618;
assign addr[6186] = -2144908484;
assign addr[6187] = -2143887273;
assign addr[6188] = -2142696065;
assign addr[6189] = -2141334954;
assign addr[6190] = -2139804048;
assign addr[6191] = -2138103468;
assign addr[6192] = -2136233350;
assign addr[6193] = -2134193842;
assign addr[6194] = -2131985106;
assign addr[6195] = -2129607316;
assign addr[6196] = -2127060661;
assign addr[6197] = -2124345343;
assign addr[6198] = -2121461578;
assign addr[6199] = -2118409593;
assign addr[6200] = -2115189632;
assign addr[6201] = -2111801949;
assign addr[6202] = -2108246813;
assign addr[6203] = -2104524506;
assign addr[6204] = -2100635323;
assign addr[6205] = -2096579573;
assign addr[6206] = -2092357577;
assign addr[6207] = -2087969669;
assign addr[6208] = -2083416198;
assign addr[6209] = -2078697525;
assign addr[6210] = -2073814024;
assign addr[6211] = -2068766083;
assign addr[6212] = -2063554100;
assign addr[6213] = -2058178491;
assign addr[6214] = -2052639680;
assign addr[6215] = -2046938108;
assign addr[6216] = -2041074226;
assign addr[6217] = -2035048499;
assign addr[6218] = -2028861406;
assign addr[6219] = -2022513436;
assign addr[6220] = -2016005093;
assign addr[6221] = -2009336893;
assign addr[6222] = -2002509365;
assign addr[6223] = -1995523051;
assign addr[6224] = -1988378503;
assign addr[6225] = -1981076290;
assign addr[6226] = -1973616989;
assign addr[6227] = -1966001192;
assign addr[6228] = -1958229503;
assign addr[6229] = -1950302539;
assign addr[6230] = -1942220928;
assign addr[6231] = -1933985310;
assign addr[6232] = -1925596340;
assign addr[6233] = -1917054681;
assign addr[6234] = -1908361011;
assign addr[6235] = -1899516021;
assign addr[6236] = -1890520410;
assign addr[6237] = -1881374892;
assign addr[6238] = -1872080193;
assign addr[6239] = -1862637049;
assign addr[6240] = -1853046210;
assign addr[6241] = -1843308435;
assign addr[6242] = -1833424497;
assign addr[6243] = -1823395180;
assign addr[6244] = -1813221279;
assign addr[6245] = -1802903601;
assign addr[6246] = -1792442963;
assign addr[6247] = -1781840195;
assign addr[6248] = -1771096139;
assign addr[6249] = -1760211645;
assign addr[6250] = -1749187577;
assign addr[6251] = -1738024810;
assign addr[6252] = -1726724227;
assign addr[6253] = -1715286726;
assign addr[6254] = -1703713213;
assign addr[6255] = -1692004606;
assign addr[6256] = -1680161834;
assign addr[6257] = -1668185835;
assign addr[6258] = -1656077559;
assign addr[6259] = -1643837966;
assign addr[6260] = -1631468027;
assign addr[6261] = -1618968722;
assign addr[6262] = -1606341043;
assign addr[6263] = -1593585992;
assign addr[6264] = -1580704578;
assign addr[6265] = -1567697824;
assign addr[6266] = -1554566762;
assign addr[6267] = -1541312431;
assign addr[6268] = -1527935884;
assign addr[6269] = -1514438181;
assign addr[6270] = -1500820393;
assign addr[6271] = -1487083598;
assign addr[6272] = -1473228887;
assign addr[6273] = -1459257358;
assign addr[6274] = -1445170118;
assign addr[6275] = -1430968286;
assign addr[6276] = -1416652986;
assign addr[6277] = -1402225355;
assign addr[6278] = -1387686535;
assign addr[6279] = -1373037681;
assign addr[6280] = -1358279953;
assign addr[6281] = -1343414522;
assign addr[6282] = -1328442566;
assign addr[6283] = -1313365273;
assign addr[6284] = -1298183838;
assign addr[6285] = -1282899464;
assign addr[6286] = -1267513365;
assign addr[6287] = -1252026760;
assign addr[6288] = -1236440877;
assign addr[6289] = -1220756951;
assign addr[6290] = -1204976227;
assign addr[6291] = -1189099956;
assign addr[6292] = -1173129396;
assign addr[6293] = -1157065814;
assign addr[6294] = -1140910484;
assign addr[6295] = -1124664687;
assign addr[6296] = -1108329711;
assign addr[6297] = -1091906851;
assign addr[6298] = -1075397409;
assign addr[6299] = -1058802695;
assign addr[6300] = -1042124025;
assign addr[6301] = -1025362720;
assign addr[6302] = -1008520110;
assign addr[6303] = -991597531;
assign addr[6304] = -974596324;
assign addr[6305] = -957517838;
assign addr[6306] = -940363427;
assign addr[6307] = -923134450;
assign addr[6308] = -905832274;
assign addr[6309] = -888458272;
assign addr[6310] = -871013820;
assign addr[6311] = -853500302;
assign addr[6312] = -835919107;
assign addr[6313] = -818271628;
assign addr[6314] = -800559266;
assign addr[6315] = -782783424;
assign addr[6316] = -764945512;
assign addr[6317] = -747046944;
assign addr[6318] = -729089140;
assign addr[6319] = -711073524;
assign addr[6320] = -693001525;
assign addr[6321] = -674874574;
assign addr[6322] = -656694110;
assign addr[6323] = -638461574;
assign addr[6324] = -620178412;
assign addr[6325] = -601846074;
assign addr[6326] = -583466013;
assign addr[6327] = -565039687;
assign addr[6328] = -546568556;
assign addr[6329] = -528054086;
assign addr[6330] = -509497745;
assign addr[6331] = -490901003;
assign addr[6332] = -472265336;
assign addr[6333] = -453592221;
assign addr[6334] = -434883140;
assign addr[6335] = -416139574;
assign addr[6336] = -397363011;
assign addr[6337] = -378554940;
assign addr[6338] = -359716852;
assign addr[6339] = -340850240;
assign addr[6340] = -321956601;
assign addr[6341] = -303037433;
assign addr[6342] = -284094236;
assign addr[6343] = -265128512;
assign addr[6344] = -246141764;
assign addr[6345] = -227135500;
assign addr[6346] = -208111224;
assign addr[6347] = -189070447;
assign addr[6348] = -170014678;
assign addr[6349] = -150945428;
assign addr[6350] = -131864208;
assign addr[6351] = -112772533;
assign addr[6352] = -93671915;
assign addr[6353] = -74563870;
assign addr[6354] = -55449912;
assign addr[6355] = -36331557;
assign addr[6356] = -17210322;
assign addr[6357] = 1912278;
assign addr[6358] = 21034727;
assign addr[6359] = 40155507;
assign addr[6360] = 59273104;
assign addr[6361] = 78386000;
assign addr[6362] = 97492681;
assign addr[6363] = 116591632;
assign addr[6364] = 135681337;
assign addr[6365] = 154760284;
assign addr[6366] = 173826959;
assign addr[6367] = 192879850;
assign addr[6368] = 211917448;
assign addr[6369] = 230938242;
assign addr[6370] = 249940723;
assign addr[6371] = 268923386;
assign addr[6372] = 287884725;
assign addr[6373] = 306823237;
assign addr[6374] = 325737419;
assign addr[6375] = 344625773;
assign addr[6376] = 363486799;
assign addr[6377] = 382319004;
assign addr[6378] = 401120892;
assign addr[6379] = 419890975;
assign addr[6380] = 438627762;
assign addr[6381] = 457329769;
assign addr[6382] = 475995513;
assign addr[6383] = 494623513;
assign addr[6384] = 513212292;
assign addr[6385] = 531760377;
assign addr[6386] = 550266296;
assign addr[6387] = 568728583;
assign addr[6388] = 587145773;
assign addr[6389] = 605516406;
assign addr[6390] = 623839025;
assign addr[6391] = 642112178;
assign addr[6392] = 660334415;
assign addr[6393] = 678504291;
assign addr[6394] = 696620367;
assign addr[6395] = 714681204;
assign addr[6396] = 732685372;
assign addr[6397] = 750631442;
assign addr[6398] = 768517992;
assign addr[6399] = 786343603;
assign addr[6400] = 804106861;
assign addr[6401] = 821806359;
assign addr[6402] = 839440693;
assign addr[6403] = 857008464;
assign addr[6404] = 874508280;
assign addr[6405] = 891938752;
assign addr[6406] = 909298500;
assign addr[6407] = 926586145;
assign addr[6408] = 943800318;
assign addr[6409] = 960939653;
assign addr[6410] = 978002791;
assign addr[6411] = 994988380;
assign addr[6412] = 1011895073;
assign addr[6413] = 1028721528;
assign addr[6414] = 1045466412;
assign addr[6415] = 1062128397;
assign addr[6416] = 1078706161;
assign addr[6417] = 1095198391;
assign addr[6418] = 1111603778;
assign addr[6419] = 1127921022;
assign addr[6420] = 1144148829;
assign addr[6421] = 1160285911;
assign addr[6422] = 1176330990;
assign addr[6423] = 1192282793;
assign addr[6424] = 1208140056;
assign addr[6425] = 1223901520;
assign addr[6426] = 1239565936;
assign addr[6427] = 1255132063;
assign addr[6428] = 1270598665;
assign addr[6429] = 1285964516;
assign addr[6430] = 1301228398;
assign addr[6431] = 1316389101;
assign addr[6432] = 1331445422;
assign addr[6433] = 1346396168;
assign addr[6434] = 1361240152;
assign addr[6435] = 1375976199;
assign addr[6436] = 1390603139;
assign addr[6437] = 1405119813;
assign addr[6438] = 1419525069;
assign addr[6439] = 1433817766;
assign addr[6440] = 1447996770;
assign addr[6441] = 1462060956;
assign addr[6442] = 1476009210;
assign addr[6443] = 1489840425;
assign addr[6444] = 1503553506;
assign addr[6445] = 1517147363;
assign addr[6446] = 1530620920;
assign addr[6447] = 1543973108;
assign addr[6448] = 1557202869;
assign addr[6449] = 1570309153;
assign addr[6450] = 1583290921;
assign addr[6451] = 1596147143;
assign addr[6452] = 1608876801;
assign addr[6453] = 1621478885;
assign addr[6454] = 1633952396;
assign addr[6455] = 1646296344;
assign addr[6456] = 1658509750;
assign addr[6457] = 1670591647;
assign addr[6458] = 1682541077;
assign addr[6459] = 1694357091;
assign addr[6460] = 1706038753;
assign addr[6461] = 1717585136;
assign addr[6462] = 1728995326;
assign addr[6463] = 1740268417;
assign addr[6464] = 1751403515;
assign addr[6465] = 1762399737;
assign addr[6466] = 1773256212;
assign addr[6467] = 1783972079;
assign addr[6468] = 1794546487;
assign addr[6469] = 1804978599;
assign addr[6470] = 1815267588;
assign addr[6471] = 1825412636;
assign addr[6472] = 1835412941;
assign addr[6473] = 1845267708;
assign addr[6474] = 1854976157;
assign addr[6475] = 1864537518;
assign addr[6476] = 1873951032;
assign addr[6477] = 1883215953;
assign addr[6478] = 1892331547;
assign addr[6479] = 1901297091;
assign addr[6480] = 1910111873;
assign addr[6481] = 1918775195;
assign addr[6482] = 1927286370;
assign addr[6483] = 1935644723;
assign addr[6484] = 1943849591;
assign addr[6485] = 1951900324;
assign addr[6486] = 1959796283;
assign addr[6487] = 1967536842;
assign addr[6488] = 1975121388;
assign addr[6489] = 1982549318;
assign addr[6490] = 1989820044;
assign addr[6491] = 1996932990;
assign addr[6492] = 2003887591;
assign addr[6493] = 2010683297;
assign addr[6494] = 2017319567;
assign addr[6495] = 2023795876;
assign addr[6496] = 2030111710;
assign addr[6497] = 2036266570;
assign addr[6498] = 2042259965;
assign addr[6499] = 2048091422;
assign addr[6500] = 2053760478;
assign addr[6501] = 2059266683;
assign addr[6502] = 2064609600;
assign addr[6503] = 2069788807;
assign addr[6504] = 2074803892;
assign addr[6505] = 2079654458;
assign addr[6506] = 2084340120;
assign addr[6507] = 2088860507;
assign addr[6508] = 2093215260;
assign addr[6509] = 2097404033;
assign addr[6510] = 2101426496;
assign addr[6511] = 2105282327;
assign addr[6512] = 2108971223;
assign addr[6513] = 2112492891;
assign addr[6514] = 2115847050;
assign addr[6515] = 2119033436;
assign addr[6516] = 2122051796;
assign addr[6517] = 2124901890;
assign addr[6518] = 2127583492;
assign addr[6519] = 2130096389;
assign addr[6520] = 2132440383;
assign addr[6521] = 2134615288;
assign addr[6522] = 2136620930;
assign addr[6523] = 2138457152;
assign addr[6524] = 2140123807;
assign addr[6525] = 2141620763;
assign addr[6526] = 2142947902;
assign addr[6527] = 2144105118;
assign addr[6528] = 2145092320;
assign addr[6529] = 2145909429;
assign addr[6530] = 2146556380;
assign addr[6531] = 2147033123;
assign addr[6532] = 2147339619;
assign addr[6533] = 2147475844;
assign addr[6534] = 2147441787;
assign addr[6535] = 2147237452;
assign addr[6536] = 2146862854;
assign addr[6537] = 2146318022;
assign addr[6538] = 2145603001;
assign addr[6539] = 2144717846;
assign addr[6540] = 2143662628;
assign addr[6541] = 2142437431;
assign addr[6542] = 2141042352;
assign addr[6543] = 2139477502;
assign addr[6544] = 2137743003;
assign addr[6545] = 2135838995;
assign addr[6546] = 2133765628;
assign addr[6547] = 2131523066;
assign addr[6548] = 2129111488;
assign addr[6549] = 2126531084;
assign addr[6550] = 2123782059;
assign addr[6551] = 2120864631;
assign addr[6552] = 2117779031;
assign addr[6553] = 2114525505;
assign addr[6554] = 2111104309;
assign addr[6555] = 2107515716;
assign addr[6556] = 2103760010;
assign addr[6557] = 2099837489;
assign addr[6558] = 2095748463;
assign addr[6559] = 2091493257;
assign addr[6560] = 2087072209;
assign addr[6561] = 2082485668;
assign addr[6562] = 2077733999;
assign addr[6563] = 2072817579;
assign addr[6564] = 2067736796;
assign addr[6565] = 2062492055;
assign addr[6566] = 2057083771;
assign addr[6567] = 2051512372;
assign addr[6568] = 2045778302;
assign addr[6569] = 2039882013;
assign addr[6570] = 2033823974;
assign addr[6571] = 2027604666;
assign addr[6572] = 2021224581;
assign addr[6573] = 2014684225;
assign addr[6574] = 2007984117;
assign addr[6575] = 2001124788;
assign addr[6576] = 1994106782;
assign addr[6577] = 1986930656;
assign addr[6578] = 1979596978;
assign addr[6579] = 1972106330;
assign addr[6580] = 1964459306;
assign addr[6581] = 1956656513;
assign addr[6582] = 1948698568;
assign addr[6583] = 1940586104;
assign addr[6584] = 1932319763;
assign addr[6585] = 1923900201;
assign addr[6586] = 1915328086;
assign addr[6587] = 1906604097;
assign addr[6588] = 1897728925;
assign addr[6589] = 1888703276;
assign addr[6590] = 1879527863;
assign addr[6591] = 1870203416;
assign addr[6592] = 1860730673;
assign addr[6593] = 1851110385;
assign addr[6594] = 1841343316;
assign addr[6595] = 1831430239;
assign addr[6596] = 1821371941;
assign addr[6597] = 1811169220;
assign addr[6598] = 1800822883;
assign addr[6599] = 1790333753;
assign addr[6600] = 1779702660;
assign addr[6601] = 1768930447;
assign addr[6602] = 1758017969;
assign addr[6603] = 1746966091;
assign addr[6604] = 1735775690;
assign addr[6605] = 1724447652;
assign addr[6606] = 1712982875;
assign addr[6607] = 1701382270;
assign addr[6608] = 1689646755;
assign addr[6609] = 1677777262;
assign addr[6610] = 1665774731;
assign addr[6611] = 1653640115;
assign addr[6612] = 1641374375;
assign addr[6613] = 1628978484;
assign addr[6614] = 1616453425;
assign addr[6615] = 1603800191;
assign addr[6616] = 1591019785;
assign addr[6617] = 1578113222;
assign addr[6618] = 1565081523;
assign addr[6619] = 1551925723;
assign addr[6620] = 1538646865;
assign addr[6621] = 1525246002;
assign addr[6622] = 1511724196;
assign addr[6623] = 1498082520;
assign addr[6624] = 1484322054;
assign addr[6625] = 1470443891;
assign addr[6626] = 1456449131;
assign addr[6627] = 1442338884;
assign addr[6628] = 1428114267;
assign addr[6629] = 1413776410;
assign addr[6630] = 1399326449;
assign addr[6631] = 1384765530;
assign addr[6632] = 1370094808;
assign addr[6633] = 1355315445;
assign addr[6634] = 1340428615;
assign addr[6635] = 1325435496;
assign addr[6636] = 1310337279;
assign addr[6637] = 1295135159;
assign addr[6638] = 1279830344;
assign addr[6639] = 1264424045;
assign addr[6640] = 1248917486;
assign addr[6641] = 1233311895;
assign addr[6642] = 1217608510;
assign addr[6643] = 1201808576;
assign addr[6644] = 1185913346;
assign addr[6645] = 1169924081;
assign addr[6646] = 1153842047;
assign addr[6647] = 1137668521;
assign addr[6648] = 1121404785;
assign addr[6649] = 1105052128;
assign addr[6650] = 1088611847;
assign addr[6651] = 1072085246;
assign addr[6652] = 1055473635;
assign addr[6653] = 1038778332;
assign addr[6654] = 1022000660;
assign addr[6655] = 1005141949;
assign addr[6656] = 988203537;
assign addr[6657] = 971186766;
assign addr[6658] = 954092986;
assign addr[6659] = 936923553;
assign addr[6660] = 919679827;
assign addr[6661] = 902363176;
assign addr[6662] = 884974973;
assign addr[6663] = 867516597;
assign addr[6664] = 849989433;
assign addr[6665] = 832394869;
assign addr[6666] = 814734301;
assign addr[6667] = 797009130;
assign addr[6668] = 779220762;
assign addr[6669] = 761370605;
assign addr[6670] = 743460077;
assign addr[6671] = 725490597;
assign addr[6672] = 707463589;
assign addr[6673] = 689380485;
assign addr[6674] = 671242716;
assign addr[6675] = 653051723;
assign addr[6676] = 634808946;
assign addr[6677] = 616515832;
assign addr[6678] = 598173833;
assign addr[6679] = 579784402;
assign addr[6680] = 561348998;
assign addr[6681] = 542869083;
assign addr[6682] = 524346121;
assign addr[6683] = 505781581;
assign addr[6684] = 487176937;
assign addr[6685] = 468533662;
assign addr[6686] = 449853235;
assign addr[6687] = 431137138;
assign addr[6688] = 412386854;
assign addr[6689] = 393603870;
assign addr[6690] = 374789676;
assign addr[6691] = 355945764;
assign addr[6692] = 337073627;
assign addr[6693] = 318174762;
assign addr[6694] = 299250668;
assign addr[6695] = 280302845;
assign addr[6696] = 261332796;
assign addr[6697] = 242342025;
assign addr[6698] = 223332037;
assign addr[6699] = 204304341;
assign addr[6700] = 185260444;
assign addr[6701] = 166201858;
assign addr[6702] = 147130093;
assign addr[6703] = 128046661;
assign addr[6704] = 108953076;
assign addr[6705] = 89850852;
assign addr[6706] = 70741503;
assign addr[6707] = 51626544;
assign addr[6708] = 32507492;
assign addr[6709] = 13385863;
assign addr[6710] = -5736829;
assign addr[6711] = -24859065;
assign addr[6712] = -43979330;
assign addr[6713] = -63096108;
assign addr[6714] = -82207882;
assign addr[6715] = -101313138;
assign addr[6716] = -120410361;
assign addr[6717] = -139498035;
assign addr[6718] = -158574649;
assign addr[6719] = -177638688;
assign addr[6720] = -196688642;
assign addr[6721] = -215722999;
assign addr[6722] = -234740251;
assign addr[6723] = -253738890;
assign addr[6724] = -272717408;
assign addr[6725] = -291674302;
assign addr[6726] = -310608068;
assign addr[6727] = -329517204;
assign addr[6728] = -348400212;
assign addr[6729] = -367255594;
assign addr[6730] = -386081854;
assign addr[6731] = -404877501;
assign addr[6732] = -423641043;
assign addr[6733] = -442370993;
assign addr[6734] = -461065866;
assign addr[6735] = -479724180;
assign addr[6736] = -498344454;
assign addr[6737] = -516925212;
assign addr[6738] = -535464981;
assign addr[6739] = -553962291;
assign addr[6740] = -572415676;
assign addr[6741] = -590823671;
assign addr[6742] = -609184818;
assign addr[6743] = -627497660;
assign addr[6744] = -645760745;
assign addr[6745] = -663972625;
assign addr[6746] = -682131857;
assign addr[6747] = -700236999;
assign addr[6748] = -718286617;
assign addr[6749] = -736279279;
assign addr[6750] = -754213559;
assign addr[6751] = -772088034;
assign addr[6752] = -789901288;
assign addr[6753] = -807651907;
assign addr[6754] = -825338484;
assign addr[6755] = -842959617;
assign addr[6756] = -860513908;
assign addr[6757] = -877999966;
assign addr[6758] = -895416404;
assign addr[6759] = -912761841;
assign addr[6760] = -930034901;
assign addr[6761] = -947234215;
assign addr[6762] = -964358420;
assign addr[6763] = -981406156;
assign addr[6764] = -998376073;
assign addr[6765] = -1015266825;
assign addr[6766] = -1032077073;
assign addr[6767] = -1048805483;
assign addr[6768] = -1065450729;
assign addr[6769] = -1082011492;
assign addr[6770] = -1098486458;
assign addr[6771] = -1114874320;
assign addr[6772] = -1131173780;
assign addr[6773] = -1147383544;
assign addr[6774] = -1163502328;
assign addr[6775] = -1179528853;
assign addr[6776] = -1195461849;
assign addr[6777] = -1211300053;
assign addr[6778] = -1227042207;
assign addr[6779] = -1242687064;
assign addr[6780] = -1258233384;
assign addr[6781] = -1273679934;
assign addr[6782] = -1289025489;
assign addr[6783] = -1304268832;
assign addr[6784] = -1319408754;
assign addr[6785] = -1334444055;
assign addr[6786] = -1349373543;
assign addr[6787] = -1364196034;
assign addr[6788] = -1378910353;
assign addr[6789] = -1393515332;
assign addr[6790] = -1408009814;
assign addr[6791] = -1422392650;
assign addr[6792] = -1436662698;
assign addr[6793] = -1450818828;
assign addr[6794] = -1464859917;
assign addr[6795] = -1478784851;
assign addr[6796] = -1492592527;
assign addr[6797] = -1506281850;
assign addr[6798] = -1519851733;
assign addr[6799] = -1533301101;
assign addr[6800] = -1546628888;
assign addr[6801] = -1559834037;
assign addr[6802] = -1572915501;
assign addr[6803] = -1585872242;
assign addr[6804] = -1598703233;
assign addr[6805] = -1611407456;
assign addr[6806] = -1623983905;
assign addr[6807] = -1636431582;
assign addr[6808] = -1648749499;
assign addr[6809] = -1660936681;
assign addr[6810] = -1672992161;
assign addr[6811] = -1684914983;
assign addr[6812] = -1696704201;
assign addr[6813] = -1708358881;
assign addr[6814] = -1719878099;
assign addr[6815] = -1731260941;
assign addr[6816] = -1742506504;
assign addr[6817] = -1753613897;
assign addr[6818] = -1764582240;
assign addr[6819] = -1775410662;
assign addr[6820] = -1786098304;
assign addr[6821] = -1796644320;
assign addr[6822] = -1807047873;
assign addr[6823] = -1817308138;
assign addr[6824] = -1827424302;
assign addr[6825] = -1837395562;
assign addr[6826] = -1847221128;
assign addr[6827] = -1856900221;
assign addr[6828] = -1866432072;
assign addr[6829] = -1875815927;
assign addr[6830] = -1885051042;
assign addr[6831] = -1894136683;
assign addr[6832] = -1903072131;
assign addr[6833] = -1911856677;
assign addr[6834] = -1920489624;
assign addr[6835] = -1928970288;
assign addr[6836] = -1937297997;
assign addr[6837] = -1945472089;
assign addr[6838] = -1953491918;
assign addr[6839] = -1961356847;
assign addr[6840] = -1969066252;
assign addr[6841] = -1976619522;
assign addr[6842] = -1984016058;
assign addr[6843] = -1991255274;
assign addr[6844] = -1998336596;
assign addr[6845] = -2005259462;
assign addr[6846] = -2012023322;
assign addr[6847] = -2018627642;
assign addr[6848] = -2025071897;
assign addr[6849] = -2031355576;
assign addr[6850] = -2037478181;
assign addr[6851] = -2043439226;
assign addr[6852] = -2049238240;
assign addr[6853] = -2054874761;
assign addr[6854] = -2060348343;
assign addr[6855] = -2065658552;
assign addr[6856] = -2070804967;
assign addr[6857] = -2075787180;
assign addr[6858] = -2080604795;
assign addr[6859] = -2085257431;
assign addr[6860] = -2089744719;
assign addr[6861] = -2094066304;
assign addr[6862] = -2098221841;
assign addr[6863] = -2102211002;
assign addr[6864] = -2106033471;
assign addr[6865] = -2109688944;
assign addr[6866] = -2113177132;
assign addr[6867] = -2116497758;
assign addr[6868] = -2119650558;
assign addr[6869] = -2122635283;
assign addr[6870] = -2125451696;
assign addr[6871] = -2128099574;
assign addr[6872] = -2130578706;
assign addr[6873] = -2132888897;
assign addr[6874] = -2135029962;
assign addr[6875] = -2137001733;
assign addr[6876] = -2138804053;
assign addr[6877] = -2140436778;
assign addr[6878] = -2141899780;
assign addr[6879] = -2143192942;
assign addr[6880] = -2144316162;
assign addr[6881] = -2145269351;
assign addr[6882] = -2146052433;
assign addr[6883] = -2146665347;
assign addr[6884] = -2147108043;
assign addr[6885] = -2147380486;
assign addr[6886] = -2147482655;
assign addr[6887] = -2147414542;
assign addr[6888] = -2147176152;
assign addr[6889] = -2146767505;
assign addr[6890] = -2146188631;
assign addr[6891] = -2145439578;
assign addr[6892] = -2144520405;
assign addr[6893] = -2143431184;
assign addr[6894] = -2142172003;
assign addr[6895] = -2140742960;
assign addr[6896] = -2139144169;
assign addr[6897] = -2137375758;
assign addr[6898] = -2135437865;
assign addr[6899] = -2133330646;
assign addr[6900] = -2131054266;
assign addr[6901] = -2128608907;
assign addr[6902] = -2125994762;
assign addr[6903] = -2123212038;
assign addr[6904] = -2120260957;
assign addr[6905] = -2117141752;
assign addr[6906] = -2113854671;
assign addr[6907] = -2110399974;
assign addr[6908] = -2106777935;
assign addr[6909] = -2102988841;
assign addr[6910] = -2099032994;
assign addr[6911] = -2094910706;
assign addr[6912] = -2090622304;
assign addr[6913] = -2086168128;
assign addr[6914] = -2081548533;
assign addr[6915] = -2076763883;
assign addr[6916] = -2071814558;
assign addr[6917] = -2066700952;
assign addr[6918] = -2061423468;
assign addr[6919] = -2055982526;
assign addr[6920] = -2050378558;
assign addr[6921] = -2044612007;
assign addr[6922] = -2038683330;
assign addr[6923] = -2032592999;
assign addr[6924] = -2026341495;
assign addr[6925] = -2019929315;
assign addr[6926] = -2013356967;
assign addr[6927] = -2006624971;
assign addr[6928] = -1999733863;
assign addr[6929] = -1992684188;
assign addr[6930] = -1985476506;
assign addr[6931] = -1978111387;
assign addr[6932] = -1970589416;
assign addr[6933] = -1962911189;
assign addr[6934] = -1955077316;
assign addr[6935] = -1947088417;
assign addr[6936] = -1938945125;
assign addr[6937] = -1930648088;
assign addr[6938] = -1922197961;
assign addr[6939] = -1913595416;
assign addr[6940] = -1904841135;
assign addr[6941] = -1895935811;
assign addr[6942] = -1886880151;
assign addr[6943] = -1877674873;
assign addr[6944] = -1868320707;
assign addr[6945] = -1858818395;
assign addr[6946] = -1849168689;
assign addr[6947] = -1839372356;
assign addr[6948] = -1829430172;
assign addr[6949] = -1819342925;
assign addr[6950] = -1809111415;
assign addr[6951] = -1798736454;
assign addr[6952] = -1788218865;
assign addr[6953] = -1777559480;
assign addr[6954] = -1766759146;
assign addr[6955] = -1755818718;
assign addr[6956] = -1744739065;
assign addr[6957] = -1733521064;
assign addr[6958] = -1722165606;
assign addr[6959] = -1710673591;
assign addr[6960] = -1699045930;
assign addr[6961] = -1687283545;
assign addr[6962] = -1675387369;
assign addr[6963] = -1663358344;
assign addr[6964] = -1651197426;
assign addr[6965] = -1638905577;
assign addr[6966] = -1626483774;
assign addr[6967] = -1613933000;
assign addr[6968] = -1601254251;
assign addr[6969] = -1588448533;
assign addr[6970] = -1575516860;
assign addr[6971] = -1562460258;
assign addr[6972] = -1549279763;
assign addr[6973] = -1535976419;
assign addr[6974] = -1522551282;
assign addr[6975] = -1509005416;
assign addr[6976] = -1495339895;
assign addr[6977] = -1481555802;
assign addr[6978] = -1467654232;
assign addr[6979] = -1453636285;
assign addr[6980] = -1439503074;
assign addr[6981] = -1425255719;
assign addr[6982] = -1410895350;
assign addr[6983] = -1396423105;
assign addr[6984] = -1381840133;
assign addr[6985] = -1367147589;
assign addr[6986] = -1352346639;
assign addr[6987] = -1337438456;
assign addr[6988] = -1322424222;
assign addr[6989] = -1307305128;
assign addr[6990] = -1292082373;
assign addr[6991] = -1276757164;
assign addr[6992] = -1261330715;
assign addr[6993] = -1245804251;
assign addr[6994] = -1230179002;
assign addr[6995] = -1214456207;
assign addr[6996] = -1198637114;
assign addr[6997] = -1182722976;
assign addr[6998] = -1166715055;
assign addr[6999] = -1150614620;
assign addr[7000] = -1134422949;
assign addr[7001] = -1118141326;
assign addr[7002] = -1101771040;
assign addr[7003] = -1085313391;
assign addr[7004] = -1068769683;
assign addr[7005] = -1052141228;
assign addr[7006] = -1035429345;
assign addr[7007] = -1018635358;
assign addr[7008] = -1001760600;
assign addr[7009] = -984806408;
assign addr[7010] = -967774128;
assign addr[7011] = -950665109;
assign addr[7012] = -933480707;
assign addr[7013] = -916222287;
assign addr[7014] = -898891215;
assign addr[7015] = -881488868;
assign addr[7016] = -864016623;
assign addr[7017] = -846475867;
assign addr[7018] = -828867991;
assign addr[7019] = -811194391;
assign addr[7020] = -793456467;
assign addr[7021] = -775655628;
assign addr[7022] = -757793284;
assign addr[7023] = -739870851;
assign addr[7024] = -721889752;
assign addr[7025] = -703851410;
assign addr[7026] = -685757258;
assign addr[7027] = -667608730;
assign addr[7028] = -649407264;
assign addr[7029] = -631154304;
assign addr[7030] = -612851297;
assign addr[7031] = -594499695;
assign addr[7032] = -576100953;
assign addr[7033] = -557656529;
assign addr[7034] = -539167887;
assign addr[7035] = -520636492;
assign addr[7036] = -502063814;
assign addr[7037] = -483451325;
assign addr[7038] = -464800501;
assign addr[7039] = -446112822;
assign addr[7040] = -427389768;
assign addr[7041] = -408632825;
assign addr[7042] = -389843480;
assign addr[7043] = -371023223;
assign addr[7044] = -352173546;
assign addr[7045] = -333295944;
assign addr[7046] = -314391913;
assign addr[7047] = -295462954;
assign addr[7048] = -276510565;
assign addr[7049] = -257536251;
assign addr[7050] = -238541516;
assign addr[7051] = -219527866;
assign addr[7052] = -200496809;
assign addr[7053] = -181449854;
assign addr[7054] = -162388511;
assign addr[7055] = -143314291;
assign addr[7056] = -124228708;
assign addr[7057] = -105133274;
assign addr[7058] = -86029503;
assign addr[7059] = -66918911;
assign addr[7060] = -47803013;
assign addr[7061] = -28683324;
assign addr[7062] = -9561361;
assign addr[7063] = 9561361;
assign addr[7064] = 28683324;
assign addr[7065] = 47803013;
assign addr[7066] = 66918911;
assign addr[7067] = 86029503;
assign addr[7068] = 105133274;
assign addr[7069] = 124228708;
assign addr[7070] = 143314291;
assign addr[7071] = 162388511;
assign addr[7072] = 181449854;
assign addr[7073] = 200496809;
assign addr[7074] = 219527866;
assign addr[7075] = 238541516;
assign addr[7076] = 257536251;
assign addr[7077] = 276510565;
assign addr[7078] = 295462954;
assign addr[7079] = 314391913;
assign addr[7080] = 333295944;
assign addr[7081] = 352173546;
assign addr[7082] = 371023223;
assign addr[7083] = 389843480;
assign addr[7084] = 408632825;
assign addr[7085] = 427389768;
assign addr[7086] = 446112822;
assign addr[7087] = 464800501;
assign addr[7088] = 483451325;
assign addr[7089] = 502063814;
assign addr[7090] = 520636492;
assign addr[7091] = 539167887;
assign addr[7092] = 557656529;
assign addr[7093] = 576100953;
assign addr[7094] = 594499695;
assign addr[7095] = 612851297;
assign addr[7096] = 631154304;
assign addr[7097] = 649407264;
assign addr[7098] = 667608730;
assign addr[7099] = 685757258;
assign addr[7100] = 703851410;
assign addr[7101] = 721889752;
assign addr[7102] = 739870851;
assign addr[7103] = 757793284;
assign addr[7104] = 775655628;
assign addr[7105] = 793456467;
assign addr[7106] = 811194391;
assign addr[7107] = 828867991;
assign addr[7108] = 846475867;
assign addr[7109] = 864016623;
assign addr[7110] = 881488868;
assign addr[7111] = 898891215;
assign addr[7112] = 916222287;
assign addr[7113] = 933480707;
assign addr[7114] = 950665109;
assign addr[7115] = 967774128;
assign addr[7116] = 984806408;
assign addr[7117] = 1001760600;
assign addr[7118] = 1018635358;
assign addr[7119] = 1035429345;
assign addr[7120] = 1052141228;
assign addr[7121] = 1068769683;
assign addr[7122] = 1085313391;
assign addr[7123] = 1101771040;
assign addr[7124] = 1118141326;
assign addr[7125] = 1134422949;
assign addr[7126] = 1150614620;
assign addr[7127] = 1166715055;
assign addr[7128] = 1182722976;
assign addr[7129] = 1198637114;
assign addr[7130] = 1214456207;
assign addr[7131] = 1230179002;
assign addr[7132] = 1245804251;
assign addr[7133] = 1261330715;
assign addr[7134] = 1276757164;
assign addr[7135] = 1292082373;
assign addr[7136] = 1307305128;
assign addr[7137] = 1322424222;
assign addr[7138] = 1337438456;
assign addr[7139] = 1352346639;
assign addr[7140] = 1367147589;
assign addr[7141] = 1381840133;
assign addr[7142] = 1396423105;
assign addr[7143] = 1410895350;
assign addr[7144] = 1425255719;
assign addr[7145] = 1439503074;
assign addr[7146] = 1453636285;
assign addr[7147] = 1467654232;
assign addr[7148] = 1481555802;
assign addr[7149] = 1495339895;
assign addr[7150] = 1509005416;
assign addr[7151] = 1522551282;
assign addr[7152] = 1535976419;
assign addr[7153] = 1549279763;
assign addr[7154] = 1562460258;
assign addr[7155] = 1575516860;
assign addr[7156] = 1588448533;
assign addr[7157] = 1601254251;
assign addr[7158] = 1613933000;
assign addr[7159] = 1626483774;
assign addr[7160] = 1638905577;
assign addr[7161] = 1651197426;
assign addr[7162] = 1663358344;
assign addr[7163] = 1675387369;
assign addr[7164] = 1687283545;
assign addr[7165] = 1699045930;
assign addr[7166] = 1710673591;
assign addr[7167] = 1722165606;
assign addr[7168] = 1733521064;
assign addr[7169] = 1744739065;
assign addr[7170] = 1755818718;
assign addr[7171] = 1766759146;
assign addr[7172] = 1777559480;
assign addr[7173] = 1788218865;
assign addr[7174] = 1798736454;
assign addr[7175] = 1809111415;
assign addr[7176] = 1819342925;
assign addr[7177] = 1829430172;
assign addr[7178] = 1839372356;
assign addr[7179] = 1849168689;
assign addr[7180] = 1858818395;
assign addr[7181] = 1868320707;
assign addr[7182] = 1877674873;
assign addr[7183] = 1886880151;
assign addr[7184] = 1895935811;
assign addr[7185] = 1904841135;
assign addr[7186] = 1913595416;
assign addr[7187] = 1922197961;
assign addr[7188] = 1930648088;
assign addr[7189] = 1938945125;
assign addr[7190] = 1947088417;
assign addr[7191] = 1955077316;
assign addr[7192] = 1962911189;
assign addr[7193] = 1970589416;
assign addr[7194] = 1978111387;
assign addr[7195] = 1985476506;
assign addr[7196] = 1992684188;
assign addr[7197] = 1999733863;
assign addr[7198] = 2006624971;
assign addr[7199] = 2013356967;
assign addr[7200] = 2019929315;
assign addr[7201] = 2026341495;
assign addr[7202] = 2032592999;
assign addr[7203] = 2038683330;
assign addr[7204] = 2044612007;
assign addr[7205] = 2050378558;
assign addr[7206] = 2055982526;
assign addr[7207] = 2061423468;
assign addr[7208] = 2066700952;
assign addr[7209] = 2071814558;
assign addr[7210] = 2076763883;
assign addr[7211] = 2081548533;
assign addr[7212] = 2086168128;
assign addr[7213] = 2090622304;
assign addr[7214] = 2094910706;
assign addr[7215] = 2099032994;
assign addr[7216] = 2102988841;
assign addr[7217] = 2106777935;
assign addr[7218] = 2110399974;
assign addr[7219] = 2113854671;
assign addr[7220] = 2117141752;
assign addr[7221] = 2120260957;
assign addr[7222] = 2123212038;
assign addr[7223] = 2125994762;
assign addr[7224] = 2128608907;
assign addr[7225] = 2131054266;
assign addr[7226] = 2133330646;
assign addr[7227] = 2135437865;
assign addr[7228] = 2137375758;
assign addr[7229] = 2139144169;
assign addr[7230] = 2140742960;
assign addr[7231] = 2142172003;
assign addr[7232] = 2143431184;
assign addr[7233] = 2144520405;
assign addr[7234] = 2145439578;
assign addr[7235] = 2146188631;
assign addr[7236] = 2146767505;
assign addr[7237] = 2147176152;
assign addr[7238] = 2147414542;
assign addr[7239] = 2147482655;
assign addr[7240] = 2147380486;
assign addr[7241] = 2147108043;
assign addr[7242] = 2146665347;
assign addr[7243] = 2146052433;
assign addr[7244] = 2145269351;
assign addr[7245] = 2144316162;
assign addr[7246] = 2143192942;
assign addr[7247] = 2141899780;
assign addr[7248] = 2140436778;
assign addr[7249] = 2138804053;
assign addr[7250] = 2137001733;
assign addr[7251] = 2135029962;
assign addr[7252] = 2132888897;
assign addr[7253] = 2130578706;
assign addr[7254] = 2128099574;
assign addr[7255] = 2125451696;
assign addr[7256] = 2122635283;
assign addr[7257] = 2119650558;
assign addr[7258] = 2116497758;
assign addr[7259] = 2113177132;
assign addr[7260] = 2109688944;
assign addr[7261] = 2106033471;
assign addr[7262] = 2102211002;
assign addr[7263] = 2098221841;
assign addr[7264] = 2094066304;
assign addr[7265] = 2089744719;
assign addr[7266] = 2085257431;
assign addr[7267] = 2080604795;
assign addr[7268] = 2075787180;
assign addr[7269] = 2070804967;
assign addr[7270] = 2065658552;
assign addr[7271] = 2060348343;
assign addr[7272] = 2054874761;
assign addr[7273] = 2049238240;
assign addr[7274] = 2043439226;
assign addr[7275] = 2037478181;
assign addr[7276] = 2031355576;
assign addr[7277] = 2025071897;
assign addr[7278] = 2018627642;
assign addr[7279] = 2012023322;
assign addr[7280] = 2005259462;
assign addr[7281] = 1998336596;
assign addr[7282] = 1991255274;
assign addr[7283] = 1984016058;
assign addr[7284] = 1976619522;
assign addr[7285] = 1969066252;
assign addr[7286] = 1961356847;
assign addr[7287] = 1953491918;
assign addr[7288] = 1945472089;
assign addr[7289] = 1937297997;
assign addr[7290] = 1928970288;
assign addr[7291] = 1920489624;
assign addr[7292] = 1911856677;
assign addr[7293] = 1903072131;
assign addr[7294] = 1894136683;
assign addr[7295] = 1885051042;
assign addr[7296] = 1875815927;
assign addr[7297] = 1866432072;
assign addr[7298] = 1856900221;
assign addr[7299] = 1847221128;
assign addr[7300] = 1837395562;
assign addr[7301] = 1827424302;
assign addr[7302] = 1817308138;
assign addr[7303] = 1807047873;
assign addr[7304] = 1796644320;
assign addr[7305] = 1786098304;
assign addr[7306] = 1775410662;
assign addr[7307] = 1764582240;
assign addr[7308] = 1753613897;
assign addr[7309] = 1742506504;
assign addr[7310] = 1731260941;
assign addr[7311] = 1719878099;
assign addr[7312] = 1708358881;
assign addr[7313] = 1696704201;
assign addr[7314] = 1684914983;
assign addr[7315] = 1672992161;
assign addr[7316] = 1660936681;
assign addr[7317] = 1648749499;
assign addr[7318] = 1636431582;
assign addr[7319] = 1623983905;
assign addr[7320] = 1611407456;
assign addr[7321] = 1598703233;
assign addr[7322] = 1585872242;
assign addr[7323] = 1572915501;
assign addr[7324] = 1559834037;
assign addr[7325] = 1546628888;
assign addr[7326] = 1533301101;
assign addr[7327] = 1519851733;
assign addr[7328] = 1506281850;
assign addr[7329] = 1492592527;
assign addr[7330] = 1478784851;
assign addr[7331] = 1464859917;
assign addr[7332] = 1450818828;
assign addr[7333] = 1436662698;
assign addr[7334] = 1422392650;
assign addr[7335] = 1408009814;
assign addr[7336] = 1393515332;
assign addr[7337] = 1378910353;
assign addr[7338] = 1364196034;
assign addr[7339] = 1349373543;
assign addr[7340] = 1334444055;
assign addr[7341] = 1319408754;
assign addr[7342] = 1304268832;
assign addr[7343] = 1289025489;
assign addr[7344] = 1273679934;
assign addr[7345] = 1258233384;
assign addr[7346] = 1242687064;
assign addr[7347] = 1227042207;
assign addr[7348] = 1211300053;
assign addr[7349] = 1195461849;
assign addr[7350] = 1179528853;
assign addr[7351] = 1163502328;
assign addr[7352] = 1147383544;
assign addr[7353] = 1131173780;
assign addr[7354] = 1114874320;
assign addr[7355] = 1098486458;
assign addr[7356] = 1082011492;
assign addr[7357] = 1065450729;
assign addr[7358] = 1048805483;
assign addr[7359] = 1032077073;
assign addr[7360] = 1015266825;
assign addr[7361] = 998376073;
assign addr[7362] = 981406156;
assign addr[7363] = 964358420;
assign addr[7364] = 947234215;
assign addr[7365] = 930034901;
assign addr[7366] = 912761841;
assign addr[7367] = 895416404;
assign addr[7368] = 877999966;
assign addr[7369] = 860513908;
assign addr[7370] = 842959617;
assign addr[7371] = 825338484;
assign addr[7372] = 807651907;
assign addr[7373] = 789901288;
assign addr[7374] = 772088034;
assign addr[7375] = 754213559;
assign addr[7376] = 736279279;
assign addr[7377] = 718286617;
assign addr[7378] = 700236999;
assign addr[7379] = 682131857;
assign addr[7380] = 663972625;
assign addr[7381] = 645760745;
assign addr[7382] = 627497660;
assign addr[7383] = 609184818;
assign addr[7384] = 590823671;
assign addr[7385] = 572415676;
assign addr[7386] = 553962291;
assign addr[7387] = 535464981;
assign addr[7388] = 516925212;
assign addr[7389] = 498344454;
assign addr[7390] = 479724180;
assign addr[7391] = 461065866;
assign addr[7392] = 442370993;
assign addr[7393] = 423641043;
assign addr[7394] = 404877501;
assign addr[7395] = 386081854;
assign addr[7396] = 367255594;
assign addr[7397] = 348400212;
assign addr[7398] = 329517204;
assign addr[7399] = 310608068;
assign addr[7400] = 291674302;
assign addr[7401] = 272717408;
assign addr[7402] = 253738890;
assign addr[7403] = 234740251;
assign addr[7404] = 215722999;
assign addr[7405] = 196688642;
assign addr[7406] = 177638688;
assign addr[7407] = 158574649;
assign addr[7408] = 139498035;
assign addr[7409] = 120410361;
assign addr[7410] = 101313138;
assign addr[7411] = 82207882;
assign addr[7412] = 63096108;
assign addr[7413] = 43979330;
assign addr[7414] = 24859065;
assign addr[7415] = 5736829;
assign addr[7416] = -13385863;
assign addr[7417] = -32507492;
assign addr[7418] = -51626544;
assign addr[7419] = -70741503;
assign addr[7420] = -89850852;
assign addr[7421] = -108953076;
assign addr[7422] = -128046661;
assign addr[7423] = -147130093;
assign addr[7424] = -166201858;
assign addr[7425] = -185260444;
assign addr[7426] = -204304341;
assign addr[7427] = -223332037;
assign addr[7428] = -242342025;
assign addr[7429] = -261332796;
assign addr[7430] = -280302845;
assign addr[7431] = -299250668;
assign addr[7432] = -318174762;
assign addr[7433] = -337073627;
assign addr[7434] = -355945764;
assign addr[7435] = -374789676;
assign addr[7436] = -393603870;
assign addr[7437] = -412386854;
assign addr[7438] = -431137138;
assign addr[7439] = -449853235;
assign addr[7440] = -468533662;
assign addr[7441] = -487176937;
assign addr[7442] = -505781581;
assign addr[7443] = -524346121;
assign addr[7444] = -542869083;
assign addr[7445] = -561348998;
assign addr[7446] = -579784402;
assign addr[7447] = -598173833;
assign addr[7448] = -616515832;
assign addr[7449] = -634808946;
assign addr[7450] = -653051723;
assign addr[7451] = -671242716;
assign addr[7452] = -689380485;
assign addr[7453] = -707463589;
assign addr[7454] = -725490597;
assign addr[7455] = -743460077;
assign addr[7456] = -761370605;
assign addr[7457] = -779220762;
assign addr[7458] = -797009130;
assign addr[7459] = -814734301;
assign addr[7460] = -832394869;
assign addr[7461] = -849989433;
assign addr[7462] = -867516597;
assign addr[7463] = -884974973;
assign addr[7464] = -902363176;
assign addr[7465] = -919679827;
assign addr[7466] = -936923553;
assign addr[7467] = -954092986;
assign addr[7468] = -971186766;
assign addr[7469] = -988203537;
assign addr[7470] = -1005141949;
assign addr[7471] = -1022000660;
assign addr[7472] = -1038778332;
assign addr[7473] = -1055473635;
assign addr[7474] = -1072085246;
assign addr[7475] = -1088611847;
assign addr[7476] = -1105052128;
assign addr[7477] = -1121404785;
assign addr[7478] = -1137668521;
assign addr[7479] = -1153842047;
assign addr[7480] = -1169924081;
assign addr[7481] = -1185913346;
assign addr[7482] = -1201808576;
assign addr[7483] = -1217608510;
assign addr[7484] = -1233311895;
assign addr[7485] = -1248917486;
assign addr[7486] = -1264424045;
assign addr[7487] = -1279830344;
assign addr[7488] = -1295135159;
assign addr[7489] = -1310337279;
assign addr[7490] = -1325435496;
assign addr[7491] = -1340428615;
assign addr[7492] = -1355315445;
assign addr[7493] = -1370094808;
assign addr[7494] = -1384765530;
assign addr[7495] = -1399326449;
assign addr[7496] = -1413776410;
assign addr[7497] = -1428114267;
assign addr[7498] = -1442338884;
assign addr[7499] = -1456449131;
assign addr[7500] = -1470443891;
assign addr[7501] = -1484322054;
assign addr[7502] = -1498082520;
assign addr[7503] = -1511724196;
assign addr[7504] = -1525246002;
assign addr[7505] = -1538646865;
assign addr[7506] = -1551925723;
assign addr[7507] = -1565081523;
assign addr[7508] = -1578113222;
assign addr[7509] = -1591019785;
assign addr[7510] = -1603800191;
assign addr[7511] = -1616453425;
assign addr[7512] = -1628978484;
assign addr[7513] = -1641374375;
assign addr[7514] = -1653640115;
assign addr[7515] = -1665774731;
assign addr[7516] = -1677777262;
assign addr[7517] = -1689646755;
assign addr[7518] = -1701382270;
assign addr[7519] = -1712982875;
assign addr[7520] = -1724447652;
assign addr[7521] = -1735775690;
assign addr[7522] = -1746966091;
assign addr[7523] = -1758017969;
assign addr[7524] = -1768930447;
assign addr[7525] = -1779702660;
assign addr[7526] = -1790333753;
assign addr[7527] = -1800822883;
assign addr[7528] = -1811169220;
assign addr[7529] = -1821371941;
assign addr[7530] = -1831430239;
assign addr[7531] = -1841343316;
assign addr[7532] = -1851110385;
assign addr[7533] = -1860730673;
assign addr[7534] = -1870203416;
assign addr[7535] = -1879527863;
assign addr[7536] = -1888703276;
assign addr[7537] = -1897728925;
assign addr[7538] = -1906604097;
assign addr[7539] = -1915328086;
assign addr[7540] = -1923900201;
assign addr[7541] = -1932319763;
assign addr[7542] = -1940586104;
assign addr[7543] = -1948698568;
assign addr[7544] = -1956656513;
assign addr[7545] = -1964459306;
assign addr[7546] = -1972106330;
assign addr[7547] = -1979596978;
assign addr[7548] = -1986930656;
assign addr[7549] = -1994106782;
assign addr[7550] = -2001124788;
assign addr[7551] = -2007984117;
assign addr[7552] = -2014684225;
assign addr[7553] = -2021224581;
assign addr[7554] = -2027604666;
assign addr[7555] = -2033823974;
assign addr[7556] = -2039882013;
assign addr[7557] = -2045778302;
assign addr[7558] = -2051512372;
assign addr[7559] = -2057083771;
assign addr[7560] = -2062492055;
assign addr[7561] = -2067736796;
assign addr[7562] = -2072817579;
assign addr[7563] = -2077733999;
assign addr[7564] = -2082485668;
assign addr[7565] = -2087072209;
assign addr[7566] = -2091493257;
assign addr[7567] = -2095748463;
assign addr[7568] = -2099837489;
assign addr[7569] = -2103760010;
assign addr[7570] = -2107515716;
assign addr[7571] = -2111104309;
assign addr[7572] = -2114525505;
assign addr[7573] = -2117779031;
assign addr[7574] = -2120864631;
assign addr[7575] = -2123782059;
assign addr[7576] = -2126531084;
assign addr[7577] = -2129111488;
assign addr[7578] = -2131523066;
assign addr[7579] = -2133765628;
assign addr[7580] = -2135838995;
assign addr[7581] = -2137743003;
assign addr[7582] = -2139477502;
assign addr[7583] = -2141042352;
assign addr[7584] = -2142437431;
assign addr[7585] = -2143662628;
assign addr[7586] = -2144717846;
assign addr[7587] = -2145603001;
assign addr[7588] = -2146318022;
assign addr[7589] = -2146862854;
assign addr[7590] = -2147237452;
assign addr[7591] = -2147441787;
assign addr[7592] = -2147475844;
assign addr[7593] = -2147339619;
assign addr[7594] = -2147033123;
assign addr[7595] = -2146556380;
assign addr[7596] = -2145909429;
assign addr[7597] = -2145092320;
assign addr[7598] = -2144105118;
assign addr[7599] = -2142947902;
assign addr[7600] = -2141620763;
assign addr[7601] = -2140123807;
assign addr[7602] = -2138457152;
assign addr[7603] = -2136620930;
assign addr[7604] = -2134615288;
assign addr[7605] = -2132440383;
assign addr[7606] = -2130096389;
assign addr[7607] = -2127583492;
assign addr[7608] = -2124901890;
assign addr[7609] = -2122051796;
assign addr[7610] = -2119033436;
assign addr[7611] = -2115847050;
assign addr[7612] = -2112492891;
assign addr[7613] = -2108971223;
assign addr[7614] = -2105282327;
assign addr[7615] = -2101426496;
assign addr[7616] = -2097404033;
assign addr[7617] = -2093215260;
assign addr[7618] = -2088860507;
assign addr[7619] = -2084340120;
assign addr[7620] = -2079654458;
assign addr[7621] = -2074803892;
assign addr[7622] = -2069788807;
assign addr[7623] = -2064609600;
assign addr[7624] = -2059266683;
assign addr[7625] = -2053760478;
assign addr[7626] = -2048091422;
assign addr[7627] = -2042259965;
assign addr[7628] = -2036266570;
assign addr[7629] = -2030111710;
assign addr[7630] = -2023795876;
assign addr[7631] = -2017319567;
assign addr[7632] = -2010683297;
assign addr[7633] = -2003887591;
assign addr[7634] = -1996932990;
assign addr[7635] = -1989820044;
assign addr[7636] = -1982549318;
assign addr[7637] = -1975121388;
assign addr[7638] = -1967536842;
assign addr[7639] = -1959796283;
assign addr[7640] = -1951900324;
assign addr[7641] = -1943849591;
assign addr[7642] = -1935644723;
assign addr[7643] = -1927286370;
assign addr[7644] = -1918775195;
assign addr[7645] = -1910111873;
assign addr[7646] = -1901297091;
assign addr[7647] = -1892331547;
assign addr[7648] = -1883215953;
assign addr[7649] = -1873951032;
assign addr[7650] = -1864537518;
assign addr[7651] = -1854976157;
assign addr[7652] = -1845267708;
assign addr[7653] = -1835412941;
assign addr[7654] = -1825412636;
assign addr[7655] = -1815267588;
assign addr[7656] = -1804978599;
assign addr[7657] = -1794546487;
assign addr[7658] = -1783972079;
assign addr[7659] = -1773256212;
assign addr[7660] = -1762399737;
assign addr[7661] = -1751403515;
assign addr[7662] = -1740268417;
assign addr[7663] = -1728995326;
assign addr[7664] = -1717585136;
assign addr[7665] = -1706038753;
assign addr[7666] = -1694357091;
assign addr[7667] = -1682541077;
assign addr[7668] = -1670591647;
assign addr[7669] = -1658509750;
assign addr[7670] = -1646296344;
assign addr[7671] = -1633952396;
assign addr[7672] = -1621478885;
assign addr[7673] = -1608876801;
assign addr[7674] = -1596147143;
assign addr[7675] = -1583290921;
assign addr[7676] = -1570309153;
assign addr[7677] = -1557202869;
assign addr[7678] = -1543973108;
assign addr[7679] = -1530620920;
assign addr[7680] = -1517147363;
assign addr[7681] = -1503553506;
assign addr[7682] = -1489840425;
assign addr[7683] = -1476009210;
assign addr[7684] = -1462060956;
assign addr[7685] = -1447996770;
assign addr[7686] = -1433817766;
assign addr[7687] = -1419525069;
assign addr[7688] = -1405119813;
assign addr[7689] = -1390603139;
assign addr[7690] = -1375976199;
assign addr[7691] = -1361240152;
assign addr[7692] = -1346396168;
assign addr[7693] = -1331445422;
assign addr[7694] = -1316389101;
assign addr[7695] = -1301228398;
assign addr[7696] = -1285964516;
assign addr[7697] = -1270598665;
assign addr[7698] = -1255132063;
assign addr[7699] = -1239565936;
assign addr[7700] = -1223901520;
assign addr[7701] = -1208140056;
assign addr[7702] = -1192282793;
assign addr[7703] = -1176330990;
assign addr[7704] = -1160285911;
assign addr[7705] = -1144148829;
assign addr[7706] = -1127921022;
assign addr[7707] = -1111603778;
assign addr[7708] = -1095198391;
assign addr[7709] = -1078706161;
assign addr[7710] = -1062128397;
assign addr[7711] = -1045466412;
assign addr[7712] = -1028721528;
assign addr[7713] = -1011895073;
assign addr[7714] = -994988380;
assign addr[7715] = -978002791;
assign addr[7716] = -960939653;
assign addr[7717] = -943800318;
assign addr[7718] = -926586145;
assign addr[7719] = -909298500;
assign addr[7720] = -891938752;
assign addr[7721] = -874508280;
assign addr[7722] = -857008464;
assign addr[7723] = -839440693;
assign addr[7724] = -821806359;
assign addr[7725] = -804106861;
assign addr[7726] = -786343603;
assign addr[7727] = -768517992;
assign addr[7728] = -750631442;
assign addr[7729] = -732685372;
assign addr[7730] = -714681204;
assign addr[7731] = -696620367;
assign addr[7732] = -678504291;
assign addr[7733] = -660334415;
assign addr[7734] = -642112178;
assign addr[7735] = -623839025;
assign addr[7736] = -605516406;
assign addr[7737] = -587145773;
assign addr[7738] = -568728583;
assign addr[7739] = -550266296;
assign addr[7740] = -531760377;
assign addr[7741] = -513212292;
assign addr[7742] = -494623513;
assign addr[7743] = -475995513;
assign addr[7744] = -457329769;
assign addr[7745] = -438627762;
assign addr[7746] = -419890975;
assign addr[7747] = -401120892;
assign addr[7748] = -382319004;
assign addr[7749] = -363486799;
assign addr[7750] = -344625773;
assign addr[7751] = -325737419;
assign addr[7752] = -306823237;
assign addr[7753] = -287884725;
assign addr[7754] = -268923386;
assign addr[7755] = -249940723;
assign addr[7756] = -230938242;
assign addr[7757] = -211917448;
assign addr[7758] = -192879850;
assign addr[7759] = -173826959;
assign addr[7760] = -154760284;
assign addr[7761] = -135681337;
assign addr[7762] = -116591632;
assign addr[7763] = -97492681;
assign addr[7764] = -78386000;
assign addr[7765] = -59273104;
assign addr[7766] = -40155507;
assign addr[7767] = -21034727;
assign addr[7768] = -1912278;
assign addr[7769] = 17210322;
assign addr[7770] = 36331557;
assign addr[7771] = 55449912;
assign addr[7772] = 74563870;
assign addr[7773] = 93671915;
assign addr[7774] = 112772533;
assign addr[7775] = 131864208;
assign addr[7776] = 150945428;
assign addr[7777] = 170014678;
assign addr[7778] = 189070447;
assign addr[7779] = 208111224;
assign addr[7780] = 227135500;
assign addr[7781] = 246141764;
assign addr[7782] = 265128512;
assign addr[7783] = 284094236;
assign addr[7784] = 303037433;
assign addr[7785] = 321956601;
assign addr[7786] = 340850240;
assign addr[7787] = 359716852;
assign addr[7788] = 378554940;
assign addr[7789] = 397363011;
assign addr[7790] = 416139574;
assign addr[7791] = 434883140;
assign addr[7792] = 453592221;
assign addr[7793] = 472265336;
assign addr[7794] = 490901003;
assign addr[7795] = 509497745;
assign addr[7796] = 528054086;
assign addr[7797] = 546568556;
assign addr[7798] = 565039687;
assign addr[7799] = 583466013;
assign addr[7800] = 601846074;
assign addr[7801] = 620178412;
assign addr[7802] = 638461574;
assign addr[7803] = 656694110;
assign addr[7804] = 674874574;
assign addr[7805] = 693001525;
assign addr[7806] = 711073524;
assign addr[7807] = 729089140;
assign addr[7808] = 747046944;
assign addr[7809] = 764945512;
assign addr[7810] = 782783424;
assign addr[7811] = 800559266;
assign addr[7812] = 818271628;
assign addr[7813] = 835919107;
assign addr[7814] = 853500302;
assign addr[7815] = 871013820;
assign addr[7816] = 888458272;
assign addr[7817] = 905832274;
assign addr[7818] = 923134450;
assign addr[7819] = 940363427;
assign addr[7820] = 957517838;
assign addr[7821] = 974596324;
assign addr[7822] = 991597531;
assign addr[7823] = 1008520110;
assign addr[7824] = 1025362720;
assign addr[7825] = 1042124025;
assign addr[7826] = 1058802695;
assign addr[7827] = 1075397409;
assign addr[7828] = 1091906851;
assign addr[7829] = 1108329711;
assign addr[7830] = 1124664687;
assign addr[7831] = 1140910484;
assign addr[7832] = 1157065814;
assign addr[7833] = 1173129396;
assign addr[7834] = 1189099956;
assign addr[7835] = 1204976227;
assign addr[7836] = 1220756951;
assign addr[7837] = 1236440877;
assign addr[7838] = 1252026760;
assign addr[7839] = 1267513365;
assign addr[7840] = 1282899464;
assign addr[7841] = 1298183838;
assign addr[7842] = 1313365273;
assign addr[7843] = 1328442566;
assign addr[7844] = 1343414522;
assign addr[7845] = 1358279953;
assign addr[7846] = 1373037681;
assign addr[7847] = 1387686535;
assign addr[7848] = 1402225355;
assign addr[7849] = 1416652986;
assign addr[7850] = 1430968286;
assign addr[7851] = 1445170118;
assign addr[7852] = 1459257358;
assign addr[7853] = 1473228887;
assign addr[7854] = 1487083598;
assign addr[7855] = 1500820393;
assign addr[7856] = 1514438181;
assign addr[7857] = 1527935884;
assign addr[7858] = 1541312431;
assign addr[7859] = 1554566762;
assign addr[7860] = 1567697824;
assign addr[7861] = 1580704578;
assign addr[7862] = 1593585992;
assign addr[7863] = 1606341043;
assign addr[7864] = 1618968722;
assign addr[7865] = 1631468027;
assign addr[7866] = 1643837966;
assign addr[7867] = 1656077559;
assign addr[7868] = 1668185835;
assign addr[7869] = 1680161834;
assign addr[7870] = 1692004606;
assign addr[7871] = 1703713213;
assign addr[7872] = 1715286726;
assign addr[7873] = 1726724227;
assign addr[7874] = 1738024810;
assign addr[7875] = 1749187577;
assign addr[7876] = 1760211645;
assign addr[7877] = 1771096139;
assign addr[7878] = 1781840195;
assign addr[7879] = 1792442963;
assign addr[7880] = 1802903601;
assign addr[7881] = 1813221279;
assign addr[7882] = 1823395180;
assign addr[7883] = 1833424497;
assign addr[7884] = 1843308435;
assign addr[7885] = 1853046210;
assign addr[7886] = 1862637049;
assign addr[7887] = 1872080193;
assign addr[7888] = 1881374892;
assign addr[7889] = 1890520410;
assign addr[7890] = 1899516021;
assign addr[7891] = 1908361011;
assign addr[7892] = 1917054681;
assign addr[7893] = 1925596340;
assign addr[7894] = 1933985310;
assign addr[7895] = 1942220928;
assign addr[7896] = 1950302539;
assign addr[7897] = 1958229503;
assign addr[7898] = 1966001192;
assign addr[7899] = 1973616989;
assign addr[7900] = 1981076290;
assign addr[7901] = 1988378503;
assign addr[7902] = 1995523051;
assign addr[7903] = 2002509365;
assign addr[7904] = 2009336893;
assign addr[7905] = 2016005093;
assign addr[7906] = 2022513436;
assign addr[7907] = 2028861406;
assign addr[7908] = 2035048499;
assign addr[7909] = 2041074226;
assign addr[7910] = 2046938108;
assign addr[7911] = 2052639680;
assign addr[7912] = 2058178491;
assign addr[7913] = 2063554100;
assign addr[7914] = 2068766083;
assign addr[7915] = 2073814024;
assign addr[7916] = 2078697525;
assign addr[7917] = 2083416198;
assign addr[7918] = 2087969669;
assign addr[7919] = 2092357577;
assign addr[7920] = 2096579573;
assign addr[7921] = 2100635323;
assign addr[7922] = 2104524506;
assign addr[7923] = 2108246813;
assign addr[7924] = 2111801949;
assign addr[7925] = 2115189632;
assign addr[7926] = 2118409593;
assign addr[7927] = 2121461578;
assign addr[7928] = 2124345343;
assign addr[7929] = 2127060661;
assign addr[7930] = 2129607316;
assign addr[7931] = 2131985106;
assign addr[7932] = 2134193842;
assign addr[7933] = 2136233350;
assign addr[7934] = 2138103468;
assign addr[7935] = 2139804048;
assign addr[7936] = 2141334954;
assign addr[7937] = 2142696065;
assign addr[7938] = 2143887273;
assign addr[7939] = 2144908484;
assign addr[7940] = 2145759618;
assign addr[7941] = 2146440605;
assign addr[7942] = 2146951393;
assign addr[7943] = 2147291941;
assign addr[7944] = 2147462221;
assign addr[7945] = 2147462221;
assign addr[7946] = 2147291941;
assign addr[7947] = 2146951393;
assign addr[7948] = 2146440605;
assign addr[7949] = 2145759618;
assign addr[7950] = 2144908484;
assign addr[7951] = 2143887273;
assign addr[7952] = 2142696065;
assign addr[7953] = 2141334954;
assign addr[7954] = 2139804048;
assign addr[7955] = 2138103468;
assign addr[7956] = 2136233350;
assign addr[7957] = 2134193842;
assign addr[7958] = 2131985106;
assign addr[7959] = 2129607316;
assign addr[7960] = 2127060661;
assign addr[7961] = 2124345343;
assign addr[7962] = 2121461578;
assign addr[7963] = 2118409593;
assign addr[7964] = 2115189632;
assign addr[7965] = 2111801949;
assign addr[7966] = 2108246813;
assign addr[7967] = 2104524506;
assign addr[7968] = 2100635323;
assign addr[7969] = 2096579573;
assign addr[7970] = 2092357577;
assign addr[7971] = 2087969669;
assign addr[7972] = 2083416198;
assign addr[7973] = 2078697525;
assign addr[7974] = 2073814024;
assign addr[7975] = 2068766083;
assign addr[7976] = 2063554100;
assign addr[7977] = 2058178491;
assign addr[7978] = 2052639680;
assign addr[7979] = 2046938108;
assign addr[7980] = 2041074226;
assign addr[7981] = 2035048499;
assign addr[7982] = 2028861406;
assign addr[7983] = 2022513436;
assign addr[7984] = 2016005093;
assign addr[7985] = 2009336893;
assign addr[7986] = 2002509365;
assign addr[7987] = 1995523051;
assign addr[7988] = 1988378503;
assign addr[7989] = 1981076290;
assign addr[7990] = 1973616989;
assign addr[7991] = 1966001192;
assign addr[7992] = 1958229503;
assign addr[7993] = 1950302539;
assign addr[7994] = 1942220928;
assign addr[7995] = 1933985310;
assign addr[7996] = 1925596340;
assign addr[7997] = 1917054681;
assign addr[7998] = 1908361011;
assign addr[7999] = 1899516021;
assign addr[8000] = 1890520410;
assign addr[8001] = 1881374892;
assign addr[8002] = 1872080193;
assign addr[8003] = 1862637049;
assign addr[8004] = 1853046210;
assign addr[8005] = 1843308435;
assign addr[8006] = 1833424497;
assign addr[8007] = 1823395180;
assign addr[8008] = 1813221279;
assign addr[8009] = 1802903601;
assign addr[8010] = 1792442963;
assign addr[8011] = 1781840195;
assign addr[8012] = 1771096139;
assign addr[8013] = 1760211645;
assign addr[8014] = 1749187577;
assign addr[8015] = 1738024810;
assign addr[8016] = 1726724227;
assign addr[8017] = 1715286726;
assign addr[8018] = 1703713213;
assign addr[8019] = 1692004606;
assign addr[8020] = 1680161834;
assign addr[8021] = 1668185835;
assign addr[8022] = 1656077559;
assign addr[8023] = 1643837966;
assign addr[8024] = 1631468027;
assign addr[8025] = 1618968722;
assign addr[8026] = 1606341043;
assign addr[8027] = 1593585992;
assign addr[8028] = 1580704578;
assign addr[8029] = 1567697824;
assign addr[8030] = 1554566762;
assign addr[8031] = 1541312431;
assign addr[8032] = 1527935884;
assign addr[8033] = 1514438181;
assign addr[8034] = 1500820393;
assign addr[8035] = 1487083598;
assign addr[8036] = 1473228887;
assign addr[8037] = 1459257358;
assign addr[8038] = 1445170118;
assign addr[8039] = 1430968286;
assign addr[8040] = 1416652986;
assign addr[8041] = 1402225355;
assign addr[8042] = 1387686535;
assign addr[8043] = 1373037681;
assign addr[8044] = 1358279953;
assign addr[8045] = 1343414522;
assign addr[8046] = 1328442566;
assign addr[8047] = 1313365273;
assign addr[8048] = 1298183838;
assign addr[8049] = 1282899464;
assign addr[8050] = 1267513365;
assign addr[8051] = 1252026760;
assign addr[8052] = 1236440877;
assign addr[8053] = 1220756951;
assign addr[8054] = 1204976227;
assign addr[8055] = 1189099956;
assign addr[8056] = 1173129396;
assign addr[8057] = 1157065814;
assign addr[8058] = 1140910484;
assign addr[8059] = 1124664687;
assign addr[8060] = 1108329711;
assign addr[8061] = 1091906851;
assign addr[8062] = 1075397409;
assign addr[8063] = 1058802695;
assign addr[8064] = 1042124025;
assign addr[8065] = 1025362720;
assign addr[8066] = 1008520110;
assign addr[8067] = 991597531;
assign addr[8068] = 974596324;
assign addr[8069] = 957517838;
assign addr[8070] = 940363427;
assign addr[8071] = 923134450;
assign addr[8072] = 905832274;
assign addr[8073] = 888458272;
assign addr[8074] = 871013820;
assign addr[8075] = 853500302;
assign addr[8076] = 835919107;
assign addr[8077] = 818271628;
assign addr[8078] = 800559266;
assign addr[8079] = 782783424;
assign addr[8080] = 764945512;
assign addr[8081] = 747046944;
assign addr[8082] = 729089140;
assign addr[8083] = 711073524;
assign addr[8084] = 693001525;
assign addr[8085] = 674874574;
assign addr[8086] = 656694110;
assign addr[8087] = 638461574;
assign addr[8088] = 620178412;
assign addr[8089] = 601846074;
assign addr[8090] = 583466013;
assign addr[8091] = 565039687;
assign addr[8092] = 546568556;
assign addr[8093] = 528054086;
assign addr[8094] = 509497745;
assign addr[8095] = 490901003;
assign addr[8096] = 472265336;
assign addr[8097] = 453592221;
assign addr[8098] = 434883140;
assign addr[8099] = 416139574;
assign addr[8100] = 397363011;
assign addr[8101] = 378554940;
assign addr[8102] = 359716852;
assign addr[8103] = 340850240;
assign addr[8104] = 321956601;
assign addr[8105] = 303037433;
assign addr[8106] = 284094236;
assign addr[8107] = 265128512;
assign addr[8108] = 246141764;
assign addr[8109] = 227135500;
assign addr[8110] = 208111224;
assign addr[8111] = 189070447;
assign addr[8112] = 170014678;
assign addr[8113] = 150945428;
assign addr[8114] = 131864208;
assign addr[8115] = 112772533;
assign addr[8116] = 93671915;
assign addr[8117] = 74563870;
assign addr[8118] = 55449912;
assign addr[8119] = 36331557;
assign addr[8120] = 17210322;
assign addr[8121] = -1912278;
assign addr[8122] = -21034727;
assign addr[8123] = -40155507;
assign addr[8124] = -59273104;
assign addr[8125] = -78386000;
assign addr[8126] = -97492681;
assign addr[8127] = -116591632;
assign addr[8128] = -135681337;
assign addr[8129] = -154760284;
assign addr[8130] = -173826959;
assign addr[8131] = -192879850;
assign addr[8132] = -211917448;
assign addr[8133] = -230938242;
assign addr[8134] = -249940723;
assign addr[8135] = -268923386;
assign addr[8136] = -287884725;
assign addr[8137] = -306823237;
assign addr[8138] = -325737419;
assign addr[8139] = -344625773;
assign addr[8140] = -363486799;
assign addr[8141] = -382319004;
assign addr[8142] = -401120892;
assign addr[8143] = -419890975;
assign addr[8144] = -438627762;
assign addr[8145] = -457329769;
assign addr[8146] = -475995513;
assign addr[8147] = -494623513;
assign addr[8148] = -513212292;
assign addr[8149] = -531760377;
assign addr[8150] = -550266296;
assign addr[8151] = -568728583;
assign addr[8152] = -587145773;
assign addr[8153] = -605516406;
assign addr[8154] = -623839025;
assign addr[8155] = -642112178;
assign addr[8156] = -660334415;
assign addr[8157] = -678504291;
assign addr[8158] = -696620367;
assign addr[8159] = -714681204;
assign addr[8160] = -732685372;
assign addr[8161] = -750631442;
assign addr[8162] = -768517992;
assign addr[8163] = -786343603;
assign addr[8164] = -804106861;
assign addr[8165] = -821806359;
assign addr[8166] = -839440693;
assign addr[8167] = -857008464;
assign addr[8168] = -874508280;
assign addr[8169] = -891938752;
assign addr[8170] = -909298500;
assign addr[8171] = -926586145;
assign addr[8172] = -943800318;
assign addr[8173] = -960939653;
assign addr[8174] = -978002791;
assign addr[8175] = -994988380;
assign addr[8176] = -1011895073;
assign addr[8177] = -1028721528;
assign addr[8178] = -1045466412;
assign addr[8179] = -1062128397;
assign addr[8180] = -1078706161;
assign addr[8181] = -1095198391;
assign addr[8182] = -1111603778;
assign addr[8183] = -1127921022;
assign addr[8184] = -1144148829;
assign addr[8185] = -1160285911;
assign addr[8186] = -1176330990;
assign addr[8187] = -1192282793;
assign addr[8188] = -1208140056;
assign addr[8189] = -1223901520;
assign addr[8190] = -1239565936;
assign addr[8191] = -1255132063;
assign addr[8192] = -1270598665;
assign addr[8193] = -1285964516;
assign addr[8194] = -1301228398;
assign addr[8195] = -1316389101;
assign addr[8196] = -1331445422;
assign addr[8197] = -1346396168;
assign addr[8198] = -1361240152;
assign addr[8199] = -1375976199;
assign addr[8200] = -1390603139;
assign addr[8201] = -1405119813;
assign addr[8202] = -1419525069;
assign addr[8203] = -1433817766;
assign addr[8204] = -1447996770;
assign addr[8205] = -1462060956;
assign addr[8206] = -1476009210;
assign addr[8207] = -1489840425;
assign addr[8208] = -1503553506;
assign addr[8209] = -1517147363;
assign addr[8210] = -1530620920;
assign addr[8211] = -1543973108;
assign addr[8212] = -1557202869;
assign addr[8213] = -1570309153;
assign addr[8214] = -1583290921;
assign addr[8215] = -1596147143;
assign addr[8216] = -1608876801;
assign addr[8217] = -1621478885;
assign addr[8218] = -1633952396;
assign addr[8219] = -1646296344;
assign addr[8220] = -1658509750;
assign addr[8221] = -1670591647;
assign addr[8222] = -1682541077;
assign addr[8223] = -1694357091;
assign addr[8224] = -1706038753;
assign addr[8225] = -1717585136;
assign addr[8226] = -1728995326;
assign addr[8227] = -1740268417;
assign addr[8228] = -1751403515;
assign addr[8229] = -1762399737;
assign addr[8230] = -1773256212;
assign addr[8231] = -1783972079;
assign addr[8232] = -1794546487;
assign addr[8233] = -1804978599;
assign addr[8234] = -1815267588;
assign addr[8235] = -1825412636;
assign addr[8236] = -1835412941;
assign addr[8237] = -1845267708;
assign addr[8238] = -1854976157;
assign addr[8239] = -1864537518;
assign addr[8240] = -1873951032;
assign addr[8241] = -1883215953;
assign addr[8242] = -1892331547;
assign addr[8243] = -1901297091;
assign addr[8244] = -1910111873;
assign addr[8245] = -1918775195;
assign addr[8246] = -1927286370;
assign addr[8247] = -1935644723;
assign addr[8248] = -1943849591;
assign addr[8249] = -1951900324;
assign addr[8250] = -1959796283;
assign addr[8251] = -1967536842;
assign addr[8252] = -1975121388;
assign addr[8253] = -1982549318;
assign addr[8254] = -1989820044;
assign addr[8255] = -1996932990;
assign addr[8256] = -2003887591;
assign addr[8257] = -2010683297;
assign addr[8258] = -2017319567;
assign addr[8259] = -2023795876;
assign addr[8260] = -2030111710;
assign addr[8261] = -2036266570;
assign addr[8262] = -2042259965;
assign addr[8263] = -2048091422;
assign addr[8264] = -2053760478;
assign addr[8265] = -2059266683;
assign addr[8266] = -2064609600;
assign addr[8267] = -2069788807;
assign addr[8268] = -2074803892;
assign addr[8269] = -2079654458;
assign addr[8270] = -2084340120;
assign addr[8271] = -2088860507;
assign addr[8272] = -2093215260;
assign addr[8273] = -2097404033;
assign addr[8274] = -2101426496;
assign addr[8275] = -2105282327;
assign addr[8276] = -2108971223;
assign addr[8277] = -2112492891;
assign addr[8278] = -2115847050;
assign addr[8279] = -2119033436;
assign addr[8280] = -2122051796;
assign addr[8281] = -2124901890;
assign addr[8282] = -2127583492;
assign addr[8283] = -2130096389;
assign addr[8284] = -2132440383;
assign addr[8285] = -2134615288;
assign addr[8286] = -2136620930;
assign addr[8287] = -2138457152;
assign addr[8288] = -2140123807;
assign addr[8289] = -2141620763;
assign addr[8290] = -2142947902;
assign addr[8291] = -2144105118;
assign addr[8292] = -2145092320;
assign addr[8293] = -2145909429;
assign addr[8294] = -2146556380;
assign addr[8295] = -2147033123;
assign addr[8296] = -2147339619;
assign addr[8297] = -2147475844;
assign addr[8298] = -2147441787;
assign addr[8299] = -2147237452;
assign addr[8300] = -2146862854;
assign addr[8301] = -2146318022;
assign addr[8302] = -2145603001;
assign addr[8303] = -2144717846;
assign addr[8304] = -2143662628;
assign addr[8305] = -2142437431;
assign addr[8306] = -2141042352;
assign addr[8307] = -2139477502;
assign addr[8308] = -2137743003;
assign addr[8309] = -2135838995;
assign addr[8310] = -2133765628;
assign addr[8311] = -2131523066;
assign addr[8312] = -2129111488;
assign addr[8313] = -2126531084;
assign addr[8314] = -2123782059;
assign addr[8315] = -2120864631;
assign addr[8316] = -2117779031;
assign addr[8317] = -2114525505;
assign addr[8318] = -2111104309;
assign addr[8319] = -2107515716;
assign addr[8320] = -2103760010;
assign addr[8321] = -2099837489;
assign addr[8322] = -2095748463;
assign addr[8323] = -2091493257;
assign addr[8324] = -2087072209;
assign addr[8325] = -2082485668;
assign addr[8326] = -2077733999;
assign addr[8327] = -2072817579;
assign addr[8328] = -2067736796;
assign addr[8329] = -2062492055;
assign addr[8330] = -2057083771;
assign addr[8331] = -2051512372;
assign addr[8332] = -2045778302;
assign addr[8333] = -2039882013;
assign addr[8334] = -2033823974;
assign addr[8335] = -2027604666;
assign addr[8336] = -2021224581;
assign addr[8337] = -2014684225;
assign addr[8338] = -2007984117;
assign addr[8339] = -2001124788;
assign addr[8340] = -1994106782;
assign addr[8341] = -1986930656;
assign addr[8342] = -1979596978;
assign addr[8343] = -1972106330;
assign addr[8344] = -1964459306;
assign addr[8345] = -1956656513;
assign addr[8346] = -1948698568;
assign addr[8347] = -1940586104;
assign addr[8348] = -1932319763;
assign addr[8349] = -1923900201;
assign addr[8350] = -1915328086;
assign addr[8351] = -1906604097;
assign addr[8352] = -1897728925;
assign addr[8353] = -1888703276;
assign addr[8354] = -1879527863;
assign addr[8355] = -1870203416;
assign addr[8356] = -1860730673;
assign addr[8357] = -1851110385;
assign addr[8358] = -1841343316;
assign addr[8359] = -1831430239;
assign addr[8360] = -1821371941;
assign addr[8361] = -1811169220;
assign addr[8362] = -1800822883;
assign addr[8363] = -1790333753;
assign addr[8364] = -1779702660;
assign addr[8365] = -1768930447;
assign addr[8366] = -1758017969;
assign addr[8367] = -1746966091;
assign addr[8368] = -1735775690;
assign addr[8369] = -1724447652;
assign addr[8370] = -1712982875;
assign addr[8371] = -1701382270;
assign addr[8372] = -1689646755;
assign addr[8373] = -1677777262;
assign addr[8374] = -1665774731;
assign addr[8375] = -1653640115;
assign addr[8376] = -1641374375;
assign addr[8377] = -1628978484;
assign addr[8378] = -1616453425;
assign addr[8379] = -1603800191;
assign addr[8380] = -1591019785;
assign addr[8381] = -1578113222;
assign addr[8382] = -1565081523;
assign addr[8383] = -1551925723;
assign addr[8384] = -1538646865;
assign addr[8385] = -1525246002;
assign addr[8386] = -1511724196;
assign addr[8387] = -1498082520;
assign addr[8388] = -1484322054;
assign addr[8389] = -1470443891;
assign addr[8390] = -1456449131;
assign addr[8391] = -1442338884;
assign addr[8392] = -1428114267;
assign addr[8393] = -1413776410;
assign addr[8394] = -1399326449;
assign addr[8395] = -1384765530;
assign addr[8396] = -1370094808;
assign addr[8397] = -1355315445;
assign addr[8398] = -1340428615;
assign addr[8399] = -1325435496;
assign addr[8400] = -1310337279;
assign addr[8401] = -1295135159;
assign addr[8402] = -1279830344;
assign addr[8403] = -1264424045;
assign addr[8404] = -1248917486;
assign addr[8405] = -1233311895;
assign addr[8406] = -1217608510;
assign addr[8407] = -1201808576;
assign addr[8408] = -1185913346;
assign addr[8409] = -1169924081;
assign addr[8410] = -1153842047;
assign addr[8411] = -1137668521;
assign addr[8412] = -1121404785;
assign addr[8413] = -1105052128;
assign addr[8414] = -1088611847;
assign addr[8415] = -1072085246;
assign addr[8416] = -1055473635;
assign addr[8417] = -1038778332;
assign addr[8418] = -1022000660;
assign addr[8419] = -1005141949;
assign addr[8420] = -988203537;
assign addr[8421] = -971186766;
assign addr[8422] = -954092986;
assign addr[8423] = -936923553;
assign addr[8424] = -919679827;
assign addr[8425] = -902363176;
assign addr[8426] = -884974973;
assign addr[8427] = -867516597;
assign addr[8428] = -849989433;
assign addr[8429] = -832394869;
assign addr[8430] = -814734301;
assign addr[8431] = -797009130;
assign addr[8432] = -779220762;
assign addr[8433] = -761370605;
assign addr[8434] = -743460077;
assign addr[8435] = -725490597;
assign addr[8436] = -707463589;
assign addr[8437] = -689380485;
assign addr[8438] = -671242716;
assign addr[8439] = -653051723;
assign addr[8440] = -634808946;
assign addr[8441] = -616515832;
assign addr[8442] = -598173833;
assign addr[8443] = -579784402;
assign addr[8444] = -561348998;
assign addr[8445] = -542869083;
assign addr[8446] = -524346121;
assign addr[8447] = -505781581;
assign addr[8448] = -487176937;
assign addr[8449] = -468533662;
assign addr[8450] = -449853235;
assign addr[8451] = -431137138;
assign addr[8452] = -412386854;
assign addr[8453] = -393603870;
assign addr[8454] = -374789676;
assign addr[8455] = -355945764;
assign addr[8456] = -337073627;
assign addr[8457] = -318174762;
assign addr[8458] = -299250668;
assign addr[8459] = -280302845;
assign addr[8460] = -261332796;
assign addr[8461] = -242342025;
assign addr[8462] = -223332037;
assign addr[8463] = -204304341;
assign addr[8464] = -185260444;
assign addr[8465] = -166201858;
assign addr[8466] = -147130093;
assign addr[8467] = -128046661;
assign addr[8468] = -108953076;
assign addr[8469] = -89850852;
assign addr[8470] = -70741503;
assign addr[8471] = -51626544;
assign addr[8472] = -32507492;
assign addr[8473] = -13385863;
assign addr[8474] = 5736829;
assign addr[8475] = 24859065;
assign addr[8476] = 43979330;
assign addr[8477] = 63096108;
assign addr[8478] = 82207882;
assign addr[8479] = 101313138;
assign addr[8480] = 120410361;
assign addr[8481] = 139498035;
assign addr[8482] = 158574649;
assign addr[8483] = 177638688;
assign addr[8484] = 196688642;
assign addr[8485] = 215722999;
assign addr[8486] = 234740251;
assign addr[8487] = 253738890;
assign addr[8488] = 272717408;
assign addr[8489] = 291674302;
assign addr[8490] = 310608068;
assign addr[8491] = 329517204;
assign addr[8492] = 348400212;
assign addr[8493] = 367255594;
assign addr[8494] = 386081854;
assign addr[8495] = 404877501;
assign addr[8496] = 423641043;
assign addr[8497] = 442370993;
assign addr[8498] = 461065866;
assign addr[8499] = 479724180;
assign addr[8500] = 498344454;
assign addr[8501] = 516925212;
assign addr[8502] = 535464981;
assign addr[8503] = 553962291;
assign addr[8504] = 572415676;
assign addr[8505] = 590823671;
assign addr[8506] = 609184818;
assign addr[8507] = 627497660;
assign addr[8508] = 645760745;
assign addr[8509] = 663972625;
assign addr[8510] = 682131857;
assign addr[8511] = 700236999;
assign addr[8512] = 718286617;
assign addr[8513] = 736279279;
assign addr[8514] = 754213559;
assign addr[8515] = 772088034;
assign addr[8516] = 789901288;
assign addr[8517] = 807651907;
assign addr[8518] = 825338484;
assign addr[8519] = 842959617;
assign addr[8520] = 860513908;
assign addr[8521] = 877999966;
assign addr[8522] = 895416404;
assign addr[8523] = 912761841;
assign addr[8524] = 930034901;
assign addr[8525] = 947234215;
assign addr[8526] = 964358420;
assign addr[8527] = 981406156;
assign addr[8528] = 998376073;
assign addr[8529] = 1015266825;
assign addr[8530] = 1032077073;
assign addr[8531] = 1048805483;
assign addr[8532] = 1065450729;
assign addr[8533] = 1082011492;
assign addr[8534] = 1098486458;
assign addr[8535] = 1114874320;
assign addr[8536] = 1131173780;
assign addr[8537] = 1147383544;
assign addr[8538] = 1163502328;
assign addr[8539] = 1179528853;
assign addr[8540] = 1195461849;
assign addr[8541] = 1211300053;
assign addr[8542] = 1227042207;
assign addr[8543] = 1242687064;
assign addr[8544] = 1258233384;
assign addr[8545] = 1273679934;
assign addr[8546] = 1289025489;
assign addr[8547] = 1304268832;
assign addr[8548] = 1319408754;
assign addr[8549] = 1334444055;
assign addr[8550] = 1349373543;
assign addr[8551] = 1364196034;
assign addr[8552] = 1378910353;
assign addr[8553] = 1393515332;
assign addr[8554] = 1408009814;
assign addr[8555] = 1422392650;
assign addr[8556] = 1436662698;
assign addr[8557] = 1450818828;
assign addr[8558] = 1464859917;
assign addr[8559] = 1478784851;
assign addr[8560] = 1492592527;
assign addr[8561] = 1506281850;
assign addr[8562] = 1519851733;
assign addr[8563] = 1533301101;
assign addr[8564] = 1546628888;
assign addr[8565] = 1559834037;
assign addr[8566] = 1572915501;
assign addr[8567] = 1585872242;
assign addr[8568] = 1598703233;
assign addr[8569] = 1611407456;
assign addr[8570] = 1623983905;
assign addr[8571] = 1636431582;
assign addr[8572] = 1648749499;
assign addr[8573] = 1660936681;
assign addr[8574] = 1672992161;
assign addr[8575] = 1684914983;
assign addr[8576] = 1696704201;
assign addr[8577] = 1708358881;
assign addr[8578] = 1719878099;
assign addr[8579] = 1731260941;
assign addr[8580] = 1742506504;
assign addr[8581] = 1753613897;
assign addr[8582] = 1764582240;
assign addr[8583] = 1775410662;
assign addr[8584] = 1786098304;
assign addr[8585] = 1796644320;
assign addr[8586] = 1807047873;
assign addr[8587] = 1817308138;
assign addr[8588] = 1827424302;
assign addr[8589] = 1837395562;
assign addr[8590] = 1847221128;
assign addr[8591] = 1856900221;
assign addr[8592] = 1866432072;
assign addr[8593] = 1875815927;
assign addr[8594] = 1885051042;
assign addr[8595] = 1894136683;
assign addr[8596] = 1903072131;
assign addr[8597] = 1911856677;
assign addr[8598] = 1920489624;
assign addr[8599] = 1928970288;
assign addr[8600] = 1937297997;
assign addr[8601] = 1945472089;
assign addr[8602] = 1953491918;
assign addr[8603] = 1961356847;
assign addr[8604] = 1969066252;
assign addr[8605] = 1976619522;
assign addr[8606] = 1984016058;
assign addr[8607] = 1991255274;
assign addr[8608] = 1998336596;
assign addr[8609] = 2005259462;
assign addr[8610] = 2012023322;
assign addr[8611] = 2018627642;
assign addr[8612] = 2025071897;
assign addr[8613] = 2031355576;
assign addr[8614] = 2037478181;
assign addr[8615] = 2043439226;
assign addr[8616] = 2049238240;
assign addr[8617] = 2054874761;
assign addr[8618] = 2060348343;
assign addr[8619] = 2065658552;
assign addr[8620] = 2070804967;
assign addr[8621] = 2075787180;
assign addr[8622] = 2080604795;
assign addr[8623] = 2085257431;
assign addr[8624] = 2089744719;
assign addr[8625] = 2094066304;
assign addr[8626] = 2098221841;
assign addr[8627] = 2102211002;
assign addr[8628] = 2106033471;
assign addr[8629] = 2109688944;
assign addr[8630] = 2113177132;
assign addr[8631] = 2116497758;
assign addr[8632] = 2119650558;
assign addr[8633] = 2122635283;
assign addr[8634] = 2125451696;
assign addr[8635] = 2128099574;
assign addr[8636] = 2130578706;
assign addr[8637] = 2132888897;
assign addr[8638] = 2135029962;
assign addr[8639] = 2137001733;
assign addr[8640] = 2138804053;
assign addr[8641] = 2140436778;
assign addr[8642] = 2141899780;
assign addr[8643] = 2143192942;
assign addr[8644] = 2144316162;
assign addr[8645] = 2145269351;
assign addr[8646] = 2146052433;
assign addr[8647] = 2146665347;
assign addr[8648] = 2147108043;
assign addr[8649] = 2147380486;
assign addr[8650] = 2147482655;
assign addr[8651] = 2147414542;
assign addr[8652] = 2147176152;
assign addr[8653] = 2146767505;
assign addr[8654] = 2146188631;
assign addr[8655] = 2145439578;
assign addr[8656] = 2144520405;
assign addr[8657] = 2143431184;
assign addr[8658] = 2142172003;
assign addr[8659] = 2140742960;
assign addr[8660] = 2139144169;
assign addr[8661] = 2137375758;
assign addr[8662] = 2135437865;
assign addr[8663] = 2133330646;
assign addr[8664] = 2131054266;
assign addr[8665] = 2128608907;
assign addr[8666] = 2125994762;
assign addr[8667] = 2123212038;
assign addr[8668] = 2120260957;
assign addr[8669] = 2117141752;
assign addr[8670] = 2113854671;
assign addr[8671] = 2110399974;
assign addr[8672] = 2106777935;
assign addr[8673] = 2102988841;
assign addr[8674] = 2099032994;
assign addr[8675] = 2094910706;
assign addr[8676] = 2090622304;
assign addr[8677] = 2086168128;
assign addr[8678] = 2081548533;
assign addr[8679] = 2076763883;
assign addr[8680] = 2071814558;
assign addr[8681] = 2066700952;
assign addr[8682] = 2061423468;
assign addr[8683] = 2055982526;
assign addr[8684] = 2050378558;
assign addr[8685] = 2044612007;
assign addr[8686] = 2038683330;
assign addr[8687] = 2032592999;
assign addr[8688] = 2026341495;
assign addr[8689] = 2019929315;
assign addr[8690] = 2013356967;
assign addr[8691] = 2006624971;
assign addr[8692] = 1999733863;
assign addr[8693] = 1992684188;
assign addr[8694] = 1985476506;
assign addr[8695] = 1978111387;
assign addr[8696] = 1970589416;
assign addr[8697] = 1962911189;
assign addr[8698] = 1955077316;
assign addr[8699] = 1947088417;
assign addr[8700] = 1938945125;
assign addr[8701] = 1930648088;
assign addr[8702] = 1922197961;
assign addr[8703] = 1913595416;
assign addr[8704] = 1904841135;
assign addr[8705] = 1895935811;
assign addr[8706] = 1886880151;
assign addr[8707] = 1877674873;
assign addr[8708] = 1868320707;
assign addr[8709] = 1858818395;
assign addr[8710] = 1849168689;
assign addr[8711] = 1839372356;
assign addr[8712] = 1829430172;
assign addr[8713] = 1819342925;
assign addr[8714] = 1809111415;
assign addr[8715] = 1798736454;
assign addr[8716] = 1788218865;
assign addr[8717] = 1777559480;
assign addr[8718] = 1766759146;
assign addr[8719] = 1755818718;
assign addr[8720] = 1744739065;
assign addr[8721] = 1733521064;
assign addr[8722] = 1722165606;
assign addr[8723] = 1710673591;
assign addr[8724] = 1699045930;
assign addr[8725] = 1687283545;
assign addr[8726] = 1675387369;
assign addr[8727] = 1663358344;
assign addr[8728] = 1651197426;
assign addr[8729] = 1638905577;
assign addr[8730] = 1626483774;
assign addr[8731] = 1613933000;
assign addr[8732] = 1601254251;
assign addr[8733] = 1588448533;
assign addr[8734] = 1575516860;
assign addr[8735] = 1562460258;
assign addr[8736] = 1549279763;
assign addr[8737] = 1535976419;
assign addr[8738] = 1522551282;
assign addr[8739] = 1509005416;
assign addr[8740] = 1495339895;
assign addr[8741] = 1481555802;
assign addr[8742] = 1467654232;
assign addr[8743] = 1453636285;
assign addr[8744] = 1439503074;
assign addr[8745] = 1425255719;
assign addr[8746] = 1410895350;
assign addr[8747] = 1396423105;
assign addr[8748] = 1381840133;
assign addr[8749] = 1367147589;
assign addr[8750] = 1352346639;
assign addr[8751] = 1337438456;
assign addr[8752] = 1322424222;
assign addr[8753] = 1307305128;
assign addr[8754] = 1292082373;
assign addr[8755] = 1276757164;
assign addr[8756] = 1261330715;
assign addr[8757] = 1245804251;
assign addr[8758] = 1230179002;
assign addr[8759] = 1214456207;
assign addr[8760] = 1198637114;
assign addr[8761] = 1182722976;
assign addr[8762] = 1166715055;
assign addr[8763] = 1150614620;
assign addr[8764] = 1134422949;
assign addr[8765] = 1118141326;
assign addr[8766] = 1101771040;
assign addr[8767] = 1085313391;
assign addr[8768] = 1068769683;
assign addr[8769] = 1052141228;
assign addr[8770] = 1035429345;
assign addr[8771] = 1018635358;
assign addr[8772] = 1001760600;
assign addr[8773] = 984806408;
assign addr[8774] = 967774128;
assign addr[8775] = 950665109;
assign addr[8776] = 933480707;
assign addr[8777] = 916222287;
assign addr[8778] = 898891215;
assign addr[8779] = 881488868;
assign addr[8780] = 864016623;
assign addr[8781] = 846475867;
assign addr[8782] = 828867991;
assign addr[8783] = 811194391;
assign addr[8784] = 793456467;
assign addr[8785] = 775655628;
assign addr[8786] = 757793284;
assign addr[8787] = 739870851;
assign addr[8788] = 721889752;
assign addr[8789] = 703851410;
assign addr[8790] = 685757258;
assign addr[8791] = 667608730;
assign addr[8792] = 649407264;
assign addr[8793] = 631154304;
assign addr[8794] = 612851297;
assign addr[8795] = 594499695;
assign addr[8796] = 576100953;
assign addr[8797] = 557656529;
assign addr[8798] = 539167887;
assign addr[8799] = 520636492;
assign addr[8800] = 502063814;
assign addr[8801] = 483451325;
assign addr[8802] = 464800501;
assign addr[8803] = 446112822;
assign addr[8804] = 427389768;
assign addr[8805] = 408632825;
assign addr[8806] = 389843480;
assign addr[8807] = 371023223;
assign addr[8808] = 352173546;
assign addr[8809] = 333295944;
assign addr[8810] = 314391913;
assign addr[8811] = 295462954;
assign addr[8812] = 276510565;
assign addr[8813] = 257536251;
assign addr[8814] = 238541516;
assign addr[8815] = 219527866;
assign addr[8816] = 200496809;
assign addr[8817] = 181449854;
assign addr[8818] = 162388511;
assign addr[8819] = 143314291;
assign addr[8820] = 124228708;
assign addr[8821] = 105133274;
assign addr[8822] = 86029503;
assign addr[8823] = 66918911;
assign addr[8824] = 47803013;
assign addr[8825] = 28683324;
assign addr[8826] = 9561361;
assign addr[8827] = -9561361;
assign addr[8828] = -28683324;
assign addr[8829] = -47803013;
assign addr[8830] = -66918911;
assign addr[8831] = -86029503;
assign addr[8832] = -105133274;
assign addr[8833] = -124228708;
assign addr[8834] = -143314291;
assign addr[8835] = -162388511;
assign addr[8836] = -181449854;
assign addr[8837] = -200496809;
assign addr[8838] = -219527866;
assign addr[8839] = -238541516;
assign addr[8840] = -257536251;
assign addr[8841] = -276510565;
assign addr[8842] = -295462954;
assign addr[8843] = -314391913;
assign addr[8844] = -333295944;
assign addr[8845] = -352173546;
assign addr[8846] = -371023223;
assign addr[8847] = -389843480;
assign addr[8848] = -408632825;
assign addr[8849] = -427389768;
assign addr[8850] = -446112822;
assign addr[8851] = -464800501;
assign addr[8852] = -483451325;
assign addr[8853] = -502063814;
assign addr[8854] = -520636492;
assign addr[8855] = -539167887;
assign addr[8856] = -557656529;
assign addr[8857] = -576100953;
assign addr[8858] = -594499695;
assign addr[8859] = -612851297;
assign addr[8860] = -631154304;
assign addr[8861] = -649407264;
assign addr[8862] = -667608730;
assign addr[8863] = -685757258;
assign addr[8864] = -703851410;
assign addr[8865] = -721889752;
assign addr[8866] = -739870851;
assign addr[8867] = -757793284;
assign addr[8868] = -775655628;
assign addr[8869] = -793456467;
assign addr[8870] = -811194391;
assign addr[8871] = -828867991;
assign addr[8872] = -846475867;
assign addr[8873] = -864016623;
assign addr[8874] = -881488868;
assign addr[8875] = -898891215;
assign addr[8876] = -916222287;
assign addr[8877] = -933480707;
assign addr[8878] = -950665109;
assign addr[8879] = -967774128;
assign addr[8880] = -984806408;
assign addr[8881] = -1001760600;
assign addr[8882] = -1018635358;
assign addr[8883] = -1035429345;
assign addr[8884] = -1052141228;
assign addr[8885] = -1068769683;
assign addr[8886] = -1085313391;
assign addr[8887] = -1101771040;
assign addr[8888] = -1118141326;
assign addr[8889] = -1134422949;
assign addr[8890] = -1150614620;
assign addr[8891] = -1166715055;
assign addr[8892] = -1182722976;
assign addr[8893] = -1198637114;
assign addr[8894] = -1214456207;
assign addr[8895] = -1230179002;
assign addr[8896] = -1245804251;
assign addr[8897] = -1261330715;
assign addr[8898] = -1276757164;
assign addr[8899] = -1292082373;
assign addr[8900] = -1307305128;
assign addr[8901] = -1322424222;
assign addr[8902] = -1337438456;
assign addr[8903] = -1352346639;
assign addr[8904] = -1367147589;
assign addr[8905] = -1381840133;
assign addr[8906] = -1396423105;
assign addr[8907] = -1410895350;
assign addr[8908] = -1425255719;
assign addr[8909] = -1439503074;
assign addr[8910] = -1453636285;
assign addr[8911] = -1467654232;
assign addr[8912] = -1481555802;
assign addr[8913] = -1495339895;
assign addr[8914] = -1509005416;
assign addr[8915] = -1522551282;
assign addr[8916] = -1535976419;
assign addr[8917] = -1549279763;
assign addr[8918] = -1562460258;
assign addr[8919] = -1575516860;
assign addr[8920] = -1588448533;
assign addr[8921] = -1601254251;
assign addr[8922] = -1613933000;
assign addr[8923] = -1626483774;
assign addr[8924] = -1638905577;
assign addr[8925] = -1651197426;
assign addr[8926] = -1663358344;
assign addr[8927] = -1675387369;
assign addr[8928] = -1687283545;
assign addr[8929] = -1699045930;
assign addr[8930] = -1710673591;
assign addr[8931] = -1722165606;
assign addr[8932] = -1733521064;
assign addr[8933] = -1744739065;
assign addr[8934] = -1755818718;
assign addr[8935] = -1766759146;
assign addr[8936] = -1777559480;
assign addr[8937] = -1788218865;
assign addr[8938] = -1798736454;
assign addr[8939] = -1809111415;
assign addr[8940] = -1819342925;
assign addr[8941] = -1829430172;
assign addr[8942] = -1839372356;
assign addr[8943] = -1849168689;
assign addr[8944] = -1858818395;
assign addr[8945] = -1868320707;
assign addr[8946] = -1877674873;
assign addr[8947] = -1886880151;
assign addr[8948] = -1895935811;
assign addr[8949] = -1904841135;
assign addr[8950] = -1913595416;
assign addr[8951] = -1922197961;
assign addr[8952] = -1930648088;
assign addr[8953] = -1938945125;
assign addr[8954] = -1947088417;
assign addr[8955] = -1955077316;
assign addr[8956] = -1962911189;
assign addr[8957] = -1970589416;
assign addr[8958] = -1978111387;
assign addr[8959] = -1985476506;
assign addr[8960] = -1992684188;
assign addr[8961] = -1999733863;
assign addr[8962] = -2006624971;
assign addr[8963] = -2013356967;
assign addr[8964] = -2019929315;
assign addr[8965] = -2026341495;
assign addr[8966] = -2032592999;
assign addr[8967] = -2038683330;
assign addr[8968] = -2044612007;
assign addr[8969] = -2050378558;
assign addr[8970] = -2055982526;
assign addr[8971] = -2061423468;
assign addr[8972] = -2066700952;
assign addr[8973] = -2071814558;
assign addr[8974] = -2076763883;
assign addr[8975] = -2081548533;
assign addr[8976] = -2086168128;
assign addr[8977] = -2090622304;
assign addr[8978] = -2094910706;
assign addr[8979] = -2099032994;
assign addr[8980] = -2102988841;
assign addr[8981] = -2106777935;
assign addr[8982] = -2110399974;
assign addr[8983] = -2113854671;
assign addr[8984] = -2117141752;
assign addr[8985] = -2120260957;
assign addr[8986] = -2123212038;
assign addr[8987] = -2125994762;
assign addr[8988] = -2128608907;
assign addr[8989] = -2131054266;
assign addr[8990] = -2133330646;
assign addr[8991] = -2135437865;
assign addr[8992] = -2137375758;
assign addr[8993] = -2139144169;
assign addr[8994] = -2140742960;
assign addr[8995] = -2142172003;
assign addr[8996] = -2143431184;
assign addr[8997] = -2144520405;
assign addr[8998] = -2145439578;
assign addr[8999] = -2146188631;
assign addr[9000] = -2146767505;
assign addr[9001] = -2147176152;
assign addr[9002] = -2147414542;
assign addr[9003] = -2147482655;
assign addr[9004] = -2147380486;
assign addr[9005] = -2147108043;
assign addr[9006] = -2146665347;
assign addr[9007] = -2146052433;
assign addr[9008] = -2145269351;
assign addr[9009] = -2144316162;
assign addr[9010] = -2143192942;
assign addr[9011] = -2141899780;
assign addr[9012] = -2140436778;
assign addr[9013] = -2138804053;
assign addr[9014] = -2137001733;
assign addr[9015] = -2135029962;
assign addr[9016] = -2132888897;
assign addr[9017] = -2130578706;
assign addr[9018] = -2128099574;
assign addr[9019] = -2125451696;
assign addr[9020] = -2122635283;
assign addr[9021] = -2119650558;
assign addr[9022] = -2116497758;
assign addr[9023] = -2113177132;
assign addr[9024] = -2109688944;
assign addr[9025] = -2106033471;
assign addr[9026] = -2102211002;
assign addr[9027] = -2098221841;
assign addr[9028] = -2094066304;
assign addr[9029] = -2089744719;
assign addr[9030] = -2085257431;
assign addr[9031] = -2080604795;
assign addr[9032] = -2075787180;
assign addr[9033] = -2070804967;
assign addr[9034] = -2065658552;
assign addr[9035] = -2060348343;
assign addr[9036] = -2054874761;
assign addr[9037] = -2049238240;
assign addr[9038] = -2043439226;
assign addr[9039] = -2037478181;
assign addr[9040] = -2031355576;
assign addr[9041] = -2025071897;
assign addr[9042] = -2018627642;
assign addr[9043] = -2012023322;
assign addr[9044] = -2005259462;
assign addr[9045] = -1998336596;
assign addr[9046] = -1991255274;
assign addr[9047] = -1984016058;
assign addr[9048] = -1976619522;
assign addr[9049] = -1969066252;
assign addr[9050] = -1961356847;
assign addr[9051] = -1953491918;
assign addr[9052] = -1945472089;
assign addr[9053] = -1937297997;
assign addr[9054] = -1928970288;
assign addr[9055] = -1920489624;
assign addr[9056] = -1911856677;
assign addr[9057] = -1903072131;
assign addr[9058] = -1894136683;
assign addr[9059] = -1885051042;
assign addr[9060] = -1875815927;
assign addr[9061] = -1866432072;
assign addr[9062] = -1856900221;
assign addr[9063] = -1847221128;
assign addr[9064] = -1837395562;
assign addr[9065] = -1827424302;
assign addr[9066] = -1817308138;
assign addr[9067] = -1807047873;
assign addr[9068] = -1796644320;
assign addr[9069] = -1786098304;
assign addr[9070] = -1775410662;
assign addr[9071] = -1764582240;
assign addr[9072] = -1753613897;
assign addr[9073] = -1742506504;
assign addr[9074] = -1731260941;
assign addr[9075] = -1719878099;
assign addr[9076] = -1708358881;
assign addr[9077] = -1696704201;
assign addr[9078] = -1684914983;
assign addr[9079] = -1672992161;
assign addr[9080] = -1660936681;
assign addr[9081] = -1648749499;
assign addr[9082] = -1636431582;
assign addr[9083] = -1623983905;
assign addr[9084] = -1611407456;
assign addr[9085] = -1598703233;
assign addr[9086] = -1585872242;
assign addr[9087] = -1572915501;
assign addr[9088] = -1559834037;
assign addr[9089] = -1546628888;
assign addr[9090] = -1533301101;
assign addr[9091] = -1519851733;
assign addr[9092] = -1506281850;
assign addr[9093] = -1492592527;
assign addr[9094] = -1478784851;
assign addr[9095] = -1464859917;
assign addr[9096] = -1450818828;
assign addr[9097] = -1436662698;
assign addr[9098] = -1422392650;
assign addr[9099] = -1408009814;
assign addr[9100] = -1393515332;
assign addr[9101] = -1378910353;
assign addr[9102] = -1364196034;
assign addr[9103] = -1349373543;
assign addr[9104] = -1334444055;
assign addr[9105] = -1319408754;
assign addr[9106] = -1304268832;
assign addr[9107] = -1289025489;
assign addr[9108] = -1273679934;
assign addr[9109] = -1258233384;
assign addr[9110] = -1242687064;
assign addr[9111] = -1227042207;
assign addr[9112] = -1211300053;
assign addr[9113] = -1195461849;
assign addr[9114] = -1179528853;
assign addr[9115] = -1163502328;
assign addr[9116] = -1147383544;
assign addr[9117] = -1131173780;
assign addr[9118] = -1114874320;
assign addr[9119] = -1098486458;
assign addr[9120] = -1082011492;
assign addr[9121] = -1065450729;
assign addr[9122] = -1048805483;
assign addr[9123] = -1032077073;
assign addr[9124] = -1015266825;
assign addr[9125] = -998376073;
assign addr[9126] = -981406156;
assign addr[9127] = -964358420;
assign addr[9128] = -947234215;
assign addr[9129] = -930034901;
assign addr[9130] = -912761841;
assign addr[9131] = -895416404;
assign addr[9132] = -877999966;
assign addr[9133] = -860513908;
assign addr[9134] = -842959617;
assign addr[9135] = -825338484;
assign addr[9136] = -807651907;
assign addr[9137] = -789901288;
assign addr[9138] = -772088034;
assign addr[9139] = -754213559;
assign addr[9140] = -736279279;
assign addr[9141] = -718286617;
assign addr[9142] = -700236999;
assign addr[9143] = -682131857;
assign addr[9144] = -663972625;
assign addr[9145] = -645760745;
assign addr[9146] = -627497660;
assign addr[9147] = -609184818;
assign addr[9148] = -590823671;
assign addr[9149] = -572415676;
assign addr[9150] = -553962291;
assign addr[9151] = -535464981;
assign addr[9152] = -516925212;
assign addr[9153] = -498344454;
assign addr[9154] = -479724180;
assign addr[9155] = -461065866;
assign addr[9156] = -442370993;
assign addr[9157] = -423641043;
assign addr[9158] = -404877501;
assign addr[9159] = -386081854;
assign addr[9160] = -367255594;
assign addr[9161] = -348400212;
assign addr[9162] = -329517204;
assign addr[9163] = -310608068;
assign addr[9164] = -291674302;
assign addr[9165] = -272717408;
assign addr[9166] = -253738890;
assign addr[9167] = -234740251;
assign addr[9168] = -215722999;
assign addr[9169] = -196688642;
assign addr[9170] = -177638688;
assign addr[9171] = -158574649;
assign addr[9172] = -139498035;
assign addr[9173] = -120410361;
assign addr[9174] = -101313138;
assign addr[9175] = -82207882;
assign addr[9176] = -63096108;
assign addr[9177] = -43979330;
assign addr[9178] = -24859065;
assign addr[9179] = -5736829;
assign addr[9180] = 13385863;
assign addr[9181] = 32507492;
assign addr[9182] = 51626544;
assign addr[9183] = 70741503;
assign addr[9184] = 89850852;
assign addr[9185] = 108953076;
assign addr[9186] = 128046661;
assign addr[9187] = 147130093;
assign addr[9188] = 166201858;
assign addr[9189] = 185260444;
assign addr[9190] = 204304341;
assign addr[9191] = 223332037;
assign addr[9192] = 242342025;
assign addr[9193] = 261332796;
assign addr[9194] = 280302845;
assign addr[9195] = 299250668;
assign addr[9196] = 318174762;
assign addr[9197] = 337073627;
assign addr[9198] = 355945764;
assign addr[9199] = 374789676;
assign addr[9200] = 393603870;
assign addr[9201] = 412386854;
assign addr[9202] = 431137138;
assign addr[9203] = 449853235;
assign addr[9204] = 468533662;
assign addr[9205] = 487176937;
assign addr[9206] = 505781581;
assign addr[9207] = 524346121;
assign addr[9208] = 542869083;
assign addr[9209] = 561348998;
assign addr[9210] = 579784402;
assign addr[9211] = 598173833;
assign addr[9212] = 616515832;
assign addr[9213] = 634808946;
assign addr[9214] = 653051723;
assign addr[9215] = 671242716;
assign addr[9216] = 689380485;
assign addr[9217] = 707463589;
assign addr[9218] = 725490597;
assign addr[9219] = 743460077;
assign addr[9220] = 761370605;
assign addr[9221] = 779220762;
assign addr[9222] = 797009130;
assign addr[9223] = 814734301;
assign addr[9224] = 832394869;
assign addr[9225] = 849989433;
assign addr[9226] = 867516597;
assign addr[9227] = 884974973;
assign addr[9228] = 902363176;
assign addr[9229] = 919679827;
assign addr[9230] = 936923553;
assign addr[9231] = 954092986;
assign addr[9232] = 971186766;
assign addr[9233] = 988203537;
assign addr[9234] = 1005141949;
assign addr[9235] = 1022000660;
assign addr[9236] = 1038778332;
assign addr[9237] = 1055473635;
assign addr[9238] = 1072085246;
assign addr[9239] = 1088611847;
assign addr[9240] = 1105052128;
assign addr[9241] = 1121404785;
assign addr[9242] = 1137668521;
assign addr[9243] = 1153842047;
assign addr[9244] = 1169924081;
assign addr[9245] = 1185913346;
assign addr[9246] = 1201808576;
assign addr[9247] = 1217608510;
assign addr[9248] = 1233311895;
assign addr[9249] = 1248917486;
assign addr[9250] = 1264424045;
assign addr[9251] = 1279830344;
assign addr[9252] = 1295135159;
assign addr[9253] = 1310337279;
assign addr[9254] = 1325435496;
assign addr[9255] = 1340428615;
assign addr[9256] = 1355315445;
assign addr[9257] = 1370094808;
assign addr[9258] = 1384765530;
assign addr[9259] = 1399326449;
assign addr[9260] = 1413776410;
assign addr[9261] = 1428114267;
assign addr[9262] = 1442338884;
assign addr[9263] = 1456449131;
assign addr[9264] = 1470443891;
assign addr[9265] = 1484322054;
assign addr[9266] = 1498082520;
assign addr[9267] = 1511724196;
assign addr[9268] = 1525246002;
assign addr[9269] = 1538646865;
assign addr[9270] = 1551925723;
assign addr[9271] = 1565081523;
assign addr[9272] = 1578113222;
assign addr[9273] = 1591019785;
assign addr[9274] = 1603800191;
assign addr[9275] = 1616453425;
assign addr[9276] = 1628978484;
assign addr[9277] = 1641374375;
assign addr[9278] = 1653640115;
assign addr[9279] = 1665774731;
assign addr[9280] = 1677777262;
assign addr[9281] = 1689646755;
assign addr[9282] = 1701382270;
assign addr[9283] = 1712982875;
assign addr[9284] = 1724447652;
assign addr[9285] = 1735775690;
assign addr[9286] = 1746966091;
assign addr[9287] = 1758017969;
assign addr[9288] = 1768930447;
assign addr[9289] = 1779702660;
assign addr[9290] = 1790333753;
assign addr[9291] = 1800822883;
assign addr[9292] = 1811169220;
assign addr[9293] = 1821371941;
assign addr[9294] = 1831430239;
assign addr[9295] = 1841343316;
assign addr[9296] = 1851110385;
assign addr[9297] = 1860730673;
assign addr[9298] = 1870203416;
assign addr[9299] = 1879527863;
assign addr[9300] = 1888703276;
assign addr[9301] = 1897728925;
assign addr[9302] = 1906604097;
assign addr[9303] = 1915328086;
assign addr[9304] = 1923900201;
assign addr[9305] = 1932319763;
assign addr[9306] = 1940586104;
assign addr[9307] = 1948698568;
assign addr[9308] = 1956656513;
assign addr[9309] = 1964459306;
assign addr[9310] = 1972106330;
assign addr[9311] = 1979596978;
assign addr[9312] = 1986930656;
assign addr[9313] = 1994106782;
assign addr[9314] = 2001124788;
assign addr[9315] = 2007984117;
assign addr[9316] = 2014684225;
assign addr[9317] = 2021224581;
assign addr[9318] = 2027604666;
assign addr[9319] = 2033823974;
assign addr[9320] = 2039882013;
assign addr[9321] = 2045778302;
assign addr[9322] = 2051512372;
assign addr[9323] = 2057083771;
assign addr[9324] = 2062492055;
assign addr[9325] = 2067736796;
assign addr[9326] = 2072817579;
assign addr[9327] = 2077733999;
assign addr[9328] = 2082485668;
assign addr[9329] = 2087072209;
assign addr[9330] = 2091493257;
assign addr[9331] = 2095748463;
assign addr[9332] = 2099837489;
assign addr[9333] = 2103760010;
assign addr[9334] = 2107515716;
assign addr[9335] = 2111104309;
assign addr[9336] = 2114525505;
assign addr[9337] = 2117779031;
assign addr[9338] = 2120864631;
assign addr[9339] = 2123782059;
assign addr[9340] = 2126531084;
assign addr[9341] = 2129111488;
assign addr[9342] = 2131523066;
assign addr[9343] = 2133765628;
assign addr[9344] = 2135838995;
assign addr[9345] = 2137743003;
assign addr[9346] = 2139477502;
assign addr[9347] = 2141042352;
assign addr[9348] = 2142437431;
assign addr[9349] = 2143662628;
assign addr[9350] = 2144717846;
assign addr[9351] = 2145603001;
assign addr[9352] = 2146318022;
assign addr[9353] = 2146862854;
assign addr[9354] = 2147237452;
assign addr[9355] = 2147441787;
assign addr[9356] = 2147475844;
assign addr[9357] = 2147339619;
assign addr[9358] = 2147033123;
assign addr[9359] = 2146556380;
assign addr[9360] = 2145909429;
assign addr[9361] = 2145092320;
assign addr[9362] = 2144105118;
assign addr[9363] = 2142947902;
assign addr[9364] = 2141620763;
assign addr[9365] = 2140123807;
assign addr[9366] = 2138457152;
assign addr[9367] = 2136620930;
assign addr[9368] = 2134615288;
assign addr[9369] = 2132440383;
assign addr[9370] = 2130096389;
assign addr[9371] = 2127583492;
assign addr[9372] = 2124901890;
assign addr[9373] = 2122051796;
assign addr[9374] = 2119033436;
assign addr[9375] = 2115847050;
assign addr[9376] = 2112492891;
assign addr[9377] = 2108971223;
assign addr[9378] = 2105282327;
assign addr[9379] = 2101426496;
assign addr[9380] = 2097404033;
assign addr[9381] = 2093215260;
assign addr[9382] = 2088860507;
assign addr[9383] = 2084340120;
assign addr[9384] = 2079654458;
assign addr[9385] = 2074803892;
assign addr[9386] = 2069788807;
assign addr[9387] = 2064609600;
assign addr[9388] = 2059266683;
assign addr[9389] = 2053760478;
assign addr[9390] = 2048091422;
assign addr[9391] = 2042259965;
assign addr[9392] = 2036266570;
assign addr[9393] = 2030111710;
assign addr[9394] = 2023795876;
assign addr[9395] = 2017319567;
assign addr[9396] = 2010683297;
assign addr[9397] = 2003887591;
assign addr[9398] = 1996932990;
assign addr[9399] = 1989820044;
assign addr[9400] = 1982549318;
assign addr[9401] = 1975121388;
assign addr[9402] = 1967536842;
assign addr[9403] = 1959796283;
assign addr[9404] = 1951900324;
assign addr[9405] = 1943849591;
assign addr[9406] = 1935644723;
assign addr[9407] = 1927286370;
assign addr[9408] = 1918775195;
assign addr[9409] = 1910111873;
assign addr[9410] = 1901297091;
assign addr[9411] = 1892331547;
assign addr[9412] = 1883215953;
assign addr[9413] = 1873951032;
assign addr[9414] = 1864537518;
assign addr[9415] = 1854976157;
assign addr[9416] = 1845267708;
assign addr[9417] = 1835412941;
assign addr[9418] = 1825412636;
assign addr[9419] = 1815267588;
assign addr[9420] = 1804978599;
assign addr[9421] = 1794546487;
assign addr[9422] = 1783972079;
assign addr[9423] = 1773256212;
assign addr[9424] = 1762399737;
assign addr[9425] = 1751403515;
assign addr[9426] = 1740268417;
assign addr[9427] = 1728995326;
assign addr[9428] = 1717585136;
assign addr[9429] = 1706038753;
assign addr[9430] = 1694357091;
assign addr[9431] = 1682541077;
assign addr[9432] = 1670591647;
assign addr[9433] = 1658509750;
assign addr[9434] = 1646296344;
assign addr[9435] = 1633952396;
assign addr[9436] = 1621478885;
assign addr[9437] = 1608876801;
assign addr[9438] = 1596147143;
assign addr[9439] = 1583290921;
assign addr[9440] = 1570309153;
assign addr[9441] = 1557202869;
assign addr[9442] = 1543973108;
assign addr[9443] = 1530620920;
assign addr[9444] = 1517147363;
assign addr[9445] = 1503553506;
assign addr[9446] = 1489840425;
assign addr[9447] = 1476009210;
assign addr[9448] = 1462060956;
assign addr[9449] = 1447996770;
assign addr[9450] = 1433817766;
assign addr[9451] = 1419525069;
assign addr[9452] = 1405119813;
assign addr[9453] = 1390603139;
assign addr[9454] = 1375976199;
assign addr[9455] = 1361240152;
assign addr[9456] = 1346396168;
assign addr[9457] = 1331445422;
assign addr[9458] = 1316389101;
assign addr[9459] = 1301228398;
assign addr[9460] = 1285964516;
assign addr[9461] = 1270598665;
assign addr[9462] = 1255132063;
assign addr[9463] = 1239565936;
assign addr[9464] = 1223901520;
assign addr[9465] = 1208140056;
assign addr[9466] = 1192282793;
assign addr[9467] = 1176330990;
assign addr[9468] = 1160285911;
assign addr[9469] = 1144148829;
assign addr[9470] = 1127921022;
assign addr[9471] = 1111603778;
assign addr[9472] = 1095198391;
assign addr[9473] = 1078706161;
assign addr[9474] = 1062128397;
assign addr[9475] = 1045466412;
assign addr[9476] = 1028721528;
assign addr[9477] = 1011895073;
assign addr[9478] = 994988380;
assign addr[9479] = 978002791;
assign addr[9480] = 960939653;
assign addr[9481] = 943800318;
assign addr[9482] = 926586145;
assign addr[9483] = 909298500;
assign addr[9484] = 891938752;
assign addr[9485] = 874508280;
assign addr[9486] = 857008464;
assign addr[9487] = 839440693;
assign addr[9488] = 821806359;
assign addr[9489] = 804106861;
assign addr[9490] = 786343603;
assign addr[9491] = 768517992;
assign addr[9492] = 750631442;
assign addr[9493] = 732685372;
assign addr[9494] = 714681204;
assign addr[9495] = 696620367;
assign addr[9496] = 678504291;
assign addr[9497] = 660334415;
assign addr[9498] = 642112178;
assign addr[9499] = 623839025;
assign addr[9500] = 605516406;
assign addr[9501] = 587145773;
assign addr[9502] = 568728583;
assign addr[9503] = 550266296;
assign addr[9504] = 531760377;
assign addr[9505] = 513212292;
assign addr[9506] = 494623513;
assign addr[9507] = 475995513;
assign addr[9508] = 457329769;
assign addr[9509] = 438627762;
assign addr[9510] = 419890975;
assign addr[9511] = 401120892;
assign addr[9512] = 382319004;
assign addr[9513] = 363486799;
assign addr[9514] = 344625773;
assign addr[9515] = 325737419;
assign addr[9516] = 306823237;
assign addr[9517] = 287884725;
assign addr[9518] = 268923386;
assign addr[9519] = 249940723;
assign addr[9520] = 230938242;
assign addr[9521] = 211917448;
assign addr[9522] = 192879850;
assign addr[9523] = 173826959;
assign addr[9524] = 154760284;
assign addr[9525] = 135681337;
assign addr[9526] = 116591632;
assign addr[9527] = 97492681;
assign addr[9528] = 78386000;
assign addr[9529] = 59273104;
assign addr[9530] = 40155507;
assign addr[9531] = 21034727;
assign addr[9532] = 1912278;
assign addr[9533] = -17210322;
assign addr[9534] = -36331557;
assign addr[9535] = -55449912;
assign addr[9536] = -74563870;
assign addr[9537] = -93671915;
assign addr[9538] = -112772533;
assign addr[9539] = -131864208;
assign addr[9540] = -150945428;
assign addr[9541] = -170014678;
assign addr[9542] = -189070447;
assign addr[9543] = -208111224;
assign addr[9544] = -227135500;
assign addr[9545] = -246141764;
assign addr[9546] = -265128512;
assign addr[9547] = -284094236;
assign addr[9548] = -303037433;
assign addr[9549] = -321956601;
assign addr[9550] = -340850240;
assign addr[9551] = -359716852;
assign addr[9552] = -378554940;
assign addr[9553] = -397363011;
assign addr[9554] = -416139574;
assign addr[9555] = -434883140;
assign addr[9556] = -453592221;
assign addr[9557] = -472265336;
assign addr[9558] = -490901003;
assign addr[9559] = -509497745;
assign addr[9560] = -528054086;
assign addr[9561] = -546568556;
assign addr[9562] = -565039687;
assign addr[9563] = -583466013;
assign addr[9564] = -601846074;
assign addr[9565] = -620178412;
assign addr[9566] = -638461574;
assign addr[9567] = -656694110;
assign addr[9568] = -674874574;
assign addr[9569] = -693001525;
assign addr[9570] = -711073524;
assign addr[9571] = -729089140;
assign addr[9572] = -747046944;
assign addr[9573] = -764945512;
assign addr[9574] = -782783424;
assign addr[9575] = -800559266;
assign addr[9576] = -818271628;
assign addr[9577] = -835919107;
assign addr[9578] = -853500302;
assign addr[9579] = -871013820;
assign addr[9580] = -888458272;
assign addr[9581] = -905832274;
assign addr[9582] = -923134450;
assign addr[9583] = -940363427;
assign addr[9584] = -957517838;
assign addr[9585] = -974596324;
assign addr[9586] = -991597531;
assign addr[9587] = -1008520110;
assign addr[9588] = -1025362720;
assign addr[9589] = -1042124025;
assign addr[9590] = -1058802695;
assign addr[9591] = -1075397409;
assign addr[9592] = -1091906851;
assign addr[9593] = -1108329711;
assign addr[9594] = -1124664687;
assign addr[9595] = -1140910484;
assign addr[9596] = -1157065814;
assign addr[9597] = -1173129396;
assign addr[9598] = -1189099956;
assign addr[9599] = -1204976227;
assign addr[9600] = -1220756951;
assign addr[9601] = -1236440877;
assign addr[9602] = -1252026760;
assign addr[9603] = -1267513365;
assign addr[9604] = -1282899464;
assign addr[9605] = -1298183838;
assign addr[9606] = -1313365273;
assign addr[9607] = -1328442566;
assign addr[9608] = -1343414522;
assign addr[9609] = -1358279953;
assign addr[9610] = -1373037681;
assign addr[9611] = -1387686535;
assign addr[9612] = -1402225355;
assign addr[9613] = -1416652986;
assign addr[9614] = -1430968286;
assign addr[9615] = -1445170118;
assign addr[9616] = -1459257358;
assign addr[9617] = -1473228887;
assign addr[9618] = -1487083598;
assign addr[9619] = -1500820393;
assign addr[9620] = -1514438181;
assign addr[9621] = -1527935884;
assign addr[9622] = -1541312431;
assign addr[9623] = -1554566762;
assign addr[9624] = -1567697824;
assign addr[9625] = -1580704578;
assign addr[9626] = -1593585992;
assign addr[9627] = -1606341043;
assign addr[9628] = -1618968722;
assign addr[9629] = -1631468027;
assign addr[9630] = -1643837966;
assign addr[9631] = -1656077559;
assign addr[9632] = -1668185835;
assign addr[9633] = -1680161834;
assign addr[9634] = -1692004606;
assign addr[9635] = -1703713213;
assign addr[9636] = -1715286726;
assign addr[9637] = -1726724227;
assign addr[9638] = -1738024810;
assign addr[9639] = -1749187577;
assign addr[9640] = -1760211645;
assign addr[9641] = -1771096139;
assign addr[9642] = -1781840195;
assign addr[9643] = -1792442963;
assign addr[9644] = -1802903601;
assign addr[9645] = -1813221279;
assign addr[9646] = -1823395180;
assign addr[9647] = -1833424497;
assign addr[9648] = -1843308435;
assign addr[9649] = -1853046210;
assign addr[9650] = -1862637049;
assign addr[9651] = -1872080193;
assign addr[9652] = -1881374892;
assign addr[9653] = -1890520410;
assign addr[9654] = -1899516021;
assign addr[9655] = -1908361011;
assign addr[9656] = -1917054681;
assign addr[9657] = -1925596340;
assign addr[9658] = -1933985310;
assign addr[9659] = -1942220928;
assign addr[9660] = -1950302539;
assign addr[9661] = -1958229503;
assign addr[9662] = -1966001192;
assign addr[9663] = -1973616989;
assign addr[9664] = -1981076290;
assign addr[9665] = -1988378503;
assign addr[9666] = -1995523051;
assign addr[9667] = -2002509365;
assign addr[9668] = -2009336893;
assign addr[9669] = -2016005093;
assign addr[9670] = -2022513436;
assign addr[9671] = -2028861406;
assign addr[9672] = -2035048499;
assign addr[9673] = -2041074226;
assign addr[9674] = -2046938108;
assign addr[9675] = -2052639680;
assign addr[9676] = -2058178491;
assign addr[9677] = -2063554100;
assign addr[9678] = -2068766083;
assign addr[9679] = -2073814024;
assign addr[9680] = -2078697525;
assign addr[9681] = -2083416198;
assign addr[9682] = -2087969669;
assign addr[9683] = -2092357577;
assign addr[9684] = -2096579573;
assign addr[9685] = -2100635323;
assign addr[9686] = -2104524506;
assign addr[9687] = -2108246813;
assign addr[9688] = -2111801949;
assign addr[9689] = -2115189632;
assign addr[9690] = -2118409593;
assign addr[9691] = -2121461578;
assign addr[9692] = -2124345343;
assign addr[9693] = -2127060661;
assign addr[9694] = -2129607316;
assign addr[9695] = -2131985106;
assign addr[9696] = -2134193842;
assign addr[9697] = -2136233350;
assign addr[9698] = -2138103468;
assign addr[9699] = -2139804048;
assign addr[9700] = -2141334954;
assign addr[9701] = -2142696065;
assign addr[9702] = -2143887273;
assign addr[9703] = -2144908484;
assign addr[9704] = -2145759618;
assign addr[9705] = -2146440605;
assign addr[9706] = -2146951393;
assign addr[9707] = -2147291941;
assign addr[9708] = -2147462221;
assign addr[9709] = -2147462221;
assign addr[9710] = -2147291941;
assign addr[9711] = -2146951393;
assign addr[9712] = -2146440605;
assign addr[9713] = -2145759618;
assign addr[9714] = -2144908484;
assign addr[9715] = -2143887273;
assign addr[9716] = -2142696065;
assign addr[9717] = -2141334954;
assign addr[9718] = -2139804048;
assign addr[9719] = -2138103468;
assign addr[9720] = -2136233350;
assign addr[9721] = -2134193842;
assign addr[9722] = -2131985106;
assign addr[9723] = -2129607316;
assign addr[9724] = -2127060661;
assign addr[9725] = -2124345343;
assign addr[9726] = -2121461578;
assign addr[9727] = -2118409593;
assign addr[9728] = -2115189632;
assign addr[9729] = -2111801949;
assign addr[9730] = -2108246813;
assign addr[9731] = -2104524506;
assign addr[9732] = -2100635323;
assign addr[9733] = -2096579573;
assign addr[9734] = -2092357577;
assign addr[9735] = -2087969669;
assign addr[9736] = -2083416198;
assign addr[9737] = -2078697525;
assign addr[9738] = -2073814024;
assign addr[9739] = -2068766083;
assign addr[9740] = -2063554100;
assign addr[9741] = -2058178491;
assign addr[9742] = -2052639680;
assign addr[9743] = -2046938108;
assign addr[9744] = -2041074226;
assign addr[9745] = -2035048499;
assign addr[9746] = -2028861406;
assign addr[9747] = -2022513436;
assign addr[9748] = -2016005093;
assign addr[9749] = -2009336893;
assign addr[9750] = -2002509365;
assign addr[9751] = -1995523051;
assign addr[9752] = -1988378503;
assign addr[9753] = -1981076290;
assign addr[9754] = -1973616989;
assign addr[9755] = -1966001192;
assign addr[9756] = -1958229503;
assign addr[9757] = -1950302539;
assign addr[9758] = -1942220928;
assign addr[9759] = -1933985310;
assign addr[9760] = -1925596340;
assign addr[9761] = -1917054681;
assign addr[9762] = -1908361011;
assign addr[9763] = -1899516021;
assign addr[9764] = -1890520410;
assign addr[9765] = -1881374892;
assign addr[9766] = -1872080193;
assign addr[9767] = -1862637049;
assign addr[9768] = -1853046210;
assign addr[9769] = -1843308435;
assign addr[9770] = -1833424497;
assign addr[9771] = -1823395180;
assign addr[9772] = -1813221279;
assign addr[9773] = -1802903601;
assign addr[9774] = -1792442963;
assign addr[9775] = -1781840195;
assign addr[9776] = -1771096139;
assign addr[9777] = -1760211645;
assign addr[9778] = -1749187577;
assign addr[9779] = -1738024810;
assign addr[9780] = -1726724227;
assign addr[9781] = -1715286726;
assign addr[9782] = -1703713213;
assign addr[9783] = -1692004606;
assign addr[9784] = -1680161834;
assign addr[9785] = -1668185835;
assign addr[9786] = -1656077559;
assign addr[9787] = -1643837966;
assign addr[9788] = -1631468027;
assign addr[9789] = -1618968722;
assign addr[9790] = -1606341043;
assign addr[9791] = -1593585992;
assign addr[9792] = -1580704578;
assign addr[9793] = -1567697824;
assign addr[9794] = -1554566762;
assign addr[9795] = -1541312431;
assign addr[9796] = -1527935884;
assign addr[9797] = -1514438181;
assign addr[9798] = -1500820393;
assign addr[9799] = -1487083598;
assign addr[9800] = -1473228887;
assign addr[9801] = -1459257358;
assign addr[9802] = -1445170118;
assign addr[9803] = -1430968286;
assign addr[9804] = -1416652986;
assign addr[9805] = -1402225355;
assign addr[9806] = -1387686535;
assign addr[9807] = -1373037681;
assign addr[9808] = -1358279953;
assign addr[9809] = -1343414522;
assign addr[9810] = -1328442566;
assign addr[9811] = -1313365273;
assign addr[9812] = -1298183838;
assign addr[9813] = -1282899464;
assign addr[9814] = -1267513365;
assign addr[9815] = -1252026760;
assign addr[9816] = -1236440877;
assign addr[9817] = -1220756951;
assign addr[9818] = -1204976227;
assign addr[9819] = -1189099956;
assign addr[9820] = -1173129396;
assign addr[9821] = -1157065814;
assign addr[9822] = -1140910484;
assign addr[9823] = -1124664687;
assign addr[9824] = -1108329711;
assign addr[9825] = -1091906851;
assign addr[9826] = -1075397409;
assign addr[9827] = -1058802695;
assign addr[9828] = -1042124025;
assign addr[9829] = -1025362720;
assign addr[9830] = -1008520110;
assign addr[9831] = -991597531;
assign addr[9832] = -974596324;
assign addr[9833] = -957517838;
assign addr[9834] = -940363427;
assign addr[9835] = -923134450;
assign addr[9836] = -905832274;
assign addr[9837] = -888458272;
assign addr[9838] = -871013820;
assign addr[9839] = -853500302;
assign addr[9840] = -835919107;
assign addr[9841] = -818271628;
assign addr[9842] = -800559266;
assign addr[9843] = -782783424;
assign addr[9844] = -764945512;
assign addr[9845] = -747046944;
assign addr[9846] = -729089140;
assign addr[9847] = -711073524;
assign addr[9848] = -693001525;
assign addr[9849] = -674874574;
assign addr[9850] = -656694110;
assign addr[9851] = -638461574;
assign addr[9852] = -620178412;
assign addr[9853] = -601846074;
assign addr[9854] = -583466013;
assign addr[9855] = -565039687;
assign addr[9856] = -546568556;
assign addr[9857] = -528054086;
assign addr[9858] = -509497745;
assign addr[9859] = -490901003;
assign addr[9860] = -472265336;
assign addr[9861] = -453592221;
assign addr[9862] = -434883140;
assign addr[9863] = -416139574;
assign addr[9864] = -397363011;
assign addr[9865] = -378554940;
assign addr[9866] = -359716852;
assign addr[9867] = -340850240;
assign addr[9868] = -321956601;
assign addr[9869] = -303037433;
assign addr[9870] = -284094236;
assign addr[9871] = -265128512;
assign addr[9872] = -246141764;
assign addr[9873] = -227135500;
assign addr[9874] = -208111224;
assign addr[9875] = -189070447;
assign addr[9876] = -170014678;
assign addr[9877] = -150945428;
assign addr[9878] = -131864208;
assign addr[9879] = -112772533;
assign addr[9880] = -93671915;
assign addr[9881] = -74563870;
assign addr[9882] = -55449912;
assign addr[9883] = -36331557;
assign addr[9884] = -17210322;
assign addr[9885] = 1912278;
assign addr[9886] = 21034727;
assign addr[9887] = 40155507;
assign addr[9888] = 59273104;
assign addr[9889] = 78386000;
assign addr[9890] = 97492681;
assign addr[9891] = 116591632;
assign addr[9892] = 135681337;
assign addr[9893] = 154760284;
assign addr[9894] = 173826959;
assign addr[9895] = 192879850;
assign addr[9896] = 211917448;
assign addr[9897] = 230938242;
assign addr[9898] = 249940723;
assign addr[9899] = 268923386;
assign addr[9900] = 287884725;
assign addr[9901] = 306823237;
assign addr[9902] = 325737419;
assign addr[9903] = 344625773;
assign addr[9904] = 363486799;
assign addr[9905] = 382319004;
assign addr[9906] = 401120892;
assign addr[9907] = 419890975;
assign addr[9908] = 438627762;
assign addr[9909] = 457329769;
assign addr[9910] = 475995513;
assign addr[9911] = 494623513;
assign addr[9912] = 513212292;
assign addr[9913] = 531760377;
assign addr[9914] = 550266296;
assign addr[9915] = 568728583;
assign addr[9916] = 587145773;
assign addr[9917] = 605516406;
assign addr[9918] = 623839025;
assign addr[9919] = 642112178;
assign addr[9920] = 660334415;
assign addr[9921] = 678504291;
assign addr[9922] = 696620367;
assign addr[9923] = 714681204;
assign addr[9924] = 732685372;
assign addr[9925] = 750631442;
assign addr[9926] = 768517992;
assign addr[9927] = 786343603;
assign addr[9928] = 804106861;
assign addr[9929] = 821806359;
assign addr[9930] = 839440693;
assign addr[9931] = 857008464;
assign addr[9932] = 874508280;
assign addr[9933] = 891938752;
assign addr[9934] = 909298500;
assign addr[9935] = 926586145;
assign addr[9936] = 943800318;
assign addr[9937] = 960939653;
assign addr[9938] = 978002791;
assign addr[9939] = 994988380;
assign addr[9940] = 1011895073;
assign addr[9941] = 1028721528;
assign addr[9942] = 1045466412;
assign addr[9943] = 1062128397;
assign addr[9944] = 1078706161;
assign addr[9945] = 1095198391;
assign addr[9946] = 1111603778;
assign addr[9947] = 1127921022;
assign addr[9948] = 1144148829;
assign addr[9949] = 1160285911;
assign addr[9950] = 1176330990;
assign addr[9951] = 1192282793;
assign addr[9952] = 1208140056;
assign addr[9953] = 1223901520;
assign addr[9954] = 1239565936;
assign addr[9955] = 1255132063;
assign addr[9956] = 1270598665;
assign addr[9957] = 1285964516;
assign addr[9958] = 1301228398;
assign addr[9959] = 1316389101;
assign addr[9960] = 1331445422;
assign addr[9961] = 1346396168;
assign addr[9962] = 1361240152;
assign addr[9963] = 1375976199;
assign addr[9964] = 1390603139;
assign addr[9965] = 1405119813;
assign addr[9966] = 1419525069;
assign addr[9967] = 1433817766;
assign addr[9968] = 1447996770;
assign addr[9969] = 1462060956;
assign addr[9970] = 1476009210;
assign addr[9971] = 1489840425;
assign addr[9972] = 1503553506;
assign addr[9973] = 1517147363;
assign addr[9974] = 1530620920;
assign addr[9975] = 1543973108;
assign addr[9976] = 1557202869;
assign addr[9977] = 1570309153;
assign addr[9978] = 1583290921;
assign addr[9979] = 1596147143;
assign addr[9980] = 1608876801;
assign addr[9981] = 1621478885;
assign addr[9982] = 1633952396;
assign addr[9983] = 1646296344;
assign addr[9984] = 1658509750;
assign addr[9985] = 1670591647;
assign addr[9986] = 1682541077;
assign addr[9987] = 1694357091;
assign addr[9988] = 1706038753;
assign addr[9989] = 1717585136;
assign addr[9990] = 1728995326;
assign addr[9991] = 1740268417;
assign addr[9992] = 1751403515;
assign addr[9993] = 1762399737;
assign addr[9994] = 1773256212;
assign addr[9995] = 1783972079;
assign addr[9996] = 1794546487;
assign addr[9997] = 1804978599;
assign addr[9998] = 1815267588;
assign addr[9999] = 1825412636;
assign addr[10000] = 1835412941;
assign addr[10001] = 1845267708;
assign addr[10002] = 1854976157;
assign addr[10003] = 1864537518;
assign addr[10004] = 1873951032;
assign addr[10005] = 1883215953;
assign addr[10006] = 1892331547;
assign addr[10007] = 1901297091;
assign addr[10008] = 1910111873;
assign addr[10009] = 1918775195;
assign addr[10010] = 1927286370;
assign addr[10011] = 1935644723;
assign addr[10012] = 1943849591;
assign addr[10013] = 1951900324;
assign addr[10014] = 1959796283;
assign addr[10015] = 1967536842;
assign addr[10016] = 1975121388;
assign addr[10017] = 1982549318;
assign addr[10018] = 1989820044;
assign addr[10019] = 1996932990;
assign addr[10020] = 2003887591;
assign addr[10021] = 2010683297;
assign addr[10022] = 2017319567;
assign addr[10023] = 2023795876;
assign addr[10024] = 2030111710;
assign addr[10025] = 2036266570;
assign addr[10026] = 2042259965;
assign addr[10027] = 2048091422;
assign addr[10028] = 2053760478;
assign addr[10029] = 2059266683;
assign addr[10030] = 2064609600;
assign addr[10031] = 2069788807;
assign addr[10032] = 2074803892;
assign addr[10033] = 2079654458;
assign addr[10034] = 2084340120;
assign addr[10035] = 2088860507;
assign addr[10036] = 2093215260;
assign addr[10037] = 2097404033;
assign addr[10038] = 2101426496;
assign addr[10039] = 2105282327;
assign addr[10040] = 2108971223;
assign addr[10041] = 2112492891;
assign addr[10042] = 2115847050;
assign addr[10043] = 2119033436;
assign addr[10044] = 2122051796;
assign addr[10045] = 2124901890;
assign addr[10046] = 2127583492;
assign addr[10047] = 2130096389;
assign addr[10048] = 2132440383;
assign addr[10049] = 2134615288;
assign addr[10050] = 2136620930;
assign addr[10051] = 2138457152;
assign addr[10052] = 2140123807;
assign addr[10053] = 2141620763;
assign addr[10054] = 2142947902;
assign addr[10055] = 2144105118;
assign addr[10056] = 2145092320;
assign addr[10057] = 2145909429;
assign addr[10058] = 2146556380;
assign addr[10059] = 2147033123;
assign addr[10060] = 2147339619;
assign addr[10061] = 2147475844;
assign addr[10062] = 2147441787;
assign addr[10063] = 2147237452;
assign addr[10064] = 2146862854;
assign addr[10065] = 2146318022;
assign addr[10066] = 2145603001;
assign addr[10067] = 2144717846;
assign addr[10068] = 2143662628;
assign addr[10069] = 2142437431;
assign addr[10070] = 2141042352;
assign addr[10071] = 2139477502;
assign addr[10072] = 2137743003;
assign addr[10073] = 2135838995;
assign addr[10074] = 2133765628;
assign addr[10075] = 2131523066;
assign addr[10076] = 2129111488;
assign addr[10077] = 2126531084;
assign addr[10078] = 2123782059;
assign addr[10079] = 2120864631;
assign addr[10080] = 2117779031;
assign addr[10081] = 2114525505;
assign addr[10082] = 2111104309;
assign addr[10083] = 2107515716;
assign addr[10084] = 2103760010;
assign addr[10085] = 2099837489;
assign addr[10086] = 2095748463;
assign addr[10087] = 2091493257;
assign addr[10088] = 2087072209;
assign addr[10089] = 2082485668;
assign addr[10090] = 2077733999;
assign addr[10091] = 2072817579;
assign addr[10092] = 2067736796;
assign addr[10093] = 2062492055;
assign addr[10094] = 2057083771;
assign addr[10095] = 2051512372;
assign addr[10096] = 2045778302;
assign addr[10097] = 2039882013;
assign addr[10098] = 2033823974;
assign addr[10099] = 2027604666;
assign addr[10100] = 2021224581;
assign addr[10101] = 2014684225;
assign addr[10102] = 2007984117;
assign addr[10103] = 2001124788;
assign addr[10104] = 1994106782;
assign addr[10105] = 1986930656;
assign addr[10106] = 1979596978;
assign addr[10107] = 1972106330;
assign addr[10108] = 1964459306;
assign addr[10109] = 1956656513;
assign addr[10110] = 1948698568;
assign addr[10111] = 1940586104;
assign addr[10112] = 1932319763;
assign addr[10113] = 1923900201;
assign addr[10114] = 1915328086;
assign addr[10115] = 1906604097;
assign addr[10116] = 1897728925;
assign addr[10117] = 1888703276;
assign addr[10118] = 1879527863;
assign addr[10119] = 1870203416;
assign addr[10120] = 1860730673;
assign addr[10121] = 1851110385;
assign addr[10122] = 1841343316;
assign addr[10123] = 1831430239;
assign addr[10124] = 1821371941;
assign addr[10125] = 1811169220;
assign addr[10126] = 1800822883;
assign addr[10127] = 1790333753;
assign addr[10128] = 1779702660;
assign addr[10129] = 1768930447;
assign addr[10130] = 1758017969;
assign addr[10131] = 1746966091;
assign addr[10132] = 1735775690;
assign addr[10133] = 1724447652;
assign addr[10134] = 1712982875;
assign addr[10135] = 1701382270;
assign addr[10136] = 1689646755;
assign addr[10137] = 1677777262;
assign addr[10138] = 1665774731;
assign addr[10139] = 1653640115;
assign addr[10140] = 1641374375;
assign addr[10141] = 1628978484;
assign addr[10142] = 1616453425;
assign addr[10143] = 1603800191;
assign addr[10144] = 1591019785;
assign addr[10145] = 1578113222;
assign addr[10146] = 1565081523;
assign addr[10147] = 1551925723;
assign addr[10148] = 1538646865;
assign addr[10149] = 1525246002;
assign addr[10150] = 1511724196;
assign addr[10151] = 1498082520;
assign addr[10152] = 1484322054;
assign addr[10153] = 1470443891;
assign addr[10154] = 1456449131;
assign addr[10155] = 1442338884;
assign addr[10156] = 1428114267;
assign addr[10157] = 1413776410;
assign addr[10158] = 1399326449;
assign addr[10159] = 1384765530;
assign addr[10160] = 1370094808;
assign addr[10161] = 1355315445;
assign addr[10162] = 1340428615;
assign addr[10163] = 1325435496;
assign addr[10164] = 1310337279;
assign addr[10165] = 1295135159;
assign addr[10166] = 1279830344;
assign addr[10167] = 1264424045;
assign addr[10168] = 1248917486;
assign addr[10169] = 1233311895;
assign addr[10170] = 1217608510;
assign addr[10171] = 1201808576;
assign addr[10172] = 1185913346;
assign addr[10173] = 1169924081;
assign addr[10174] = 1153842047;
assign addr[10175] = 1137668521;
assign addr[10176] = 1121404785;
assign addr[10177] = 1105052128;
assign addr[10178] = 1088611847;
assign addr[10179] = 1072085246;
assign addr[10180] = 1055473635;
assign addr[10181] = 1038778332;
assign addr[10182] = 1022000660;
assign addr[10183] = 1005141949;
assign addr[10184] = 988203537;
assign addr[10185] = 971186766;
assign addr[10186] = 954092986;
assign addr[10187] = 936923553;
assign addr[10188] = 919679827;
assign addr[10189] = 902363176;
assign addr[10190] = 884974973;
assign addr[10191] = 867516597;
assign addr[10192] = 849989433;
assign addr[10193] = 832394869;
assign addr[10194] = 814734301;
assign addr[10195] = 797009130;
assign addr[10196] = 779220762;
assign addr[10197] = 761370605;
assign addr[10198] = 743460077;
assign addr[10199] = 725490597;
assign addr[10200] = 707463589;
assign addr[10201] = 689380485;
assign addr[10202] = 671242716;
assign addr[10203] = 653051723;
assign addr[10204] = 634808946;
assign addr[10205] = 616515832;
assign addr[10206] = 598173833;
assign addr[10207] = 579784402;
assign addr[10208] = 561348998;
assign addr[10209] = 542869083;
assign addr[10210] = 524346121;
assign addr[10211] = 505781581;
assign addr[10212] = 487176937;
assign addr[10213] = 468533662;
assign addr[10214] = 449853235;
assign addr[10215] = 431137138;
assign addr[10216] = 412386854;
assign addr[10217] = 393603870;
assign addr[10218] = 374789676;
assign addr[10219] = 355945764;
assign addr[10220] = 337073627;
assign addr[10221] = 318174762;
assign addr[10222] = 299250668;
assign addr[10223] = 280302845;
assign addr[10224] = 261332796;
assign addr[10225] = 242342025;
assign addr[10226] = 223332037;
assign addr[10227] = 204304341;
assign addr[10228] = 185260444;
assign addr[10229] = 166201858;
assign addr[10230] = 147130093;
assign addr[10231] = 128046661;
assign addr[10232] = 108953076;
assign addr[10233] = 89850852;
assign addr[10234] = 70741503;
assign addr[10235] = 51626544;
assign addr[10236] = 32507492;
assign addr[10237] = 13385863;
assign addr[10238] = -5736829;
assign addr[10239] = -24859065;
assign addr[10240] = -43979330;
assign addr[10241] = -63096108;
assign addr[10242] = -82207882;
assign addr[10243] = -101313138;
assign addr[10244] = -120410361;
assign addr[10245] = -139498035;
assign addr[10246] = -158574649;
assign addr[10247] = -177638688;
assign addr[10248] = -196688642;
assign addr[10249] = -215722999;
assign addr[10250] = -234740251;
assign addr[10251] = -253738890;
assign addr[10252] = -272717408;
assign addr[10253] = -291674302;
assign addr[10254] = -310608068;
assign addr[10255] = -329517204;
assign addr[10256] = -348400212;
assign addr[10257] = -367255594;
assign addr[10258] = -386081854;
assign addr[10259] = -404877501;
assign addr[10260] = -423641043;
assign addr[10261] = -442370993;
assign addr[10262] = -461065866;
assign addr[10263] = -479724180;
assign addr[10264] = -498344454;
assign addr[10265] = -516925212;
assign addr[10266] = -535464981;
assign addr[10267] = -553962291;
assign addr[10268] = -572415676;
assign addr[10269] = -590823671;
assign addr[10270] = -609184818;
assign addr[10271] = -627497660;
assign addr[10272] = -645760745;
assign addr[10273] = -663972625;
assign addr[10274] = -682131857;
assign addr[10275] = -700236999;
assign addr[10276] = -718286617;
assign addr[10277] = -736279279;
assign addr[10278] = -754213559;
assign addr[10279] = -772088034;
assign addr[10280] = -789901288;
assign addr[10281] = -807651907;
assign addr[10282] = -825338484;
assign addr[10283] = -842959617;
assign addr[10284] = -860513908;
assign addr[10285] = -877999966;
assign addr[10286] = -895416404;
assign addr[10287] = -912761841;
assign addr[10288] = -930034901;
assign addr[10289] = -947234215;
assign addr[10290] = -964358420;
assign addr[10291] = -981406156;
assign addr[10292] = -998376073;
assign addr[10293] = -1015266825;
assign addr[10294] = -1032077073;
assign addr[10295] = -1048805483;
assign addr[10296] = -1065450729;
assign addr[10297] = -1082011492;
assign addr[10298] = -1098486458;
assign addr[10299] = -1114874320;
assign addr[10300] = -1131173780;
assign addr[10301] = -1147383544;
assign addr[10302] = -1163502328;
assign addr[10303] = -1179528853;
assign addr[10304] = -1195461849;
assign addr[10305] = -1211300053;
assign addr[10306] = -1227042207;
assign addr[10307] = -1242687064;
assign addr[10308] = -1258233384;
assign addr[10309] = -1273679934;
assign addr[10310] = -1289025489;
assign addr[10311] = -1304268832;
assign addr[10312] = -1319408754;
assign addr[10313] = -1334444055;
assign addr[10314] = -1349373543;
assign addr[10315] = -1364196034;
assign addr[10316] = -1378910353;
assign addr[10317] = -1393515332;
assign addr[10318] = -1408009814;
assign addr[10319] = -1422392650;
assign addr[10320] = -1436662698;
assign addr[10321] = -1450818828;
assign addr[10322] = -1464859917;
assign addr[10323] = -1478784851;
assign addr[10324] = -1492592527;
assign addr[10325] = -1506281850;
assign addr[10326] = -1519851733;
assign addr[10327] = -1533301101;
assign addr[10328] = -1546628888;
assign addr[10329] = -1559834037;
assign addr[10330] = -1572915501;
assign addr[10331] = -1585872242;
assign addr[10332] = -1598703233;
assign addr[10333] = -1611407456;
assign addr[10334] = -1623983905;
assign addr[10335] = -1636431582;
assign addr[10336] = -1648749499;
assign addr[10337] = -1660936681;
assign addr[10338] = -1672992161;
assign addr[10339] = -1684914983;
assign addr[10340] = -1696704201;
assign addr[10341] = -1708358881;
assign addr[10342] = -1719878099;
assign addr[10343] = -1731260941;
assign addr[10344] = -1742506504;
assign addr[10345] = -1753613897;
assign addr[10346] = -1764582240;
assign addr[10347] = -1775410662;
assign addr[10348] = -1786098304;
assign addr[10349] = -1796644320;
assign addr[10350] = -1807047873;
assign addr[10351] = -1817308138;
assign addr[10352] = -1827424302;
assign addr[10353] = -1837395562;
assign addr[10354] = -1847221128;
assign addr[10355] = -1856900221;
assign addr[10356] = -1866432072;
assign addr[10357] = -1875815927;
assign addr[10358] = -1885051042;
assign addr[10359] = -1894136683;
assign addr[10360] = -1903072131;
assign addr[10361] = -1911856677;
assign addr[10362] = -1920489624;
assign addr[10363] = -1928970288;
assign addr[10364] = -1937297997;
assign addr[10365] = -1945472089;
assign addr[10366] = -1953491918;
assign addr[10367] = -1961356847;
assign addr[10368] = -1969066252;
assign addr[10369] = -1976619522;
assign addr[10370] = -1984016058;
assign addr[10371] = -1991255274;
assign addr[10372] = -1998336596;
assign addr[10373] = -2005259462;
assign addr[10374] = -2012023322;
assign addr[10375] = -2018627642;
assign addr[10376] = -2025071897;
assign addr[10377] = -2031355576;
assign addr[10378] = -2037478181;
assign addr[10379] = -2043439226;
assign addr[10380] = -2049238240;
assign addr[10381] = -2054874761;
assign addr[10382] = -2060348343;
assign addr[10383] = -2065658552;
assign addr[10384] = -2070804967;
assign addr[10385] = -2075787180;
assign addr[10386] = -2080604795;
assign addr[10387] = -2085257431;
assign addr[10388] = -2089744719;
assign addr[10389] = -2094066304;
assign addr[10390] = -2098221841;
assign addr[10391] = -2102211002;
assign addr[10392] = -2106033471;
assign addr[10393] = -2109688944;
assign addr[10394] = -2113177132;
assign addr[10395] = -2116497758;
assign addr[10396] = -2119650558;
assign addr[10397] = -2122635283;
assign addr[10398] = -2125451696;
assign addr[10399] = -2128099574;
assign addr[10400] = -2130578706;
assign addr[10401] = -2132888897;
assign addr[10402] = -2135029962;
assign addr[10403] = -2137001733;
assign addr[10404] = -2138804053;
assign addr[10405] = -2140436778;
assign addr[10406] = -2141899780;
assign addr[10407] = -2143192942;
assign addr[10408] = -2144316162;
assign addr[10409] = -2145269351;
assign addr[10410] = -2146052433;
assign addr[10411] = -2146665347;
assign addr[10412] = -2147108043;
assign addr[10413] = -2147380486;
assign addr[10414] = -2147482655;
assign addr[10415] = -2147414542;
assign addr[10416] = -2147176152;
assign addr[10417] = -2146767505;
assign addr[10418] = -2146188631;
assign addr[10419] = -2145439578;
assign addr[10420] = -2144520405;
assign addr[10421] = -2143431184;
assign addr[10422] = -2142172003;
assign addr[10423] = -2140742960;
assign addr[10424] = -2139144169;
assign addr[10425] = -2137375758;
assign addr[10426] = -2135437865;
assign addr[10427] = -2133330646;
assign addr[10428] = -2131054266;
assign addr[10429] = -2128608907;
assign addr[10430] = -2125994762;
assign addr[10431] = -2123212038;
assign addr[10432] = -2120260957;
assign addr[10433] = -2117141752;
assign addr[10434] = -2113854671;
assign addr[10435] = -2110399974;
assign addr[10436] = -2106777935;
assign addr[10437] = -2102988841;
assign addr[10438] = -2099032994;
assign addr[10439] = -2094910706;
assign addr[10440] = -2090622304;
assign addr[10441] = -2086168128;
assign addr[10442] = -2081548533;
assign addr[10443] = -2076763883;
assign addr[10444] = -2071814558;
assign addr[10445] = -2066700952;
assign addr[10446] = -2061423468;
assign addr[10447] = -2055982526;
assign addr[10448] = -2050378558;
assign addr[10449] = -2044612007;
assign addr[10450] = -2038683330;
assign addr[10451] = -2032592999;
assign addr[10452] = -2026341495;
assign addr[10453] = -2019929315;
assign addr[10454] = -2013356967;
assign addr[10455] = -2006624971;
assign addr[10456] = -1999733863;
assign addr[10457] = -1992684188;
assign addr[10458] = -1985476506;
assign addr[10459] = -1978111387;
assign addr[10460] = -1970589416;
assign addr[10461] = -1962911189;
assign addr[10462] = -1955077316;
assign addr[10463] = -1947088417;
assign addr[10464] = -1938945125;
assign addr[10465] = -1930648088;
assign addr[10466] = -1922197961;
assign addr[10467] = -1913595416;
assign addr[10468] = -1904841135;
assign addr[10469] = -1895935811;
assign addr[10470] = -1886880151;
assign addr[10471] = -1877674873;
assign addr[10472] = -1868320707;
assign addr[10473] = -1858818395;
assign addr[10474] = -1849168689;
assign addr[10475] = -1839372356;
assign addr[10476] = -1829430172;
assign addr[10477] = -1819342925;
assign addr[10478] = -1809111415;
assign addr[10479] = -1798736454;
assign addr[10480] = -1788218865;
assign addr[10481] = -1777559480;
assign addr[10482] = -1766759146;
assign addr[10483] = -1755818718;
assign addr[10484] = -1744739065;
assign addr[10485] = -1733521064;
assign addr[10486] = -1722165606;
assign addr[10487] = -1710673591;
assign addr[10488] = -1699045930;
assign addr[10489] = -1687283545;
assign addr[10490] = -1675387369;
assign addr[10491] = -1663358344;
assign addr[10492] = -1651197426;
assign addr[10493] = -1638905577;
assign addr[10494] = -1626483774;
assign addr[10495] = -1613933000;
assign addr[10496] = -1601254251;
assign addr[10497] = -1588448533;
assign addr[10498] = -1575516860;
assign addr[10499] = -1562460258;
assign addr[10500] = -1549279763;
assign addr[10501] = -1535976419;
assign addr[10502] = -1522551282;
assign addr[10503] = -1509005416;
assign addr[10504] = -1495339895;
assign addr[10505] = -1481555802;
assign addr[10506] = -1467654232;
assign addr[10507] = -1453636285;
assign addr[10508] = -1439503074;
assign addr[10509] = -1425255719;
assign addr[10510] = -1410895350;
assign addr[10511] = -1396423105;
assign addr[10512] = -1381840133;
assign addr[10513] = -1367147589;
assign addr[10514] = -1352346639;
assign addr[10515] = -1337438456;
assign addr[10516] = -1322424222;
assign addr[10517] = -1307305128;
assign addr[10518] = -1292082373;
assign addr[10519] = -1276757164;
assign addr[10520] = -1261330715;
assign addr[10521] = -1245804251;
assign addr[10522] = -1230179002;
assign addr[10523] = -1214456207;
assign addr[10524] = -1198637114;
assign addr[10525] = -1182722976;
assign addr[10526] = -1166715055;
assign addr[10527] = -1150614620;
assign addr[10528] = -1134422949;
assign addr[10529] = -1118141326;
assign addr[10530] = -1101771040;
assign addr[10531] = -1085313391;
assign addr[10532] = -1068769683;
assign addr[10533] = -1052141228;
assign addr[10534] = -1035429345;
assign addr[10535] = -1018635358;
assign addr[10536] = -1001760600;
assign addr[10537] = -984806408;
assign addr[10538] = -967774128;
assign addr[10539] = -950665109;
assign addr[10540] = -933480707;
assign addr[10541] = -916222287;
assign addr[10542] = -898891215;
assign addr[10543] = -881488868;
assign addr[10544] = -864016623;
assign addr[10545] = -846475867;
assign addr[10546] = -828867991;
assign addr[10547] = -811194391;
assign addr[10548] = -793456467;
assign addr[10549] = -775655628;
assign addr[10550] = -757793284;
assign addr[10551] = -739870851;
assign addr[10552] = -721889752;
assign addr[10553] = -703851410;
assign addr[10554] = -685757258;
assign addr[10555] = -667608730;
assign addr[10556] = -649407264;
assign addr[10557] = -631154304;
assign addr[10558] = -612851297;
assign addr[10559] = -594499695;
assign addr[10560] = -576100953;
assign addr[10561] = -557656529;
assign addr[10562] = -539167887;
assign addr[10563] = -520636492;
assign addr[10564] = -502063814;
assign addr[10565] = -483451325;
assign addr[10566] = -464800501;
assign addr[10567] = -446112822;
assign addr[10568] = -427389768;
assign addr[10569] = -408632825;
assign addr[10570] = -389843480;
assign addr[10571] = -371023223;
assign addr[10572] = -352173546;
assign addr[10573] = -333295944;
assign addr[10574] = -314391913;
assign addr[10575] = -295462954;
assign addr[10576] = -276510565;
assign addr[10577] = -257536251;
assign addr[10578] = -238541516;
assign addr[10579] = -219527866;
assign addr[10580] = -200496809;
assign addr[10581] = -181449854;
assign addr[10582] = -162388511;
assign addr[10583] = -143314291;
assign addr[10584] = -124228708;
assign addr[10585] = -105133274;
assign addr[10586] = -86029503;
assign addr[10587] = -66918911;
assign addr[10588] = -47803013;
assign addr[10589] = -28683324;
assign addr[10590] = -9561361;
assign addr[10591] = 9561361;
assign addr[10592] = 28683324;
assign addr[10593] = 47803013;
assign addr[10594] = 66918911;
assign addr[10595] = 86029503;
assign addr[10596] = 105133274;
assign addr[10597] = 124228708;
assign addr[10598] = 143314291;
assign addr[10599] = 162388511;
assign addr[10600] = 181449854;
assign addr[10601] = 200496809;
assign addr[10602] = 219527866;
assign addr[10603] = 238541516;
assign addr[10604] = 257536251;
assign addr[10605] = 276510565;
assign addr[10606] = 295462954;
assign addr[10607] = 314391913;
assign addr[10608] = 333295944;
assign addr[10609] = 352173546;
assign addr[10610] = 371023223;
assign addr[10611] = 389843480;
assign addr[10612] = 408632825;
assign addr[10613] = 427389768;
assign addr[10614] = 446112822;
assign addr[10615] = 464800501;
assign addr[10616] = 483451325;
assign addr[10617] = 502063814;
assign addr[10618] = 520636492;
assign addr[10619] = 539167887;
assign addr[10620] = 557656529;
assign addr[10621] = 576100953;
assign addr[10622] = 594499695;
assign addr[10623] = 612851297;
assign addr[10624] = 631154304;
assign addr[10625] = 649407264;
assign addr[10626] = 667608730;
assign addr[10627] = 685757258;
assign addr[10628] = 703851410;
assign addr[10629] = 721889752;
assign addr[10630] = 739870851;
assign addr[10631] = 757793284;
assign addr[10632] = 775655628;
assign addr[10633] = 793456467;
assign addr[10634] = 811194391;
assign addr[10635] = 828867991;
assign addr[10636] = 846475867;
assign addr[10637] = 864016623;
assign addr[10638] = 881488868;
assign addr[10639] = 898891215;
assign addr[10640] = 916222287;
assign addr[10641] = 933480707;
assign addr[10642] = 950665109;
assign addr[10643] = 967774128;
assign addr[10644] = 984806408;
assign addr[10645] = 1001760600;
assign addr[10646] = 1018635358;
assign addr[10647] = 1035429345;
assign addr[10648] = 1052141228;
assign addr[10649] = 1068769683;
assign addr[10650] = 1085313391;
assign addr[10651] = 1101771040;
assign addr[10652] = 1118141326;
assign addr[10653] = 1134422949;
assign addr[10654] = 1150614620;
assign addr[10655] = 1166715055;
assign addr[10656] = 1182722976;
assign addr[10657] = 1198637114;
assign addr[10658] = 1214456207;
assign addr[10659] = 1230179002;
assign addr[10660] = 1245804251;
assign addr[10661] = 1261330715;
assign addr[10662] = 1276757164;
assign addr[10663] = 1292082373;
assign addr[10664] = 1307305128;
assign addr[10665] = 1322424222;
assign addr[10666] = 1337438456;
assign addr[10667] = 1352346639;
assign addr[10668] = 1367147589;
assign addr[10669] = 1381840133;
assign addr[10670] = 1396423105;
assign addr[10671] = 1410895350;
assign addr[10672] = 1425255719;
assign addr[10673] = 1439503074;
assign addr[10674] = 1453636285;
assign addr[10675] = 1467654232;
assign addr[10676] = 1481555802;
assign addr[10677] = 1495339895;
assign addr[10678] = 1509005416;
assign addr[10679] = 1522551282;
assign addr[10680] = 1535976419;
assign addr[10681] = 1549279763;
assign addr[10682] = 1562460258;
assign addr[10683] = 1575516860;
assign addr[10684] = 1588448533;
assign addr[10685] = 1601254251;
assign addr[10686] = 1613933000;
assign addr[10687] = 1626483774;
assign addr[10688] = 1638905577;
assign addr[10689] = 1651197426;
assign addr[10690] = 1663358344;
assign addr[10691] = 1675387369;
assign addr[10692] = 1687283545;
assign addr[10693] = 1699045930;
assign addr[10694] = 1710673591;
assign addr[10695] = 1722165606;
assign addr[10696] = 1733521064;
assign addr[10697] = 1744739065;
assign addr[10698] = 1755818718;
assign addr[10699] = 1766759146;
assign addr[10700] = 1777559480;
assign addr[10701] = 1788218865;
assign addr[10702] = 1798736454;
assign addr[10703] = 1809111415;
assign addr[10704] = 1819342925;
assign addr[10705] = 1829430172;
assign addr[10706] = 1839372356;
assign addr[10707] = 1849168689;
assign addr[10708] = 1858818395;
assign addr[10709] = 1868320707;
assign addr[10710] = 1877674873;
assign addr[10711] = 1886880151;
assign addr[10712] = 1895935811;
assign addr[10713] = 1904841135;
assign addr[10714] = 1913595416;
assign addr[10715] = 1922197961;
assign addr[10716] = 1930648088;
assign addr[10717] = 1938945125;
assign addr[10718] = 1947088417;
assign addr[10719] = 1955077316;
assign addr[10720] = 1962911189;
assign addr[10721] = 1970589416;
assign addr[10722] = 1978111387;
assign addr[10723] = 1985476506;
assign addr[10724] = 1992684188;
assign addr[10725] = 1999733863;
assign addr[10726] = 2006624971;
assign addr[10727] = 2013356967;
assign addr[10728] = 2019929315;
assign addr[10729] = 2026341495;
assign addr[10730] = 2032592999;
assign addr[10731] = 2038683330;
assign addr[10732] = 2044612007;
assign addr[10733] = 2050378558;
assign addr[10734] = 2055982526;
assign addr[10735] = 2061423468;
assign addr[10736] = 2066700952;
assign addr[10737] = 2071814558;
assign addr[10738] = 2076763883;
assign addr[10739] = 2081548533;
assign addr[10740] = 2086168128;
assign addr[10741] = 2090622304;
assign addr[10742] = 2094910706;
assign addr[10743] = 2099032994;
assign addr[10744] = 2102988841;
assign addr[10745] = 2106777935;
assign addr[10746] = 2110399974;
assign addr[10747] = 2113854671;
assign addr[10748] = 2117141752;
assign addr[10749] = 2120260957;
assign addr[10750] = 2123212038;
assign addr[10751] = 2125994762;
assign addr[10752] = 2128608907;
assign addr[10753] = 2131054266;
assign addr[10754] = 2133330646;
assign addr[10755] = 2135437865;
assign addr[10756] = 2137375758;
assign addr[10757] = 2139144169;
assign addr[10758] = 2140742960;
assign addr[10759] = 2142172003;
assign addr[10760] = 2143431184;
assign addr[10761] = 2144520405;
assign addr[10762] = 2145439578;
assign addr[10763] = 2146188631;
assign addr[10764] = 2146767505;
assign addr[10765] = 2147176152;
assign addr[10766] = 2147414542;
assign addr[10767] = 2147482655;
assign addr[10768] = 2147380486;
assign addr[10769] = 2147108043;
assign addr[10770] = 2146665347;
assign addr[10771] = 2146052433;
assign addr[10772] = 2145269351;
assign addr[10773] = 2144316162;
assign addr[10774] = 2143192942;
assign addr[10775] = 2141899780;
assign addr[10776] = 2140436778;
assign addr[10777] = 2138804053;
assign addr[10778] = 2137001733;
assign addr[10779] = 2135029962;
assign addr[10780] = 2132888897;
assign addr[10781] = 2130578706;
assign addr[10782] = 2128099574;
assign addr[10783] = 2125451696;
assign addr[10784] = 2122635283;
assign addr[10785] = 2119650558;
assign addr[10786] = 2116497758;
assign addr[10787] = 2113177132;
assign addr[10788] = 2109688944;
assign addr[10789] = 2106033471;
assign addr[10790] = 2102211002;
assign addr[10791] = 2098221841;
assign addr[10792] = 2094066304;
assign addr[10793] = 2089744719;
assign addr[10794] = 2085257431;
assign addr[10795] = 2080604795;
assign addr[10796] = 2075787180;
assign addr[10797] = 2070804967;
assign addr[10798] = 2065658552;
assign addr[10799] = 2060348343;
assign addr[10800] = 2054874761;
assign addr[10801] = 2049238240;
assign addr[10802] = 2043439226;
assign addr[10803] = 2037478181;
assign addr[10804] = 2031355576;
assign addr[10805] = 2025071897;
assign addr[10806] = 2018627642;
assign addr[10807] = 2012023322;
assign addr[10808] = 2005259462;
assign addr[10809] = 1998336596;
assign addr[10810] = 1991255274;
assign addr[10811] = 1984016058;
assign addr[10812] = 1976619522;
assign addr[10813] = 1969066252;
assign addr[10814] = 1961356847;
assign addr[10815] = 1953491918;
assign addr[10816] = 1945472089;
assign addr[10817] = 1937297997;
assign addr[10818] = 1928970288;
assign addr[10819] = 1920489624;
assign addr[10820] = 1911856677;
assign addr[10821] = 1903072131;
assign addr[10822] = 1894136683;
assign addr[10823] = 1885051042;
assign addr[10824] = 1875815927;
assign addr[10825] = 1866432072;
assign addr[10826] = 1856900221;
assign addr[10827] = 1847221128;
assign addr[10828] = 1837395562;
assign addr[10829] = 1827424302;
assign addr[10830] = 1817308138;
assign addr[10831] = 1807047873;
assign addr[10832] = 1796644320;
assign addr[10833] = 1786098304;
assign addr[10834] = 1775410662;
assign addr[10835] = 1764582240;
assign addr[10836] = 1753613897;
assign addr[10837] = 1742506504;
assign addr[10838] = 1731260941;
assign addr[10839] = 1719878099;
assign addr[10840] = 1708358881;
assign addr[10841] = 1696704201;
assign addr[10842] = 1684914983;
assign addr[10843] = 1672992161;
assign addr[10844] = 1660936681;
assign addr[10845] = 1648749499;
assign addr[10846] = 1636431582;
assign addr[10847] = 1623983905;
assign addr[10848] = 1611407456;
assign addr[10849] = 1598703233;
assign addr[10850] = 1585872242;
assign addr[10851] = 1572915501;
assign addr[10852] = 1559834037;
assign addr[10853] = 1546628888;
assign addr[10854] = 1533301101;
assign addr[10855] = 1519851733;
assign addr[10856] = 1506281850;
assign addr[10857] = 1492592527;
assign addr[10858] = 1478784851;
assign addr[10859] = 1464859917;
assign addr[10860] = 1450818828;
assign addr[10861] = 1436662698;
assign addr[10862] = 1422392650;
assign addr[10863] = 1408009814;
assign addr[10864] = 1393515332;
assign addr[10865] = 1378910353;
assign addr[10866] = 1364196034;
assign addr[10867] = 1349373543;
assign addr[10868] = 1334444055;
assign addr[10869] = 1319408754;
assign addr[10870] = 1304268832;
assign addr[10871] = 1289025489;
assign addr[10872] = 1273679934;
assign addr[10873] = 1258233384;
assign addr[10874] = 1242687064;
assign addr[10875] = 1227042207;
assign addr[10876] = 1211300053;
assign addr[10877] = 1195461849;
assign addr[10878] = 1179528853;
assign addr[10879] = 1163502328;
assign addr[10880] = 1147383544;
assign addr[10881] = 1131173780;
assign addr[10882] = 1114874320;
assign addr[10883] = 1098486458;
assign addr[10884] = 1082011492;
assign addr[10885] = 1065450729;
assign addr[10886] = 1048805483;
assign addr[10887] = 1032077073;
assign addr[10888] = 1015266825;
assign addr[10889] = 998376073;
assign addr[10890] = 981406156;
assign addr[10891] = 964358420;
assign addr[10892] = 947234215;
assign addr[10893] = 930034901;
assign addr[10894] = 912761841;
assign addr[10895] = 895416404;
assign addr[10896] = 877999966;
assign addr[10897] = 860513908;
assign addr[10898] = 842959617;
assign addr[10899] = 825338484;
assign addr[10900] = 807651907;
assign addr[10901] = 789901288;
assign addr[10902] = 772088034;
assign addr[10903] = 754213559;
assign addr[10904] = 736279279;
assign addr[10905] = 718286617;
assign addr[10906] = 700236999;
assign addr[10907] = 682131857;
assign addr[10908] = 663972625;
assign addr[10909] = 645760745;
assign addr[10910] = 627497660;
assign addr[10911] = 609184818;
assign addr[10912] = 590823671;
assign addr[10913] = 572415676;
assign addr[10914] = 553962291;
assign addr[10915] = 535464981;
assign addr[10916] = 516925212;
assign addr[10917] = 498344454;
assign addr[10918] = 479724180;
assign addr[10919] = 461065866;
assign addr[10920] = 442370993;
assign addr[10921] = 423641043;
assign addr[10922] = 404877501;
assign addr[10923] = 386081854;
assign addr[10924] = 367255594;
assign addr[10925] = 348400212;
assign addr[10926] = 329517204;
assign addr[10927] = 310608068;
assign addr[10928] = 291674302;
assign addr[10929] = 272717408;
assign addr[10930] = 253738890;
assign addr[10931] = 234740251;
assign addr[10932] = 215722999;
assign addr[10933] = 196688642;
assign addr[10934] = 177638688;
assign addr[10935] = 158574649;
assign addr[10936] = 139498035;
assign addr[10937] = 120410361;
assign addr[10938] = 101313138;
assign addr[10939] = 82207882;
assign addr[10940] = 63096108;
assign addr[10941] = 43979330;
assign addr[10942] = 24859065;
assign addr[10943] = 5736829;
assign addr[10944] = -13385863;
assign addr[10945] = -32507492;
assign addr[10946] = -51626544;
assign addr[10947] = -70741503;
assign addr[10948] = -89850852;
assign addr[10949] = -108953076;
assign addr[10950] = -128046661;
assign addr[10951] = -147130093;
assign addr[10952] = -166201858;
assign addr[10953] = -185260444;
assign addr[10954] = -204304341;
assign addr[10955] = -223332037;
assign addr[10956] = -242342025;
assign addr[10957] = -261332796;
assign addr[10958] = -280302845;
assign addr[10959] = -299250668;
assign addr[10960] = -318174762;
assign addr[10961] = -337073627;
assign addr[10962] = -355945764;
assign addr[10963] = -374789676;
assign addr[10964] = -393603870;
assign addr[10965] = -412386854;
assign addr[10966] = -431137138;
assign addr[10967] = -449853235;
assign addr[10968] = -468533662;
assign addr[10969] = -487176937;
assign addr[10970] = -505781581;
assign addr[10971] = -524346121;
assign addr[10972] = -542869083;
assign addr[10973] = -561348998;
assign addr[10974] = -579784402;
assign addr[10975] = -598173833;
assign addr[10976] = -616515832;
assign addr[10977] = -634808946;
assign addr[10978] = -653051723;
assign addr[10979] = -671242716;
assign addr[10980] = -689380485;
assign addr[10981] = -707463589;
assign addr[10982] = -725490597;
assign addr[10983] = -743460077;
assign addr[10984] = -761370605;
assign addr[10985] = -779220762;
assign addr[10986] = -797009130;
assign addr[10987] = -814734301;
assign addr[10988] = -832394869;
assign addr[10989] = -849989433;
assign addr[10990] = -867516597;
assign addr[10991] = -884974973;
assign addr[10992] = -902363176;
assign addr[10993] = -919679827;
assign addr[10994] = -936923553;
assign addr[10995] = -954092986;
assign addr[10996] = -971186766;
assign addr[10997] = -988203537;
assign addr[10998] = -1005141949;
assign addr[10999] = -1022000660;
assign addr[11000] = -1038778332;
assign addr[11001] = -1055473635;
assign addr[11002] = -1072085246;
assign addr[11003] = -1088611847;
assign addr[11004] = -1105052128;
assign addr[11005] = -1121404785;
assign addr[11006] = -1137668521;
assign addr[11007] = -1153842047;
assign addr[11008] = -1169924081;
assign addr[11009] = -1185913346;
assign addr[11010] = -1201808576;
assign addr[11011] = -1217608510;
assign addr[11012] = -1233311895;
assign addr[11013] = -1248917486;
assign addr[11014] = -1264424045;
assign addr[11015] = -1279830344;
assign addr[11016] = -1295135159;
assign addr[11017] = -1310337279;
assign addr[11018] = -1325435496;
assign addr[11019] = -1340428615;
assign addr[11020] = -1355315445;
assign addr[11021] = -1370094808;
assign addr[11022] = -1384765530;
assign addr[11023] = -1399326449;
assign addr[11024] = -1413776410;
assign addr[11025] = -1428114267;
assign addr[11026] = -1442338884;
assign addr[11027] = -1456449131;
assign addr[11028] = -1470443891;
assign addr[11029] = -1484322054;
assign addr[11030] = -1498082520;
assign addr[11031] = -1511724196;
assign addr[11032] = -1525246002;
assign addr[11033] = -1538646865;
assign addr[11034] = -1551925723;
assign addr[11035] = -1565081523;
assign addr[11036] = -1578113222;
assign addr[11037] = -1591019785;
assign addr[11038] = -1603800191;
assign addr[11039] = -1616453425;
assign addr[11040] = -1628978484;
assign addr[11041] = -1641374375;
assign addr[11042] = -1653640115;
assign addr[11043] = -1665774731;
assign addr[11044] = -1677777262;
assign addr[11045] = -1689646755;
assign addr[11046] = -1701382270;
assign addr[11047] = -1712982875;
assign addr[11048] = -1724447652;
assign addr[11049] = -1735775690;
assign addr[11050] = -1746966091;
assign addr[11051] = -1758017969;
assign addr[11052] = -1768930447;
assign addr[11053] = -1779702660;
assign addr[11054] = -1790333753;
assign addr[11055] = -1800822883;
assign addr[11056] = -1811169220;
assign addr[11057] = -1821371941;
assign addr[11058] = -1831430239;
assign addr[11059] = -1841343316;
assign addr[11060] = -1851110385;
assign addr[11061] = -1860730673;
assign addr[11062] = -1870203416;
assign addr[11063] = -1879527863;
assign addr[11064] = -1888703276;
assign addr[11065] = -1897728925;
assign addr[11066] = -1906604097;
assign addr[11067] = -1915328086;
assign addr[11068] = -1923900201;
assign addr[11069] = -1932319763;
assign addr[11070] = -1940586104;
assign addr[11071] = -1948698568;
assign addr[11072] = -1956656513;
assign addr[11073] = -1964459306;
assign addr[11074] = -1972106330;
assign addr[11075] = -1979596978;
assign addr[11076] = -1986930656;
assign addr[11077] = -1994106782;
assign addr[11078] = -2001124788;
assign addr[11079] = -2007984117;
assign addr[11080] = -2014684225;
assign addr[11081] = -2021224581;
assign addr[11082] = -2027604666;
assign addr[11083] = -2033823974;
assign addr[11084] = -2039882013;
assign addr[11085] = -2045778302;
assign addr[11086] = -2051512372;
assign addr[11087] = -2057083771;
assign addr[11088] = -2062492055;
assign addr[11089] = -2067736796;
assign addr[11090] = -2072817579;
assign addr[11091] = -2077733999;
assign addr[11092] = -2082485668;
assign addr[11093] = -2087072209;
assign addr[11094] = -2091493257;
assign addr[11095] = -2095748463;
assign addr[11096] = -2099837489;
assign addr[11097] = -2103760010;
assign addr[11098] = -2107515716;
assign addr[11099] = -2111104309;
assign addr[11100] = -2114525505;
assign addr[11101] = -2117779031;
assign addr[11102] = -2120864631;
assign addr[11103] = -2123782059;
assign addr[11104] = -2126531084;
assign addr[11105] = -2129111488;
assign addr[11106] = -2131523066;
assign addr[11107] = -2133765628;
assign addr[11108] = -2135838995;
assign addr[11109] = -2137743003;
assign addr[11110] = -2139477502;
assign addr[11111] = -2141042352;
assign addr[11112] = -2142437431;
assign addr[11113] = -2143662628;
assign addr[11114] = -2144717846;
assign addr[11115] = -2145603001;
assign addr[11116] = -2146318022;
assign addr[11117] = -2146862854;
assign addr[11118] = -2147237452;
assign addr[11119] = -2147441787;
assign addr[11120] = -2147475844;
assign addr[11121] = -2147339619;
assign addr[11122] = -2147033123;
assign addr[11123] = -2146556380;
assign addr[11124] = -2145909429;
assign addr[11125] = -2145092320;
assign addr[11126] = -2144105118;
assign addr[11127] = -2142947902;
assign addr[11128] = -2141620763;
assign addr[11129] = -2140123807;
assign addr[11130] = -2138457152;
assign addr[11131] = -2136620930;
assign addr[11132] = -2134615288;
assign addr[11133] = -2132440383;
assign addr[11134] = -2130096389;
assign addr[11135] = -2127583492;
assign addr[11136] = -2124901890;
assign addr[11137] = -2122051796;
assign addr[11138] = -2119033436;
assign addr[11139] = -2115847050;
assign addr[11140] = -2112492891;
assign addr[11141] = -2108971223;
assign addr[11142] = -2105282327;
assign addr[11143] = -2101426496;
assign addr[11144] = -2097404033;
assign addr[11145] = -2093215260;
assign addr[11146] = -2088860507;
assign addr[11147] = -2084340120;
assign addr[11148] = -2079654458;
assign addr[11149] = -2074803892;
assign addr[11150] = -2069788807;
assign addr[11151] = -2064609600;
assign addr[11152] = -2059266683;
assign addr[11153] = -2053760478;
assign addr[11154] = -2048091422;
assign addr[11155] = -2042259965;
assign addr[11156] = -2036266570;
assign addr[11157] = -2030111710;
assign addr[11158] = -2023795876;
assign addr[11159] = -2017319567;
assign addr[11160] = -2010683297;
assign addr[11161] = -2003887591;
assign addr[11162] = -1996932990;
assign addr[11163] = -1989820044;
assign addr[11164] = -1982549318;
assign addr[11165] = -1975121388;
assign addr[11166] = -1967536842;
assign addr[11167] = -1959796283;
assign addr[11168] = -1951900324;
assign addr[11169] = -1943849591;
assign addr[11170] = -1935644723;
assign addr[11171] = -1927286370;
assign addr[11172] = -1918775195;
assign addr[11173] = -1910111873;
assign addr[11174] = -1901297091;
assign addr[11175] = -1892331547;
assign addr[11176] = -1883215953;
assign addr[11177] = -1873951032;
assign addr[11178] = -1864537518;
assign addr[11179] = -1854976157;
assign addr[11180] = -1845267708;
assign addr[11181] = -1835412941;
assign addr[11182] = -1825412636;
assign addr[11183] = -1815267588;
assign addr[11184] = -1804978599;
assign addr[11185] = -1794546487;
assign addr[11186] = -1783972079;
assign addr[11187] = -1773256212;
assign addr[11188] = -1762399737;
assign addr[11189] = -1751403515;
assign addr[11190] = -1740268417;
assign addr[11191] = -1728995326;
assign addr[11192] = -1717585136;
assign addr[11193] = -1706038753;
assign addr[11194] = -1694357091;
assign addr[11195] = -1682541077;
assign addr[11196] = -1670591647;
assign addr[11197] = -1658509750;
assign addr[11198] = -1646296344;
assign addr[11199] = -1633952396;
assign addr[11200] = -1621478885;
assign addr[11201] = -1608876801;
assign addr[11202] = -1596147143;
assign addr[11203] = -1583290921;
assign addr[11204] = -1570309153;
assign addr[11205] = -1557202869;
assign addr[11206] = -1543973108;
assign addr[11207] = -1530620920;
assign addr[11208] = -1517147363;
assign addr[11209] = -1503553506;
assign addr[11210] = -1489840425;
assign addr[11211] = -1476009210;
assign addr[11212] = -1462060956;
assign addr[11213] = -1447996770;
assign addr[11214] = -1433817766;
assign addr[11215] = -1419525069;
assign addr[11216] = -1405119813;
assign addr[11217] = -1390603139;
assign addr[11218] = -1375976199;
assign addr[11219] = -1361240152;
assign addr[11220] = -1346396168;
assign addr[11221] = -1331445422;
assign addr[11222] = -1316389101;
assign addr[11223] = -1301228398;
assign addr[11224] = -1285964516;
assign addr[11225] = -1270598665;
assign addr[11226] = -1255132063;
assign addr[11227] = -1239565936;
assign addr[11228] = -1223901520;
assign addr[11229] = -1208140056;
assign addr[11230] = -1192282793;
assign addr[11231] = -1176330990;
assign addr[11232] = -1160285911;
assign addr[11233] = -1144148829;
assign addr[11234] = -1127921022;
assign addr[11235] = -1111603778;
assign addr[11236] = -1095198391;
assign addr[11237] = -1078706161;
assign addr[11238] = -1062128397;
assign addr[11239] = -1045466412;
assign addr[11240] = -1028721528;
assign addr[11241] = -1011895073;
assign addr[11242] = -994988380;
assign addr[11243] = -978002791;
assign addr[11244] = -960939653;
assign addr[11245] = -943800318;
assign addr[11246] = -926586145;
assign addr[11247] = -909298500;
assign addr[11248] = -891938752;
assign addr[11249] = -874508280;
assign addr[11250] = -857008464;
assign addr[11251] = -839440693;
assign addr[11252] = -821806359;
assign addr[11253] = -804106861;
assign addr[11254] = -786343603;
assign addr[11255] = -768517992;
assign addr[11256] = -750631442;
assign addr[11257] = -732685372;
assign addr[11258] = -714681204;
assign addr[11259] = -696620367;
assign addr[11260] = -678504291;
assign addr[11261] = -660334415;
assign addr[11262] = -642112178;
assign addr[11263] = -623839025;
assign addr[11264] = -605516406;
assign addr[11265] = -587145773;
assign addr[11266] = -568728583;
assign addr[11267] = -550266296;
assign addr[11268] = -531760377;
assign addr[11269] = -513212292;
assign addr[11270] = -494623513;
assign addr[11271] = -475995513;
assign addr[11272] = -457329769;
assign addr[11273] = -438627762;
assign addr[11274] = -419890975;
assign addr[11275] = -401120892;
assign addr[11276] = -382319004;
assign addr[11277] = -363486799;
assign addr[11278] = -344625773;
assign addr[11279] = -325737419;
assign addr[11280] = -306823237;
assign addr[11281] = -287884725;
assign addr[11282] = -268923386;
assign addr[11283] = -249940723;
assign addr[11284] = -230938242;
assign addr[11285] = -211917448;
assign addr[11286] = -192879850;
assign addr[11287] = -173826959;
assign addr[11288] = -154760284;
assign addr[11289] = -135681337;
assign addr[11290] = -116591632;
assign addr[11291] = -97492681;
assign addr[11292] = -78386000;
assign addr[11293] = -59273104;
assign addr[11294] = -40155507;
assign addr[11295] = -21034727;
assign addr[11296] = -1912278;
assign addr[11297] = 17210322;
assign addr[11298] = 36331557;
assign addr[11299] = 55449912;
assign addr[11300] = 74563870;
assign addr[11301] = 93671915;
assign addr[11302] = 112772533;
assign addr[11303] = 131864208;
assign addr[11304] = 150945428;
assign addr[11305] = 170014678;
assign addr[11306] = 189070447;
assign addr[11307] = 208111224;
assign addr[11308] = 227135500;
assign addr[11309] = 246141764;
assign addr[11310] = 265128512;
assign addr[11311] = 284094236;
assign addr[11312] = 303037433;
assign addr[11313] = 321956601;
assign addr[11314] = 340850240;
assign addr[11315] = 359716852;
assign addr[11316] = 378554940;
assign addr[11317] = 397363011;
assign addr[11318] = 416139574;
assign addr[11319] = 434883140;
assign addr[11320] = 453592221;
assign addr[11321] = 472265336;
assign addr[11322] = 490901003;
assign addr[11323] = 509497745;
assign addr[11324] = 528054086;
assign addr[11325] = 546568556;
assign addr[11326] = 565039687;
assign addr[11327] = 583466013;
assign addr[11328] = 601846074;
assign addr[11329] = 620178412;
assign addr[11330] = 638461574;
assign addr[11331] = 656694110;
assign addr[11332] = 674874574;
assign addr[11333] = 693001525;
assign addr[11334] = 711073524;
assign addr[11335] = 729089140;
assign addr[11336] = 747046944;
assign addr[11337] = 764945512;
assign addr[11338] = 782783424;
assign addr[11339] = 800559266;
assign addr[11340] = 818271628;
assign addr[11341] = 835919107;
assign addr[11342] = 853500302;
assign addr[11343] = 871013820;
assign addr[11344] = 888458272;
assign addr[11345] = 905832274;
assign addr[11346] = 923134450;
assign addr[11347] = 940363427;
assign addr[11348] = 957517838;
assign addr[11349] = 974596324;
assign addr[11350] = 991597531;
assign addr[11351] = 1008520110;
assign addr[11352] = 1025362720;
assign addr[11353] = 1042124025;
assign addr[11354] = 1058802695;
assign addr[11355] = 1075397409;
assign addr[11356] = 1091906851;
assign addr[11357] = 1108329711;
assign addr[11358] = 1124664687;
assign addr[11359] = 1140910484;
assign addr[11360] = 1157065814;
assign addr[11361] = 1173129396;
assign addr[11362] = 1189099956;
assign addr[11363] = 1204976227;
assign addr[11364] = 1220756951;
assign addr[11365] = 1236440877;
assign addr[11366] = 1252026760;
assign addr[11367] = 1267513365;
assign addr[11368] = 1282899464;
assign addr[11369] = 1298183838;
assign addr[11370] = 1313365273;
assign addr[11371] = 1328442566;
assign addr[11372] = 1343414522;
assign addr[11373] = 1358279953;
assign addr[11374] = 1373037681;
assign addr[11375] = 1387686535;
assign addr[11376] = 1402225355;
assign addr[11377] = 1416652986;
assign addr[11378] = 1430968286;
assign addr[11379] = 1445170118;
assign addr[11380] = 1459257358;
assign addr[11381] = 1473228887;
assign addr[11382] = 1487083598;
assign addr[11383] = 1500820393;
assign addr[11384] = 1514438181;
assign addr[11385] = 1527935884;
assign addr[11386] = 1541312431;
assign addr[11387] = 1554566762;
assign addr[11388] = 1567697824;
assign addr[11389] = 1580704578;
assign addr[11390] = 1593585992;
assign addr[11391] = 1606341043;
assign addr[11392] = 1618968722;
assign addr[11393] = 1631468027;
assign addr[11394] = 1643837966;
assign addr[11395] = 1656077559;
assign addr[11396] = 1668185835;
assign addr[11397] = 1680161834;
assign addr[11398] = 1692004606;
assign addr[11399] = 1703713213;
assign addr[11400] = 1715286726;
assign addr[11401] = 1726724227;
assign addr[11402] = 1738024810;
assign addr[11403] = 1749187577;
assign addr[11404] = 1760211645;
assign addr[11405] = 1771096139;
assign addr[11406] = 1781840195;
assign addr[11407] = 1792442963;
assign addr[11408] = 1802903601;
assign addr[11409] = 1813221279;
assign addr[11410] = 1823395180;
assign addr[11411] = 1833424497;
assign addr[11412] = 1843308435;
assign addr[11413] = 1853046210;
assign addr[11414] = 1862637049;
assign addr[11415] = 1872080193;
assign addr[11416] = 1881374892;
assign addr[11417] = 1890520410;
assign addr[11418] = 1899516021;
assign addr[11419] = 1908361011;
assign addr[11420] = 1917054681;
assign addr[11421] = 1925596340;
assign addr[11422] = 1933985310;
assign addr[11423] = 1942220928;
assign addr[11424] = 1950302539;
assign addr[11425] = 1958229503;
assign addr[11426] = 1966001192;
assign addr[11427] = 1973616989;
assign addr[11428] = 1981076290;
assign addr[11429] = 1988378503;
assign addr[11430] = 1995523051;
assign addr[11431] = 2002509365;
assign addr[11432] = 2009336893;
assign addr[11433] = 2016005093;
assign addr[11434] = 2022513436;
assign addr[11435] = 2028861406;
assign addr[11436] = 2035048499;
assign addr[11437] = 2041074226;
assign addr[11438] = 2046938108;
assign addr[11439] = 2052639680;
assign addr[11440] = 2058178491;
assign addr[11441] = 2063554100;
assign addr[11442] = 2068766083;
assign addr[11443] = 2073814024;
assign addr[11444] = 2078697525;
assign addr[11445] = 2083416198;
assign addr[11446] = 2087969669;
assign addr[11447] = 2092357577;
assign addr[11448] = 2096579573;
assign addr[11449] = 2100635323;
assign addr[11450] = 2104524506;
assign addr[11451] = 2108246813;
assign addr[11452] = 2111801949;
assign addr[11453] = 2115189632;
assign addr[11454] = 2118409593;
assign addr[11455] = 2121461578;
assign addr[11456] = 2124345343;
assign addr[11457] = 2127060661;
assign addr[11458] = 2129607316;
assign addr[11459] = 2131985106;
assign addr[11460] = 2134193842;
assign addr[11461] = 2136233350;
assign addr[11462] = 2138103468;
assign addr[11463] = 2139804048;
assign addr[11464] = 2141334954;
assign addr[11465] = 2142696065;
assign addr[11466] = 2143887273;
assign addr[11467] = 2144908484;
assign addr[11468] = 2145759618;
assign addr[11469] = 2146440605;
assign addr[11470] = 2146951393;
assign addr[11471] = 2147291941;
assign addr[11472] = 2147462221;
assign addr[11473] = 2147462221;
assign addr[11474] = 2147291941;
assign addr[11475] = 2146951393;
assign addr[11476] = 2146440605;
assign addr[11477] = 2145759618;
assign addr[11478] = 2144908484;
assign addr[11479] = 2143887273;
assign addr[11480] = 2142696065;
assign addr[11481] = 2141334954;
assign addr[11482] = 2139804048;
assign addr[11483] = 2138103468;
assign addr[11484] = 2136233350;
assign addr[11485] = 2134193842;
assign addr[11486] = 2131985106;
assign addr[11487] = 2129607316;
assign addr[11488] = 2127060661;
assign addr[11489] = 2124345343;
assign addr[11490] = 2121461578;
assign addr[11491] = 2118409593;
assign addr[11492] = 2115189632;
assign addr[11493] = 2111801949;
assign addr[11494] = 2108246813;
assign addr[11495] = 2104524506;
assign addr[11496] = 2100635323;
assign addr[11497] = 2096579573;
assign addr[11498] = 2092357577;
assign addr[11499] = 2087969669;
assign addr[11500] = 2083416198;
assign addr[11501] = 2078697525;
assign addr[11502] = 2073814024;
assign addr[11503] = 2068766083;
assign addr[11504] = 2063554100;
assign addr[11505] = 2058178491;
assign addr[11506] = 2052639680;
assign addr[11507] = 2046938108;
assign addr[11508] = 2041074226;
assign addr[11509] = 2035048499;
assign addr[11510] = 2028861406;
assign addr[11511] = 2022513436;
assign addr[11512] = 2016005093;
assign addr[11513] = 2009336893;
assign addr[11514] = 2002509365;
assign addr[11515] = 1995523051;
assign addr[11516] = 1988378503;
assign addr[11517] = 1981076290;
assign addr[11518] = 1973616989;
assign addr[11519] = 1966001192;
assign addr[11520] = 1958229503;
assign addr[11521] = 1950302539;
assign addr[11522] = 1942220928;
assign addr[11523] = 1933985310;
assign addr[11524] = 1925596340;
assign addr[11525] = 1917054681;
assign addr[11526] = 1908361011;
assign addr[11527] = 1899516021;
assign addr[11528] = 1890520410;
assign addr[11529] = 1881374892;
assign addr[11530] = 1872080193;
assign addr[11531] = 1862637049;
assign addr[11532] = 1853046210;
assign addr[11533] = 1843308435;
assign addr[11534] = 1833424497;
assign addr[11535] = 1823395180;
assign addr[11536] = 1813221279;
assign addr[11537] = 1802903601;
assign addr[11538] = 1792442963;
assign addr[11539] = 1781840195;
assign addr[11540] = 1771096139;
assign addr[11541] = 1760211645;
assign addr[11542] = 1749187577;
assign addr[11543] = 1738024810;
assign addr[11544] = 1726724227;
assign addr[11545] = 1715286726;
assign addr[11546] = 1703713213;
assign addr[11547] = 1692004606;
assign addr[11548] = 1680161834;
assign addr[11549] = 1668185835;
assign addr[11550] = 1656077559;
assign addr[11551] = 1643837966;
assign addr[11552] = 1631468027;
assign addr[11553] = 1618968722;
assign addr[11554] = 1606341043;
assign addr[11555] = 1593585992;
assign addr[11556] = 1580704578;
assign addr[11557] = 1567697824;
assign addr[11558] = 1554566762;
assign addr[11559] = 1541312431;
assign addr[11560] = 1527935884;
assign addr[11561] = 1514438181;
assign addr[11562] = 1500820393;
assign addr[11563] = 1487083598;
assign addr[11564] = 1473228887;
assign addr[11565] = 1459257358;
assign addr[11566] = 1445170118;
assign addr[11567] = 1430968286;
assign addr[11568] = 1416652986;
assign addr[11569] = 1402225355;
assign addr[11570] = 1387686535;
assign addr[11571] = 1373037681;
assign addr[11572] = 1358279953;
assign addr[11573] = 1343414522;
assign addr[11574] = 1328442566;
assign addr[11575] = 1313365273;
assign addr[11576] = 1298183838;
assign addr[11577] = 1282899464;
assign addr[11578] = 1267513365;
assign addr[11579] = 1252026760;
assign addr[11580] = 1236440877;
assign addr[11581] = 1220756951;
assign addr[11582] = 1204976227;
assign addr[11583] = 1189099956;
assign addr[11584] = 1173129396;
assign addr[11585] = 1157065814;
assign addr[11586] = 1140910484;
assign addr[11587] = 1124664687;
assign addr[11588] = 1108329711;
assign addr[11589] = 1091906851;
assign addr[11590] = 1075397409;
assign addr[11591] = 1058802695;
assign addr[11592] = 1042124025;
assign addr[11593] = 1025362720;
assign addr[11594] = 1008520110;
assign addr[11595] = 991597531;
assign addr[11596] = 974596324;
assign addr[11597] = 957517838;
assign addr[11598] = 940363427;
assign addr[11599] = 923134450;
assign addr[11600] = 905832274;
assign addr[11601] = 888458272;
assign addr[11602] = 871013820;
assign addr[11603] = 853500302;
assign addr[11604] = 835919107;
assign addr[11605] = 818271628;
assign addr[11606] = 800559266;
assign addr[11607] = 782783424;
assign addr[11608] = 764945512;
assign addr[11609] = 747046944;
assign addr[11610] = 729089140;
assign addr[11611] = 711073524;
assign addr[11612] = 693001525;
assign addr[11613] = 674874574;
assign addr[11614] = 656694110;
assign addr[11615] = 638461574;
assign addr[11616] = 620178412;
assign addr[11617] = 601846074;
assign addr[11618] = 583466013;
assign addr[11619] = 565039687;
assign addr[11620] = 546568556;
assign addr[11621] = 528054086;
assign addr[11622] = 509497745;
assign addr[11623] = 490901003;
assign addr[11624] = 472265336;
assign addr[11625] = 453592221;
assign addr[11626] = 434883140;
assign addr[11627] = 416139574;
assign addr[11628] = 397363011;
assign addr[11629] = 378554940;
assign addr[11630] = 359716852;
assign addr[11631] = 340850240;
assign addr[11632] = 321956601;
assign addr[11633] = 303037433;
assign addr[11634] = 284094236;
assign addr[11635] = 265128512;
assign addr[11636] = 246141764;
assign addr[11637] = 227135500;
assign addr[11638] = 208111224;
assign addr[11639] = 189070447;
assign addr[11640] = 170014678;
assign addr[11641] = 150945428;
assign addr[11642] = 131864208;
assign addr[11643] = 112772533;
assign addr[11644] = 93671915;
assign addr[11645] = 74563870;
assign addr[11646] = 55449912;
assign addr[11647] = 36331557;
assign addr[11648] = 17210322;
assign addr[11649] = -1912278;
assign addr[11650] = -21034727;
assign addr[11651] = -40155507;
assign addr[11652] = -59273104;
assign addr[11653] = -78386000;
assign addr[11654] = -97492681;
assign addr[11655] = -116591632;
assign addr[11656] = -135681337;
assign addr[11657] = -154760284;
assign addr[11658] = -173826959;
assign addr[11659] = -192879850;
assign addr[11660] = -211917448;
assign addr[11661] = -230938242;
assign addr[11662] = -249940723;
assign addr[11663] = -268923386;
assign addr[11664] = -287884725;
assign addr[11665] = -306823237;
assign addr[11666] = -325737419;
assign addr[11667] = -344625773;
assign addr[11668] = -363486799;
assign addr[11669] = -382319004;
assign addr[11670] = -401120892;
assign addr[11671] = -419890975;
assign addr[11672] = -438627762;
assign addr[11673] = -457329769;
assign addr[11674] = -475995513;
assign addr[11675] = -494623513;
assign addr[11676] = -513212292;
assign addr[11677] = -531760377;
assign addr[11678] = -550266296;
assign addr[11679] = -568728583;
assign addr[11680] = -587145773;
assign addr[11681] = -605516406;
assign addr[11682] = -623839025;
assign addr[11683] = -642112178;
assign addr[11684] = -660334415;
assign addr[11685] = -678504291;
assign addr[11686] = -696620367;
assign addr[11687] = -714681204;
assign addr[11688] = -732685372;
assign addr[11689] = -750631442;
assign addr[11690] = -768517992;
assign addr[11691] = -786343603;
assign addr[11692] = -804106861;
assign addr[11693] = -821806359;
assign addr[11694] = -839440693;
assign addr[11695] = -857008464;
assign addr[11696] = -874508280;
assign addr[11697] = -891938752;
assign addr[11698] = -909298500;
assign addr[11699] = -926586145;
assign addr[11700] = -943800318;
assign addr[11701] = -960939653;
assign addr[11702] = -978002791;
assign addr[11703] = -994988380;
assign addr[11704] = -1011895073;
assign addr[11705] = -1028721528;
assign addr[11706] = -1045466412;
assign addr[11707] = -1062128397;
assign addr[11708] = -1078706161;
assign addr[11709] = -1095198391;
assign addr[11710] = -1111603778;
assign addr[11711] = -1127921022;
assign addr[11712] = -1144148829;
assign addr[11713] = -1160285911;
assign addr[11714] = -1176330990;
assign addr[11715] = -1192282793;
assign addr[11716] = -1208140056;
assign addr[11717] = -1223901520;
assign addr[11718] = -1239565936;
assign addr[11719] = -1255132063;
assign addr[11720] = -1270598665;
assign addr[11721] = -1285964516;
assign addr[11722] = -1301228398;
assign addr[11723] = -1316389101;
assign addr[11724] = -1331445422;
assign addr[11725] = -1346396168;
assign addr[11726] = -1361240152;
assign addr[11727] = -1375976199;
assign addr[11728] = -1390603139;
assign addr[11729] = -1405119813;
assign addr[11730] = -1419525069;
assign addr[11731] = -1433817766;
assign addr[11732] = -1447996770;
assign addr[11733] = -1462060956;
assign addr[11734] = -1476009210;
assign addr[11735] = -1489840425;
assign addr[11736] = -1503553506;
assign addr[11737] = -1517147363;
assign addr[11738] = -1530620920;
assign addr[11739] = -1543973108;
assign addr[11740] = -1557202869;
assign addr[11741] = -1570309153;
assign addr[11742] = -1583290921;
assign addr[11743] = -1596147143;
assign addr[11744] = -1608876801;
assign addr[11745] = -1621478885;
assign addr[11746] = -1633952396;
assign addr[11747] = -1646296344;
assign addr[11748] = -1658509750;
assign addr[11749] = -1670591647;
assign addr[11750] = -1682541077;
assign addr[11751] = -1694357091;
assign addr[11752] = -1706038753;
assign addr[11753] = -1717585136;
assign addr[11754] = -1728995326;
assign addr[11755] = -1740268417;
assign addr[11756] = -1751403515;
assign addr[11757] = -1762399737;
assign addr[11758] = -1773256212;
assign addr[11759] = -1783972079;
assign addr[11760] = -1794546487;
assign addr[11761] = -1804978599;
assign addr[11762] = -1815267588;
assign addr[11763] = -1825412636;
assign addr[11764] = -1835412941;
assign addr[11765] = -1845267708;
assign addr[11766] = -1854976157;
assign addr[11767] = -1864537518;
assign addr[11768] = -1873951032;
assign addr[11769] = -1883215953;
assign addr[11770] = -1892331547;
assign addr[11771] = -1901297091;
assign addr[11772] = -1910111873;
assign addr[11773] = -1918775195;
assign addr[11774] = -1927286370;
assign addr[11775] = -1935644723;
assign addr[11776] = -1943849591;
assign addr[11777] = -1951900324;
assign addr[11778] = -1959796283;
assign addr[11779] = -1967536842;
assign addr[11780] = -1975121388;
assign addr[11781] = -1982549318;
assign addr[11782] = -1989820044;
assign addr[11783] = -1996932990;
assign addr[11784] = -2003887591;
assign addr[11785] = -2010683297;
assign addr[11786] = -2017319567;
assign addr[11787] = -2023795876;
assign addr[11788] = -2030111710;
assign addr[11789] = -2036266570;
assign addr[11790] = -2042259965;
assign addr[11791] = -2048091422;
assign addr[11792] = -2053760478;
assign addr[11793] = -2059266683;
assign addr[11794] = -2064609600;
assign addr[11795] = -2069788807;
assign addr[11796] = -2074803892;
assign addr[11797] = -2079654458;
assign addr[11798] = -2084340120;
assign addr[11799] = -2088860507;
assign addr[11800] = -2093215260;
assign addr[11801] = -2097404033;
assign addr[11802] = -2101426496;
assign addr[11803] = -2105282327;
assign addr[11804] = -2108971223;
assign addr[11805] = -2112492891;
assign addr[11806] = -2115847050;
assign addr[11807] = -2119033436;
assign addr[11808] = -2122051796;
assign addr[11809] = -2124901890;
assign addr[11810] = -2127583492;
assign addr[11811] = -2130096389;
assign addr[11812] = -2132440383;
assign addr[11813] = -2134615288;
assign addr[11814] = -2136620930;
assign addr[11815] = -2138457152;
assign addr[11816] = -2140123807;
assign addr[11817] = -2141620763;
assign addr[11818] = -2142947902;
assign addr[11819] = -2144105118;
assign addr[11820] = -2145092320;
assign addr[11821] = -2145909429;
assign addr[11822] = -2146556380;
assign addr[11823] = -2147033123;
assign addr[11824] = -2147339619;
assign addr[11825] = -2147475844;
assign addr[11826] = -2147441787;
assign addr[11827] = -2147237452;
assign addr[11828] = -2146862854;
assign addr[11829] = -2146318022;
assign addr[11830] = -2145603001;
assign addr[11831] = -2144717846;
assign addr[11832] = -2143662628;
assign addr[11833] = -2142437431;
assign addr[11834] = -2141042352;
assign addr[11835] = -2139477502;
assign addr[11836] = -2137743003;
assign addr[11837] = -2135838995;
assign addr[11838] = -2133765628;
assign addr[11839] = -2131523066;
assign addr[11840] = -2129111488;
assign addr[11841] = -2126531084;
assign addr[11842] = -2123782059;
assign addr[11843] = -2120864631;
assign addr[11844] = -2117779031;
assign addr[11845] = -2114525505;
assign addr[11846] = -2111104309;
assign addr[11847] = -2107515716;
assign addr[11848] = -2103760010;
assign addr[11849] = -2099837489;
assign addr[11850] = -2095748463;
assign addr[11851] = -2091493257;
assign addr[11852] = -2087072209;
assign addr[11853] = -2082485668;
assign addr[11854] = -2077733999;
assign addr[11855] = -2072817579;
assign addr[11856] = -2067736796;
assign addr[11857] = -2062492055;
assign addr[11858] = -2057083771;
assign addr[11859] = -2051512372;
assign addr[11860] = -2045778302;
assign addr[11861] = -2039882013;
assign addr[11862] = -2033823974;
assign addr[11863] = -2027604666;
assign addr[11864] = -2021224581;
assign addr[11865] = -2014684225;
assign addr[11866] = -2007984117;
assign addr[11867] = -2001124788;
assign addr[11868] = -1994106782;
assign addr[11869] = -1986930656;
assign addr[11870] = -1979596978;
assign addr[11871] = -1972106330;
assign addr[11872] = -1964459306;
assign addr[11873] = -1956656513;
assign addr[11874] = -1948698568;
assign addr[11875] = -1940586104;
assign addr[11876] = -1932319763;
assign addr[11877] = -1923900201;
assign addr[11878] = -1915328086;
assign addr[11879] = -1906604097;
assign addr[11880] = -1897728925;
assign addr[11881] = -1888703276;
assign addr[11882] = -1879527863;
assign addr[11883] = -1870203416;
assign addr[11884] = -1860730673;
assign addr[11885] = -1851110385;
assign addr[11886] = -1841343316;
assign addr[11887] = -1831430239;
assign addr[11888] = -1821371941;
assign addr[11889] = -1811169220;
assign addr[11890] = -1800822883;
assign addr[11891] = -1790333753;
assign addr[11892] = -1779702660;
assign addr[11893] = -1768930447;
assign addr[11894] = -1758017969;
assign addr[11895] = -1746966091;
assign addr[11896] = -1735775690;
assign addr[11897] = -1724447652;
assign addr[11898] = -1712982875;
assign addr[11899] = -1701382270;
assign addr[11900] = -1689646755;
assign addr[11901] = -1677777262;
assign addr[11902] = -1665774731;
assign addr[11903] = -1653640115;
assign addr[11904] = -1641374375;
assign addr[11905] = -1628978484;
assign addr[11906] = -1616453425;
assign addr[11907] = -1603800191;
assign addr[11908] = -1591019785;
assign addr[11909] = -1578113222;
assign addr[11910] = -1565081523;
assign addr[11911] = -1551925723;
assign addr[11912] = -1538646865;
assign addr[11913] = -1525246002;
assign addr[11914] = -1511724196;
assign addr[11915] = -1498082520;
assign addr[11916] = -1484322054;
assign addr[11917] = -1470443891;
assign addr[11918] = -1456449131;
assign addr[11919] = -1442338884;
assign addr[11920] = -1428114267;
assign addr[11921] = -1413776410;
assign addr[11922] = -1399326449;
assign addr[11923] = -1384765530;
assign addr[11924] = -1370094808;
assign addr[11925] = -1355315445;
assign addr[11926] = -1340428615;
assign addr[11927] = -1325435496;
assign addr[11928] = -1310337279;
assign addr[11929] = -1295135159;
assign addr[11930] = -1279830344;
assign addr[11931] = -1264424045;
assign addr[11932] = -1248917486;
assign addr[11933] = -1233311895;
assign addr[11934] = -1217608510;
assign addr[11935] = -1201808576;
assign addr[11936] = -1185913346;
assign addr[11937] = -1169924081;
assign addr[11938] = -1153842047;
assign addr[11939] = -1137668521;
assign addr[11940] = -1121404785;
assign addr[11941] = -1105052128;
assign addr[11942] = -1088611847;
assign addr[11943] = -1072085246;
assign addr[11944] = -1055473635;
assign addr[11945] = -1038778332;
assign addr[11946] = -1022000660;
assign addr[11947] = -1005141949;
assign addr[11948] = -988203537;
assign addr[11949] = -971186766;
assign addr[11950] = -954092986;
assign addr[11951] = -936923553;
assign addr[11952] = -919679827;
assign addr[11953] = -902363176;
assign addr[11954] = -884974973;
assign addr[11955] = -867516597;
assign addr[11956] = -849989433;
assign addr[11957] = -832394869;
assign addr[11958] = -814734301;
assign addr[11959] = -797009130;
assign addr[11960] = -779220762;
assign addr[11961] = -761370605;
assign addr[11962] = -743460077;
assign addr[11963] = -725490597;
assign addr[11964] = -707463589;
assign addr[11965] = -689380485;
assign addr[11966] = -671242716;
assign addr[11967] = -653051723;
assign addr[11968] = -634808946;
assign addr[11969] = -616515832;
assign addr[11970] = -598173833;
assign addr[11971] = -579784402;
assign addr[11972] = -561348998;
assign addr[11973] = -542869083;
assign addr[11974] = -524346121;
assign addr[11975] = -505781581;
assign addr[11976] = -487176937;
assign addr[11977] = -468533662;
assign addr[11978] = -449853235;
assign addr[11979] = -431137138;
assign addr[11980] = -412386854;
assign addr[11981] = -393603870;
assign addr[11982] = -374789676;
assign addr[11983] = -355945764;
assign addr[11984] = -337073627;
assign addr[11985] = -318174762;
assign addr[11986] = -299250668;
assign addr[11987] = -280302845;
assign addr[11988] = -261332796;
assign addr[11989] = -242342025;
assign addr[11990] = -223332037;
assign addr[11991] = -204304341;
assign addr[11992] = -185260444;
assign addr[11993] = -166201858;
assign addr[11994] = -147130093;
assign addr[11995] = -128046661;
assign addr[11996] = -108953076;
assign addr[11997] = -89850852;
assign addr[11998] = -70741503;
assign addr[11999] = -51626544;
assign addr[12000] = -32507492;
assign addr[12001] = -13385863;
assign addr[12002] = 5736829;
assign addr[12003] = 24859065;
assign addr[12004] = 43979330;
assign addr[12005] = 63096108;
assign addr[12006] = 82207882;
assign addr[12007] = 101313138;
assign addr[12008] = 120410361;
assign addr[12009] = 139498035;
assign addr[12010] = 158574649;
assign addr[12011] = 177638688;
assign addr[12012] = 196688642;
assign addr[12013] = 215722999;
assign addr[12014] = 234740251;
assign addr[12015] = 253738890;
assign addr[12016] = 272717408;
assign addr[12017] = 291674302;
assign addr[12018] = 310608068;
assign addr[12019] = 329517204;
assign addr[12020] = 348400212;
assign addr[12021] = 367255594;
assign addr[12022] = 386081854;
assign addr[12023] = 404877501;
assign addr[12024] = 423641043;
assign addr[12025] = 442370993;
assign addr[12026] = 461065866;
assign addr[12027] = 479724180;
assign addr[12028] = 498344454;
assign addr[12029] = 516925212;
assign addr[12030] = 535464981;
assign addr[12031] = 553962291;
assign addr[12032] = 572415676;
assign addr[12033] = 590823671;
assign addr[12034] = 609184818;
assign addr[12035] = 627497660;
assign addr[12036] = 645760745;
assign addr[12037] = 663972625;
assign addr[12038] = 682131857;
assign addr[12039] = 700236999;
assign addr[12040] = 718286617;
assign addr[12041] = 736279279;
assign addr[12042] = 754213559;
assign addr[12043] = 772088034;
assign addr[12044] = 789901288;
assign addr[12045] = 807651907;
assign addr[12046] = 825338484;
assign addr[12047] = 842959617;
assign addr[12048] = 860513908;
assign addr[12049] = 877999966;
assign addr[12050] = 895416404;
assign addr[12051] = 912761841;
assign addr[12052] = 930034901;
assign addr[12053] = 947234215;
assign addr[12054] = 964358420;
assign addr[12055] = 981406156;
assign addr[12056] = 998376073;
assign addr[12057] = 1015266825;
assign addr[12058] = 1032077073;
assign addr[12059] = 1048805483;
assign addr[12060] = 1065450729;
assign addr[12061] = 1082011492;
assign addr[12062] = 1098486458;
assign addr[12063] = 1114874320;
assign addr[12064] = 1131173780;
assign addr[12065] = 1147383544;
assign addr[12066] = 1163502328;
assign addr[12067] = 1179528853;
assign addr[12068] = 1195461849;
assign addr[12069] = 1211300053;
assign addr[12070] = 1227042207;
assign addr[12071] = 1242687064;
assign addr[12072] = 1258233384;
assign addr[12073] = 1273679934;
assign addr[12074] = 1289025489;
assign addr[12075] = 1304268832;
assign addr[12076] = 1319408754;
assign addr[12077] = 1334444055;
assign addr[12078] = 1349373543;
assign addr[12079] = 1364196034;
assign addr[12080] = 1378910353;
assign addr[12081] = 1393515332;
assign addr[12082] = 1408009814;
assign addr[12083] = 1422392650;
assign addr[12084] = 1436662698;
assign addr[12085] = 1450818828;
assign addr[12086] = 1464859917;
assign addr[12087] = 1478784851;
assign addr[12088] = 1492592527;
assign addr[12089] = 1506281850;
assign addr[12090] = 1519851733;
assign addr[12091] = 1533301101;
assign addr[12092] = 1546628888;
assign addr[12093] = 1559834037;
assign addr[12094] = 1572915501;
assign addr[12095] = 1585872242;
assign addr[12096] = 1598703233;
assign addr[12097] = 1611407456;
assign addr[12098] = 1623983905;
assign addr[12099] = 1636431582;
assign addr[12100] = 1648749499;
assign addr[12101] = 1660936681;
assign addr[12102] = 1672992161;
assign addr[12103] = 1684914983;
assign addr[12104] = 1696704201;
assign addr[12105] = 1708358881;
assign addr[12106] = 1719878099;
assign addr[12107] = 1731260941;
assign addr[12108] = 1742506504;
assign addr[12109] = 1753613897;
assign addr[12110] = 1764582240;
assign addr[12111] = 1775410662;
assign addr[12112] = 1786098304;
assign addr[12113] = 1796644320;
assign addr[12114] = 1807047873;
assign addr[12115] = 1817308138;
assign addr[12116] = 1827424302;
assign addr[12117] = 1837395562;
assign addr[12118] = 1847221128;
assign addr[12119] = 1856900221;
assign addr[12120] = 1866432072;
assign addr[12121] = 1875815927;
assign addr[12122] = 1885051042;
assign addr[12123] = 1894136683;
assign addr[12124] = 1903072131;
assign addr[12125] = 1911856677;
assign addr[12126] = 1920489624;
assign addr[12127] = 1928970288;
assign addr[12128] = 1937297997;
assign addr[12129] = 1945472089;
assign addr[12130] = 1953491918;
assign addr[12131] = 1961356847;
assign addr[12132] = 1969066252;
assign addr[12133] = 1976619522;
assign addr[12134] = 1984016058;
assign addr[12135] = 1991255274;
assign addr[12136] = 1998336596;
assign addr[12137] = 2005259462;
assign addr[12138] = 2012023322;
assign addr[12139] = 2018627642;
assign addr[12140] = 2025071897;
assign addr[12141] = 2031355576;
assign addr[12142] = 2037478181;
assign addr[12143] = 2043439226;
assign addr[12144] = 2049238240;
assign addr[12145] = 2054874761;
assign addr[12146] = 2060348343;
assign addr[12147] = 2065658552;
assign addr[12148] = 2070804967;
assign addr[12149] = 2075787180;
assign addr[12150] = 2080604795;
assign addr[12151] = 2085257431;
assign addr[12152] = 2089744719;
assign addr[12153] = 2094066304;
assign addr[12154] = 2098221841;
assign addr[12155] = 2102211002;
assign addr[12156] = 2106033471;
assign addr[12157] = 2109688944;
assign addr[12158] = 2113177132;
assign addr[12159] = 2116497758;
assign addr[12160] = 2119650558;
assign addr[12161] = 2122635283;
assign addr[12162] = 2125451696;
assign addr[12163] = 2128099574;
assign addr[12164] = 2130578706;
assign addr[12165] = 2132888897;
assign addr[12166] = 2135029962;
assign addr[12167] = 2137001733;
assign addr[12168] = 2138804053;
assign addr[12169] = 2140436778;
assign addr[12170] = 2141899780;
assign addr[12171] = 2143192942;
assign addr[12172] = 2144316162;
assign addr[12173] = 2145269351;
assign addr[12174] = 2146052433;
assign addr[12175] = 2146665347;
assign addr[12176] = 2147108043;
assign addr[12177] = 2147380486;
assign addr[12178] = 2147482655;
assign addr[12179] = 2147414542;
assign addr[12180] = 2147176152;
assign addr[12181] = 2146767505;
assign addr[12182] = 2146188631;
assign addr[12183] = 2145439578;
assign addr[12184] = 2144520405;
assign addr[12185] = 2143431184;
assign addr[12186] = 2142172003;
assign addr[12187] = 2140742960;
assign addr[12188] = 2139144169;
assign addr[12189] = 2137375758;
assign addr[12190] = 2135437865;
assign addr[12191] = 2133330646;
assign addr[12192] = 2131054266;
assign addr[12193] = 2128608907;
assign addr[12194] = 2125994762;
assign addr[12195] = 2123212038;
assign addr[12196] = 2120260957;
assign addr[12197] = 2117141752;
assign addr[12198] = 2113854671;
assign addr[12199] = 2110399974;
assign addr[12200] = 2106777935;
assign addr[12201] = 2102988841;
assign addr[12202] = 2099032994;
assign addr[12203] = 2094910706;
assign addr[12204] = 2090622304;
assign addr[12205] = 2086168128;
assign addr[12206] = 2081548533;
assign addr[12207] = 2076763883;
assign addr[12208] = 2071814558;
assign addr[12209] = 2066700952;
assign addr[12210] = 2061423468;
assign addr[12211] = 2055982526;
assign addr[12212] = 2050378558;
assign addr[12213] = 2044612007;
assign addr[12214] = 2038683330;
assign addr[12215] = 2032592999;
assign addr[12216] = 2026341495;
assign addr[12217] = 2019929315;
assign addr[12218] = 2013356967;
assign addr[12219] = 2006624971;
assign addr[12220] = 1999733863;
assign addr[12221] = 1992684188;
assign addr[12222] = 1985476506;
assign addr[12223] = 1978111387;
assign addr[12224] = 1970589416;
assign addr[12225] = 1962911189;
assign addr[12226] = 1955077316;
assign addr[12227] = 1947088417;
assign addr[12228] = 1938945125;
assign addr[12229] = 1930648088;
assign addr[12230] = 1922197961;
assign addr[12231] = 1913595416;
assign addr[12232] = 1904841135;
assign addr[12233] = 1895935811;
assign addr[12234] = 1886880151;
assign addr[12235] = 1877674873;
assign addr[12236] = 1868320707;
assign addr[12237] = 1858818395;
assign addr[12238] = 1849168689;
assign addr[12239] = 1839372356;
assign addr[12240] = 1829430172;
assign addr[12241] = 1819342925;
assign addr[12242] = 1809111415;
assign addr[12243] = 1798736454;
assign addr[12244] = 1788218865;
assign addr[12245] = 1777559480;
assign addr[12246] = 1766759146;
assign addr[12247] = 1755818718;
assign addr[12248] = 1744739065;
assign addr[12249] = 1733521064;
assign addr[12250] = 1722165606;
assign addr[12251] = 1710673591;
assign addr[12252] = 1699045930;
assign addr[12253] = 1687283545;
assign addr[12254] = 1675387369;
assign addr[12255] = 1663358344;
assign addr[12256] = 1651197426;
assign addr[12257] = 1638905577;
assign addr[12258] = 1626483774;
assign addr[12259] = 1613933000;
assign addr[12260] = 1601254251;
assign addr[12261] = 1588448533;
assign addr[12262] = 1575516860;
assign addr[12263] = 1562460258;
assign addr[12264] = 1549279763;
assign addr[12265] = 1535976419;
assign addr[12266] = 1522551282;
assign addr[12267] = 1509005416;
assign addr[12268] = 1495339895;
assign addr[12269] = 1481555802;
assign addr[12270] = 1467654232;
assign addr[12271] = 1453636285;
assign addr[12272] = 1439503074;
assign addr[12273] = 1425255719;
assign addr[12274] = 1410895350;
assign addr[12275] = 1396423105;
assign addr[12276] = 1381840133;
assign addr[12277] = 1367147589;
assign addr[12278] = 1352346639;
assign addr[12279] = 1337438456;
assign addr[12280] = 1322424222;
assign addr[12281] = 1307305128;
assign addr[12282] = 1292082373;
assign addr[12283] = 1276757164;
assign addr[12284] = 1261330715;
assign addr[12285] = 1245804251;
assign addr[12286] = 1230179002;
assign addr[12287] = 1214456207;
assign addr[12288] = 1198637114;
assign addr[12289] = 1182722976;
assign addr[12290] = 1166715055;
assign addr[12291] = 1150614620;
assign addr[12292] = 1134422949;
assign addr[12293] = 1118141326;
assign addr[12294] = 1101771040;
assign addr[12295] = 1085313391;
assign addr[12296] = 1068769683;
assign addr[12297] = 1052141228;
assign addr[12298] = 1035429345;
assign addr[12299] = 1018635358;
assign addr[12300] = 1001760600;
assign addr[12301] = 984806408;
assign addr[12302] = 967774128;
assign addr[12303] = 950665109;
assign addr[12304] = 933480707;
assign addr[12305] = 916222287;
assign addr[12306] = 898891215;
assign addr[12307] = 881488868;
assign addr[12308] = 864016623;
assign addr[12309] = 846475867;
assign addr[12310] = 828867991;
assign addr[12311] = 811194391;
assign addr[12312] = 793456467;
assign addr[12313] = 775655628;
assign addr[12314] = 757793284;
assign addr[12315] = 739870851;
assign addr[12316] = 721889752;
assign addr[12317] = 703851410;
assign addr[12318] = 685757258;
assign addr[12319] = 667608730;
assign addr[12320] = 649407264;
assign addr[12321] = 631154304;
assign addr[12322] = 612851297;
assign addr[12323] = 594499695;
assign addr[12324] = 576100953;
assign addr[12325] = 557656529;
assign addr[12326] = 539167887;
assign addr[12327] = 520636492;
assign addr[12328] = 502063814;
assign addr[12329] = 483451325;
assign addr[12330] = 464800501;
assign addr[12331] = 446112822;
assign addr[12332] = 427389768;
assign addr[12333] = 408632825;
assign addr[12334] = 389843480;
assign addr[12335] = 371023223;
assign addr[12336] = 352173546;
assign addr[12337] = 333295944;
assign addr[12338] = 314391913;
assign addr[12339] = 295462954;
assign addr[12340] = 276510565;
assign addr[12341] = 257536251;
assign addr[12342] = 238541516;
assign addr[12343] = 219527866;
assign addr[12344] = 200496809;
assign addr[12345] = 181449854;
assign addr[12346] = 162388511;
assign addr[12347] = 143314291;
assign addr[12348] = 124228708;
assign addr[12349] = 105133274;
assign addr[12350] = 86029503;
assign addr[12351] = 66918911;
assign addr[12352] = 47803013;
assign addr[12353] = 28683324;
assign addr[12354] = 9561361;
assign addr[12355] = -9561361;
assign addr[12356] = -28683324;
assign addr[12357] = -47803013;
assign addr[12358] = -66918911;
assign addr[12359] = -86029503;
assign addr[12360] = -105133274;
assign addr[12361] = -124228708;
assign addr[12362] = -143314291;
assign addr[12363] = -162388511;
assign addr[12364] = -181449854;
assign addr[12365] = -200496809;
assign addr[12366] = -219527866;
assign addr[12367] = -238541516;
assign addr[12368] = -257536251;
assign addr[12369] = -276510565;
assign addr[12370] = -295462954;
assign addr[12371] = -314391913;
assign addr[12372] = -333295944;
assign addr[12373] = -352173546;
assign addr[12374] = -371023223;
assign addr[12375] = -389843480;
assign addr[12376] = -408632825;
assign addr[12377] = -427389768;
assign addr[12378] = -446112822;
assign addr[12379] = -464800501;
assign addr[12380] = -483451325;
assign addr[12381] = -502063814;
assign addr[12382] = -520636492;
assign addr[12383] = -539167887;
assign addr[12384] = -557656529;
assign addr[12385] = -576100953;
assign addr[12386] = -594499695;
assign addr[12387] = -612851297;
assign addr[12388] = -631154304;
assign addr[12389] = -649407264;
assign addr[12390] = -667608730;
assign addr[12391] = -685757258;
assign addr[12392] = -703851410;
assign addr[12393] = -721889752;
assign addr[12394] = -739870851;
assign addr[12395] = -757793284;
assign addr[12396] = -775655628;
assign addr[12397] = -793456467;
assign addr[12398] = -811194391;
assign addr[12399] = -828867991;
assign addr[12400] = -846475867;
assign addr[12401] = -864016623;
assign addr[12402] = -881488868;
assign addr[12403] = -898891215;
assign addr[12404] = -916222287;
assign addr[12405] = -933480707;
assign addr[12406] = -950665109;
assign addr[12407] = -967774128;
assign addr[12408] = -984806408;
assign addr[12409] = -1001760600;
assign addr[12410] = -1018635358;
assign addr[12411] = -1035429345;
assign addr[12412] = -1052141228;
assign addr[12413] = -1068769683;
assign addr[12414] = -1085313391;
assign addr[12415] = -1101771040;
assign addr[12416] = -1118141326;
assign addr[12417] = -1134422949;
assign addr[12418] = -1150614620;
assign addr[12419] = -1166715055;
assign addr[12420] = -1182722976;
assign addr[12421] = -1198637114;
assign addr[12422] = -1214456207;
assign addr[12423] = -1230179002;
assign addr[12424] = -1245804251;
assign addr[12425] = -1261330715;
assign addr[12426] = -1276757164;
assign addr[12427] = -1292082373;
assign addr[12428] = -1307305128;
assign addr[12429] = -1322424222;
assign addr[12430] = -1337438456;
assign addr[12431] = -1352346639;
assign addr[12432] = -1367147589;
assign addr[12433] = -1381840133;
assign addr[12434] = -1396423105;
assign addr[12435] = -1410895350;
assign addr[12436] = -1425255719;
assign addr[12437] = -1439503074;
assign addr[12438] = -1453636285;
assign addr[12439] = -1467654232;
assign addr[12440] = -1481555802;
assign addr[12441] = -1495339895;
assign addr[12442] = -1509005416;
assign addr[12443] = -1522551282;
assign addr[12444] = -1535976419;
assign addr[12445] = -1549279763;
assign addr[12446] = -1562460258;
assign addr[12447] = -1575516860;
assign addr[12448] = -1588448533;
assign addr[12449] = -1601254251;
assign addr[12450] = -1613933000;
assign addr[12451] = -1626483774;
assign addr[12452] = -1638905577;
assign addr[12453] = -1651197426;
assign addr[12454] = -1663358344;
assign addr[12455] = -1675387369;
assign addr[12456] = -1687283545;
assign addr[12457] = -1699045930;
assign addr[12458] = -1710673591;
assign addr[12459] = -1722165606;
assign addr[12460] = -1733521064;
assign addr[12461] = -1744739065;
assign addr[12462] = -1755818718;
assign addr[12463] = -1766759146;
assign addr[12464] = -1777559480;
assign addr[12465] = -1788218865;
assign addr[12466] = -1798736454;
assign addr[12467] = -1809111415;
assign addr[12468] = -1819342925;
assign addr[12469] = -1829430172;
assign addr[12470] = -1839372356;
assign addr[12471] = -1849168689;
assign addr[12472] = -1858818395;
assign addr[12473] = -1868320707;
assign addr[12474] = -1877674873;
assign addr[12475] = -1886880151;
assign addr[12476] = -1895935811;
assign addr[12477] = -1904841135;
assign addr[12478] = -1913595416;
assign addr[12479] = -1922197961;
assign addr[12480] = -1930648088;
assign addr[12481] = -1938945125;
assign addr[12482] = -1947088417;
assign addr[12483] = -1955077316;
assign addr[12484] = -1962911189;
assign addr[12485] = -1970589416;
assign addr[12486] = -1978111387;
assign addr[12487] = -1985476506;
assign addr[12488] = -1992684188;
assign addr[12489] = -1999733863;
assign addr[12490] = -2006624971;
assign addr[12491] = -2013356967;
assign addr[12492] = -2019929315;
assign addr[12493] = -2026341495;
assign addr[12494] = -2032592999;
assign addr[12495] = -2038683330;
assign addr[12496] = -2044612007;
assign addr[12497] = -2050378558;
assign addr[12498] = -2055982526;
assign addr[12499] = -2061423468;
assign addr[12500] = -2066700952;
assign addr[12501] = -2071814558;
assign addr[12502] = -2076763883;
assign addr[12503] = -2081548533;
assign addr[12504] = -2086168128;
assign addr[12505] = -2090622304;
assign addr[12506] = -2094910706;
assign addr[12507] = -2099032994;
assign addr[12508] = -2102988841;
assign addr[12509] = -2106777935;
assign addr[12510] = -2110399974;
assign addr[12511] = -2113854671;
assign addr[12512] = -2117141752;
assign addr[12513] = -2120260957;
assign addr[12514] = -2123212038;
assign addr[12515] = -2125994762;
assign addr[12516] = -2128608907;
assign addr[12517] = -2131054266;
assign addr[12518] = -2133330646;
assign addr[12519] = -2135437865;
assign addr[12520] = -2137375758;
assign addr[12521] = -2139144169;
assign addr[12522] = -2140742960;
assign addr[12523] = -2142172003;
assign addr[12524] = -2143431184;
assign addr[12525] = -2144520405;
assign addr[12526] = -2145439578;
assign addr[12527] = -2146188631;
assign addr[12528] = -2146767505;
assign addr[12529] = -2147176152;
assign addr[12530] = -2147414542;
assign addr[12531] = -2147482655;
assign addr[12532] = -2147380486;
assign addr[12533] = -2147108043;
assign addr[12534] = -2146665347;
assign addr[12535] = -2146052433;
assign addr[12536] = -2145269351;
assign addr[12537] = -2144316162;
assign addr[12538] = -2143192942;
assign addr[12539] = -2141899780;
assign addr[12540] = -2140436778;
assign addr[12541] = -2138804053;
assign addr[12542] = -2137001733;
assign addr[12543] = -2135029962;
assign addr[12544] = -2132888897;
assign addr[12545] = -2130578706;
assign addr[12546] = -2128099574;
assign addr[12547] = -2125451696;
assign addr[12548] = -2122635283;
assign addr[12549] = -2119650558;
assign addr[12550] = -2116497758;
assign addr[12551] = -2113177132;
assign addr[12552] = -2109688944;
assign addr[12553] = -2106033471;
assign addr[12554] = -2102211002;
assign addr[12555] = -2098221841;
assign addr[12556] = -2094066304;
assign addr[12557] = -2089744719;
assign addr[12558] = -2085257431;
assign addr[12559] = -2080604795;
assign addr[12560] = -2075787180;
assign addr[12561] = -2070804967;
assign addr[12562] = -2065658552;
assign addr[12563] = -2060348343;
assign addr[12564] = -2054874761;
assign addr[12565] = -2049238240;
assign addr[12566] = -2043439226;
assign addr[12567] = -2037478181;
assign addr[12568] = -2031355576;
assign addr[12569] = -2025071897;
assign addr[12570] = -2018627642;
assign addr[12571] = -2012023322;
assign addr[12572] = -2005259462;
assign addr[12573] = -1998336596;
assign addr[12574] = -1991255274;
assign addr[12575] = -1984016058;
assign addr[12576] = -1976619522;
assign addr[12577] = -1969066252;
assign addr[12578] = -1961356847;
assign addr[12579] = -1953491918;
assign addr[12580] = -1945472089;
assign addr[12581] = -1937297997;
assign addr[12582] = -1928970288;
assign addr[12583] = -1920489624;
assign addr[12584] = -1911856677;
assign addr[12585] = -1903072131;
assign addr[12586] = -1894136683;
assign addr[12587] = -1885051042;
assign addr[12588] = -1875815927;
assign addr[12589] = -1866432072;
assign addr[12590] = -1856900221;
assign addr[12591] = -1847221128;
assign addr[12592] = -1837395562;
assign addr[12593] = -1827424302;
assign addr[12594] = -1817308138;
assign addr[12595] = -1807047873;
assign addr[12596] = -1796644320;
assign addr[12597] = -1786098304;
assign addr[12598] = -1775410662;
assign addr[12599] = -1764582240;
assign addr[12600] = -1753613897;
assign addr[12601] = -1742506504;
assign addr[12602] = -1731260941;
assign addr[12603] = -1719878099;
assign addr[12604] = -1708358881;
assign addr[12605] = -1696704201;
assign addr[12606] = -1684914983;
assign addr[12607] = -1672992161;
assign addr[12608] = -1660936681;
assign addr[12609] = -1648749499;
assign addr[12610] = -1636431582;
assign addr[12611] = -1623983905;
assign addr[12612] = -1611407456;
assign addr[12613] = -1598703233;
assign addr[12614] = -1585872242;
assign addr[12615] = -1572915501;
assign addr[12616] = -1559834037;
assign addr[12617] = -1546628888;
assign addr[12618] = -1533301101;
assign addr[12619] = -1519851733;
assign addr[12620] = -1506281850;
assign addr[12621] = -1492592527;
assign addr[12622] = -1478784851;
assign addr[12623] = -1464859917;
assign addr[12624] = -1450818828;
assign addr[12625] = -1436662698;
assign addr[12626] = -1422392650;
assign addr[12627] = -1408009814;
assign addr[12628] = -1393515332;
assign addr[12629] = -1378910353;
assign addr[12630] = -1364196034;
assign addr[12631] = -1349373543;
assign addr[12632] = -1334444055;
assign addr[12633] = -1319408754;
assign addr[12634] = -1304268832;
assign addr[12635] = -1289025489;
assign addr[12636] = -1273679934;
assign addr[12637] = -1258233384;
assign addr[12638] = -1242687064;
assign addr[12639] = -1227042207;
assign addr[12640] = -1211300053;
assign addr[12641] = -1195461849;
assign addr[12642] = -1179528853;
assign addr[12643] = -1163502328;
assign addr[12644] = -1147383544;
assign addr[12645] = -1131173780;
assign addr[12646] = -1114874320;
assign addr[12647] = -1098486458;
assign addr[12648] = -1082011492;
assign addr[12649] = -1065450729;
assign addr[12650] = -1048805483;
assign addr[12651] = -1032077073;
assign addr[12652] = -1015266825;
assign addr[12653] = -998376073;
assign addr[12654] = -981406156;
assign addr[12655] = -964358420;
assign addr[12656] = -947234215;
assign addr[12657] = -930034901;
assign addr[12658] = -912761841;
assign addr[12659] = -895416404;
assign addr[12660] = -877999966;
assign addr[12661] = -860513908;
assign addr[12662] = -842959617;
assign addr[12663] = -825338484;
assign addr[12664] = -807651907;
assign addr[12665] = -789901288;
assign addr[12666] = -772088034;
assign addr[12667] = -754213559;
assign addr[12668] = -736279279;
assign addr[12669] = -718286617;
assign addr[12670] = -700236999;
assign addr[12671] = -682131857;
assign addr[12672] = -663972625;
assign addr[12673] = -645760745;
assign addr[12674] = -627497660;
assign addr[12675] = -609184818;
assign addr[12676] = -590823671;
assign addr[12677] = -572415676;
assign addr[12678] = -553962291;
assign addr[12679] = -535464981;
assign addr[12680] = -516925212;
assign addr[12681] = -498344454;
assign addr[12682] = -479724180;
assign addr[12683] = -461065866;
assign addr[12684] = -442370993;
assign addr[12685] = -423641043;
assign addr[12686] = -404877501;
assign addr[12687] = -386081854;
assign addr[12688] = -367255594;
assign addr[12689] = -348400212;
assign addr[12690] = -329517204;
assign addr[12691] = -310608068;
assign addr[12692] = -291674302;
assign addr[12693] = -272717408;
assign addr[12694] = -253738890;
assign addr[12695] = -234740251;
assign addr[12696] = -215722999;
assign addr[12697] = -196688642;
assign addr[12698] = -177638688;
assign addr[12699] = -158574649;
assign addr[12700] = -139498035;
assign addr[12701] = -120410361;
assign addr[12702] = -101313138;
assign addr[12703] = -82207882;
assign addr[12704] = -63096108;
assign addr[12705] = -43979330;
assign addr[12706] = -24859065;
assign addr[12707] = -5736829;
assign addr[12708] = 13385863;
assign addr[12709] = 32507492;
assign addr[12710] = 51626544;
assign addr[12711] = 70741503;
assign addr[12712] = 89850852;
assign addr[12713] = 108953076;
assign addr[12714] = 128046661;
assign addr[12715] = 147130093;
assign addr[12716] = 166201858;
assign addr[12717] = 185260444;
assign addr[12718] = 204304341;
assign addr[12719] = 223332037;
assign addr[12720] = 242342025;
assign addr[12721] = 261332796;
assign addr[12722] = 280302845;
assign addr[12723] = 299250668;
assign addr[12724] = 318174762;
assign addr[12725] = 337073627;
assign addr[12726] = 355945764;
assign addr[12727] = 374789676;
assign addr[12728] = 393603870;
assign addr[12729] = 412386854;
assign addr[12730] = 431137138;
assign addr[12731] = 449853235;
assign addr[12732] = 468533662;
assign addr[12733] = 487176937;
assign addr[12734] = 505781581;
assign addr[12735] = 524346121;
assign addr[12736] = 542869083;
assign addr[12737] = 561348998;
assign addr[12738] = 579784402;
assign addr[12739] = 598173833;
assign addr[12740] = 616515832;
assign addr[12741] = 634808946;
assign addr[12742] = 653051723;
assign addr[12743] = 671242716;
assign addr[12744] = 689380485;
assign addr[12745] = 707463589;
assign addr[12746] = 725490597;
assign addr[12747] = 743460077;
assign addr[12748] = 761370605;
assign addr[12749] = 779220762;
assign addr[12750] = 797009130;
assign addr[12751] = 814734301;
assign addr[12752] = 832394869;
assign addr[12753] = 849989433;
assign addr[12754] = 867516597;
assign addr[12755] = 884974973;
assign addr[12756] = 902363176;
assign addr[12757] = 919679827;
assign addr[12758] = 936923553;
assign addr[12759] = 954092986;
assign addr[12760] = 971186766;
assign addr[12761] = 988203537;
assign addr[12762] = 1005141949;
assign addr[12763] = 1022000660;
assign addr[12764] = 1038778332;
assign addr[12765] = 1055473635;
assign addr[12766] = 1072085246;
assign addr[12767] = 1088611847;
assign addr[12768] = 1105052128;
assign addr[12769] = 1121404785;
assign addr[12770] = 1137668521;
assign addr[12771] = 1153842047;
assign addr[12772] = 1169924081;
assign addr[12773] = 1185913346;
assign addr[12774] = 1201808576;
assign addr[12775] = 1217608510;
assign addr[12776] = 1233311895;
assign addr[12777] = 1248917486;
assign addr[12778] = 1264424045;
assign addr[12779] = 1279830344;
assign addr[12780] = 1295135159;
assign addr[12781] = 1310337279;
assign addr[12782] = 1325435496;
assign addr[12783] = 1340428615;
assign addr[12784] = 1355315445;
assign addr[12785] = 1370094808;
assign addr[12786] = 1384765530;
assign addr[12787] = 1399326449;
assign addr[12788] = 1413776410;
assign addr[12789] = 1428114267;
assign addr[12790] = 1442338884;
assign addr[12791] = 1456449131;
assign addr[12792] = 1470443891;
assign addr[12793] = 1484322054;
assign addr[12794] = 1498082520;
assign addr[12795] = 1511724196;
assign addr[12796] = 1525246002;
assign addr[12797] = 1538646865;
assign addr[12798] = 1551925723;
assign addr[12799] = 1565081523;
assign addr[12800] = 1578113222;
assign addr[12801] = 1591019785;
assign addr[12802] = 1603800191;
assign addr[12803] = 1616453425;
assign addr[12804] = 1628978484;
assign addr[12805] = 1641374375;
assign addr[12806] = 1653640115;
assign addr[12807] = 1665774731;
assign addr[12808] = 1677777262;
assign addr[12809] = 1689646755;
assign addr[12810] = 1701382270;
assign addr[12811] = 1712982875;
assign addr[12812] = 1724447652;
assign addr[12813] = 1735775690;
assign addr[12814] = 1746966091;
assign addr[12815] = 1758017969;
assign addr[12816] = 1768930447;
assign addr[12817] = 1779702660;
assign addr[12818] = 1790333753;
assign addr[12819] = 1800822883;
assign addr[12820] = 1811169220;
assign addr[12821] = 1821371941;
assign addr[12822] = 1831430239;
assign addr[12823] = 1841343316;
assign addr[12824] = 1851110385;
assign addr[12825] = 1860730673;
assign addr[12826] = 1870203416;
assign addr[12827] = 1879527863;
assign addr[12828] = 1888703276;
assign addr[12829] = 1897728925;
assign addr[12830] = 1906604097;
assign addr[12831] = 1915328086;
assign addr[12832] = 1923900201;
assign addr[12833] = 1932319763;
assign addr[12834] = 1940586104;
assign addr[12835] = 1948698568;
assign addr[12836] = 1956656513;
assign addr[12837] = 1964459306;
assign addr[12838] = 1972106330;
assign addr[12839] = 1979596978;
assign addr[12840] = 1986930656;
assign addr[12841] = 1994106782;
assign addr[12842] = 2001124788;
assign addr[12843] = 2007984117;
assign addr[12844] = 2014684225;
assign addr[12845] = 2021224581;
assign addr[12846] = 2027604666;
assign addr[12847] = 2033823974;
assign addr[12848] = 2039882013;
assign addr[12849] = 2045778302;
assign addr[12850] = 2051512372;
assign addr[12851] = 2057083771;
assign addr[12852] = 2062492055;
assign addr[12853] = 2067736796;
assign addr[12854] = 2072817579;
assign addr[12855] = 2077733999;
assign addr[12856] = 2082485668;
assign addr[12857] = 2087072209;
assign addr[12858] = 2091493257;
assign addr[12859] = 2095748463;
assign addr[12860] = 2099837489;
assign addr[12861] = 2103760010;
assign addr[12862] = 2107515716;
assign addr[12863] = 2111104309;
assign addr[12864] = 2114525505;
assign addr[12865] = 2117779031;
assign addr[12866] = 2120864631;
assign addr[12867] = 2123782059;
assign addr[12868] = 2126531084;
assign addr[12869] = 2129111488;
assign addr[12870] = 2131523066;
assign addr[12871] = 2133765628;
assign addr[12872] = 2135838995;
assign addr[12873] = 2137743003;
assign addr[12874] = 2139477502;
assign addr[12875] = 2141042352;
assign addr[12876] = 2142437431;
assign addr[12877] = 2143662628;
assign addr[12878] = 2144717846;
assign addr[12879] = 2145603001;
assign addr[12880] = 2146318022;
assign addr[12881] = 2146862854;
assign addr[12882] = 2147237452;
assign addr[12883] = 2147441787;
assign addr[12884] = 2147475844;
assign addr[12885] = 2147339619;
assign addr[12886] = 2147033123;
assign addr[12887] = 2146556380;
assign addr[12888] = 2145909429;
assign addr[12889] = 2145092320;
assign addr[12890] = 2144105118;
assign addr[12891] = 2142947902;
assign addr[12892] = 2141620763;
assign addr[12893] = 2140123807;
assign addr[12894] = 2138457152;
assign addr[12895] = 2136620930;
assign addr[12896] = 2134615288;
assign addr[12897] = 2132440383;
assign addr[12898] = 2130096389;
assign addr[12899] = 2127583492;
assign addr[12900] = 2124901890;
assign addr[12901] = 2122051796;
assign addr[12902] = 2119033436;
assign addr[12903] = 2115847050;
assign addr[12904] = 2112492891;
assign addr[12905] = 2108971223;
assign addr[12906] = 2105282327;
assign addr[12907] = 2101426496;
assign addr[12908] = 2097404033;
assign addr[12909] = 2093215260;
assign addr[12910] = 2088860507;
assign addr[12911] = 2084340120;
assign addr[12912] = 2079654458;
assign addr[12913] = 2074803892;
assign addr[12914] = 2069788807;
assign addr[12915] = 2064609600;
assign addr[12916] = 2059266683;
assign addr[12917] = 2053760478;
assign addr[12918] = 2048091422;
assign addr[12919] = 2042259965;
assign addr[12920] = 2036266570;
assign addr[12921] = 2030111710;
assign addr[12922] = 2023795876;
assign addr[12923] = 2017319567;
assign addr[12924] = 2010683297;
assign addr[12925] = 2003887591;
assign addr[12926] = 1996932990;
assign addr[12927] = 1989820044;
assign addr[12928] = 1982549318;
assign addr[12929] = 1975121388;
assign addr[12930] = 1967536842;
assign addr[12931] = 1959796283;
assign addr[12932] = 1951900324;
assign addr[12933] = 1943849591;
assign addr[12934] = 1935644723;
assign addr[12935] = 1927286370;
assign addr[12936] = 1918775195;
assign addr[12937] = 1910111873;
assign addr[12938] = 1901297091;
assign addr[12939] = 1892331547;
assign addr[12940] = 1883215953;
assign addr[12941] = 1873951032;
assign addr[12942] = 1864537518;
assign addr[12943] = 1854976157;
assign addr[12944] = 1845267708;
assign addr[12945] = 1835412941;
assign addr[12946] = 1825412636;
assign addr[12947] = 1815267588;
assign addr[12948] = 1804978599;
assign addr[12949] = 1794546487;
assign addr[12950] = 1783972079;
assign addr[12951] = 1773256212;
assign addr[12952] = 1762399737;
assign addr[12953] = 1751403515;
assign addr[12954] = 1740268417;
assign addr[12955] = 1728995326;
assign addr[12956] = 1717585136;
assign addr[12957] = 1706038753;
assign addr[12958] = 1694357091;
assign addr[12959] = 1682541077;
assign addr[12960] = 1670591647;
assign addr[12961] = 1658509750;
assign addr[12962] = 1646296344;
assign addr[12963] = 1633952396;
assign addr[12964] = 1621478885;
assign addr[12965] = 1608876801;
assign addr[12966] = 1596147143;
assign addr[12967] = 1583290921;
assign addr[12968] = 1570309153;
assign addr[12969] = 1557202869;
assign addr[12970] = 1543973108;
assign addr[12971] = 1530620920;
assign addr[12972] = 1517147363;
assign addr[12973] = 1503553506;
assign addr[12974] = 1489840425;
assign addr[12975] = 1476009210;
assign addr[12976] = 1462060956;
assign addr[12977] = 1447996770;
assign addr[12978] = 1433817766;
assign addr[12979] = 1419525069;
assign addr[12980] = 1405119813;
assign addr[12981] = 1390603139;
assign addr[12982] = 1375976199;
assign addr[12983] = 1361240152;
assign addr[12984] = 1346396168;
assign addr[12985] = 1331445422;
assign addr[12986] = 1316389101;
assign addr[12987] = 1301228398;
assign addr[12988] = 1285964516;
assign addr[12989] = 1270598665;
assign addr[12990] = 1255132063;
assign addr[12991] = 1239565936;
assign addr[12992] = 1223901520;
assign addr[12993] = 1208140056;
assign addr[12994] = 1192282793;
assign addr[12995] = 1176330990;
assign addr[12996] = 1160285911;
assign addr[12997] = 1144148829;
assign addr[12998] = 1127921022;
assign addr[12999] = 1111603778;
assign addr[13000] = 1095198391;
assign addr[13001] = 1078706161;
assign addr[13002] = 1062128397;
assign addr[13003] = 1045466412;
assign addr[13004] = 1028721528;
assign addr[13005] = 1011895073;
assign addr[13006] = 994988380;
assign addr[13007] = 978002791;
assign addr[13008] = 960939653;
assign addr[13009] = 943800318;
assign addr[13010] = 926586145;
assign addr[13011] = 909298500;
assign addr[13012] = 891938752;
assign addr[13013] = 874508280;
assign addr[13014] = 857008464;
assign addr[13015] = 839440693;
assign addr[13016] = 821806359;
assign addr[13017] = 804106861;
assign addr[13018] = 786343603;
assign addr[13019] = 768517992;
assign addr[13020] = 750631442;
assign addr[13021] = 732685372;
assign addr[13022] = 714681204;
assign addr[13023] = 696620367;
assign addr[13024] = 678504291;
assign addr[13025] = 660334415;
assign addr[13026] = 642112178;
assign addr[13027] = 623839025;
assign addr[13028] = 605516406;
assign addr[13029] = 587145773;
assign addr[13030] = 568728583;
assign addr[13031] = 550266296;
assign addr[13032] = 531760377;
assign addr[13033] = 513212292;
assign addr[13034] = 494623513;
assign addr[13035] = 475995513;
assign addr[13036] = 457329769;
assign addr[13037] = 438627762;
assign addr[13038] = 419890975;
assign addr[13039] = 401120892;
assign addr[13040] = 382319004;
assign addr[13041] = 363486799;
assign addr[13042] = 344625773;
assign addr[13043] = 325737419;
assign addr[13044] = 306823237;
assign addr[13045] = 287884725;
assign addr[13046] = 268923386;
assign addr[13047] = 249940723;
assign addr[13048] = 230938242;
assign addr[13049] = 211917448;
assign addr[13050] = 192879850;
assign addr[13051] = 173826959;
assign addr[13052] = 154760284;
assign addr[13053] = 135681337;
assign addr[13054] = 116591632;
assign addr[13055] = 97492681;
assign addr[13056] = 78386000;
assign addr[13057] = 59273104;
assign addr[13058] = 40155507;
assign addr[13059] = 21034727;
assign addr[13060] = 1912278;
assign addr[13061] = -17210322;
assign addr[13062] = -36331557;
assign addr[13063] = -55449912;
assign addr[13064] = -74563870;
assign addr[13065] = -93671915;
assign addr[13066] = -112772533;
assign addr[13067] = -131864208;
assign addr[13068] = -150945428;
assign addr[13069] = -170014678;
assign addr[13070] = -189070447;
assign addr[13071] = -208111224;
assign addr[13072] = -227135500;
assign addr[13073] = -246141764;
assign addr[13074] = -265128512;
assign addr[13075] = -284094236;
assign addr[13076] = -303037433;
assign addr[13077] = -321956601;
assign addr[13078] = -340850240;
assign addr[13079] = -359716852;
assign addr[13080] = -378554940;
assign addr[13081] = -397363011;
assign addr[13082] = -416139574;
assign addr[13083] = -434883140;
assign addr[13084] = -453592221;
assign addr[13085] = -472265336;
assign addr[13086] = -490901003;
assign addr[13087] = -509497745;
assign addr[13088] = -528054086;
assign addr[13089] = -546568556;
assign addr[13090] = -565039687;
assign addr[13091] = -583466013;
assign addr[13092] = -601846074;
assign addr[13093] = -620178412;
assign addr[13094] = -638461574;
assign addr[13095] = -656694110;
assign addr[13096] = -674874574;
assign addr[13097] = -693001525;
assign addr[13098] = -711073524;
assign addr[13099] = -729089140;
assign addr[13100] = -747046944;
assign addr[13101] = -764945512;
assign addr[13102] = -782783424;
assign addr[13103] = -800559266;
assign addr[13104] = -818271628;
assign addr[13105] = -835919107;
assign addr[13106] = -853500302;
assign addr[13107] = -871013820;
assign addr[13108] = -888458272;
assign addr[13109] = -905832274;
assign addr[13110] = -923134450;
assign addr[13111] = -940363427;
assign addr[13112] = -957517838;
assign addr[13113] = -974596324;
assign addr[13114] = -991597531;
assign addr[13115] = -1008520110;
assign addr[13116] = -1025362720;
assign addr[13117] = -1042124025;
assign addr[13118] = -1058802695;
assign addr[13119] = -1075397409;
assign addr[13120] = -1091906851;
assign addr[13121] = -1108329711;
assign addr[13122] = -1124664687;
assign addr[13123] = -1140910484;
assign addr[13124] = -1157065814;
assign addr[13125] = -1173129396;
assign addr[13126] = -1189099956;
assign addr[13127] = -1204976227;
assign addr[13128] = -1220756951;
assign addr[13129] = -1236440877;
assign addr[13130] = -1252026760;
assign addr[13131] = -1267513365;
assign addr[13132] = -1282899464;
assign addr[13133] = -1298183838;
assign addr[13134] = -1313365273;
assign addr[13135] = -1328442566;
assign addr[13136] = -1343414522;
assign addr[13137] = -1358279953;
assign addr[13138] = -1373037681;
assign addr[13139] = -1387686535;
assign addr[13140] = -1402225355;
assign addr[13141] = -1416652986;
assign addr[13142] = -1430968286;
assign addr[13143] = -1445170118;
assign addr[13144] = -1459257358;
assign addr[13145] = -1473228887;
assign addr[13146] = -1487083598;
assign addr[13147] = -1500820393;
assign addr[13148] = -1514438181;
assign addr[13149] = -1527935884;
assign addr[13150] = -1541312431;
assign addr[13151] = -1554566762;
assign addr[13152] = -1567697824;
assign addr[13153] = -1580704578;
assign addr[13154] = -1593585992;
assign addr[13155] = -1606341043;
assign addr[13156] = -1618968722;
assign addr[13157] = -1631468027;
assign addr[13158] = -1643837966;
assign addr[13159] = -1656077559;
assign addr[13160] = -1668185835;
assign addr[13161] = -1680161834;
assign addr[13162] = -1692004606;
assign addr[13163] = -1703713213;
assign addr[13164] = -1715286726;
assign addr[13165] = -1726724227;
assign addr[13166] = -1738024810;
assign addr[13167] = -1749187577;
assign addr[13168] = -1760211645;
assign addr[13169] = -1771096139;
assign addr[13170] = -1781840195;
assign addr[13171] = -1792442963;
assign addr[13172] = -1802903601;
assign addr[13173] = -1813221279;
assign addr[13174] = -1823395180;
assign addr[13175] = -1833424497;
assign addr[13176] = -1843308435;
assign addr[13177] = -1853046210;
assign addr[13178] = -1862637049;
assign addr[13179] = -1872080193;
assign addr[13180] = -1881374892;
assign addr[13181] = -1890520410;
assign addr[13182] = -1899516021;
assign addr[13183] = -1908361011;
assign addr[13184] = -1917054681;
assign addr[13185] = -1925596340;
assign addr[13186] = -1933985310;
assign addr[13187] = -1942220928;
assign addr[13188] = -1950302539;
assign addr[13189] = -1958229503;
assign addr[13190] = -1966001192;
assign addr[13191] = -1973616989;
assign addr[13192] = -1981076290;
assign addr[13193] = -1988378503;
assign addr[13194] = -1995523051;
assign addr[13195] = -2002509365;
assign addr[13196] = -2009336893;
assign addr[13197] = -2016005093;
assign addr[13198] = -2022513436;
assign addr[13199] = -2028861406;
assign addr[13200] = -2035048499;
assign addr[13201] = -2041074226;
assign addr[13202] = -2046938108;
assign addr[13203] = -2052639680;
assign addr[13204] = -2058178491;
assign addr[13205] = -2063554100;
assign addr[13206] = -2068766083;
assign addr[13207] = -2073814024;
assign addr[13208] = -2078697525;
assign addr[13209] = -2083416198;
assign addr[13210] = -2087969669;
assign addr[13211] = -2092357577;
assign addr[13212] = -2096579573;
assign addr[13213] = -2100635323;
assign addr[13214] = -2104524506;
assign addr[13215] = -2108246813;
assign addr[13216] = -2111801949;
assign addr[13217] = -2115189632;
assign addr[13218] = -2118409593;
assign addr[13219] = -2121461578;
assign addr[13220] = -2124345343;
assign addr[13221] = -2127060661;
assign addr[13222] = -2129607316;
assign addr[13223] = -2131985106;
assign addr[13224] = -2134193842;
assign addr[13225] = -2136233350;
assign addr[13226] = -2138103468;
assign addr[13227] = -2139804048;
assign addr[13228] = -2141334954;
assign addr[13229] = -2142696065;
assign addr[13230] = -2143887273;
assign addr[13231] = -2144908484;
assign addr[13232] = -2145759618;
assign addr[13233] = -2146440605;
assign addr[13234] = -2146951393;
assign addr[13235] = -2147291941;
assign addr[13236] = -2147462221;
assign addr[13237] = -2147462221;
assign addr[13238] = -2147291941;
assign addr[13239] = -2146951393;
assign addr[13240] = -2146440605;
assign addr[13241] = -2145759618;
assign addr[13242] = -2144908484;
assign addr[13243] = -2143887273;
assign addr[13244] = -2142696065;
assign addr[13245] = -2141334954;
assign addr[13246] = -2139804048;
assign addr[13247] = -2138103468;
assign addr[13248] = -2136233350;
assign addr[13249] = -2134193842;
assign addr[13250] = -2131985106;
assign addr[13251] = -2129607316;
assign addr[13252] = -2127060661;
assign addr[13253] = -2124345343;
assign addr[13254] = -2121461578;
assign addr[13255] = -2118409593;
assign addr[13256] = -2115189632;
assign addr[13257] = -2111801949;
assign addr[13258] = -2108246813;
assign addr[13259] = -2104524506;
assign addr[13260] = -2100635323;
assign addr[13261] = -2096579573;
assign addr[13262] = -2092357577;
assign addr[13263] = -2087969669;
assign addr[13264] = -2083416198;
assign addr[13265] = -2078697525;
assign addr[13266] = -2073814024;
assign addr[13267] = -2068766083;
assign addr[13268] = -2063554100;
assign addr[13269] = -2058178491;
assign addr[13270] = -2052639680;
assign addr[13271] = -2046938108;
assign addr[13272] = -2041074226;
assign addr[13273] = -2035048499;
assign addr[13274] = -2028861406;
assign addr[13275] = -2022513436;
assign addr[13276] = -2016005093;
assign addr[13277] = -2009336893;
assign addr[13278] = -2002509365;
assign addr[13279] = -1995523051;
assign addr[13280] = -1988378503;
assign addr[13281] = -1981076290;
assign addr[13282] = -1973616989;
assign addr[13283] = -1966001192;
assign addr[13284] = -1958229503;
assign addr[13285] = -1950302539;
assign addr[13286] = -1942220928;
assign addr[13287] = -1933985310;
assign addr[13288] = -1925596340;
assign addr[13289] = -1917054681;
assign addr[13290] = -1908361011;
assign addr[13291] = -1899516021;
assign addr[13292] = -1890520410;
assign addr[13293] = -1881374892;
assign addr[13294] = -1872080193;
assign addr[13295] = -1862637049;
assign addr[13296] = -1853046210;
assign addr[13297] = -1843308435;
assign addr[13298] = -1833424497;
assign addr[13299] = -1823395180;
assign addr[13300] = -1813221279;
assign addr[13301] = -1802903601;
assign addr[13302] = -1792442963;
assign addr[13303] = -1781840195;
assign addr[13304] = -1771096139;
assign addr[13305] = -1760211645;
assign addr[13306] = -1749187577;
assign addr[13307] = -1738024810;
assign addr[13308] = -1726724227;
assign addr[13309] = -1715286726;
assign addr[13310] = -1703713213;
assign addr[13311] = -1692004606;
assign addr[13312] = -1680161834;
assign addr[13313] = -1668185835;
assign addr[13314] = -1656077559;
assign addr[13315] = -1643837966;
assign addr[13316] = -1631468027;
assign addr[13317] = -1618968722;
assign addr[13318] = -1606341043;
assign addr[13319] = -1593585992;
assign addr[13320] = -1580704578;
assign addr[13321] = -1567697824;
assign addr[13322] = -1554566762;
assign addr[13323] = -1541312431;
assign addr[13324] = -1527935884;
assign addr[13325] = -1514438181;
assign addr[13326] = -1500820393;
assign addr[13327] = -1487083598;
assign addr[13328] = -1473228887;
assign addr[13329] = -1459257358;
assign addr[13330] = -1445170118;
assign addr[13331] = -1430968286;
assign addr[13332] = -1416652986;
assign addr[13333] = -1402225355;
assign addr[13334] = -1387686535;
assign addr[13335] = -1373037681;
assign addr[13336] = -1358279953;
assign addr[13337] = -1343414522;
assign addr[13338] = -1328442566;
assign addr[13339] = -1313365273;
assign addr[13340] = -1298183838;
assign addr[13341] = -1282899464;
assign addr[13342] = -1267513365;
assign addr[13343] = -1252026760;
assign addr[13344] = -1236440877;
assign addr[13345] = -1220756951;
assign addr[13346] = -1204976227;
assign addr[13347] = -1189099956;
assign addr[13348] = -1173129396;
assign addr[13349] = -1157065814;
assign addr[13350] = -1140910484;
assign addr[13351] = -1124664687;
assign addr[13352] = -1108329711;
assign addr[13353] = -1091906851;
assign addr[13354] = -1075397409;
assign addr[13355] = -1058802695;
assign addr[13356] = -1042124025;
assign addr[13357] = -1025362720;
assign addr[13358] = -1008520110;
assign addr[13359] = -991597531;
assign addr[13360] = -974596324;
assign addr[13361] = -957517838;
assign addr[13362] = -940363427;
assign addr[13363] = -923134450;
assign addr[13364] = -905832274;
assign addr[13365] = -888458272;
assign addr[13366] = -871013820;
assign addr[13367] = -853500302;
assign addr[13368] = -835919107;
assign addr[13369] = -818271628;
assign addr[13370] = -800559266;
assign addr[13371] = -782783424;
assign addr[13372] = -764945512;
assign addr[13373] = -747046944;
assign addr[13374] = -729089140;
assign addr[13375] = -711073524;
assign addr[13376] = -693001525;
assign addr[13377] = -674874574;
assign addr[13378] = -656694110;
assign addr[13379] = -638461574;
assign addr[13380] = -620178412;
assign addr[13381] = -601846074;
assign addr[13382] = -583466013;
assign addr[13383] = -565039687;
assign addr[13384] = -546568556;
assign addr[13385] = -528054086;
assign addr[13386] = -509497745;
assign addr[13387] = -490901003;
assign addr[13388] = -472265336;
assign addr[13389] = -453592221;
assign addr[13390] = -434883140;
assign addr[13391] = -416139574;
assign addr[13392] = -397363011;
assign addr[13393] = -378554940;
assign addr[13394] = -359716852;
assign addr[13395] = -340850240;
assign addr[13396] = -321956601;
assign addr[13397] = -303037433;
assign addr[13398] = -284094236;
assign addr[13399] = -265128512;
assign addr[13400] = -246141764;
assign addr[13401] = -227135500;
assign addr[13402] = -208111224;
assign addr[13403] = -189070447;
assign addr[13404] = -170014678;
assign addr[13405] = -150945428;
assign addr[13406] = -131864208;
assign addr[13407] = -112772533;
assign addr[13408] = -93671915;
assign addr[13409] = -74563870;
assign addr[13410] = -55449912;
assign addr[13411] = -36331557;
assign addr[13412] = -17210322;
assign addr[13413] = 1912278;
assign addr[13414] = 21034727;
assign addr[13415] = 40155507;
assign addr[13416] = 59273104;
assign addr[13417] = 78386000;
assign addr[13418] = 97492681;
assign addr[13419] = 116591632;
assign addr[13420] = 135681337;
assign addr[13421] = 154760284;
assign addr[13422] = 173826959;
assign addr[13423] = 192879850;
assign addr[13424] = 211917448;
assign addr[13425] = 230938242;
assign addr[13426] = 249940723;
assign addr[13427] = 268923386;
assign addr[13428] = 287884725;
assign addr[13429] = 306823237;
assign addr[13430] = 325737419;
assign addr[13431] = 344625773;
assign addr[13432] = 363486799;
assign addr[13433] = 382319004;
assign addr[13434] = 401120892;
assign addr[13435] = 419890975;
assign addr[13436] = 438627762;
assign addr[13437] = 457329769;
assign addr[13438] = 475995513;
assign addr[13439] = 494623513;
assign addr[13440] = 513212292;
assign addr[13441] = 531760377;
assign addr[13442] = 550266296;
assign addr[13443] = 568728583;
assign addr[13444] = 587145773;
assign addr[13445] = 605516406;
assign addr[13446] = 623839025;
assign addr[13447] = 642112178;
assign addr[13448] = 660334415;
assign addr[13449] = 678504291;
assign addr[13450] = 696620367;
assign addr[13451] = 714681204;
assign addr[13452] = 732685372;
assign addr[13453] = 750631442;
assign addr[13454] = 768517992;
assign addr[13455] = 786343603;
assign addr[13456] = 804106861;
assign addr[13457] = 821806359;
assign addr[13458] = 839440693;
assign addr[13459] = 857008464;
assign addr[13460] = 874508280;
assign addr[13461] = 891938752;
assign addr[13462] = 909298500;
assign addr[13463] = 926586145;
assign addr[13464] = 943800318;
assign addr[13465] = 960939653;
assign addr[13466] = 978002791;
assign addr[13467] = 994988380;
assign addr[13468] = 1011895073;
assign addr[13469] = 1028721528;
assign addr[13470] = 1045466412;
assign addr[13471] = 1062128397;
assign addr[13472] = 1078706161;
assign addr[13473] = 1095198391;
assign addr[13474] = 1111603778;
assign addr[13475] = 1127921022;
assign addr[13476] = 1144148829;
assign addr[13477] = 1160285911;
assign addr[13478] = 1176330990;
assign addr[13479] = 1192282793;
assign addr[13480] = 1208140056;
assign addr[13481] = 1223901520;
assign addr[13482] = 1239565936;
assign addr[13483] = 1255132063;
assign addr[13484] = 1270598665;
assign addr[13485] = 1285964516;
assign addr[13486] = 1301228398;
assign addr[13487] = 1316389101;
assign addr[13488] = 1331445422;
assign addr[13489] = 1346396168;
assign addr[13490] = 1361240152;
assign addr[13491] = 1375976199;
assign addr[13492] = 1390603139;
assign addr[13493] = 1405119813;
assign addr[13494] = 1419525069;
assign addr[13495] = 1433817766;
assign addr[13496] = 1447996770;
assign addr[13497] = 1462060956;
assign addr[13498] = 1476009210;
assign addr[13499] = 1489840425;
assign addr[13500] = 1503553506;
assign addr[13501] = 1517147363;
assign addr[13502] = 1530620920;
assign addr[13503] = 1543973108;
assign addr[13504] = 1557202869;
assign addr[13505] = 1570309153;
assign addr[13506] = 1583290921;
assign addr[13507] = 1596147143;
assign addr[13508] = 1608876801;
assign addr[13509] = 1621478885;
assign addr[13510] = 1633952396;
assign addr[13511] = 1646296344;
assign addr[13512] = 1658509750;
assign addr[13513] = 1670591647;
assign addr[13514] = 1682541077;
assign addr[13515] = 1694357091;
assign addr[13516] = 1706038753;
assign addr[13517] = 1717585136;
assign addr[13518] = 1728995326;
assign addr[13519] = 1740268417;
assign addr[13520] = 1751403515;
assign addr[13521] = 1762399737;
assign addr[13522] = 1773256212;
assign addr[13523] = 1783972079;
assign addr[13524] = 1794546487;
assign addr[13525] = 1804978599;
assign addr[13526] = 1815267588;
assign addr[13527] = 1825412636;
assign addr[13528] = 1835412941;
assign addr[13529] = 1845267708;
assign addr[13530] = 1854976157;
assign addr[13531] = 1864537518;
assign addr[13532] = 1873951032;
assign addr[13533] = 1883215953;
assign addr[13534] = 1892331547;
assign addr[13535] = 1901297091;
assign addr[13536] = 1910111873;
assign addr[13537] = 1918775195;
assign addr[13538] = 1927286370;
assign addr[13539] = 1935644723;
assign addr[13540] = 1943849591;
assign addr[13541] = 1951900324;
assign addr[13542] = 1959796283;
assign addr[13543] = 1967536842;
assign addr[13544] = 1975121388;
assign addr[13545] = 1982549318;
assign addr[13546] = 1989820044;
assign addr[13547] = 1996932990;
assign addr[13548] = 2003887591;
assign addr[13549] = 2010683297;
assign addr[13550] = 2017319567;
assign addr[13551] = 2023795876;
assign addr[13552] = 2030111710;
assign addr[13553] = 2036266570;
assign addr[13554] = 2042259965;
assign addr[13555] = 2048091422;
assign addr[13556] = 2053760478;
assign addr[13557] = 2059266683;
assign addr[13558] = 2064609600;
assign addr[13559] = 2069788807;
assign addr[13560] = 2074803892;
assign addr[13561] = 2079654458;
assign addr[13562] = 2084340120;
assign addr[13563] = 2088860507;
assign addr[13564] = 2093215260;
assign addr[13565] = 2097404033;
assign addr[13566] = 2101426496;
assign addr[13567] = 2105282327;
assign addr[13568] = 2108971223;
assign addr[13569] = 2112492891;
assign addr[13570] = 2115847050;
assign addr[13571] = 2119033436;
assign addr[13572] = 2122051796;
assign addr[13573] = 2124901890;
assign addr[13574] = 2127583492;
assign addr[13575] = 2130096389;
assign addr[13576] = 2132440383;
assign addr[13577] = 2134615288;
assign addr[13578] = 2136620930;
assign addr[13579] = 2138457152;
assign addr[13580] = 2140123807;
assign addr[13581] = 2141620763;
assign addr[13582] = 2142947902;
assign addr[13583] = 2144105118;
assign addr[13584] = 2145092320;
assign addr[13585] = 2145909429;
assign addr[13586] = 2146556380;
assign addr[13587] = 2147033123;
assign addr[13588] = 2147339619;
assign addr[13589] = 2147475844;
assign addr[13590] = 2147441787;
assign addr[13591] = 2147237452;
assign addr[13592] = 2146862854;
assign addr[13593] = 2146318022;
assign addr[13594] = 2145603001;
assign addr[13595] = 2144717846;
assign addr[13596] = 2143662628;
assign addr[13597] = 2142437431;
assign addr[13598] = 2141042352;
assign addr[13599] = 2139477502;
assign addr[13600] = 2137743003;
assign addr[13601] = 2135838995;
assign addr[13602] = 2133765628;
assign addr[13603] = 2131523066;
assign addr[13604] = 2129111488;
assign addr[13605] = 2126531084;
assign addr[13606] = 2123782059;
assign addr[13607] = 2120864631;
assign addr[13608] = 2117779031;
assign addr[13609] = 2114525505;
assign addr[13610] = 2111104309;
assign addr[13611] = 2107515716;
assign addr[13612] = 2103760010;
assign addr[13613] = 2099837489;
assign addr[13614] = 2095748463;
assign addr[13615] = 2091493257;
assign addr[13616] = 2087072209;
assign addr[13617] = 2082485668;
assign addr[13618] = 2077733999;
assign addr[13619] = 2072817579;
assign addr[13620] = 2067736796;
assign addr[13621] = 2062492055;
assign addr[13622] = 2057083771;
assign addr[13623] = 2051512372;
assign addr[13624] = 2045778302;
assign addr[13625] = 2039882013;
assign addr[13626] = 2033823974;
assign addr[13627] = 2027604666;
assign addr[13628] = 2021224581;
assign addr[13629] = 2014684225;
assign addr[13630] = 2007984117;
assign addr[13631] = 2001124788;
assign addr[13632] = 1994106782;
assign addr[13633] = 1986930656;
assign addr[13634] = 1979596978;
assign addr[13635] = 1972106330;
assign addr[13636] = 1964459306;
assign addr[13637] = 1956656513;
assign addr[13638] = 1948698568;
assign addr[13639] = 1940586104;
assign addr[13640] = 1932319763;
assign addr[13641] = 1923900201;
assign addr[13642] = 1915328086;
assign addr[13643] = 1906604097;
assign addr[13644] = 1897728925;
assign addr[13645] = 1888703276;
assign addr[13646] = 1879527863;
assign addr[13647] = 1870203416;
assign addr[13648] = 1860730673;
assign addr[13649] = 1851110385;
assign addr[13650] = 1841343316;
assign addr[13651] = 1831430239;
assign addr[13652] = 1821371941;
assign addr[13653] = 1811169220;
assign addr[13654] = 1800822883;
assign addr[13655] = 1790333753;
assign addr[13656] = 1779702660;
assign addr[13657] = 1768930447;
assign addr[13658] = 1758017969;
assign addr[13659] = 1746966091;
assign addr[13660] = 1735775690;
assign addr[13661] = 1724447652;
assign addr[13662] = 1712982875;
assign addr[13663] = 1701382270;
assign addr[13664] = 1689646755;
assign addr[13665] = 1677777262;
assign addr[13666] = 1665774731;
assign addr[13667] = 1653640115;
assign addr[13668] = 1641374375;
assign addr[13669] = 1628978484;
assign addr[13670] = 1616453425;
assign addr[13671] = 1603800191;
assign addr[13672] = 1591019785;
assign addr[13673] = 1578113222;
assign addr[13674] = 1565081523;
assign addr[13675] = 1551925723;
assign addr[13676] = 1538646865;
assign addr[13677] = 1525246002;
assign addr[13678] = 1511724196;
assign addr[13679] = 1498082520;
assign addr[13680] = 1484322054;
assign addr[13681] = 1470443891;
assign addr[13682] = 1456449131;
assign addr[13683] = 1442338884;
assign addr[13684] = 1428114267;
assign addr[13685] = 1413776410;
assign addr[13686] = 1399326449;
assign addr[13687] = 1384765530;
assign addr[13688] = 1370094808;
assign addr[13689] = 1355315445;
assign addr[13690] = 1340428615;
assign addr[13691] = 1325435496;
assign addr[13692] = 1310337279;
assign addr[13693] = 1295135159;
assign addr[13694] = 1279830344;
assign addr[13695] = 1264424045;
assign addr[13696] = 1248917486;
assign addr[13697] = 1233311895;
assign addr[13698] = 1217608510;
assign addr[13699] = 1201808576;
assign addr[13700] = 1185913346;
assign addr[13701] = 1169924081;
assign addr[13702] = 1153842047;
assign addr[13703] = 1137668521;
assign addr[13704] = 1121404785;
assign addr[13705] = 1105052128;
assign addr[13706] = 1088611847;
assign addr[13707] = 1072085246;
assign addr[13708] = 1055473635;
assign addr[13709] = 1038778332;
assign addr[13710] = 1022000660;
assign addr[13711] = 1005141949;
assign addr[13712] = 988203537;
assign addr[13713] = 971186766;
assign addr[13714] = 954092986;
assign addr[13715] = 936923553;
assign addr[13716] = 919679827;
assign addr[13717] = 902363176;
assign addr[13718] = 884974973;
assign addr[13719] = 867516597;
assign addr[13720] = 849989433;
assign addr[13721] = 832394869;
assign addr[13722] = 814734301;
assign addr[13723] = 797009130;
assign addr[13724] = 779220762;
assign addr[13725] = 761370605;
assign addr[13726] = 743460077;
assign addr[13727] = 725490597;
assign addr[13728] = 707463589;
assign addr[13729] = 689380485;
assign addr[13730] = 671242716;
assign addr[13731] = 653051723;
assign addr[13732] = 634808946;
assign addr[13733] = 616515832;
assign addr[13734] = 598173833;
assign addr[13735] = 579784402;
assign addr[13736] = 561348998;
assign addr[13737] = 542869083;
assign addr[13738] = 524346121;
assign addr[13739] = 505781581;
assign addr[13740] = 487176937;
assign addr[13741] = 468533662;
assign addr[13742] = 449853235;
assign addr[13743] = 431137138;
assign addr[13744] = 412386854;
assign addr[13745] = 393603870;
assign addr[13746] = 374789676;
assign addr[13747] = 355945764;
assign addr[13748] = 337073627;
assign addr[13749] = 318174762;
assign addr[13750] = 299250668;
assign addr[13751] = 280302845;
assign addr[13752] = 261332796;
assign addr[13753] = 242342025;
assign addr[13754] = 223332037;
assign addr[13755] = 204304341;
assign addr[13756] = 185260444;
assign addr[13757] = 166201858;
assign addr[13758] = 147130093;
assign addr[13759] = 128046661;
assign addr[13760] = 108953076;
assign addr[13761] = 89850852;
assign addr[13762] = 70741503;
assign addr[13763] = 51626544;
assign addr[13764] = 32507492;
assign addr[13765] = 13385863;
assign addr[13766] = -5736829;
assign addr[13767] = -24859065;
assign addr[13768] = -43979330;
assign addr[13769] = -63096108;
assign addr[13770] = -82207882;
assign addr[13771] = -101313138;
assign addr[13772] = -120410361;
assign addr[13773] = -139498035;
assign addr[13774] = -158574649;
assign addr[13775] = -177638688;
assign addr[13776] = -196688642;
assign addr[13777] = -215722999;
assign addr[13778] = -234740251;
assign addr[13779] = -253738890;
assign addr[13780] = -272717408;
assign addr[13781] = -291674302;
assign addr[13782] = -310608068;
assign addr[13783] = -329517204;
assign addr[13784] = -348400212;
assign addr[13785] = -367255594;
assign addr[13786] = -386081854;
assign addr[13787] = -404877501;
assign addr[13788] = -423641043;
assign addr[13789] = -442370993;
assign addr[13790] = -461065866;
assign addr[13791] = -479724180;
assign addr[13792] = -498344454;
assign addr[13793] = -516925212;
assign addr[13794] = -535464981;
assign addr[13795] = -553962291;
assign addr[13796] = -572415676;
assign addr[13797] = -590823671;
assign addr[13798] = -609184818;
assign addr[13799] = -627497660;
assign addr[13800] = -645760745;
assign addr[13801] = -663972625;
assign addr[13802] = -682131857;
assign addr[13803] = -700236999;
assign addr[13804] = -718286617;
assign addr[13805] = -736279279;
assign addr[13806] = -754213559;
assign addr[13807] = -772088034;
assign addr[13808] = -789901288;
assign addr[13809] = -807651907;
assign addr[13810] = -825338484;
assign addr[13811] = -842959617;
assign addr[13812] = -860513908;
assign addr[13813] = -877999966;
assign addr[13814] = -895416404;
assign addr[13815] = -912761841;
assign addr[13816] = -930034901;
assign addr[13817] = -947234215;
assign addr[13818] = -964358420;
assign addr[13819] = -981406156;
assign addr[13820] = -998376073;
assign addr[13821] = -1015266825;
assign addr[13822] = -1032077073;
assign addr[13823] = -1048805483;
assign addr[13824] = -1065450729;
assign addr[13825] = -1082011492;
assign addr[13826] = -1098486458;
assign addr[13827] = -1114874320;
assign addr[13828] = -1131173780;
assign addr[13829] = -1147383544;
assign addr[13830] = -1163502328;
assign addr[13831] = -1179528853;
assign addr[13832] = -1195461849;
assign addr[13833] = -1211300053;
assign addr[13834] = -1227042207;
assign addr[13835] = -1242687064;
assign addr[13836] = -1258233384;
assign addr[13837] = -1273679934;
assign addr[13838] = -1289025489;
assign addr[13839] = -1304268832;
assign addr[13840] = -1319408754;
assign addr[13841] = -1334444055;
assign addr[13842] = -1349373543;
assign addr[13843] = -1364196034;
assign addr[13844] = -1378910353;
assign addr[13845] = -1393515332;
assign addr[13846] = -1408009814;
assign addr[13847] = -1422392650;
assign addr[13848] = -1436662698;
assign addr[13849] = -1450818828;
assign addr[13850] = -1464859917;
assign addr[13851] = -1478784851;
assign addr[13852] = -1492592527;
assign addr[13853] = -1506281850;
assign addr[13854] = -1519851733;
assign addr[13855] = -1533301101;
assign addr[13856] = -1546628888;
assign addr[13857] = -1559834037;
assign addr[13858] = -1572915501;
assign addr[13859] = -1585872242;
assign addr[13860] = -1598703233;
assign addr[13861] = -1611407456;
assign addr[13862] = -1623983905;
assign addr[13863] = -1636431582;
assign addr[13864] = -1648749499;
assign addr[13865] = -1660936681;
assign addr[13866] = -1672992161;
assign addr[13867] = -1684914983;
assign addr[13868] = -1696704201;
assign addr[13869] = -1708358881;
assign addr[13870] = -1719878099;
assign addr[13871] = -1731260941;
assign addr[13872] = -1742506504;
assign addr[13873] = -1753613897;
assign addr[13874] = -1764582240;
assign addr[13875] = -1775410662;
assign addr[13876] = -1786098304;
assign addr[13877] = -1796644320;
assign addr[13878] = -1807047873;
assign addr[13879] = -1817308138;
assign addr[13880] = -1827424302;
assign addr[13881] = -1837395562;
assign addr[13882] = -1847221128;
assign addr[13883] = -1856900221;
assign addr[13884] = -1866432072;
assign addr[13885] = -1875815927;
assign addr[13886] = -1885051042;
assign addr[13887] = -1894136683;
assign addr[13888] = -1903072131;
assign addr[13889] = -1911856677;
assign addr[13890] = -1920489624;
assign addr[13891] = -1928970288;
assign addr[13892] = -1937297997;
assign addr[13893] = -1945472089;
assign addr[13894] = -1953491918;
assign addr[13895] = -1961356847;
assign addr[13896] = -1969066252;
assign addr[13897] = -1976619522;
assign addr[13898] = -1984016058;
assign addr[13899] = -1991255274;
assign addr[13900] = -1998336596;
assign addr[13901] = -2005259462;
assign addr[13902] = -2012023322;
assign addr[13903] = -2018627642;
assign addr[13904] = -2025071897;
assign addr[13905] = -2031355576;
assign addr[13906] = -2037478181;
assign addr[13907] = -2043439226;
assign addr[13908] = -2049238240;
assign addr[13909] = -2054874761;
assign addr[13910] = -2060348343;
assign addr[13911] = -2065658552;
assign addr[13912] = -2070804967;
assign addr[13913] = -2075787180;
assign addr[13914] = -2080604795;
assign addr[13915] = -2085257431;
assign addr[13916] = -2089744719;
assign addr[13917] = -2094066304;
assign addr[13918] = -2098221841;
assign addr[13919] = -2102211002;
assign addr[13920] = -2106033471;
assign addr[13921] = -2109688944;
assign addr[13922] = -2113177132;
assign addr[13923] = -2116497758;
assign addr[13924] = -2119650558;
assign addr[13925] = -2122635283;
assign addr[13926] = -2125451696;
assign addr[13927] = -2128099574;
assign addr[13928] = -2130578706;
assign addr[13929] = -2132888897;
assign addr[13930] = -2135029962;
assign addr[13931] = -2137001733;
assign addr[13932] = -2138804053;
assign addr[13933] = -2140436778;
assign addr[13934] = -2141899780;
assign addr[13935] = -2143192942;
assign addr[13936] = -2144316162;
assign addr[13937] = -2145269351;
assign addr[13938] = -2146052433;
assign addr[13939] = -2146665347;
assign addr[13940] = -2147108043;
assign addr[13941] = -2147380486;
assign addr[13942] = -2147482655;
assign addr[13943] = -2147414542;
assign addr[13944] = -2147176152;
assign addr[13945] = -2146767505;
assign addr[13946] = -2146188631;
assign addr[13947] = -2145439578;
assign addr[13948] = -2144520405;
assign addr[13949] = -2143431184;
assign addr[13950] = -2142172003;
assign addr[13951] = -2140742960;
assign addr[13952] = -2139144169;
assign addr[13953] = -2137375758;
assign addr[13954] = -2135437865;
assign addr[13955] = -2133330646;
assign addr[13956] = -2131054266;
assign addr[13957] = -2128608907;
assign addr[13958] = -2125994762;
assign addr[13959] = -2123212038;
assign addr[13960] = -2120260957;
assign addr[13961] = -2117141752;
assign addr[13962] = -2113854671;
assign addr[13963] = -2110399974;
assign addr[13964] = -2106777935;
assign addr[13965] = -2102988841;
assign addr[13966] = -2099032994;
assign addr[13967] = -2094910706;
assign addr[13968] = -2090622304;
assign addr[13969] = -2086168128;
assign addr[13970] = -2081548533;
assign addr[13971] = -2076763883;
assign addr[13972] = -2071814558;
assign addr[13973] = -2066700952;
assign addr[13974] = -2061423468;
assign addr[13975] = -2055982526;
assign addr[13976] = -2050378558;
assign addr[13977] = -2044612007;
assign addr[13978] = -2038683330;
assign addr[13979] = -2032592999;
assign addr[13980] = -2026341495;
assign addr[13981] = -2019929315;
assign addr[13982] = -2013356967;
assign addr[13983] = -2006624971;
assign addr[13984] = -1999733863;
assign addr[13985] = -1992684188;
assign addr[13986] = -1985476506;
assign addr[13987] = -1978111387;
assign addr[13988] = -1970589416;
assign addr[13989] = -1962911189;
assign addr[13990] = -1955077316;
assign addr[13991] = -1947088417;
assign addr[13992] = -1938945125;
assign addr[13993] = -1930648088;
assign addr[13994] = -1922197961;
assign addr[13995] = -1913595416;
assign addr[13996] = -1904841135;
assign addr[13997] = -1895935811;
assign addr[13998] = -1886880151;
assign addr[13999] = -1877674873;
assign addr[14000] = -1868320707;
assign addr[14001] = -1858818395;
assign addr[14002] = -1849168689;
assign addr[14003] = -1839372356;
assign addr[14004] = -1829430172;
assign addr[14005] = -1819342925;
assign addr[14006] = -1809111415;
assign addr[14007] = -1798736454;
assign addr[14008] = -1788218865;
assign addr[14009] = -1777559480;
assign addr[14010] = -1766759146;
assign addr[14011] = -1755818718;
assign addr[14012] = -1744739065;
assign addr[14013] = -1733521064;
assign addr[14014] = -1722165606;
assign addr[14015] = -1710673591;
assign addr[14016] = -1699045930;
assign addr[14017] = -1687283545;
assign addr[14018] = -1675387369;
assign addr[14019] = -1663358344;
assign addr[14020] = -1651197426;
assign addr[14021] = -1638905577;
assign addr[14022] = -1626483774;
assign addr[14023] = -1613933000;
assign addr[14024] = -1601254251;
assign addr[14025] = -1588448533;
assign addr[14026] = -1575516860;
assign addr[14027] = -1562460258;
assign addr[14028] = -1549279763;
assign addr[14029] = -1535976419;
assign addr[14030] = -1522551282;
assign addr[14031] = -1509005416;
assign addr[14032] = -1495339895;
assign addr[14033] = -1481555802;
assign addr[14034] = -1467654232;
assign addr[14035] = -1453636285;
assign addr[14036] = -1439503074;
assign addr[14037] = -1425255719;
assign addr[14038] = -1410895350;
assign addr[14039] = -1396423105;
assign addr[14040] = -1381840133;
assign addr[14041] = -1367147589;
assign addr[14042] = -1352346639;
assign addr[14043] = -1337438456;
assign addr[14044] = -1322424222;
assign addr[14045] = -1307305128;
assign addr[14046] = -1292082373;
assign addr[14047] = -1276757164;
assign addr[14048] = -1261330715;
assign addr[14049] = -1245804251;
assign addr[14050] = -1230179002;
assign addr[14051] = -1214456207;
assign addr[14052] = -1198637114;
assign addr[14053] = -1182722976;
assign addr[14054] = -1166715055;
assign addr[14055] = -1150614620;
assign addr[14056] = -1134422949;
assign addr[14057] = -1118141326;
assign addr[14058] = -1101771040;
assign addr[14059] = -1085313391;
assign addr[14060] = -1068769683;
assign addr[14061] = -1052141228;
assign addr[14062] = -1035429345;
assign addr[14063] = -1018635358;
assign addr[14064] = -1001760600;
assign addr[14065] = -984806408;
assign addr[14066] = -967774128;
assign addr[14067] = -950665109;
assign addr[14068] = -933480707;
assign addr[14069] = -916222287;
assign addr[14070] = -898891215;
assign addr[14071] = -881488868;
assign addr[14072] = -864016623;
assign addr[14073] = -846475867;
assign addr[14074] = -828867991;
assign addr[14075] = -811194391;
assign addr[14076] = -793456467;
assign addr[14077] = -775655628;
assign addr[14078] = -757793284;
assign addr[14079] = -739870851;
assign addr[14080] = -721889752;
assign addr[14081] = -703851410;
assign addr[14082] = -685757258;
assign addr[14083] = -667608730;
assign addr[14084] = -649407264;
assign addr[14085] = -631154304;
assign addr[14086] = -612851297;
assign addr[14087] = -594499695;
assign addr[14088] = -576100953;
assign addr[14089] = -557656529;
assign addr[14090] = -539167887;
assign addr[14091] = -520636492;
assign addr[14092] = -502063814;
assign addr[14093] = -483451325;
assign addr[14094] = -464800501;
assign addr[14095] = -446112822;
assign addr[14096] = -427389768;
assign addr[14097] = -408632825;
assign addr[14098] = -389843480;
assign addr[14099] = -371023223;
assign addr[14100] = -352173546;
assign addr[14101] = -333295944;
assign addr[14102] = -314391913;
assign addr[14103] = -295462954;
assign addr[14104] = -276510565;
assign addr[14105] = -257536251;
assign addr[14106] = -238541516;
assign addr[14107] = -219527866;
assign addr[14108] = -200496809;
assign addr[14109] = -181449854;
assign addr[14110] = -162388511;
assign addr[14111] = -143314291;
assign addr[14112] = -124228708;
assign addr[14113] = -105133274;
assign addr[14114] = -86029503;
assign addr[14115] = -66918911;
assign addr[14116] = -47803013;
assign addr[14117] = -28683324;
assign addr[14118] = -9561361;
assign addr[14119] = 9561361;
assign addr[14120] = 28683324;
assign addr[14121] = 47803013;
assign addr[14122] = 66918911;
assign addr[14123] = 86029503;
assign addr[14124] = 105133274;
assign addr[14125] = 124228708;
assign addr[14126] = 143314291;
assign addr[14127] = 162388511;
assign addr[14128] = 181449854;
assign addr[14129] = 200496809;
assign addr[14130] = 219527866;
assign addr[14131] = 238541516;
assign addr[14132] = 257536251;
assign addr[14133] = 276510565;
assign addr[14134] = 295462954;
assign addr[14135] = 314391913;
assign addr[14136] = 333295944;
assign addr[14137] = 352173546;
assign addr[14138] = 371023223;
assign addr[14139] = 389843480;
assign addr[14140] = 408632825;
assign addr[14141] = 427389768;
assign addr[14142] = 446112822;
assign addr[14143] = 464800501;
assign addr[14144] = 483451325;
assign addr[14145] = 502063814;
assign addr[14146] = 520636492;
assign addr[14147] = 539167887;
assign addr[14148] = 557656529;
assign addr[14149] = 576100953;
assign addr[14150] = 594499695;
assign addr[14151] = 612851297;
assign addr[14152] = 631154304;
assign addr[14153] = 649407264;
assign addr[14154] = 667608730;
assign addr[14155] = 685757258;
assign addr[14156] = 703851410;
assign addr[14157] = 721889752;
assign addr[14158] = 739870851;
assign addr[14159] = 757793284;
assign addr[14160] = 775655628;
assign addr[14161] = 793456467;
assign addr[14162] = 811194391;
assign addr[14163] = 828867991;
assign addr[14164] = 846475867;
assign addr[14165] = 864016623;
assign addr[14166] = 881488868;
assign addr[14167] = 898891215;
assign addr[14168] = 916222287;
assign addr[14169] = 933480707;
assign addr[14170] = 950665109;
assign addr[14171] = 967774128;
assign addr[14172] = 984806408;
assign addr[14173] = 1001760600;
assign addr[14174] = 1018635358;
assign addr[14175] = 1035429345;
assign addr[14176] = 1052141228;
assign addr[14177] = 1068769683;
assign addr[14178] = 1085313391;
assign addr[14179] = 1101771040;
assign addr[14180] = 1118141326;
assign addr[14181] = 1134422949;
assign addr[14182] = 1150614620;
assign addr[14183] = 1166715055;
assign addr[14184] = 1182722976;
assign addr[14185] = 1198637114;
assign addr[14186] = 1214456207;
assign addr[14187] = 1230179002;
assign addr[14188] = 1245804251;
assign addr[14189] = 1261330715;
assign addr[14190] = 1276757164;
assign addr[14191] = 1292082373;
assign addr[14192] = 1307305128;
assign addr[14193] = 1322424222;
assign addr[14194] = 1337438456;
assign addr[14195] = 1352346639;
assign addr[14196] = 1367147589;
assign addr[14197] = 1381840133;
assign addr[14198] = 1396423105;
assign addr[14199] = 1410895350;
assign addr[14200] = 1425255719;
assign addr[14201] = 1439503074;
assign addr[14202] = 1453636285;
assign addr[14203] = 1467654232;
assign addr[14204] = 1481555802;
assign addr[14205] = 1495339895;
assign addr[14206] = 1509005416;
assign addr[14207] = 1522551282;
assign addr[14208] = 1535976419;
assign addr[14209] = 1549279763;
assign addr[14210] = 1562460258;
assign addr[14211] = 1575516860;
assign addr[14212] = 1588448533;
assign addr[14213] = 1601254251;
assign addr[14214] = 1613933000;
assign addr[14215] = 1626483774;
assign addr[14216] = 1638905577;
assign addr[14217] = 1651197426;
assign addr[14218] = 1663358344;
assign addr[14219] = 1675387369;
assign addr[14220] = 1687283545;
assign addr[14221] = 1699045930;
assign addr[14222] = 1710673591;
assign addr[14223] = 1722165606;
assign addr[14224] = 1733521064;
assign addr[14225] = 1744739065;
assign addr[14226] = 1755818718;
assign addr[14227] = 1766759146;
assign addr[14228] = 1777559480;
assign addr[14229] = 1788218865;
assign addr[14230] = 1798736454;
assign addr[14231] = 1809111415;
assign addr[14232] = 1819342925;
assign addr[14233] = 1829430172;
assign addr[14234] = 1839372356;
assign addr[14235] = 1849168689;
assign addr[14236] = 1858818395;
assign addr[14237] = 1868320707;
assign addr[14238] = 1877674873;
assign addr[14239] = 1886880151;
assign addr[14240] = 1895935811;
assign addr[14241] = 1904841135;
assign addr[14242] = 1913595416;
assign addr[14243] = 1922197961;
assign addr[14244] = 1930648088;
assign addr[14245] = 1938945125;
assign addr[14246] = 1947088417;
assign addr[14247] = 1955077316;
assign addr[14248] = 1962911189;
assign addr[14249] = 1970589416;
assign addr[14250] = 1978111387;
assign addr[14251] = 1985476506;
assign addr[14252] = 1992684188;
assign addr[14253] = 1999733863;
assign addr[14254] = 2006624971;
assign addr[14255] = 2013356967;
assign addr[14256] = 2019929315;
assign addr[14257] = 2026341495;
assign addr[14258] = 2032592999;
assign addr[14259] = 2038683330;
assign addr[14260] = 2044612007;
assign addr[14261] = 2050378558;
assign addr[14262] = 2055982526;
assign addr[14263] = 2061423468;
assign addr[14264] = 2066700952;
assign addr[14265] = 2071814558;
assign addr[14266] = 2076763883;
assign addr[14267] = 2081548533;
assign addr[14268] = 2086168128;
assign addr[14269] = 2090622304;
assign addr[14270] = 2094910706;
assign addr[14271] = 2099032994;
assign addr[14272] = 2102988841;
assign addr[14273] = 2106777935;
assign addr[14274] = 2110399974;
assign addr[14275] = 2113854671;
assign addr[14276] = 2117141752;
assign addr[14277] = 2120260957;
assign addr[14278] = 2123212038;
assign addr[14279] = 2125994762;
assign addr[14280] = 2128608907;
assign addr[14281] = 2131054266;
assign addr[14282] = 2133330646;
assign addr[14283] = 2135437865;
assign addr[14284] = 2137375758;
assign addr[14285] = 2139144169;
assign addr[14286] = 2140742960;
assign addr[14287] = 2142172003;
assign addr[14288] = 2143431184;
assign addr[14289] = 2144520405;
assign addr[14290] = 2145439578;
assign addr[14291] = 2146188631;
assign addr[14292] = 2146767505;
assign addr[14293] = 2147176152;
assign addr[14294] = 2147414542;
assign addr[14295] = 2147482655;
assign addr[14296] = 2147380486;
assign addr[14297] = 2147108043;
assign addr[14298] = 2146665347;
assign addr[14299] = 2146052433;
assign addr[14300] = 2145269351;
assign addr[14301] = 2144316162;
assign addr[14302] = 2143192942;
assign addr[14303] = 2141899780;
assign addr[14304] = 2140436778;
assign addr[14305] = 2138804053;
assign addr[14306] = 2137001733;
assign addr[14307] = 2135029962;
assign addr[14308] = 2132888897;
assign addr[14309] = 2130578706;
assign addr[14310] = 2128099574;
assign addr[14311] = 2125451696;
assign addr[14312] = 2122635283;
assign addr[14313] = 2119650558;
assign addr[14314] = 2116497758;
assign addr[14315] = 2113177132;
assign addr[14316] = 2109688944;
assign addr[14317] = 2106033471;
assign addr[14318] = 2102211002;
assign addr[14319] = 2098221841;
assign addr[14320] = 2094066304;
assign addr[14321] = 2089744719;
assign addr[14322] = 2085257431;
assign addr[14323] = 2080604795;
assign addr[14324] = 2075787180;
assign addr[14325] = 2070804967;
assign addr[14326] = 2065658552;
assign addr[14327] = 2060348343;
assign addr[14328] = 2054874761;
assign addr[14329] = 2049238240;
assign addr[14330] = 2043439226;
assign addr[14331] = 2037478181;
assign addr[14332] = 2031355576;
assign addr[14333] = 2025071897;
assign addr[14334] = 2018627642;
assign addr[14335] = 2012023322;
assign addr[14336] = 2005259462;
assign addr[14337] = 1998336596;
assign addr[14338] = 1991255274;
assign addr[14339] = 1984016058;
assign addr[14340] = 1976619522;
assign addr[14341] = 1969066252;
assign addr[14342] = 1961356847;
assign addr[14343] = 1953491918;
assign addr[14344] = 1945472089;
assign addr[14345] = 1937297997;
assign addr[14346] = 1928970288;
assign addr[14347] = 1920489624;
assign addr[14348] = 1911856677;
assign addr[14349] = 1903072131;
assign addr[14350] = 1894136683;
assign addr[14351] = 1885051042;
assign addr[14352] = 1875815927;
assign addr[14353] = 1866432072;
assign addr[14354] = 1856900221;
assign addr[14355] = 1847221128;
assign addr[14356] = 1837395562;
assign addr[14357] = 1827424302;
assign addr[14358] = 1817308138;
assign addr[14359] = 1807047873;
assign addr[14360] = 1796644320;
assign addr[14361] = 1786098304;
assign addr[14362] = 1775410662;
assign addr[14363] = 1764582240;
assign addr[14364] = 1753613897;
assign addr[14365] = 1742506504;
assign addr[14366] = 1731260941;
assign addr[14367] = 1719878099;
assign addr[14368] = 1708358881;
assign addr[14369] = 1696704201;
assign addr[14370] = 1684914983;
assign addr[14371] = 1672992161;
assign addr[14372] = 1660936681;
assign addr[14373] = 1648749499;
assign addr[14374] = 1636431582;
assign addr[14375] = 1623983905;
assign addr[14376] = 1611407456;
assign addr[14377] = 1598703233;
assign addr[14378] = 1585872242;
assign addr[14379] = 1572915501;
assign addr[14380] = 1559834037;
assign addr[14381] = 1546628888;
assign addr[14382] = 1533301101;
assign addr[14383] = 1519851733;
assign addr[14384] = 1506281850;
assign addr[14385] = 1492592527;
assign addr[14386] = 1478784851;
assign addr[14387] = 1464859917;
assign addr[14388] = 1450818828;
assign addr[14389] = 1436662698;
assign addr[14390] = 1422392650;
assign addr[14391] = 1408009814;
assign addr[14392] = 1393515332;
assign addr[14393] = 1378910353;
assign addr[14394] = 1364196034;
assign addr[14395] = 1349373543;
assign addr[14396] = 1334444055;
assign addr[14397] = 1319408754;
assign addr[14398] = 1304268832;
assign addr[14399] = 1289025489;
assign addr[14400] = 1273679934;
assign addr[14401] = 1258233384;
assign addr[14402] = 1242687064;
assign addr[14403] = 1227042207;
assign addr[14404] = 1211300053;
assign addr[14405] = 1195461849;
assign addr[14406] = 1179528853;
assign addr[14407] = 1163502328;
assign addr[14408] = 1147383544;
assign addr[14409] = 1131173780;
assign addr[14410] = 1114874320;
assign addr[14411] = 1098486458;
assign addr[14412] = 1082011492;
assign addr[14413] = 1065450729;
assign addr[14414] = 1048805483;
assign addr[14415] = 1032077073;
assign addr[14416] = 1015266825;
assign addr[14417] = 998376073;
assign addr[14418] = 981406156;
assign addr[14419] = 964358420;
assign addr[14420] = 947234215;
assign addr[14421] = 930034901;
assign addr[14422] = 912761841;
assign addr[14423] = 895416404;
assign addr[14424] = 877999966;
assign addr[14425] = 860513908;
assign addr[14426] = 842959617;
assign addr[14427] = 825338484;
assign addr[14428] = 807651907;
assign addr[14429] = 789901288;
assign addr[14430] = 772088034;
assign addr[14431] = 754213559;
assign addr[14432] = 736279279;
assign addr[14433] = 718286617;
assign addr[14434] = 700236999;
assign addr[14435] = 682131857;
assign addr[14436] = 663972625;
assign addr[14437] = 645760745;
assign addr[14438] = 627497660;
assign addr[14439] = 609184818;
assign addr[14440] = 590823671;
assign addr[14441] = 572415676;
assign addr[14442] = 553962291;
assign addr[14443] = 535464981;
assign addr[14444] = 516925212;
assign addr[14445] = 498344454;
assign addr[14446] = 479724180;
assign addr[14447] = 461065866;
assign addr[14448] = 442370993;
assign addr[14449] = 423641043;
assign addr[14450] = 404877501;
assign addr[14451] = 386081854;
assign addr[14452] = 367255594;
assign addr[14453] = 348400212;
assign addr[14454] = 329517204;
assign addr[14455] = 310608068;
assign addr[14456] = 291674302;
assign addr[14457] = 272717408;
assign addr[14458] = 253738890;
assign addr[14459] = 234740251;
assign addr[14460] = 215722999;
assign addr[14461] = 196688642;
assign addr[14462] = 177638688;
assign addr[14463] = 158574649;
assign addr[14464] = 139498035;
assign addr[14465] = 120410361;
assign addr[14466] = 101313138;
assign addr[14467] = 82207882;
assign addr[14468] = 63096108;
assign addr[14469] = 43979330;
assign addr[14470] = 24859065;
assign addr[14471] = 5736829;
assign addr[14472] = -13385863;
assign addr[14473] = -32507492;
assign addr[14474] = -51626544;
assign addr[14475] = -70741503;
assign addr[14476] = -89850852;
assign addr[14477] = -108953076;
assign addr[14478] = -128046661;
assign addr[14479] = -147130093;
assign addr[14480] = -166201858;
assign addr[14481] = -185260444;
assign addr[14482] = -204304341;
assign addr[14483] = -223332037;
assign addr[14484] = -242342025;
assign addr[14485] = -261332796;
assign addr[14486] = -280302845;
assign addr[14487] = -299250668;
assign addr[14488] = -318174762;
assign addr[14489] = -337073627;
assign addr[14490] = -355945764;
assign addr[14491] = -374789676;
assign addr[14492] = -393603870;
assign addr[14493] = -412386854;
assign addr[14494] = -431137138;
assign addr[14495] = -449853235;
assign addr[14496] = -468533662;
assign addr[14497] = -487176937;
assign addr[14498] = -505781581;
assign addr[14499] = -524346121;
assign addr[14500] = -542869083;
assign addr[14501] = -561348998;
assign addr[14502] = -579784402;
assign addr[14503] = -598173833;
assign addr[14504] = -616515832;
assign addr[14505] = -634808946;
assign addr[14506] = -653051723;
assign addr[14507] = -671242716;
assign addr[14508] = -689380485;
assign addr[14509] = -707463589;
assign addr[14510] = -725490597;
assign addr[14511] = -743460077;
assign addr[14512] = -761370605;
assign addr[14513] = -779220762;
assign addr[14514] = -797009130;
assign addr[14515] = -814734301;
assign addr[14516] = -832394869;
assign addr[14517] = -849989433;
assign addr[14518] = -867516597;
assign addr[14519] = -884974973;
assign addr[14520] = -902363176;
assign addr[14521] = -919679827;
assign addr[14522] = -936923553;
assign addr[14523] = -954092986;
assign addr[14524] = -971186766;
assign addr[14525] = -988203537;
assign addr[14526] = -1005141949;
assign addr[14527] = -1022000660;
assign addr[14528] = -1038778332;
assign addr[14529] = -1055473635;
assign addr[14530] = -1072085246;
assign addr[14531] = -1088611847;
assign addr[14532] = -1105052128;
assign addr[14533] = -1121404785;
assign addr[14534] = -1137668521;
assign addr[14535] = -1153842047;
assign addr[14536] = -1169924081;
assign addr[14537] = -1185913346;
assign addr[14538] = -1201808576;
assign addr[14539] = -1217608510;
assign addr[14540] = -1233311895;
assign addr[14541] = -1248917486;
assign addr[14542] = -1264424045;
assign addr[14543] = -1279830344;
assign addr[14544] = -1295135159;
assign addr[14545] = -1310337279;
assign addr[14546] = -1325435496;
assign addr[14547] = -1340428615;
assign addr[14548] = -1355315445;
assign addr[14549] = -1370094808;
assign addr[14550] = -1384765530;
assign addr[14551] = -1399326449;
assign addr[14552] = -1413776410;
assign addr[14553] = -1428114267;
assign addr[14554] = -1442338884;
assign addr[14555] = -1456449131;
assign addr[14556] = -1470443891;
assign addr[14557] = -1484322054;
assign addr[14558] = -1498082520;
assign addr[14559] = -1511724196;
assign addr[14560] = -1525246002;
assign addr[14561] = -1538646865;
assign addr[14562] = -1551925723;
assign addr[14563] = -1565081523;
assign addr[14564] = -1578113222;
assign addr[14565] = -1591019785;
assign addr[14566] = -1603800191;
assign addr[14567] = -1616453425;
assign addr[14568] = -1628978484;
assign addr[14569] = -1641374375;
assign addr[14570] = -1653640115;
assign addr[14571] = -1665774731;
assign addr[14572] = -1677777262;
assign addr[14573] = -1689646755;
assign addr[14574] = -1701382270;
assign addr[14575] = -1712982875;
assign addr[14576] = -1724447652;
assign addr[14577] = -1735775690;
assign addr[14578] = -1746966091;
assign addr[14579] = -1758017969;
assign addr[14580] = -1768930447;
assign addr[14581] = -1779702660;
assign addr[14582] = -1790333753;
assign addr[14583] = -1800822883;
assign addr[14584] = -1811169220;
assign addr[14585] = -1821371941;
assign addr[14586] = -1831430239;
assign addr[14587] = -1841343316;
assign addr[14588] = -1851110385;
assign addr[14589] = -1860730673;
assign addr[14590] = -1870203416;
assign addr[14591] = -1879527863;
assign addr[14592] = -1888703276;
assign addr[14593] = -1897728925;
assign addr[14594] = -1906604097;
assign addr[14595] = -1915328086;
assign addr[14596] = -1923900201;
assign addr[14597] = -1932319763;
assign addr[14598] = -1940586104;
assign addr[14599] = -1948698568;
assign addr[14600] = -1956656513;
assign addr[14601] = -1964459306;
assign addr[14602] = -1972106330;
assign addr[14603] = -1979596978;
assign addr[14604] = -1986930656;
assign addr[14605] = -1994106782;
assign addr[14606] = -2001124788;
assign addr[14607] = -2007984117;
assign addr[14608] = -2014684225;
assign addr[14609] = -2021224581;
assign addr[14610] = -2027604666;
assign addr[14611] = -2033823974;
assign addr[14612] = -2039882013;
assign addr[14613] = -2045778302;
assign addr[14614] = -2051512372;
assign addr[14615] = -2057083771;
assign addr[14616] = -2062492055;
assign addr[14617] = -2067736796;
assign addr[14618] = -2072817579;
assign addr[14619] = -2077733999;
assign addr[14620] = -2082485668;
assign addr[14621] = -2087072209;
assign addr[14622] = -2091493257;
assign addr[14623] = -2095748463;
assign addr[14624] = -2099837489;
assign addr[14625] = -2103760010;
assign addr[14626] = -2107515716;
assign addr[14627] = -2111104309;
assign addr[14628] = -2114525505;
assign addr[14629] = -2117779031;
assign addr[14630] = -2120864631;
assign addr[14631] = -2123782059;
assign addr[14632] = -2126531084;
assign addr[14633] = -2129111488;
assign addr[14634] = -2131523066;
assign addr[14635] = -2133765628;
assign addr[14636] = -2135838995;
assign addr[14637] = -2137743003;
assign addr[14638] = -2139477502;
assign addr[14639] = -2141042352;
assign addr[14640] = -2142437431;
assign addr[14641] = -2143662628;
assign addr[14642] = -2144717846;
assign addr[14643] = -2145603001;
assign addr[14644] = -2146318022;
assign addr[14645] = -2146862854;
assign addr[14646] = -2147237452;
assign addr[14647] = -2147441787;
assign addr[14648] = -2147475844;
assign addr[14649] = -2147339619;
assign addr[14650] = -2147033123;
assign addr[14651] = -2146556380;
assign addr[14652] = -2145909429;
assign addr[14653] = -2145092320;
assign addr[14654] = -2144105118;
assign addr[14655] = -2142947902;
assign addr[14656] = -2141620763;
assign addr[14657] = -2140123807;
assign addr[14658] = -2138457152;
assign addr[14659] = -2136620930;
assign addr[14660] = -2134615288;
assign addr[14661] = -2132440383;
assign addr[14662] = -2130096389;
assign addr[14663] = -2127583492;
assign addr[14664] = -2124901890;
assign addr[14665] = -2122051796;
assign addr[14666] = -2119033436;
assign addr[14667] = -2115847050;
assign addr[14668] = -2112492891;
assign addr[14669] = -2108971223;
assign addr[14670] = -2105282327;
assign addr[14671] = -2101426496;
assign addr[14672] = -2097404033;
assign addr[14673] = -2093215260;
assign addr[14674] = -2088860507;
assign addr[14675] = -2084340120;
assign addr[14676] = -2079654458;
assign addr[14677] = -2074803892;
assign addr[14678] = -2069788807;
assign addr[14679] = -2064609600;
assign addr[14680] = -2059266683;
assign addr[14681] = -2053760478;
assign addr[14682] = -2048091422;
assign addr[14683] = -2042259965;
assign addr[14684] = -2036266570;
assign addr[14685] = -2030111710;
assign addr[14686] = -2023795876;
assign addr[14687] = -2017319567;
assign addr[14688] = -2010683297;
assign addr[14689] = -2003887591;
assign addr[14690] = -1996932990;
assign addr[14691] = -1989820044;
assign addr[14692] = -1982549318;
assign addr[14693] = -1975121388;
assign addr[14694] = -1967536842;
assign addr[14695] = -1959796283;
assign addr[14696] = -1951900324;
assign addr[14697] = -1943849591;
assign addr[14698] = -1935644723;
assign addr[14699] = -1927286370;
assign addr[14700] = -1918775195;
assign addr[14701] = -1910111873;
assign addr[14702] = -1901297091;
assign addr[14703] = -1892331547;
assign addr[14704] = -1883215953;
assign addr[14705] = -1873951032;
assign addr[14706] = -1864537518;
assign addr[14707] = -1854976157;
assign addr[14708] = -1845267708;
assign addr[14709] = -1835412941;
assign addr[14710] = -1825412636;
assign addr[14711] = -1815267588;
assign addr[14712] = -1804978599;
assign addr[14713] = -1794546487;
assign addr[14714] = -1783972079;
assign addr[14715] = -1773256212;
assign addr[14716] = -1762399737;
assign addr[14717] = -1751403515;
assign addr[14718] = -1740268417;
assign addr[14719] = -1728995326;
assign addr[14720] = -1717585136;
assign addr[14721] = -1706038753;
assign addr[14722] = -1694357091;
assign addr[14723] = -1682541077;
assign addr[14724] = -1670591647;
assign addr[14725] = -1658509750;
assign addr[14726] = -1646296344;
assign addr[14727] = -1633952396;
assign addr[14728] = -1621478885;
assign addr[14729] = -1608876801;
assign addr[14730] = -1596147143;
assign addr[14731] = -1583290921;
assign addr[14732] = -1570309153;
assign addr[14733] = -1557202869;
assign addr[14734] = -1543973108;
assign addr[14735] = -1530620920;
assign addr[14736] = -1517147363;
assign addr[14737] = -1503553506;
assign addr[14738] = -1489840425;
assign addr[14739] = -1476009210;
assign addr[14740] = -1462060956;
assign addr[14741] = -1447996770;
assign addr[14742] = -1433817766;
assign addr[14743] = -1419525069;
assign addr[14744] = -1405119813;
assign addr[14745] = -1390603139;
assign addr[14746] = -1375976199;
assign addr[14747] = -1361240152;
assign addr[14748] = -1346396168;
assign addr[14749] = -1331445422;
assign addr[14750] = -1316389101;
assign addr[14751] = -1301228398;
assign addr[14752] = -1285964516;
assign addr[14753] = -1270598665;
assign addr[14754] = -1255132063;
assign addr[14755] = -1239565936;
assign addr[14756] = -1223901520;
assign addr[14757] = -1208140056;
assign addr[14758] = -1192282793;
assign addr[14759] = -1176330990;
assign addr[14760] = -1160285911;
assign addr[14761] = -1144148829;
assign addr[14762] = -1127921022;
assign addr[14763] = -1111603778;
assign addr[14764] = -1095198391;
assign addr[14765] = -1078706161;
assign addr[14766] = -1062128397;
assign addr[14767] = -1045466412;
assign addr[14768] = -1028721528;
assign addr[14769] = -1011895073;
assign addr[14770] = -994988380;
assign addr[14771] = -978002791;
assign addr[14772] = -960939653;
assign addr[14773] = -943800318;
assign addr[14774] = -926586145;
assign addr[14775] = -909298500;
assign addr[14776] = -891938752;
assign addr[14777] = -874508280;
assign addr[14778] = -857008464;
assign addr[14779] = -839440693;
assign addr[14780] = -821806359;
assign addr[14781] = -804106861;
assign addr[14782] = -786343603;
assign addr[14783] = -768517992;
assign addr[14784] = -750631442;
assign addr[14785] = -732685372;
assign addr[14786] = -714681204;
assign addr[14787] = -696620367;
assign addr[14788] = -678504291;
assign addr[14789] = -660334415;
assign addr[14790] = -642112178;
assign addr[14791] = -623839025;
assign addr[14792] = -605516406;
assign addr[14793] = -587145773;
assign addr[14794] = -568728583;
assign addr[14795] = -550266296;
assign addr[14796] = -531760377;
assign addr[14797] = -513212292;
assign addr[14798] = -494623513;
assign addr[14799] = -475995513;
assign addr[14800] = -457329769;
assign addr[14801] = -438627762;
assign addr[14802] = -419890975;
assign addr[14803] = -401120892;
assign addr[14804] = -382319004;
assign addr[14805] = -363486799;
assign addr[14806] = -344625773;
assign addr[14807] = -325737419;
assign addr[14808] = -306823237;
assign addr[14809] = -287884725;
assign addr[14810] = -268923386;
assign addr[14811] = -249940723;
assign addr[14812] = -230938242;
assign addr[14813] = -211917448;
assign addr[14814] = -192879850;
assign addr[14815] = -173826959;
assign addr[14816] = -154760284;
assign addr[14817] = -135681337;
assign addr[14818] = -116591632;
assign addr[14819] = -97492681;
assign addr[14820] = -78386000;
assign addr[14821] = -59273104;
assign addr[14822] = -40155507;
assign addr[14823] = -21034727;
assign addr[14824] = -1912278;
assign addr[14825] = 17210322;
assign addr[14826] = 36331557;
assign addr[14827] = 55449912;
assign addr[14828] = 74563870;
assign addr[14829] = 93671915;
assign addr[14830] = 112772533;
assign addr[14831] = 131864208;
assign addr[14832] = 150945428;
assign addr[14833] = 170014678;
assign addr[14834] = 189070447;
assign addr[14835] = 208111224;
assign addr[14836] = 227135500;
assign addr[14837] = 246141764;
assign addr[14838] = 265128512;
assign addr[14839] = 284094236;
assign addr[14840] = 303037433;
assign addr[14841] = 321956601;
assign addr[14842] = 340850240;
assign addr[14843] = 359716852;
assign addr[14844] = 378554940;
assign addr[14845] = 397363011;
assign addr[14846] = 416139574;
assign addr[14847] = 434883140;
assign addr[14848] = 453592221;
assign addr[14849] = 472265336;
assign addr[14850] = 490901003;
assign addr[14851] = 509497745;
assign addr[14852] = 528054086;
assign addr[14853] = 546568556;
assign addr[14854] = 565039687;
assign addr[14855] = 583466013;
assign addr[14856] = 601846074;
assign addr[14857] = 620178412;
assign addr[14858] = 638461574;
assign addr[14859] = 656694110;
assign addr[14860] = 674874574;
assign addr[14861] = 693001525;
assign addr[14862] = 711073524;
assign addr[14863] = 729089140;
assign addr[14864] = 747046944;
assign addr[14865] = 764945512;
assign addr[14866] = 782783424;
assign addr[14867] = 800559266;
assign addr[14868] = 818271628;
assign addr[14869] = 835919107;
assign addr[14870] = 853500302;
assign addr[14871] = 871013820;
assign addr[14872] = 888458272;
assign addr[14873] = 905832274;
assign addr[14874] = 923134450;
assign addr[14875] = 940363427;
assign addr[14876] = 957517838;
assign addr[14877] = 974596324;
assign addr[14878] = 991597531;
assign addr[14879] = 1008520110;
assign addr[14880] = 1025362720;
assign addr[14881] = 1042124025;
assign addr[14882] = 1058802695;
assign addr[14883] = 1075397409;
assign addr[14884] = 1091906851;
assign addr[14885] = 1108329711;
assign addr[14886] = 1124664687;
assign addr[14887] = 1140910484;
assign addr[14888] = 1157065814;
assign addr[14889] = 1173129396;
assign addr[14890] = 1189099956;
assign addr[14891] = 1204976227;
assign addr[14892] = 1220756951;
assign addr[14893] = 1236440877;
assign addr[14894] = 1252026760;
assign addr[14895] = 1267513365;
assign addr[14896] = 1282899464;
assign addr[14897] = 1298183838;
assign addr[14898] = 1313365273;
assign addr[14899] = 1328442566;
assign addr[14900] = 1343414522;
assign addr[14901] = 1358279953;
assign addr[14902] = 1373037681;
assign addr[14903] = 1387686535;
assign addr[14904] = 1402225355;
assign addr[14905] = 1416652986;
assign addr[14906] = 1430968286;
assign addr[14907] = 1445170118;
assign addr[14908] = 1459257358;
assign addr[14909] = 1473228887;
assign addr[14910] = 1487083598;
assign addr[14911] = 1500820393;
assign addr[14912] = 1514438181;
assign addr[14913] = 1527935884;
assign addr[14914] = 1541312431;
assign addr[14915] = 1554566762;
assign addr[14916] = 1567697824;
assign addr[14917] = 1580704578;
assign addr[14918] = 1593585992;
assign addr[14919] = 1606341043;
assign addr[14920] = 1618968722;
assign addr[14921] = 1631468027;
assign addr[14922] = 1643837966;
assign addr[14923] = 1656077559;
assign addr[14924] = 1668185835;
assign addr[14925] = 1680161834;
assign addr[14926] = 1692004606;
assign addr[14927] = 1703713213;
assign addr[14928] = 1715286726;
assign addr[14929] = 1726724227;
assign addr[14930] = 1738024810;
assign addr[14931] = 1749187577;
assign addr[14932] = 1760211645;
assign addr[14933] = 1771096139;
assign addr[14934] = 1781840195;
assign addr[14935] = 1792442963;
assign addr[14936] = 1802903601;
assign addr[14937] = 1813221279;
assign addr[14938] = 1823395180;
assign addr[14939] = 1833424497;
assign addr[14940] = 1843308435;
assign addr[14941] = 1853046210;
assign addr[14942] = 1862637049;
assign addr[14943] = 1872080193;
assign addr[14944] = 1881374892;
assign addr[14945] = 1890520410;
assign addr[14946] = 1899516021;
assign addr[14947] = 1908361011;
assign addr[14948] = 1917054681;
assign addr[14949] = 1925596340;
assign addr[14950] = 1933985310;
assign addr[14951] = 1942220928;
assign addr[14952] = 1950302539;
assign addr[14953] = 1958229503;
assign addr[14954] = 1966001192;
assign addr[14955] = 1973616989;
assign addr[14956] = 1981076290;
assign addr[14957] = 1988378503;
assign addr[14958] = 1995523051;
assign addr[14959] = 2002509365;
assign addr[14960] = 2009336893;
assign addr[14961] = 2016005093;
assign addr[14962] = 2022513436;
assign addr[14963] = 2028861406;
assign addr[14964] = 2035048499;
assign addr[14965] = 2041074226;
assign addr[14966] = 2046938108;
assign addr[14967] = 2052639680;
assign addr[14968] = 2058178491;
assign addr[14969] = 2063554100;
assign addr[14970] = 2068766083;
assign addr[14971] = 2073814024;
assign addr[14972] = 2078697525;
assign addr[14973] = 2083416198;
assign addr[14974] = 2087969669;
assign addr[14975] = 2092357577;
assign addr[14976] = 2096579573;
assign addr[14977] = 2100635323;
assign addr[14978] = 2104524506;
assign addr[14979] = 2108246813;
assign addr[14980] = 2111801949;
assign addr[14981] = 2115189632;
assign addr[14982] = 2118409593;
assign addr[14983] = 2121461578;
assign addr[14984] = 2124345343;
assign addr[14985] = 2127060661;
assign addr[14986] = 2129607316;
assign addr[14987] = 2131985106;
assign addr[14988] = 2134193842;
assign addr[14989] = 2136233350;
assign addr[14990] = 2138103468;
assign addr[14991] = 2139804048;
assign addr[14992] = 2141334954;
assign addr[14993] = 2142696065;
assign addr[14994] = 2143887273;
assign addr[14995] = 2144908484;
assign addr[14996] = 2145759618;
assign addr[14997] = 2146440605;
assign addr[14998] = 2146951393;
assign addr[14999] = 2147291941;
assign addr[15000] = 2147462221;
assign addr[15001] = 2147462221;
assign addr[15002] = 2147291941;
assign addr[15003] = 2146951393;
assign addr[15004] = 2146440605;
assign addr[15005] = 2145759618;
assign addr[15006] = 2144908484;
assign addr[15007] = 2143887273;
assign addr[15008] = 2142696065;
assign addr[15009] = 2141334954;
assign addr[15010] = 2139804048;
assign addr[15011] = 2138103468;
assign addr[15012] = 2136233350;
assign addr[15013] = 2134193842;
assign addr[15014] = 2131985106;
assign addr[15015] = 2129607316;
assign addr[15016] = 2127060661;
assign addr[15017] = 2124345343;
assign addr[15018] = 2121461578;
assign addr[15019] = 2118409593;
assign addr[15020] = 2115189632;
assign addr[15021] = 2111801949;
assign addr[15022] = 2108246813;
assign addr[15023] = 2104524506;
assign addr[15024] = 2100635323;
assign addr[15025] = 2096579573;
assign addr[15026] = 2092357577;
assign addr[15027] = 2087969669;
assign addr[15028] = 2083416198;
assign addr[15029] = 2078697525;
assign addr[15030] = 2073814024;
assign addr[15031] = 2068766083;
assign addr[15032] = 2063554100;
assign addr[15033] = 2058178491;
assign addr[15034] = 2052639680;
assign addr[15035] = 2046938108;
assign addr[15036] = 2041074226;
assign addr[15037] = 2035048499;
assign addr[15038] = 2028861406;
assign addr[15039] = 2022513436;
assign addr[15040] = 2016005093;
assign addr[15041] = 2009336893;
assign addr[15042] = 2002509365;
assign addr[15043] = 1995523051;
assign addr[15044] = 1988378503;
assign addr[15045] = 1981076290;
assign addr[15046] = 1973616989;
assign addr[15047] = 1966001192;
assign addr[15048] = 1958229503;
assign addr[15049] = 1950302539;
assign addr[15050] = 1942220928;
assign addr[15051] = 1933985310;
assign addr[15052] = 1925596340;
assign addr[15053] = 1917054681;
assign addr[15054] = 1908361011;
assign addr[15055] = 1899516021;
assign addr[15056] = 1890520410;
assign addr[15057] = 1881374892;
assign addr[15058] = 1872080193;
assign addr[15059] = 1862637049;
assign addr[15060] = 1853046210;
assign addr[15061] = 1843308435;
assign addr[15062] = 1833424497;
assign addr[15063] = 1823395180;
assign addr[15064] = 1813221279;
assign addr[15065] = 1802903601;
assign addr[15066] = 1792442963;
assign addr[15067] = 1781840195;
assign addr[15068] = 1771096139;
assign addr[15069] = 1760211645;
assign addr[15070] = 1749187577;
assign addr[15071] = 1738024810;
assign addr[15072] = 1726724227;
assign addr[15073] = 1715286726;
assign addr[15074] = 1703713213;
assign addr[15075] = 1692004606;
assign addr[15076] = 1680161834;
assign addr[15077] = 1668185835;
assign addr[15078] = 1656077559;
assign addr[15079] = 1643837966;
assign addr[15080] = 1631468027;
assign addr[15081] = 1618968722;
assign addr[15082] = 1606341043;
assign addr[15083] = 1593585992;
assign addr[15084] = 1580704578;
assign addr[15085] = 1567697824;
assign addr[15086] = 1554566762;
assign addr[15087] = 1541312431;
assign addr[15088] = 1527935884;
assign addr[15089] = 1514438181;
assign addr[15090] = 1500820393;
assign addr[15091] = 1487083598;
assign addr[15092] = 1473228887;
assign addr[15093] = 1459257358;
assign addr[15094] = 1445170118;
assign addr[15095] = 1430968286;
assign addr[15096] = 1416652986;
assign addr[15097] = 1402225355;
assign addr[15098] = 1387686535;
assign addr[15099] = 1373037681;
assign addr[15100] = 1358279953;
assign addr[15101] = 1343414522;
assign addr[15102] = 1328442566;
assign addr[15103] = 1313365273;
assign addr[15104] = 1298183838;
assign addr[15105] = 1282899464;
assign addr[15106] = 1267513365;
assign addr[15107] = 1252026760;
assign addr[15108] = 1236440877;
assign addr[15109] = 1220756951;
assign addr[15110] = 1204976227;
assign addr[15111] = 1189099956;
assign addr[15112] = 1173129396;
assign addr[15113] = 1157065814;
assign addr[15114] = 1140910484;
assign addr[15115] = 1124664687;
assign addr[15116] = 1108329711;
assign addr[15117] = 1091906851;
assign addr[15118] = 1075397409;
assign addr[15119] = 1058802695;
assign addr[15120] = 1042124025;
assign addr[15121] = 1025362720;
assign addr[15122] = 1008520110;
assign addr[15123] = 991597531;
assign addr[15124] = 974596324;
assign addr[15125] = 957517838;
assign addr[15126] = 940363427;
assign addr[15127] = 923134450;
assign addr[15128] = 905832274;
assign addr[15129] = 888458272;
assign addr[15130] = 871013820;
assign addr[15131] = 853500302;
assign addr[15132] = 835919107;
assign addr[15133] = 818271628;
assign addr[15134] = 800559266;
assign addr[15135] = 782783424;
assign addr[15136] = 764945512;
assign addr[15137] = 747046944;
assign addr[15138] = 729089140;
assign addr[15139] = 711073524;
assign addr[15140] = 693001525;
assign addr[15141] = 674874574;
assign addr[15142] = 656694110;
assign addr[15143] = 638461574;
assign addr[15144] = 620178412;
assign addr[15145] = 601846074;
assign addr[15146] = 583466013;
assign addr[15147] = 565039687;
assign addr[15148] = 546568556;
assign addr[15149] = 528054086;
assign addr[15150] = 509497745;
assign addr[15151] = 490901003;
assign addr[15152] = 472265336;
assign addr[15153] = 453592221;
assign addr[15154] = 434883140;
assign addr[15155] = 416139574;
assign addr[15156] = 397363011;
assign addr[15157] = 378554940;
assign addr[15158] = 359716852;
assign addr[15159] = 340850240;
assign addr[15160] = 321956601;
assign addr[15161] = 303037433;
assign addr[15162] = 284094236;
assign addr[15163] = 265128512;
assign addr[15164] = 246141764;
assign addr[15165] = 227135500;
assign addr[15166] = 208111224;
assign addr[15167] = 189070447;
assign addr[15168] = 170014678;
assign addr[15169] = 150945428;
assign addr[15170] = 131864208;
assign addr[15171] = 112772533;
assign addr[15172] = 93671915;
assign addr[15173] = 74563870;
assign addr[15174] = 55449912;
assign addr[15175] = 36331557;
assign addr[15176] = 17210322;
assign addr[15177] = -1912278;
assign addr[15178] = -21034727;
assign addr[15179] = -40155507;
assign addr[15180] = -59273104;
assign addr[15181] = -78386000;
assign addr[15182] = -97492681;
assign addr[15183] = -116591632;
assign addr[15184] = -135681337;
assign addr[15185] = -154760284;
assign addr[15186] = -173826959;
assign addr[15187] = -192879850;
assign addr[15188] = -211917448;
assign addr[15189] = -230938242;
assign addr[15190] = -249940723;
assign addr[15191] = -268923386;
assign addr[15192] = -287884725;
assign addr[15193] = -306823237;
assign addr[15194] = -325737419;
assign addr[15195] = -344625773;
assign addr[15196] = -363486799;
assign addr[15197] = -382319004;
assign addr[15198] = -401120892;
assign addr[15199] = -419890975;
assign addr[15200] = -438627762;
assign addr[15201] = -457329769;
assign addr[15202] = -475995513;
assign addr[15203] = -494623513;
assign addr[15204] = -513212292;
assign addr[15205] = -531760377;
assign addr[15206] = -550266296;
assign addr[15207] = -568728583;
assign addr[15208] = -587145773;
assign addr[15209] = -605516406;
assign addr[15210] = -623839025;
assign addr[15211] = -642112178;
assign addr[15212] = -660334415;
assign addr[15213] = -678504291;
assign addr[15214] = -696620367;
assign addr[15215] = -714681204;
assign addr[15216] = -732685372;
assign addr[15217] = -750631442;
assign addr[15218] = -768517992;
assign addr[15219] = -786343603;
assign addr[15220] = -804106861;
assign addr[15221] = -821806359;
assign addr[15222] = -839440693;
assign addr[15223] = -857008464;
assign addr[15224] = -874508280;
assign addr[15225] = -891938752;
assign addr[15226] = -909298500;
assign addr[15227] = -926586145;
assign addr[15228] = -943800318;
assign addr[15229] = -960939653;
assign addr[15230] = -978002791;
assign addr[15231] = -994988380;
assign addr[15232] = -1011895073;
assign addr[15233] = -1028721528;
assign addr[15234] = -1045466412;
assign addr[15235] = -1062128397;
assign addr[15236] = -1078706161;
assign addr[15237] = -1095198391;
assign addr[15238] = -1111603778;
assign addr[15239] = -1127921022;
assign addr[15240] = -1144148829;
assign addr[15241] = -1160285911;
assign addr[15242] = -1176330990;
assign addr[15243] = -1192282793;
assign addr[15244] = -1208140056;
assign addr[15245] = -1223901520;
assign addr[15246] = -1239565936;
assign addr[15247] = -1255132063;
assign addr[15248] = -1270598665;
assign addr[15249] = -1285964516;
assign addr[15250] = -1301228398;
assign addr[15251] = -1316389101;
assign addr[15252] = -1331445422;
assign addr[15253] = -1346396168;
assign addr[15254] = -1361240152;
assign addr[15255] = -1375976199;
assign addr[15256] = -1390603139;
assign addr[15257] = -1405119813;
assign addr[15258] = -1419525069;
assign addr[15259] = -1433817766;
assign addr[15260] = -1447996770;
assign addr[15261] = -1462060956;
assign addr[15262] = -1476009210;
assign addr[15263] = -1489840425;
assign addr[15264] = -1503553506;
assign addr[15265] = -1517147363;
assign addr[15266] = -1530620920;
assign addr[15267] = -1543973108;
assign addr[15268] = -1557202869;
assign addr[15269] = -1570309153;
assign addr[15270] = -1583290921;
assign addr[15271] = -1596147143;
assign addr[15272] = -1608876801;
assign addr[15273] = -1621478885;
assign addr[15274] = -1633952396;
assign addr[15275] = -1646296344;
assign addr[15276] = -1658509750;
assign addr[15277] = -1670591647;
assign addr[15278] = -1682541077;
assign addr[15279] = -1694357091;
assign addr[15280] = -1706038753;
assign addr[15281] = -1717585136;
assign addr[15282] = -1728995326;
assign addr[15283] = -1740268417;
assign addr[15284] = -1751403515;
assign addr[15285] = -1762399737;
assign addr[15286] = -1773256212;
assign addr[15287] = -1783972079;
assign addr[15288] = -1794546487;
assign addr[15289] = -1804978599;
assign addr[15290] = -1815267588;
assign addr[15291] = -1825412636;
assign addr[15292] = -1835412941;
assign addr[15293] = -1845267708;
assign addr[15294] = -1854976157;
assign addr[15295] = -1864537518;
assign addr[15296] = -1873951032;
assign addr[15297] = -1883215953;
assign addr[15298] = -1892331547;
assign addr[15299] = -1901297091;
assign addr[15300] = -1910111873;
assign addr[15301] = -1918775195;
assign addr[15302] = -1927286370;
assign addr[15303] = -1935644723;
assign addr[15304] = -1943849591;
assign addr[15305] = -1951900324;
assign addr[15306] = -1959796283;
assign addr[15307] = -1967536842;
assign addr[15308] = -1975121388;
assign addr[15309] = -1982549318;
assign addr[15310] = -1989820044;
assign addr[15311] = -1996932990;
assign addr[15312] = -2003887591;
assign addr[15313] = -2010683297;
assign addr[15314] = -2017319567;
assign addr[15315] = -2023795876;
assign addr[15316] = -2030111710;
assign addr[15317] = -2036266570;
assign addr[15318] = -2042259965;
assign addr[15319] = -2048091422;
assign addr[15320] = -2053760478;
assign addr[15321] = -2059266683;
assign addr[15322] = -2064609600;
assign addr[15323] = -2069788807;
assign addr[15324] = -2074803892;
assign addr[15325] = -2079654458;
assign addr[15326] = -2084340120;
assign addr[15327] = -2088860507;
assign addr[15328] = -2093215260;
assign addr[15329] = -2097404033;
assign addr[15330] = -2101426496;
assign addr[15331] = -2105282327;
assign addr[15332] = -2108971223;
assign addr[15333] = -2112492891;
assign addr[15334] = -2115847050;
assign addr[15335] = -2119033436;
assign addr[15336] = -2122051796;
assign addr[15337] = -2124901890;
assign addr[15338] = -2127583492;
assign addr[15339] = -2130096389;
assign addr[15340] = -2132440383;
assign addr[15341] = -2134615288;
assign addr[15342] = -2136620930;
assign addr[15343] = -2138457152;
assign addr[15344] = -2140123807;
assign addr[15345] = -2141620763;
assign addr[15346] = -2142947902;
assign addr[15347] = -2144105118;
assign addr[15348] = -2145092320;
assign addr[15349] = -2145909429;
assign addr[15350] = -2146556380;
assign addr[15351] = -2147033123;
assign addr[15352] = -2147339619;
assign addr[15353] = -2147475844;
assign addr[15354] = -2147441787;
assign addr[15355] = -2147237452;
assign addr[15356] = -2146862854;
assign addr[15357] = -2146318022;
assign addr[15358] = -2145603001;
assign addr[15359] = -2144717846;
assign addr[15360] = -2143662628;
assign addr[15361] = -2142437431;
assign addr[15362] = -2141042352;
assign addr[15363] = -2139477502;
assign addr[15364] = -2137743003;
assign addr[15365] = -2135838995;
assign addr[15366] = -2133765628;
assign addr[15367] = -2131523066;
assign addr[15368] = -2129111488;
assign addr[15369] = -2126531084;
assign addr[15370] = -2123782059;
assign addr[15371] = -2120864631;
assign addr[15372] = -2117779031;
assign addr[15373] = -2114525505;
assign addr[15374] = -2111104309;
assign addr[15375] = -2107515716;
assign addr[15376] = -2103760010;
assign addr[15377] = -2099837489;
assign addr[15378] = -2095748463;
assign addr[15379] = -2091493257;
assign addr[15380] = -2087072209;
assign addr[15381] = -2082485668;
assign addr[15382] = -2077733999;
assign addr[15383] = -2072817579;
assign addr[15384] = -2067736796;
assign addr[15385] = -2062492055;
assign addr[15386] = -2057083771;
assign addr[15387] = -2051512372;
assign addr[15388] = -2045778302;
assign addr[15389] = -2039882013;
assign addr[15390] = -2033823974;
assign addr[15391] = -2027604666;
assign addr[15392] = -2021224581;
assign addr[15393] = -2014684225;
assign addr[15394] = -2007984117;
assign addr[15395] = -2001124788;
assign addr[15396] = -1994106782;
assign addr[15397] = -1986930656;
assign addr[15398] = -1979596978;
assign addr[15399] = -1972106330;
assign addr[15400] = -1964459306;
assign addr[15401] = -1956656513;
assign addr[15402] = -1948698568;
assign addr[15403] = -1940586104;
assign addr[15404] = -1932319763;
assign addr[15405] = -1923900201;
assign addr[15406] = -1915328086;
assign addr[15407] = -1906604097;
assign addr[15408] = -1897728925;
assign addr[15409] = -1888703276;
assign addr[15410] = -1879527863;
assign addr[15411] = -1870203416;
assign addr[15412] = -1860730673;
assign addr[15413] = -1851110385;
assign addr[15414] = -1841343316;
assign addr[15415] = -1831430239;
assign addr[15416] = -1821371941;
assign addr[15417] = -1811169220;
assign addr[15418] = -1800822883;
assign addr[15419] = -1790333753;
assign addr[15420] = -1779702660;
assign addr[15421] = -1768930447;
assign addr[15422] = -1758017969;
assign addr[15423] = -1746966091;
assign addr[15424] = -1735775690;
assign addr[15425] = -1724447652;
assign addr[15426] = -1712982875;
assign addr[15427] = -1701382270;
assign addr[15428] = -1689646755;
assign addr[15429] = -1677777262;
assign addr[15430] = -1665774731;
assign addr[15431] = -1653640115;
assign addr[15432] = -1641374375;
assign addr[15433] = -1628978484;
assign addr[15434] = -1616453425;
assign addr[15435] = -1603800191;
assign addr[15436] = -1591019785;
assign addr[15437] = -1578113222;
assign addr[15438] = -1565081523;
assign addr[15439] = -1551925723;
assign addr[15440] = -1538646865;
assign addr[15441] = -1525246002;
assign addr[15442] = -1511724196;
assign addr[15443] = -1498082520;
assign addr[15444] = -1484322054;
assign addr[15445] = -1470443891;
assign addr[15446] = -1456449131;
assign addr[15447] = -1442338884;
assign addr[15448] = -1428114267;
assign addr[15449] = -1413776410;
assign addr[15450] = -1399326449;
assign addr[15451] = -1384765530;
assign addr[15452] = -1370094808;
assign addr[15453] = -1355315445;
assign addr[15454] = -1340428615;
assign addr[15455] = -1325435496;
assign addr[15456] = -1310337279;
assign addr[15457] = -1295135159;
assign addr[15458] = -1279830344;
assign addr[15459] = -1264424045;
assign addr[15460] = -1248917486;
assign addr[15461] = -1233311895;
assign addr[15462] = -1217608510;
assign addr[15463] = -1201808576;
assign addr[15464] = -1185913346;
assign addr[15465] = -1169924081;
assign addr[15466] = -1153842047;
assign addr[15467] = -1137668521;
assign addr[15468] = -1121404785;
assign addr[15469] = -1105052128;
assign addr[15470] = -1088611847;
assign addr[15471] = -1072085246;
assign addr[15472] = -1055473635;
assign addr[15473] = -1038778332;
assign addr[15474] = -1022000660;
assign addr[15475] = -1005141949;
assign addr[15476] = -988203537;
assign addr[15477] = -971186766;
assign addr[15478] = -954092986;
assign addr[15479] = -936923553;
assign addr[15480] = -919679827;
assign addr[15481] = -902363176;
assign addr[15482] = -884974973;
assign addr[15483] = -867516597;
assign addr[15484] = -849989433;
assign addr[15485] = -832394869;
assign addr[15486] = -814734301;
assign addr[15487] = -797009130;
assign addr[15488] = -779220762;
assign addr[15489] = -761370605;
assign addr[15490] = -743460077;
assign addr[15491] = -725490597;
assign addr[15492] = -707463589;
assign addr[15493] = -689380485;
assign addr[15494] = -671242716;
assign addr[15495] = -653051723;
assign addr[15496] = -634808946;
assign addr[15497] = -616515832;
assign addr[15498] = -598173833;
assign addr[15499] = -579784402;
assign addr[15500] = -561348998;
assign addr[15501] = -542869083;
assign addr[15502] = -524346121;
assign addr[15503] = -505781581;
assign addr[15504] = -487176937;
assign addr[15505] = -468533662;
assign addr[15506] = -449853235;
assign addr[15507] = -431137138;
assign addr[15508] = -412386854;
assign addr[15509] = -393603870;
assign addr[15510] = -374789676;
assign addr[15511] = -355945764;
assign addr[15512] = -337073627;
assign addr[15513] = -318174762;
assign addr[15514] = -299250668;
assign addr[15515] = -280302845;
assign addr[15516] = -261332796;
assign addr[15517] = -242342025;
assign addr[15518] = -223332037;
assign addr[15519] = -204304341;
assign addr[15520] = -185260444;
assign addr[15521] = -166201858;
assign addr[15522] = -147130093;
assign addr[15523] = -128046661;
assign addr[15524] = -108953076;
assign addr[15525] = -89850852;
assign addr[15526] = -70741503;
assign addr[15527] = -51626544;
assign addr[15528] = -32507492;
assign addr[15529] = -13385863;
assign addr[15530] = 5736829;
assign addr[15531] = 24859065;
assign addr[15532] = 43979330;
assign addr[15533] = 63096108;
assign addr[15534] = 82207882;
assign addr[15535] = 101313138;
assign addr[15536] = 120410361;
assign addr[15537] = 139498035;
assign addr[15538] = 158574649;
assign addr[15539] = 177638688;
assign addr[15540] = 196688642;
assign addr[15541] = 215722999;
assign addr[15542] = 234740251;
assign addr[15543] = 253738890;
assign addr[15544] = 272717408;
assign addr[15545] = 291674302;
assign addr[15546] = 310608068;
assign addr[15547] = 329517204;
assign addr[15548] = 348400212;
assign addr[15549] = 367255594;
assign addr[15550] = 386081854;
assign addr[15551] = 404877501;
assign addr[15552] = 423641043;
assign addr[15553] = 442370993;
assign addr[15554] = 461065866;
assign addr[15555] = 479724180;
assign addr[15556] = 498344454;
assign addr[15557] = 516925212;
assign addr[15558] = 535464981;
assign addr[15559] = 553962291;
assign addr[15560] = 572415676;
assign addr[15561] = 590823671;
assign addr[15562] = 609184818;
assign addr[15563] = 627497660;
assign addr[15564] = 645760745;
assign addr[15565] = 663972625;
assign addr[15566] = 682131857;
assign addr[15567] = 700236999;
assign addr[15568] = 718286617;
assign addr[15569] = 736279279;
assign addr[15570] = 754213559;
assign addr[15571] = 772088034;
assign addr[15572] = 789901288;
assign addr[15573] = 807651907;
assign addr[15574] = 825338484;
assign addr[15575] = 842959617;
assign addr[15576] = 860513908;
assign addr[15577] = 877999966;
assign addr[15578] = 895416404;
assign addr[15579] = 912761841;
assign addr[15580] = 930034901;
assign addr[15581] = 947234215;
assign addr[15582] = 964358420;
assign addr[15583] = 981406156;
assign addr[15584] = 998376073;
assign addr[15585] = 1015266825;
assign addr[15586] = 1032077073;
assign addr[15587] = 1048805483;
assign addr[15588] = 1065450729;
assign addr[15589] = 1082011492;
assign addr[15590] = 1098486458;
assign addr[15591] = 1114874320;
assign addr[15592] = 1131173780;
assign addr[15593] = 1147383544;
assign addr[15594] = 1163502328;
assign addr[15595] = 1179528853;
assign addr[15596] = 1195461849;
assign addr[15597] = 1211300053;
assign addr[15598] = 1227042207;
assign addr[15599] = 1242687064;
assign addr[15600] = 1258233384;
assign addr[15601] = 1273679934;
assign addr[15602] = 1289025489;
assign addr[15603] = 1304268832;
assign addr[15604] = 1319408754;
assign addr[15605] = 1334444055;
assign addr[15606] = 1349373543;
assign addr[15607] = 1364196034;
assign addr[15608] = 1378910353;
assign addr[15609] = 1393515332;
assign addr[15610] = 1408009814;
assign addr[15611] = 1422392650;
assign addr[15612] = 1436662698;
assign addr[15613] = 1450818828;
assign addr[15614] = 1464859917;
assign addr[15615] = 1478784851;
assign addr[15616] = 1492592527;
assign addr[15617] = 1506281850;
assign addr[15618] = 1519851733;
assign addr[15619] = 1533301101;
assign addr[15620] = 1546628888;
assign addr[15621] = 1559834037;
assign addr[15622] = 1572915501;
assign addr[15623] = 1585872242;
assign addr[15624] = 1598703233;
assign addr[15625] = 1611407456;
assign addr[15626] = 1623983905;
assign addr[15627] = 1636431582;
assign addr[15628] = 1648749499;
assign addr[15629] = 1660936681;
assign addr[15630] = 1672992161;
assign addr[15631] = 1684914983;
assign addr[15632] = 1696704201;
assign addr[15633] = 1708358881;
assign addr[15634] = 1719878099;
assign addr[15635] = 1731260941;
assign addr[15636] = 1742506504;
assign addr[15637] = 1753613897;
assign addr[15638] = 1764582240;
assign addr[15639] = 1775410662;
assign addr[15640] = 1786098304;
assign addr[15641] = 1796644320;
assign addr[15642] = 1807047873;
assign addr[15643] = 1817308138;
assign addr[15644] = 1827424302;
assign addr[15645] = 1837395562;
assign addr[15646] = 1847221128;
assign addr[15647] = 1856900221;
assign addr[15648] = 1866432072;
assign addr[15649] = 1875815927;
assign addr[15650] = 1885051042;
assign addr[15651] = 1894136683;
assign addr[15652] = 1903072131;
assign addr[15653] = 1911856677;
assign addr[15654] = 1920489624;
assign addr[15655] = 1928970288;
assign addr[15656] = 1937297997;
assign addr[15657] = 1945472089;
assign addr[15658] = 1953491918;
assign addr[15659] = 1961356847;
assign addr[15660] = 1969066252;
assign addr[15661] = 1976619522;
assign addr[15662] = 1984016058;
assign addr[15663] = 1991255274;
assign addr[15664] = 1998336596;
assign addr[15665] = 2005259462;
assign addr[15666] = 2012023322;
assign addr[15667] = 2018627642;
assign addr[15668] = 2025071897;
assign addr[15669] = 2031355576;
assign addr[15670] = 2037478181;
assign addr[15671] = 2043439226;
assign addr[15672] = 2049238240;
assign addr[15673] = 2054874761;
assign addr[15674] = 2060348343;
assign addr[15675] = 2065658552;
assign addr[15676] = 2070804967;
assign addr[15677] = 2075787180;
assign addr[15678] = 2080604795;
assign addr[15679] = 2085257431;
assign addr[15680] = 2089744719;
assign addr[15681] = 2094066304;
assign addr[15682] = 2098221841;
assign addr[15683] = 2102211002;
assign addr[15684] = 2106033471;
assign addr[15685] = 2109688944;
assign addr[15686] = 2113177132;
assign addr[15687] = 2116497758;
assign addr[15688] = 2119650558;
assign addr[15689] = 2122635283;
assign addr[15690] = 2125451696;
assign addr[15691] = 2128099574;
assign addr[15692] = 2130578706;
assign addr[15693] = 2132888897;
assign addr[15694] = 2135029962;
assign addr[15695] = 2137001733;
assign addr[15696] = 2138804053;
assign addr[15697] = 2140436778;
assign addr[15698] = 2141899780;
assign addr[15699] = 2143192942;
assign addr[15700] = 2144316162;
assign addr[15701] = 2145269351;
assign addr[15702] = 2146052433;
assign addr[15703] = 2146665347;
assign addr[15704] = 2147108043;
assign addr[15705] = 2147380486;
assign addr[15706] = 2147482655;
assign addr[15707] = 2147414542;
assign addr[15708] = 2147176152;
assign addr[15709] = 2146767505;
assign addr[15710] = 2146188631;
assign addr[15711] = 2145439578;
assign addr[15712] = 2144520405;
assign addr[15713] = 2143431184;
assign addr[15714] = 2142172003;
assign addr[15715] = 2140742960;
assign addr[15716] = 2139144169;
assign addr[15717] = 2137375758;
assign addr[15718] = 2135437865;
assign addr[15719] = 2133330646;
assign addr[15720] = 2131054266;
assign addr[15721] = 2128608907;
assign addr[15722] = 2125994762;
assign addr[15723] = 2123212038;
assign addr[15724] = 2120260957;
assign addr[15725] = 2117141752;
assign addr[15726] = 2113854671;
assign addr[15727] = 2110399974;
assign addr[15728] = 2106777935;
assign addr[15729] = 2102988841;
assign addr[15730] = 2099032994;
assign addr[15731] = 2094910706;
assign addr[15732] = 2090622304;
assign addr[15733] = 2086168128;
assign addr[15734] = 2081548533;
assign addr[15735] = 2076763883;
assign addr[15736] = 2071814558;
assign addr[15737] = 2066700952;
assign addr[15738] = 2061423468;
assign addr[15739] = 2055982526;
assign addr[15740] = 2050378558;
assign addr[15741] = 2044612007;
assign addr[15742] = 2038683330;
assign addr[15743] = 2032592999;
assign addr[15744] = 2026341495;
assign addr[15745] = 2019929315;
assign addr[15746] = 2013356967;
assign addr[15747] = 2006624971;
assign addr[15748] = 1999733863;
assign addr[15749] = 1992684188;
assign addr[15750] = 1985476506;
assign addr[15751] = 1978111387;
assign addr[15752] = 1970589416;
assign addr[15753] = 1962911189;
assign addr[15754] = 1955077316;
assign addr[15755] = 1947088417;
assign addr[15756] = 1938945125;
assign addr[15757] = 1930648088;
assign addr[15758] = 1922197961;
assign addr[15759] = 1913595416;
assign addr[15760] = 1904841135;
assign addr[15761] = 1895935811;
assign addr[15762] = 1886880151;
assign addr[15763] = 1877674873;
assign addr[15764] = 1868320707;
assign addr[15765] = 1858818395;
assign addr[15766] = 1849168689;
assign addr[15767] = 1839372356;
assign addr[15768] = 1829430172;
assign addr[15769] = 1819342925;
assign addr[15770] = 1809111415;
assign addr[15771] = 1798736454;
assign addr[15772] = 1788218865;
assign addr[15773] = 1777559480;
assign addr[15774] = 1766759146;
assign addr[15775] = 1755818718;
assign addr[15776] = 1744739065;
assign addr[15777] = 1733521064;
assign addr[15778] = 1722165606;
assign addr[15779] = 1710673591;
assign addr[15780] = 1699045930;
assign addr[15781] = 1687283545;
assign addr[15782] = 1675387369;
assign addr[15783] = 1663358344;
assign addr[15784] = 1651197426;
assign addr[15785] = 1638905577;
assign addr[15786] = 1626483774;
assign addr[15787] = 1613933000;
assign addr[15788] = 1601254251;
assign addr[15789] = 1588448533;
assign addr[15790] = 1575516860;
assign addr[15791] = 1562460258;
assign addr[15792] = 1549279763;
assign addr[15793] = 1535976419;
assign addr[15794] = 1522551282;
assign addr[15795] = 1509005416;
assign addr[15796] = 1495339895;
assign addr[15797] = 1481555802;
assign addr[15798] = 1467654232;
assign addr[15799] = 1453636285;
assign addr[15800] = 1439503074;
assign addr[15801] = 1425255719;
assign addr[15802] = 1410895350;
assign addr[15803] = 1396423105;
assign addr[15804] = 1381840133;
assign addr[15805] = 1367147589;
assign addr[15806] = 1352346639;
assign addr[15807] = 1337438456;
assign addr[15808] = 1322424222;
assign addr[15809] = 1307305128;
assign addr[15810] = 1292082373;
assign addr[15811] = 1276757164;
assign addr[15812] = 1261330715;
assign addr[15813] = 1245804251;
assign addr[15814] = 1230179002;
assign addr[15815] = 1214456207;
assign addr[15816] = 1198637114;
assign addr[15817] = 1182722976;
assign addr[15818] = 1166715055;
assign addr[15819] = 1150614620;
assign addr[15820] = 1134422949;
assign addr[15821] = 1118141326;
assign addr[15822] = 1101771040;
assign addr[15823] = 1085313391;
assign addr[15824] = 1068769683;
assign addr[15825] = 1052141228;
assign addr[15826] = 1035429345;
assign addr[15827] = 1018635358;
assign addr[15828] = 1001760600;
assign addr[15829] = 984806408;
assign addr[15830] = 967774128;
assign addr[15831] = 950665109;
assign addr[15832] = 933480707;
assign addr[15833] = 916222287;
assign addr[15834] = 898891215;
assign addr[15835] = 881488868;
assign addr[15836] = 864016623;
assign addr[15837] = 846475867;
assign addr[15838] = 828867991;
assign addr[15839] = 811194391;
assign addr[15840] = 793456467;
assign addr[15841] = 775655628;
assign addr[15842] = 757793284;
assign addr[15843] = 739870851;
assign addr[15844] = 721889752;
assign addr[15845] = 703851410;
assign addr[15846] = 685757258;
assign addr[15847] = 667608730;
assign addr[15848] = 649407264;
assign addr[15849] = 631154304;
assign addr[15850] = 612851297;
assign addr[15851] = 594499695;
assign addr[15852] = 576100953;
assign addr[15853] = 557656529;
assign addr[15854] = 539167887;
assign addr[15855] = 520636492;
assign addr[15856] = 502063814;
assign addr[15857] = 483451325;
assign addr[15858] = 464800501;
assign addr[15859] = 446112822;
assign addr[15860] = 427389768;
assign addr[15861] = 408632825;
assign addr[15862] = 389843480;
assign addr[15863] = 371023223;
assign addr[15864] = 352173546;
assign addr[15865] = 333295944;
assign addr[15866] = 314391913;
assign addr[15867] = 295462954;
assign addr[15868] = 276510565;
assign addr[15869] = 257536251;
assign addr[15870] = 238541516;
assign addr[15871] = 219527866;
assign addr[15872] = 200496809;
assign addr[15873] = 181449854;
assign addr[15874] = 162388511;
assign addr[15875] = 143314291;
assign addr[15876] = 124228708;
assign addr[15877] = 105133274;
assign addr[15878] = 86029503;
assign addr[15879] = 66918911;
assign addr[15880] = 47803013;
assign addr[15881] = 28683324;
assign addr[15882] = 9561361;
assign addr[15883] = -9561361;
assign addr[15884] = -28683324;
assign addr[15885] = -47803013;
assign addr[15886] = -66918911;
assign addr[15887] = -86029503;
assign addr[15888] = -105133274;
assign addr[15889] = -124228708;
assign addr[15890] = -143314291;
assign addr[15891] = -162388511;
assign addr[15892] = -181449854;
assign addr[15893] = -200496809;
assign addr[15894] = -219527866;
assign addr[15895] = -238541516;
assign addr[15896] = -257536251;
assign addr[15897] = -276510565;
assign addr[15898] = -295462954;
assign addr[15899] = -314391913;
assign addr[15900] = -333295944;
assign addr[15901] = -352173546;
assign addr[15902] = -371023223;
assign addr[15903] = -389843480;
assign addr[15904] = -408632825;
assign addr[15905] = -427389768;
assign addr[15906] = -446112822;
assign addr[15907] = -464800501;
assign addr[15908] = -483451325;
assign addr[15909] = -502063814;
assign addr[15910] = -520636492;
assign addr[15911] = -539167887;
assign addr[15912] = -557656529;
assign addr[15913] = -576100953;
assign addr[15914] = -594499695;
assign addr[15915] = -612851297;
assign addr[15916] = -631154304;
assign addr[15917] = -649407264;
assign addr[15918] = -667608730;
assign addr[15919] = -685757258;
assign addr[15920] = -703851410;
assign addr[15921] = -721889752;
assign addr[15922] = -739870851;
assign addr[15923] = -757793284;
assign addr[15924] = -775655628;
assign addr[15925] = -793456467;
assign addr[15926] = -811194391;
assign addr[15927] = -828867991;
assign addr[15928] = -846475867;
assign addr[15929] = -864016623;
assign addr[15930] = -881488868;
assign addr[15931] = -898891215;
assign addr[15932] = -916222287;
assign addr[15933] = -933480707;
assign addr[15934] = -950665109;
assign addr[15935] = -967774128;
assign addr[15936] = -984806408;
assign addr[15937] = -1001760600;
assign addr[15938] = -1018635358;
assign addr[15939] = -1035429345;
assign addr[15940] = -1052141228;
assign addr[15941] = -1068769683;
assign addr[15942] = -1085313391;
assign addr[15943] = -1101771040;
assign addr[15944] = -1118141326;
assign addr[15945] = -1134422949;
assign addr[15946] = -1150614620;
assign addr[15947] = -1166715055;
assign addr[15948] = -1182722976;
assign addr[15949] = -1198637114;
assign addr[15950] = -1214456207;
assign addr[15951] = -1230179002;
assign addr[15952] = -1245804251;
assign addr[15953] = -1261330715;
assign addr[15954] = -1276757164;
assign addr[15955] = -1292082373;
assign addr[15956] = -1307305128;
assign addr[15957] = -1322424222;
assign addr[15958] = -1337438456;
assign addr[15959] = -1352346639;
assign addr[15960] = -1367147589;
assign addr[15961] = -1381840133;
assign addr[15962] = -1396423105;
assign addr[15963] = -1410895350;
assign addr[15964] = -1425255719;
assign addr[15965] = -1439503074;
assign addr[15966] = -1453636285;
assign addr[15967] = -1467654232;
assign addr[15968] = -1481555802;
assign addr[15969] = -1495339895;
assign addr[15970] = -1509005416;
assign addr[15971] = -1522551282;
assign addr[15972] = -1535976419;
assign addr[15973] = -1549279763;
assign addr[15974] = -1562460258;
assign addr[15975] = -1575516860;
assign addr[15976] = -1588448533;
assign addr[15977] = -1601254251;
assign addr[15978] = -1613933000;
assign addr[15979] = -1626483774;
assign addr[15980] = -1638905577;
assign addr[15981] = -1651197426;
assign addr[15982] = -1663358344;
assign addr[15983] = -1675387369;
assign addr[15984] = -1687283545;
assign addr[15985] = -1699045930;
assign addr[15986] = -1710673591;
assign addr[15987] = -1722165606;
assign addr[15988] = -1733521064;
assign addr[15989] = -1744739065;
assign addr[15990] = -1755818718;
assign addr[15991] = -1766759146;
assign addr[15992] = -1777559480;
assign addr[15993] = -1788218865;
assign addr[15994] = -1798736454;
assign addr[15995] = -1809111415;
assign addr[15996] = -1819342925;
assign addr[15997] = -1829430172;
assign addr[15998] = -1839372356;
assign addr[15999] = -1849168689;
assign addr[16000] = -1858818395;
assign addr[16001] = -1868320707;
assign addr[16002] = -1877674873;
assign addr[16003] = -1886880151;
assign addr[16004] = -1895935811;
assign addr[16005] = -1904841135;
assign addr[16006] = -1913595416;
assign addr[16007] = -1922197961;
assign addr[16008] = -1930648088;
assign addr[16009] = -1938945125;
assign addr[16010] = -1947088417;
assign addr[16011] = -1955077316;
assign addr[16012] = -1962911189;
assign addr[16013] = -1970589416;
assign addr[16014] = -1978111387;
assign addr[16015] = -1985476506;
assign addr[16016] = -1992684188;
assign addr[16017] = -1999733863;
assign addr[16018] = -2006624971;
assign addr[16019] = -2013356967;
assign addr[16020] = -2019929315;
assign addr[16021] = -2026341495;
assign addr[16022] = -2032592999;
assign addr[16023] = -2038683330;
assign addr[16024] = -2044612007;
assign addr[16025] = -2050378558;
assign addr[16026] = -2055982526;
assign addr[16027] = -2061423468;
assign addr[16028] = -2066700952;
assign addr[16029] = -2071814558;
assign addr[16030] = -2076763883;
assign addr[16031] = -2081548533;
assign addr[16032] = -2086168128;
assign addr[16033] = -2090622304;
assign addr[16034] = -2094910706;
assign addr[16035] = -2099032994;
assign addr[16036] = -2102988841;
assign addr[16037] = -2106777935;
assign addr[16038] = -2110399974;
assign addr[16039] = -2113854671;
assign addr[16040] = -2117141752;
assign addr[16041] = -2120260957;
assign addr[16042] = -2123212038;
assign addr[16043] = -2125994762;
assign addr[16044] = -2128608907;
assign addr[16045] = -2131054266;
assign addr[16046] = -2133330646;
assign addr[16047] = -2135437865;
assign addr[16048] = -2137375758;
assign addr[16049] = -2139144169;
assign addr[16050] = -2140742960;
assign addr[16051] = -2142172003;
assign addr[16052] = -2143431184;
assign addr[16053] = -2144520405;
assign addr[16054] = -2145439578;
assign addr[16055] = -2146188631;
assign addr[16056] = -2146767505;
assign addr[16057] = -2147176152;
assign addr[16058] = -2147414542;
assign addr[16059] = -2147482655;
assign addr[16060] = -2147380486;
assign addr[16061] = -2147108043;
assign addr[16062] = -2146665347;
assign addr[16063] = -2146052433;
assign addr[16064] = -2145269351;
assign addr[16065] = -2144316162;
assign addr[16066] = -2143192942;
assign addr[16067] = -2141899780;
assign addr[16068] = -2140436778;
assign addr[16069] = -2138804053;
assign addr[16070] = -2137001733;
assign addr[16071] = -2135029962;
assign addr[16072] = -2132888897;
assign addr[16073] = -2130578706;
assign addr[16074] = -2128099574;
assign addr[16075] = -2125451696;
assign addr[16076] = -2122635283;
assign addr[16077] = -2119650558;
assign addr[16078] = -2116497758;
assign addr[16079] = -2113177132;
assign addr[16080] = -2109688944;
assign addr[16081] = -2106033471;
assign addr[16082] = -2102211002;
assign addr[16083] = -2098221841;
assign addr[16084] = -2094066304;
assign addr[16085] = -2089744719;
assign addr[16086] = -2085257431;
assign addr[16087] = -2080604795;
assign addr[16088] = -2075787180;
assign addr[16089] = -2070804967;
assign addr[16090] = -2065658552;
assign addr[16091] = -2060348343;
assign addr[16092] = -2054874761;
assign addr[16093] = -2049238240;
assign addr[16094] = -2043439226;
assign addr[16095] = -2037478181;
assign addr[16096] = -2031355576;
assign addr[16097] = -2025071897;
assign addr[16098] = -2018627642;
assign addr[16099] = -2012023322;
assign addr[16100] = -2005259462;
assign addr[16101] = -1998336596;
assign addr[16102] = -1991255274;
assign addr[16103] = -1984016058;
assign addr[16104] = -1976619522;
assign addr[16105] = -1969066252;
assign addr[16106] = -1961356847;
assign addr[16107] = -1953491918;
assign addr[16108] = -1945472089;
assign addr[16109] = -1937297997;
assign addr[16110] = -1928970288;
assign addr[16111] = -1920489624;
assign addr[16112] = -1911856677;
assign addr[16113] = -1903072131;
assign addr[16114] = -1894136683;
assign addr[16115] = -1885051042;
assign addr[16116] = -1875815927;
assign addr[16117] = -1866432072;
assign addr[16118] = -1856900221;
assign addr[16119] = -1847221128;
assign addr[16120] = -1837395562;
assign addr[16121] = -1827424302;
assign addr[16122] = -1817308138;
assign addr[16123] = -1807047873;
assign addr[16124] = -1796644320;
assign addr[16125] = -1786098304;
assign addr[16126] = -1775410662;
assign addr[16127] = -1764582240;
assign addr[16128] = -1753613897;
assign addr[16129] = -1742506504;
assign addr[16130] = -1731260941;
assign addr[16131] = -1719878099;
assign addr[16132] = -1708358881;
assign addr[16133] = -1696704201;
assign addr[16134] = -1684914983;
assign addr[16135] = -1672992161;
assign addr[16136] = -1660936681;
assign addr[16137] = -1648749499;
assign addr[16138] = -1636431582;
assign addr[16139] = -1623983905;
assign addr[16140] = -1611407456;
assign addr[16141] = -1598703233;
assign addr[16142] = -1585872242;
assign addr[16143] = -1572915501;
assign addr[16144] = -1559834037;
assign addr[16145] = -1546628888;
assign addr[16146] = -1533301101;
assign addr[16147] = -1519851733;
assign addr[16148] = -1506281850;
assign addr[16149] = -1492592527;
assign addr[16150] = -1478784851;
assign addr[16151] = -1464859917;
assign addr[16152] = -1450818828;
assign addr[16153] = -1436662698;
assign addr[16154] = -1422392650;
assign addr[16155] = -1408009814;
assign addr[16156] = -1393515332;
assign addr[16157] = -1378910353;
assign addr[16158] = -1364196034;
assign addr[16159] = -1349373543;
assign addr[16160] = -1334444055;
assign addr[16161] = -1319408754;
assign addr[16162] = -1304268832;
assign addr[16163] = -1289025489;
assign addr[16164] = -1273679934;
assign addr[16165] = -1258233384;
assign addr[16166] = -1242687064;
assign addr[16167] = -1227042207;
assign addr[16168] = -1211300053;
assign addr[16169] = -1195461849;
assign addr[16170] = -1179528853;
assign addr[16171] = -1163502328;
assign addr[16172] = -1147383544;
assign addr[16173] = -1131173780;
assign addr[16174] = -1114874320;
assign addr[16175] = -1098486458;
assign addr[16176] = -1082011492;
assign addr[16177] = -1065450729;
assign addr[16178] = -1048805483;
assign addr[16179] = -1032077073;
assign addr[16180] = -1015266825;
assign addr[16181] = -998376073;
assign addr[16182] = -981406156;
assign addr[16183] = -964358420;
assign addr[16184] = -947234215;
assign addr[16185] = -930034901;
assign addr[16186] = -912761841;
assign addr[16187] = -895416404;
assign addr[16188] = -877999966;
assign addr[16189] = -860513908;
assign addr[16190] = -842959617;
assign addr[16191] = -825338484;
assign addr[16192] = -807651907;
assign addr[16193] = -789901288;
assign addr[16194] = -772088034;
assign addr[16195] = -754213559;
assign addr[16196] = -736279279;
assign addr[16197] = -718286617;
assign addr[16198] = -700236999;
assign addr[16199] = -682131857;
assign addr[16200] = -663972625;
assign addr[16201] = -645760745;
assign addr[16202] = -627497660;
assign addr[16203] = -609184818;
assign addr[16204] = -590823671;
assign addr[16205] = -572415676;
assign addr[16206] = -553962291;
assign addr[16207] = -535464981;
assign addr[16208] = -516925212;
assign addr[16209] = -498344454;
assign addr[16210] = -479724180;
assign addr[16211] = -461065866;
assign addr[16212] = -442370993;
assign addr[16213] = -423641043;
assign addr[16214] = -404877501;
assign addr[16215] = -386081854;
assign addr[16216] = -367255594;
assign addr[16217] = -348400212;
assign addr[16218] = -329517204;
assign addr[16219] = -310608068;
assign addr[16220] = -291674302;
assign addr[16221] = -272717408;
assign addr[16222] = -253738890;
assign addr[16223] = -234740251;
assign addr[16224] = -215722999;
assign addr[16225] = -196688642;
assign addr[16226] = -177638688;
assign addr[16227] = -158574649;
assign addr[16228] = -139498035;
assign addr[16229] = -120410361;
assign addr[16230] = -101313138;
assign addr[16231] = -82207882;
assign addr[16232] = -63096108;
assign addr[16233] = -43979330;
assign addr[16234] = -24859065;
assign addr[16235] = -5736829;
assign addr[16236] = 13385863;
assign addr[16237] = 32507492;
assign addr[16238] = 51626544;
assign addr[16239] = 70741503;
assign addr[16240] = 89850852;
assign addr[16241] = 108953076;
assign addr[16242] = 128046661;
assign addr[16243] = 147130093;
assign addr[16244] = 166201858;
assign addr[16245] = 185260444;
assign addr[16246] = 204304341;
assign addr[16247] = 223332037;
assign addr[16248] = 242342025;
assign addr[16249] = 261332796;
assign addr[16250] = 280302845;
assign addr[16251] = 299250668;
assign addr[16252] = 318174762;
assign addr[16253] = 337073627;
assign addr[16254] = 355945764;
assign addr[16255] = 374789676;
assign addr[16256] = 393603870;
assign addr[16257] = 412386854;
assign addr[16258] = 431137138;
assign addr[16259] = 449853235;
assign addr[16260] = 468533662;
assign addr[16261] = 487176937;
assign addr[16262] = 505781581;
assign addr[16263] = 524346121;
assign addr[16264] = 542869083;
assign addr[16265] = 561348998;
assign addr[16266] = 579784402;
assign addr[16267] = 598173833;
assign addr[16268] = 616515832;
assign addr[16269] = 634808946;
assign addr[16270] = 653051723;
assign addr[16271] = 671242716;
assign addr[16272] = 689380485;
assign addr[16273] = 707463589;
assign addr[16274] = 725490597;
assign addr[16275] = 743460077;
assign addr[16276] = 761370605;
assign addr[16277] = 779220762;
assign addr[16278] = 797009130;
assign addr[16279] = 814734301;
assign addr[16280] = 832394869;
assign addr[16281] = 849989433;
assign addr[16282] = 867516597;
assign addr[16283] = 884974973;
assign addr[16284] = 902363176;
assign addr[16285] = 919679827;
assign addr[16286] = 936923553;
assign addr[16287] = 954092986;
assign addr[16288] = 971186766;
assign addr[16289] = 988203537;
assign addr[16290] = 1005141949;
assign addr[16291] = 1022000660;
assign addr[16292] = 1038778332;
assign addr[16293] = 1055473635;
assign addr[16294] = 1072085246;
assign addr[16295] = 1088611847;
assign addr[16296] = 1105052128;
assign addr[16297] = 1121404785;
assign addr[16298] = 1137668521;
assign addr[16299] = 1153842047;
assign addr[16300] = 1169924081;
assign addr[16301] = 1185913346;
assign addr[16302] = 1201808576;
assign addr[16303] = 1217608510;
assign addr[16304] = 1233311895;
assign addr[16305] = 1248917486;
assign addr[16306] = 1264424045;
assign addr[16307] = 1279830344;
assign addr[16308] = 1295135159;
assign addr[16309] = 1310337279;
assign addr[16310] = 1325435496;
assign addr[16311] = 1340428615;
assign addr[16312] = 1355315445;
assign addr[16313] = 1370094808;
assign addr[16314] = 1384765530;
assign addr[16315] = 1399326449;
assign addr[16316] = 1413776410;
assign addr[16317] = 1428114267;
assign addr[16318] = 1442338884;
assign addr[16319] = 1456449131;
assign addr[16320] = 1470443891;
assign addr[16321] = 1484322054;
assign addr[16322] = 1498082520;
assign addr[16323] = 1511724196;
assign addr[16324] = 1525246002;
assign addr[16325] = 1538646865;
assign addr[16326] = 1551925723;
assign addr[16327] = 1565081523;
assign addr[16328] = 1578113222;
assign addr[16329] = 1591019785;
assign addr[16330] = 1603800191;
assign addr[16331] = 1616453425;
assign addr[16332] = 1628978484;
assign addr[16333] = 1641374375;
assign addr[16334] = 1653640115;
assign addr[16335] = 1665774731;
assign addr[16336] = 1677777262;
assign addr[16337] = 1689646755;
assign addr[16338] = 1701382270;
assign addr[16339] = 1712982875;
assign addr[16340] = 1724447652;
assign addr[16341] = 1735775690;
assign addr[16342] = 1746966091;
assign addr[16343] = 1758017969;
assign addr[16344] = 1768930447;
assign addr[16345] = 1779702660;
assign addr[16346] = 1790333753;
assign addr[16347] = 1800822883;
assign addr[16348] = 1811169220;
assign addr[16349] = 1821371941;
assign addr[16350] = 1831430239;
assign addr[16351] = 1841343316;
assign addr[16352] = 1851110385;
assign addr[16353] = 1860730673;
assign addr[16354] = 1870203416;
assign addr[16355] = 1879527863;
assign addr[16356] = 1888703276;
assign addr[16357] = 1897728925;
assign addr[16358] = 1906604097;
assign addr[16359] = 1915328086;
assign addr[16360] = 1923900201;
assign addr[16361] = 1932319763;
assign addr[16362] = 1940586104;
assign addr[16363] = 1948698568;
assign addr[16364] = 1956656513;
assign addr[16365] = 1964459306;
assign addr[16366] = 1972106330;
assign addr[16367] = 1979596978;
assign addr[16368] = 1986930656;
assign addr[16369] = 1994106782;
assign addr[16370] = 2001124788;
assign addr[16371] = 2007984117;
assign addr[16372] = 2014684225;
assign addr[16373] = 2021224581;
assign addr[16374] = 2027604666;
assign addr[16375] = 2033823974;
assign addr[16376] = 2039882013;
assign addr[16377] = 2045778302;
assign addr[16378] = 2051512372;
assign addr[16379] = 2057083771;
assign addr[16380] = 2062492055;
assign addr[16381] = 2067736796;
assign addr[16382] = 2072817579;
assign addr[16383] = 2077733999;
assign addr[16384] = 2082485668;
assign addr[16385] = 2087072209;
assign addr[16386] = 2091493257;
assign addr[16387] = 2095748463;
assign addr[16388] = 2099837489;
assign addr[16389] = 2103760010;
assign addr[16390] = 2107515716;
assign addr[16391] = 2111104309;
assign addr[16392] = 2114525505;
assign addr[16393] = 2117779031;
assign addr[16394] = 2120864631;
assign addr[16395] = 2123782059;
assign addr[16396] = 2126531084;
assign addr[16397] = 2129111488;
assign addr[16398] = 2131523066;
assign addr[16399] = 2133765628;
assign addr[16400] = 2135838995;
assign addr[16401] = 2137743003;
assign addr[16402] = 2139477502;
assign addr[16403] = 2141042352;
assign addr[16404] = 2142437431;
assign addr[16405] = 2143662628;
assign addr[16406] = 2144717846;
assign addr[16407] = 2145603001;
assign addr[16408] = 2146318022;
assign addr[16409] = 2146862854;
assign addr[16410] = 2147237452;
assign addr[16411] = 2147441787;
assign addr[16412] = 2147475844;
assign addr[16413] = 2147339619;
assign addr[16414] = 2147033123;
assign addr[16415] = 2146556380;
assign addr[16416] = 2145909429;
assign addr[16417] = 2145092320;
assign addr[16418] = 2144105118;
assign addr[16419] = 2142947902;
assign addr[16420] = 2141620763;
assign addr[16421] = 2140123807;
assign addr[16422] = 2138457152;
assign addr[16423] = 2136620930;
assign addr[16424] = 2134615288;
assign addr[16425] = 2132440383;
assign addr[16426] = 2130096389;
assign addr[16427] = 2127583492;
assign addr[16428] = 2124901890;
assign addr[16429] = 2122051796;
assign addr[16430] = 2119033436;
assign addr[16431] = 2115847050;
assign addr[16432] = 2112492891;
assign addr[16433] = 2108971223;
assign addr[16434] = 2105282327;
assign addr[16435] = 2101426496;
assign addr[16436] = 2097404033;
assign addr[16437] = 2093215260;
assign addr[16438] = 2088860507;
assign addr[16439] = 2084340120;
assign addr[16440] = 2079654458;
assign addr[16441] = 2074803892;
assign addr[16442] = 2069788807;
assign addr[16443] = 2064609600;
assign addr[16444] = 2059266683;
assign addr[16445] = 2053760478;
assign addr[16446] = 2048091422;
assign addr[16447] = 2042259965;
assign addr[16448] = 2036266570;
assign addr[16449] = 2030111710;
assign addr[16450] = 2023795876;
assign addr[16451] = 2017319567;
assign addr[16452] = 2010683297;
assign addr[16453] = 2003887591;
assign addr[16454] = 1996932990;
assign addr[16455] = 1989820044;
assign addr[16456] = 1982549318;
assign addr[16457] = 1975121388;
assign addr[16458] = 1967536842;
assign addr[16459] = 1959796283;
assign addr[16460] = 1951900324;
assign addr[16461] = 1943849591;
assign addr[16462] = 1935644723;
assign addr[16463] = 1927286370;
assign addr[16464] = 1918775195;
assign addr[16465] = 1910111873;
assign addr[16466] = 1901297091;
assign addr[16467] = 1892331547;
assign addr[16468] = 1883215953;
assign addr[16469] = 1873951032;
assign addr[16470] = 1864537518;
assign addr[16471] = 1854976157;
assign addr[16472] = 1845267708;
assign addr[16473] = 1835412941;
assign addr[16474] = 1825412636;
assign addr[16475] = 1815267588;
assign addr[16476] = 1804978599;
assign addr[16477] = 1794546487;
assign addr[16478] = 1783972079;
assign addr[16479] = 1773256212;
assign addr[16480] = 1762399737;
assign addr[16481] = 1751403515;
assign addr[16482] = 1740268417;
assign addr[16483] = 1728995326;
assign addr[16484] = 1717585136;
assign addr[16485] = 1706038753;
assign addr[16486] = 1694357091;
assign addr[16487] = 1682541077;
assign addr[16488] = 1670591647;
assign addr[16489] = 1658509750;
assign addr[16490] = 1646296344;
assign addr[16491] = 1633952396;
assign addr[16492] = 1621478885;
assign addr[16493] = 1608876801;
assign addr[16494] = 1596147143;
assign addr[16495] = 1583290921;
assign addr[16496] = 1570309153;
assign addr[16497] = 1557202869;
assign addr[16498] = 1543973108;
assign addr[16499] = 1530620920;
assign addr[16500] = 1517147363;
assign addr[16501] = 1503553506;
assign addr[16502] = 1489840425;
assign addr[16503] = 1476009210;
assign addr[16504] = 1462060956;
assign addr[16505] = 1447996770;
assign addr[16506] = 1433817766;
assign addr[16507] = 1419525069;
assign addr[16508] = 1405119813;
assign addr[16509] = 1390603139;
assign addr[16510] = 1375976199;
assign addr[16511] = 1361240152;
assign addr[16512] = 1346396168;
assign addr[16513] = 1331445422;
assign addr[16514] = 1316389101;
assign addr[16515] = 1301228398;
assign addr[16516] = 1285964516;
assign addr[16517] = 1270598665;
assign addr[16518] = 1255132063;
assign addr[16519] = 1239565936;
assign addr[16520] = 1223901520;
assign addr[16521] = 1208140056;
assign addr[16522] = 1192282793;
assign addr[16523] = 1176330990;
assign addr[16524] = 1160285911;
assign addr[16525] = 1144148829;
assign addr[16526] = 1127921022;
assign addr[16527] = 1111603778;
assign addr[16528] = 1095198391;
assign addr[16529] = 1078706161;
assign addr[16530] = 1062128397;
assign addr[16531] = 1045466412;
assign addr[16532] = 1028721528;
assign addr[16533] = 1011895073;
assign addr[16534] = 994988380;
assign addr[16535] = 978002791;
assign addr[16536] = 960939653;
assign addr[16537] = 943800318;
assign addr[16538] = 926586145;
assign addr[16539] = 909298500;
assign addr[16540] = 891938752;
assign addr[16541] = 874508280;
assign addr[16542] = 857008464;
assign addr[16543] = 839440693;
assign addr[16544] = 821806359;
assign addr[16545] = 804106861;
assign addr[16546] = 786343603;
assign addr[16547] = 768517992;
assign addr[16548] = 750631442;
assign addr[16549] = 732685372;
assign addr[16550] = 714681204;
assign addr[16551] = 696620367;
assign addr[16552] = 678504291;
assign addr[16553] = 660334415;
assign addr[16554] = 642112178;
assign addr[16555] = 623839025;
assign addr[16556] = 605516406;
assign addr[16557] = 587145773;
assign addr[16558] = 568728583;
assign addr[16559] = 550266296;
assign addr[16560] = 531760377;
assign addr[16561] = 513212292;
assign addr[16562] = 494623513;
assign addr[16563] = 475995513;
assign addr[16564] = 457329769;
assign addr[16565] = 438627762;
assign addr[16566] = 419890975;
assign addr[16567] = 401120892;
assign addr[16568] = 382319004;
assign addr[16569] = 363486799;
assign addr[16570] = 344625773;
assign addr[16571] = 325737419;
assign addr[16572] = 306823237;
assign addr[16573] = 287884725;
assign addr[16574] = 268923386;
assign addr[16575] = 249940723;
assign addr[16576] = 230938242;
assign addr[16577] = 211917448;
assign addr[16578] = 192879850;
assign addr[16579] = 173826959;
assign addr[16580] = 154760284;
assign addr[16581] = 135681337;
assign addr[16582] = 116591632;
assign addr[16583] = 97492681;
assign addr[16584] = 78386000;
assign addr[16585] = 59273104;
assign addr[16586] = 40155507;
assign addr[16587] = 21034727;
assign addr[16588] = 1912278;
assign addr[16589] = -17210322;
assign addr[16590] = -36331557;
assign addr[16591] = -55449912;
assign addr[16592] = -74563870;
assign addr[16593] = -93671915;
assign addr[16594] = -112772533;
assign addr[16595] = -131864208;
assign addr[16596] = -150945428;
assign addr[16597] = -170014678;
assign addr[16598] = -189070447;
assign addr[16599] = -208111224;
assign addr[16600] = -227135500;
assign addr[16601] = -246141764;
assign addr[16602] = -265128512;
assign addr[16603] = -284094236;
assign addr[16604] = -303037433;
assign addr[16605] = -321956601;
assign addr[16606] = -340850240;
assign addr[16607] = -359716852;
assign addr[16608] = -378554940;
assign addr[16609] = -397363011;
assign addr[16610] = -416139574;
assign addr[16611] = -434883140;
assign addr[16612] = -453592221;
assign addr[16613] = -472265336;
assign addr[16614] = -490901003;
assign addr[16615] = -509497745;
assign addr[16616] = -528054086;
assign addr[16617] = -546568556;
assign addr[16618] = -565039687;
assign addr[16619] = -583466013;
assign addr[16620] = -601846074;
assign addr[16621] = -620178412;
assign addr[16622] = -638461574;
assign addr[16623] = -656694110;
assign addr[16624] = -674874574;
assign addr[16625] = -693001525;
assign addr[16626] = -711073524;
assign addr[16627] = -729089140;
assign addr[16628] = -747046944;
assign addr[16629] = -764945512;
assign addr[16630] = -782783424;
assign addr[16631] = -800559266;
assign addr[16632] = -818271628;
assign addr[16633] = -835919107;
assign addr[16634] = -853500302;
assign addr[16635] = -871013820;
assign addr[16636] = -888458272;
assign addr[16637] = -905832274;
assign addr[16638] = -923134450;
assign addr[16639] = -940363427;
assign addr[16640] = -957517838;
assign addr[16641] = -974596324;
assign addr[16642] = -991597531;
assign addr[16643] = -1008520110;
assign addr[16644] = -1025362720;
assign addr[16645] = -1042124025;
assign addr[16646] = -1058802695;
assign addr[16647] = -1075397409;
assign addr[16648] = -1091906851;
assign addr[16649] = -1108329711;
assign addr[16650] = -1124664687;
assign addr[16651] = -1140910484;
assign addr[16652] = -1157065814;
assign addr[16653] = -1173129396;
assign addr[16654] = -1189099956;
assign addr[16655] = -1204976227;
assign addr[16656] = -1220756951;
assign addr[16657] = -1236440877;
assign addr[16658] = -1252026760;
assign addr[16659] = -1267513365;
assign addr[16660] = -1282899464;
assign addr[16661] = -1298183838;
assign addr[16662] = -1313365273;
assign addr[16663] = -1328442566;
assign addr[16664] = -1343414522;
assign addr[16665] = -1358279953;
assign addr[16666] = -1373037681;
assign addr[16667] = -1387686535;
assign addr[16668] = -1402225355;
assign addr[16669] = -1416652986;
assign addr[16670] = -1430968286;
assign addr[16671] = -1445170118;
assign addr[16672] = -1459257358;
assign addr[16673] = -1473228887;
assign addr[16674] = -1487083598;
assign addr[16675] = -1500820393;
assign addr[16676] = -1514438181;
assign addr[16677] = -1527935884;
assign addr[16678] = -1541312431;
assign addr[16679] = -1554566762;
assign addr[16680] = -1567697824;
assign addr[16681] = -1580704578;
assign addr[16682] = -1593585992;
assign addr[16683] = -1606341043;
assign addr[16684] = -1618968722;
assign addr[16685] = -1631468027;
assign addr[16686] = -1643837966;
assign addr[16687] = -1656077559;
assign addr[16688] = -1668185835;
assign addr[16689] = -1680161834;
assign addr[16690] = -1692004606;
assign addr[16691] = -1703713213;
assign addr[16692] = -1715286726;
assign addr[16693] = -1726724227;
assign addr[16694] = -1738024810;
assign addr[16695] = -1749187577;
assign addr[16696] = -1760211645;
assign addr[16697] = -1771096139;
assign addr[16698] = -1781840195;
assign addr[16699] = -1792442963;
assign addr[16700] = -1802903601;
assign addr[16701] = -1813221279;
assign addr[16702] = -1823395180;
assign addr[16703] = -1833424497;
assign addr[16704] = -1843308435;
assign addr[16705] = -1853046210;
assign addr[16706] = -1862637049;
assign addr[16707] = -1872080193;
assign addr[16708] = -1881374892;
assign addr[16709] = -1890520410;
assign addr[16710] = -1899516021;
assign addr[16711] = -1908361011;
assign addr[16712] = -1917054681;
assign addr[16713] = -1925596340;
assign addr[16714] = -1933985310;
assign addr[16715] = -1942220928;
assign addr[16716] = -1950302539;
assign addr[16717] = -1958229503;
assign addr[16718] = -1966001192;
assign addr[16719] = -1973616989;
assign addr[16720] = -1981076290;
assign addr[16721] = -1988378503;
assign addr[16722] = -1995523051;
assign addr[16723] = -2002509365;
assign addr[16724] = -2009336893;
assign addr[16725] = -2016005093;
assign addr[16726] = -2022513436;
assign addr[16727] = -2028861406;
assign addr[16728] = -2035048499;
assign addr[16729] = -2041074226;
assign addr[16730] = -2046938108;
assign addr[16731] = -2052639680;
assign addr[16732] = -2058178491;
assign addr[16733] = -2063554100;
assign addr[16734] = -2068766083;
assign addr[16735] = -2073814024;
assign addr[16736] = -2078697525;
assign addr[16737] = -2083416198;
assign addr[16738] = -2087969669;
assign addr[16739] = -2092357577;
assign addr[16740] = -2096579573;
assign addr[16741] = -2100635323;
assign addr[16742] = -2104524506;
assign addr[16743] = -2108246813;
assign addr[16744] = -2111801949;
assign addr[16745] = -2115189632;
assign addr[16746] = -2118409593;
assign addr[16747] = -2121461578;
assign addr[16748] = -2124345343;
assign addr[16749] = -2127060661;
assign addr[16750] = -2129607316;
assign addr[16751] = -2131985106;
assign addr[16752] = -2134193842;
assign addr[16753] = -2136233350;
assign addr[16754] = -2138103468;
assign addr[16755] = -2139804048;
assign addr[16756] = -2141334954;
assign addr[16757] = -2142696065;
assign addr[16758] = -2143887273;
assign addr[16759] = -2144908484;
assign addr[16760] = -2145759618;
assign addr[16761] = -2146440605;
assign addr[16762] = -2146951393;
assign addr[16763] = -2147291941;
assign addr[16764] = -2147462221;
assign addr[16765] = -2147462221;
assign addr[16766] = -2147291941;
assign addr[16767] = -2146951393;
assign addr[16768] = -2146440605;
assign addr[16769] = -2145759618;
assign addr[16770] = -2144908484;
assign addr[16771] = -2143887273;
assign addr[16772] = -2142696065;
assign addr[16773] = -2141334954;
assign addr[16774] = -2139804048;
assign addr[16775] = -2138103468;
assign addr[16776] = -2136233350;
assign addr[16777] = -2134193842;
assign addr[16778] = -2131985106;
assign addr[16779] = -2129607316;
assign addr[16780] = -2127060661;
assign addr[16781] = -2124345343;
assign addr[16782] = -2121461578;
assign addr[16783] = -2118409593;
assign addr[16784] = -2115189632;
assign addr[16785] = -2111801949;
assign addr[16786] = -2108246813;
assign addr[16787] = -2104524506;
assign addr[16788] = -2100635323;
assign addr[16789] = -2096579573;
assign addr[16790] = -2092357577;
assign addr[16791] = -2087969669;
assign addr[16792] = -2083416198;
assign addr[16793] = -2078697525;
assign addr[16794] = -2073814024;
assign addr[16795] = -2068766083;
assign addr[16796] = -2063554100;
assign addr[16797] = -2058178491;
assign addr[16798] = -2052639680;
assign addr[16799] = -2046938108;
assign addr[16800] = -2041074226;
assign addr[16801] = -2035048499;
assign addr[16802] = -2028861406;
assign addr[16803] = -2022513436;
assign addr[16804] = -2016005093;
assign addr[16805] = -2009336893;
assign addr[16806] = -2002509365;
assign addr[16807] = -1995523051;
assign addr[16808] = -1988378503;
assign addr[16809] = -1981076290;
assign addr[16810] = -1973616989;
assign addr[16811] = -1966001192;
assign addr[16812] = -1958229503;
assign addr[16813] = -1950302539;
assign addr[16814] = -1942220928;
assign addr[16815] = -1933985310;
assign addr[16816] = -1925596340;
assign addr[16817] = -1917054681;
assign addr[16818] = -1908361011;
assign addr[16819] = -1899516021;
assign addr[16820] = -1890520410;
assign addr[16821] = -1881374892;
assign addr[16822] = -1872080193;
assign addr[16823] = -1862637049;
assign addr[16824] = -1853046210;
assign addr[16825] = -1843308435;
assign addr[16826] = -1833424497;
assign addr[16827] = -1823395180;
assign addr[16828] = -1813221279;
assign addr[16829] = -1802903601;
assign addr[16830] = -1792442963;
assign addr[16831] = -1781840195;
assign addr[16832] = -1771096139;
assign addr[16833] = -1760211645;
assign addr[16834] = -1749187577;
assign addr[16835] = -1738024810;
assign addr[16836] = -1726724227;
assign addr[16837] = -1715286726;
assign addr[16838] = -1703713213;
assign addr[16839] = -1692004606;
assign addr[16840] = -1680161834;
assign addr[16841] = -1668185835;
assign addr[16842] = -1656077559;
assign addr[16843] = -1643837966;
assign addr[16844] = -1631468027;
assign addr[16845] = -1618968722;
assign addr[16846] = -1606341043;
assign addr[16847] = -1593585992;
assign addr[16848] = -1580704578;
assign addr[16849] = -1567697824;
assign addr[16850] = -1554566762;
assign addr[16851] = -1541312431;
assign addr[16852] = -1527935884;
assign addr[16853] = -1514438181;
assign addr[16854] = -1500820393;
assign addr[16855] = -1487083598;
assign addr[16856] = -1473228887;
assign addr[16857] = -1459257358;
assign addr[16858] = -1445170118;
assign addr[16859] = -1430968286;
assign addr[16860] = -1416652986;
assign addr[16861] = -1402225355;
assign addr[16862] = -1387686535;
assign addr[16863] = -1373037681;
assign addr[16864] = -1358279953;
assign addr[16865] = -1343414522;
assign addr[16866] = -1328442566;
assign addr[16867] = -1313365273;
assign addr[16868] = -1298183838;
assign addr[16869] = -1282899464;
assign addr[16870] = -1267513365;
assign addr[16871] = -1252026760;
assign addr[16872] = -1236440877;
assign addr[16873] = -1220756951;
assign addr[16874] = -1204976227;
assign addr[16875] = -1189099956;
assign addr[16876] = -1173129396;
assign addr[16877] = -1157065814;
assign addr[16878] = -1140910484;
assign addr[16879] = -1124664687;
assign addr[16880] = -1108329711;
assign addr[16881] = -1091906851;
assign addr[16882] = -1075397409;
assign addr[16883] = -1058802695;
assign addr[16884] = -1042124025;
assign addr[16885] = -1025362720;
assign addr[16886] = -1008520110;
assign addr[16887] = -991597531;
assign addr[16888] = -974596324;
assign addr[16889] = -957517838;
assign addr[16890] = -940363427;
assign addr[16891] = -923134450;
assign addr[16892] = -905832274;
assign addr[16893] = -888458272;
assign addr[16894] = -871013820;
assign addr[16895] = -853500302;
assign addr[16896] = -835919107;
assign addr[16897] = -818271628;
assign addr[16898] = -800559266;
assign addr[16899] = -782783424;
assign addr[16900] = -764945512;
assign addr[16901] = -747046944;
assign addr[16902] = -729089140;
assign addr[16903] = -711073524;
assign addr[16904] = -693001525;
assign addr[16905] = -674874574;
assign addr[16906] = -656694110;
assign addr[16907] = -638461574;
assign addr[16908] = -620178412;
assign addr[16909] = -601846074;
assign addr[16910] = -583466013;
assign addr[16911] = -565039687;
assign addr[16912] = -546568556;
assign addr[16913] = -528054086;
assign addr[16914] = -509497745;
assign addr[16915] = -490901003;
assign addr[16916] = -472265336;
assign addr[16917] = -453592221;
assign addr[16918] = -434883140;
assign addr[16919] = -416139574;
assign addr[16920] = -397363011;
assign addr[16921] = -378554940;
assign addr[16922] = -359716852;
assign addr[16923] = -340850240;
assign addr[16924] = -321956601;
assign addr[16925] = -303037433;
assign addr[16926] = -284094236;
assign addr[16927] = -265128512;
assign addr[16928] = -246141764;
assign addr[16929] = -227135500;
assign addr[16930] = -208111224;
assign addr[16931] = -189070447;
assign addr[16932] = -170014678;
assign addr[16933] = -150945428;
assign addr[16934] = -131864208;
assign addr[16935] = -112772533;
assign addr[16936] = -93671915;
assign addr[16937] = -74563870;
assign addr[16938] = -55449912;
assign addr[16939] = -36331557;
assign addr[16940] = -17210322;
assign addr[16941] = 1912278;
assign addr[16942] = 21034727;
assign addr[16943] = 40155507;
assign addr[16944] = 59273104;
assign addr[16945] = 78386000;
assign addr[16946] = 97492681;
assign addr[16947] = 116591632;
assign addr[16948] = 135681337;
assign addr[16949] = 154760284;
assign addr[16950] = 173826959;
assign addr[16951] = 192879850;
assign addr[16952] = 211917448;
assign addr[16953] = 230938242;
assign addr[16954] = 249940723;
assign addr[16955] = 268923386;
assign addr[16956] = 287884725;
assign addr[16957] = 306823237;
assign addr[16958] = 325737419;
assign addr[16959] = 344625773;
assign addr[16960] = 363486799;
assign addr[16961] = 382319004;
assign addr[16962] = 401120892;
assign addr[16963] = 419890975;
assign addr[16964] = 438627762;
assign addr[16965] = 457329769;
assign addr[16966] = 475995513;
assign addr[16967] = 494623513;
assign addr[16968] = 513212292;
assign addr[16969] = 531760377;
assign addr[16970] = 550266296;
assign addr[16971] = 568728583;
assign addr[16972] = 587145773;
assign addr[16973] = 605516406;
assign addr[16974] = 623839025;
assign addr[16975] = 642112178;
assign addr[16976] = 660334415;
assign addr[16977] = 678504291;
assign addr[16978] = 696620367;
assign addr[16979] = 714681204;
assign addr[16980] = 732685372;
assign addr[16981] = 750631442;
assign addr[16982] = 768517992;
assign addr[16983] = 786343603;
assign addr[16984] = 804106861;
assign addr[16985] = 821806359;
assign addr[16986] = 839440693;
assign addr[16987] = 857008464;
assign addr[16988] = 874508280;
assign addr[16989] = 891938752;
assign addr[16990] = 909298500;
assign addr[16991] = 926586145;
assign addr[16992] = 943800318;
assign addr[16993] = 960939653;
assign addr[16994] = 978002791;
assign addr[16995] = 994988380;
assign addr[16996] = 1011895073;
assign addr[16997] = 1028721528;
assign addr[16998] = 1045466412;
assign addr[16999] = 1062128397;
assign addr[17000] = 1078706161;
assign addr[17001] = 1095198391;
assign addr[17002] = 1111603778;
assign addr[17003] = 1127921022;
assign addr[17004] = 1144148829;
assign addr[17005] = 1160285911;
assign addr[17006] = 1176330990;
assign addr[17007] = 1192282793;
assign addr[17008] = 1208140056;
assign addr[17009] = 1223901520;
assign addr[17010] = 1239565936;
assign addr[17011] = 1255132063;
assign addr[17012] = 1270598665;
assign addr[17013] = 1285964516;
assign addr[17014] = 1301228398;
assign addr[17015] = 1316389101;
assign addr[17016] = 1331445422;
assign addr[17017] = 1346396168;
assign addr[17018] = 1361240152;
assign addr[17019] = 1375976199;
assign addr[17020] = 1390603139;
assign addr[17021] = 1405119813;
assign addr[17022] = 1419525069;
assign addr[17023] = 1433817766;
assign addr[17024] = 1447996770;
assign addr[17025] = 1462060956;
assign addr[17026] = 1476009210;
assign addr[17027] = 1489840425;
assign addr[17028] = 1503553506;
assign addr[17029] = 1517147363;
assign addr[17030] = 1530620920;
assign addr[17031] = 1543973108;
assign addr[17032] = 1557202869;
assign addr[17033] = 1570309153;
assign addr[17034] = 1583290921;
assign addr[17035] = 1596147143;
assign addr[17036] = 1608876801;
assign addr[17037] = 1621478885;
assign addr[17038] = 1633952396;
assign addr[17039] = 1646296344;
assign addr[17040] = 1658509750;
assign addr[17041] = 1670591647;
assign addr[17042] = 1682541077;
assign addr[17043] = 1694357091;
assign addr[17044] = 1706038753;
assign addr[17045] = 1717585136;
assign addr[17046] = 1728995326;
assign addr[17047] = 1740268417;
assign addr[17048] = 1751403515;
assign addr[17049] = 1762399737;
assign addr[17050] = 1773256212;
assign addr[17051] = 1783972079;
assign addr[17052] = 1794546487;
assign addr[17053] = 1804978599;
assign addr[17054] = 1815267588;
assign addr[17055] = 1825412636;
assign addr[17056] = 1835412941;
assign addr[17057] = 1845267708;
assign addr[17058] = 1854976157;
assign addr[17059] = 1864537518;
assign addr[17060] = 1873951032;
assign addr[17061] = 1883215953;
assign addr[17062] = 1892331547;
assign addr[17063] = 1901297091;
assign addr[17064] = 1910111873;
assign addr[17065] = 1918775195;
assign addr[17066] = 1927286370;
assign addr[17067] = 1935644723;
assign addr[17068] = 1943849591;
assign addr[17069] = 1951900324;
assign addr[17070] = 1959796283;
assign addr[17071] = 1967536842;
assign addr[17072] = 1975121388;
assign addr[17073] = 1982549318;
assign addr[17074] = 1989820044;
assign addr[17075] = 1996932990;
assign addr[17076] = 2003887591;
assign addr[17077] = 2010683297;
assign addr[17078] = 2017319567;
assign addr[17079] = 2023795876;
assign addr[17080] = 2030111710;
assign addr[17081] = 2036266570;
assign addr[17082] = 2042259965;
assign addr[17083] = 2048091422;
assign addr[17084] = 2053760478;
assign addr[17085] = 2059266683;
assign addr[17086] = 2064609600;
assign addr[17087] = 2069788807;
assign addr[17088] = 2074803892;
assign addr[17089] = 2079654458;
assign addr[17090] = 2084340120;
assign addr[17091] = 2088860507;
assign addr[17092] = 2093215260;
assign addr[17093] = 2097404033;
assign addr[17094] = 2101426496;
assign addr[17095] = 2105282327;
assign addr[17096] = 2108971223;
assign addr[17097] = 2112492891;
assign addr[17098] = 2115847050;
assign addr[17099] = 2119033436;
assign addr[17100] = 2122051796;
assign addr[17101] = 2124901890;
assign addr[17102] = 2127583492;
assign addr[17103] = 2130096389;
assign addr[17104] = 2132440383;
assign addr[17105] = 2134615288;
assign addr[17106] = 2136620930;
assign addr[17107] = 2138457152;
assign addr[17108] = 2140123807;
assign addr[17109] = 2141620763;
assign addr[17110] = 2142947902;
assign addr[17111] = 2144105118;
assign addr[17112] = 2145092320;
assign addr[17113] = 2145909429;
assign addr[17114] = 2146556380;
assign addr[17115] = 2147033123;
assign addr[17116] = 2147339619;
assign addr[17117] = 2147475844;
assign addr[17118] = 2147441787;
assign addr[17119] = 2147237452;
assign addr[17120] = 2146862854;
assign addr[17121] = 2146318022;
assign addr[17122] = 2145603001;
assign addr[17123] = 2144717846;
assign addr[17124] = 2143662628;
assign addr[17125] = 2142437431;
assign addr[17126] = 2141042352;
assign addr[17127] = 2139477502;
assign addr[17128] = 2137743003;
assign addr[17129] = 2135838995;
assign addr[17130] = 2133765628;
assign addr[17131] = 2131523066;
assign addr[17132] = 2129111488;
assign addr[17133] = 2126531084;
assign addr[17134] = 2123782059;
assign addr[17135] = 2120864631;
assign addr[17136] = 2117779031;
assign addr[17137] = 2114525505;
assign addr[17138] = 2111104309;
assign addr[17139] = 2107515716;
assign addr[17140] = 2103760010;
assign addr[17141] = 2099837489;
assign addr[17142] = 2095748463;
assign addr[17143] = 2091493257;
assign addr[17144] = 2087072209;
assign addr[17145] = 2082485668;
assign addr[17146] = 2077733999;
assign addr[17147] = 2072817579;
assign addr[17148] = 2067736796;
assign addr[17149] = 2062492055;
assign addr[17150] = 2057083771;
assign addr[17151] = 2051512372;
assign addr[17152] = 2045778302;
assign addr[17153] = 2039882013;
assign addr[17154] = 2033823974;
assign addr[17155] = 2027604666;
assign addr[17156] = 2021224581;
assign addr[17157] = 2014684225;
assign addr[17158] = 2007984117;
assign addr[17159] = 2001124788;
assign addr[17160] = 1994106782;
assign addr[17161] = 1986930656;
assign addr[17162] = 1979596978;
assign addr[17163] = 1972106330;
assign addr[17164] = 1964459306;
assign addr[17165] = 1956656513;
assign addr[17166] = 1948698568;
assign addr[17167] = 1940586104;
assign addr[17168] = 1932319763;
assign addr[17169] = 1923900201;
assign addr[17170] = 1915328086;
assign addr[17171] = 1906604097;
assign addr[17172] = 1897728925;
assign addr[17173] = 1888703276;
assign addr[17174] = 1879527863;
assign addr[17175] = 1870203416;
assign addr[17176] = 1860730673;
assign addr[17177] = 1851110385;
assign addr[17178] = 1841343316;
assign addr[17179] = 1831430239;
assign addr[17180] = 1821371941;
assign addr[17181] = 1811169220;
assign addr[17182] = 1800822883;
assign addr[17183] = 1790333753;
assign addr[17184] = 1779702660;
assign addr[17185] = 1768930447;
assign addr[17186] = 1758017969;
assign addr[17187] = 1746966091;
assign addr[17188] = 1735775690;
assign addr[17189] = 1724447652;
assign addr[17190] = 1712982875;
assign addr[17191] = 1701382270;
assign addr[17192] = 1689646755;
assign addr[17193] = 1677777262;
assign addr[17194] = 1665774731;
assign addr[17195] = 1653640115;
assign addr[17196] = 1641374375;
assign addr[17197] = 1628978484;
assign addr[17198] = 1616453425;
assign addr[17199] = 1603800191;
assign addr[17200] = 1591019785;
assign addr[17201] = 1578113222;
assign addr[17202] = 1565081523;
assign addr[17203] = 1551925723;
assign addr[17204] = 1538646865;
assign addr[17205] = 1525246002;
assign addr[17206] = 1511724196;
assign addr[17207] = 1498082520;
assign addr[17208] = 1484322054;
assign addr[17209] = 1470443891;
assign addr[17210] = 1456449131;
assign addr[17211] = 1442338884;
assign addr[17212] = 1428114267;
assign addr[17213] = 1413776410;
assign addr[17214] = 1399326449;
assign addr[17215] = 1384765530;
assign addr[17216] = 1370094808;
assign addr[17217] = 1355315445;
assign addr[17218] = 1340428615;
assign addr[17219] = 1325435496;
assign addr[17220] = 1310337279;
assign addr[17221] = 1295135159;
assign addr[17222] = 1279830344;
assign addr[17223] = 1264424045;
assign addr[17224] = 1248917486;
assign addr[17225] = 1233311895;
assign addr[17226] = 1217608510;
assign addr[17227] = 1201808576;
assign addr[17228] = 1185913346;
assign addr[17229] = 1169924081;
assign addr[17230] = 1153842047;
assign addr[17231] = 1137668521;
assign addr[17232] = 1121404785;
assign addr[17233] = 1105052128;
assign addr[17234] = 1088611847;
assign addr[17235] = 1072085246;
assign addr[17236] = 1055473635;
assign addr[17237] = 1038778332;
assign addr[17238] = 1022000660;
assign addr[17239] = 1005141949;
assign addr[17240] = 988203537;
assign addr[17241] = 971186766;
assign addr[17242] = 954092986;
assign addr[17243] = 936923553;
assign addr[17244] = 919679827;
assign addr[17245] = 902363176;
assign addr[17246] = 884974973;
assign addr[17247] = 867516597;
assign addr[17248] = 849989433;
assign addr[17249] = 832394869;
assign addr[17250] = 814734301;
assign addr[17251] = 797009130;
assign addr[17252] = 779220762;
assign addr[17253] = 761370605;
assign addr[17254] = 743460077;
assign addr[17255] = 725490597;
assign addr[17256] = 707463589;
assign addr[17257] = 689380485;
assign addr[17258] = 671242716;
assign addr[17259] = 653051723;
assign addr[17260] = 634808946;
assign addr[17261] = 616515832;
assign addr[17262] = 598173833;
assign addr[17263] = 579784402;
assign addr[17264] = 561348998;
assign addr[17265] = 542869083;
assign addr[17266] = 524346121;
assign addr[17267] = 505781581;
assign addr[17268] = 487176937;
assign addr[17269] = 468533662;
assign addr[17270] = 449853235;
assign addr[17271] = 431137138;
assign addr[17272] = 412386854;
assign addr[17273] = 393603870;
assign addr[17274] = 374789676;
assign addr[17275] = 355945764;
assign addr[17276] = 337073627;
assign addr[17277] = 318174762;
assign addr[17278] = 299250668;
assign addr[17279] = 280302845;
assign addr[17280] = 261332796;
assign addr[17281] = 242342025;
assign addr[17282] = 223332037;
assign addr[17283] = 204304341;
assign addr[17284] = 185260444;
assign addr[17285] = 166201858;
assign addr[17286] = 147130093;
assign addr[17287] = 128046661;
assign addr[17288] = 108953076;
assign addr[17289] = 89850852;
assign addr[17290] = 70741503;
assign addr[17291] = 51626544;
assign addr[17292] = 32507492;
assign addr[17293] = 13385863;
assign addr[17294] = -5736829;
assign addr[17295] = -24859065;
assign addr[17296] = -43979330;
assign addr[17297] = -63096108;
assign addr[17298] = -82207882;
assign addr[17299] = -101313138;
assign addr[17300] = -120410361;
assign addr[17301] = -139498035;
assign addr[17302] = -158574649;
assign addr[17303] = -177638688;
assign addr[17304] = -196688642;
assign addr[17305] = -215722999;
assign addr[17306] = -234740251;
assign addr[17307] = -253738890;
assign addr[17308] = -272717408;
assign addr[17309] = -291674302;
assign addr[17310] = -310608068;
assign addr[17311] = -329517204;
assign addr[17312] = -348400212;
assign addr[17313] = -367255594;
assign addr[17314] = -386081854;
assign addr[17315] = -404877501;
assign addr[17316] = -423641043;
assign addr[17317] = -442370993;
assign addr[17318] = -461065866;
assign addr[17319] = -479724180;
assign addr[17320] = -498344454;
assign addr[17321] = -516925212;
assign addr[17322] = -535464981;
assign addr[17323] = -553962291;
assign addr[17324] = -572415676;
assign addr[17325] = -590823671;
assign addr[17326] = -609184818;
assign addr[17327] = -627497660;
assign addr[17328] = -645760745;
assign addr[17329] = -663972625;
assign addr[17330] = -682131857;
assign addr[17331] = -700236999;
assign addr[17332] = -718286617;
assign addr[17333] = -736279279;
assign addr[17334] = -754213559;
assign addr[17335] = -772088034;
assign addr[17336] = -789901288;
assign addr[17337] = -807651907;
assign addr[17338] = -825338484;
assign addr[17339] = -842959617;
assign addr[17340] = -860513908;
assign addr[17341] = -877999966;
assign addr[17342] = -895416404;
assign addr[17343] = -912761841;
assign addr[17344] = -930034901;
assign addr[17345] = -947234215;
assign addr[17346] = -964358420;
assign addr[17347] = -981406156;
assign addr[17348] = -998376073;
assign addr[17349] = -1015266825;
assign addr[17350] = -1032077073;
assign addr[17351] = -1048805483;
assign addr[17352] = -1065450729;
assign addr[17353] = -1082011492;
assign addr[17354] = -1098486458;
assign addr[17355] = -1114874320;
assign addr[17356] = -1131173780;
assign addr[17357] = -1147383544;
assign addr[17358] = -1163502328;
assign addr[17359] = -1179528853;
assign addr[17360] = -1195461849;
assign addr[17361] = -1211300053;
assign addr[17362] = -1227042207;
assign addr[17363] = -1242687064;
assign addr[17364] = -1258233384;
assign addr[17365] = -1273679934;
assign addr[17366] = -1289025489;
assign addr[17367] = -1304268832;
assign addr[17368] = -1319408754;
assign addr[17369] = -1334444055;
assign addr[17370] = -1349373543;
assign addr[17371] = -1364196034;
assign addr[17372] = -1378910353;
assign addr[17373] = -1393515332;
assign addr[17374] = -1408009814;
assign addr[17375] = -1422392650;
assign addr[17376] = -1436662698;
assign addr[17377] = -1450818828;
assign addr[17378] = -1464859917;
assign addr[17379] = -1478784851;
assign addr[17380] = -1492592527;
assign addr[17381] = -1506281850;
assign addr[17382] = -1519851733;
assign addr[17383] = -1533301101;
assign addr[17384] = -1546628888;
assign addr[17385] = -1559834037;
assign addr[17386] = -1572915501;
assign addr[17387] = -1585872242;
assign addr[17388] = -1598703233;
assign addr[17389] = -1611407456;
assign addr[17390] = -1623983905;
assign addr[17391] = -1636431582;
assign addr[17392] = -1648749499;
assign addr[17393] = -1660936681;
assign addr[17394] = -1672992161;
assign addr[17395] = -1684914983;
assign addr[17396] = -1696704201;
assign addr[17397] = -1708358881;
assign addr[17398] = -1719878099;
assign addr[17399] = -1731260941;
assign addr[17400] = -1742506504;
assign addr[17401] = -1753613897;
assign addr[17402] = -1764582240;
assign addr[17403] = -1775410662;
assign addr[17404] = -1786098304;
assign addr[17405] = -1796644320;
assign addr[17406] = -1807047873;
assign addr[17407] = -1817308138;
assign addr[17408] = -1827424302;
assign addr[17409] = -1837395562;
assign addr[17410] = -1847221128;
assign addr[17411] = -1856900221;
assign addr[17412] = -1866432072;
assign addr[17413] = -1875815927;
assign addr[17414] = -1885051042;
assign addr[17415] = -1894136683;
assign addr[17416] = -1903072131;
assign addr[17417] = -1911856677;
assign addr[17418] = -1920489624;
assign addr[17419] = -1928970288;
assign addr[17420] = -1937297997;
assign addr[17421] = -1945472089;
assign addr[17422] = -1953491918;
assign addr[17423] = -1961356847;
assign addr[17424] = -1969066252;
assign addr[17425] = -1976619522;
assign addr[17426] = -1984016058;
assign addr[17427] = -1991255274;
assign addr[17428] = -1998336596;
assign addr[17429] = -2005259462;
assign addr[17430] = -2012023322;
assign addr[17431] = -2018627642;
assign addr[17432] = -2025071897;
assign addr[17433] = -2031355576;
assign addr[17434] = -2037478181;
assign addr[17435] = -2043439226;
assign addr[17436] = -2049238240;
assign addr[17437] = -2054874761;
assign addr[17438] = -2060348343;
assign addr[17439] = -2065658552;
assign addr[17440] = -2070804967;
assign addr[17441] = -2075787180;
assign addr[17442] = -2080604795;
assign addr[17443] = -2085257431;
assign addr[17444] = -2089744719;
assign addr[17445] = -2094066304;
assign addr[17446] = -2098221841;
assign addr[17447] = -2102211002;
assign addr[17448] = -2106033471;
assign addr[17449] = -2109688944;
assign addr[17450] = -2113177132;
assign addr[17451] = -2116497758;
assign addr[17452] = -2119650558;
assign addr[17453] = -2122635283;
assign addr[17454] = -2125451696;
assign addr[17455] = -2128099574;
assign addr[17456] = -2130578706;
assign addr[17457] = -2132888897;
assign addr[17458] = -2135029962;
assign addr[17459] = -2137001733;
assign addr[17460] = -2138804053;
assign addr[17461] = -2140436778;
assign addr[17462] = -2141899780;
assign addr[17463] = -2143192942;
assign addr[17464] = -2144316162;
assign addr[17465] = -2145269351;
assign addr[17466] = -2146052433;
assign addr[17467] = -2146665347;
assign addr[17468] = -2147108043;
assign addr[17469] = -2147380486;
assign addr[17470] = -2147482655;
assign addr[17471] = -2147414542;
assign addr[17472] = -2147176152;
assign addr[17473] = -2146767505;
assign addr[17474] = -2146188631;
assign addr[17475] = -2145439578;
assign addr[17476] = -2144520405;
assign addr[17477] = -2143431184;
assign addr[17478] = -2142172003;
assign addr[17479] = -2140742960;
assign addr[17480] = -2139144169;
assign addr[17481] = -2137375758;
assign addr[17482] = -2135437865;
assign addr[17483] = -2133330646;
assign addr[17484] = -2131054266;
assign addr[17485] = -2128608907;
assign addr[17486] = -2125994762;
assign addr[17487] = -2123212038;
assign addr[17488] = -2120260957;
assign addr[17489] = -2117141752;
assign addr[17490] = -2113854671;
assign addr[17491] = -2110399974;
assign addr[17492] = -2106777935;
assign addr[17493] = -2102988841;
assign addr[17494] = -2099032994;
assign addr[17495] = -2094910706;
assign addr[17496] = -2090622304;
assign addr[17497] = -2086168128;
assign addr[17498] = -2081548533;
assign addr[17499] = -2076763883;
assign addr[17500] = -2071814558;
assign addr[17501] = -2066700952;
assign addr[17502] = -2061423468;
assign addr[17503] = -2055982526;
assign addr[17504] = -2050378558;
assign addr[17505] = -2044612007;
assign addr[17506] = -2038683330;
assign addr[17507] = -2032592999;
assign addr[17508] = -2026341495;
assign addr[17509] = -2019929315;
assign addr[17510] = -2013356967;
assign addr[17511] = -2006624971;
assign addr[17512] = -1999733863;
assign addr[17513] = -1992684188;
assign addr[17514] = -1985476506;
assign addr[17515] = -1978111387;
assign addr[17516] = -1970589416;
assign addr[17517] = -1962911189;
assign addr[17518] = -1955077316;
assign addr[17519] = -1947088417;
assign addr[17520] = -1938945125;
assign addr[17521] = -1930648088;
assign addr[17522] = -1922197961;
assign addr[17523] = -1913595416;
assign addr[17524] = -1904841135;
assign addr[17525] = -1895935811;
assign addr[17526] = -1886880151;
assign addr[17527] = -1877674873;
assign addr[17528] = -1868320707;
assign addr[17529] = -1858818395;
assign addr[17530] = -1849168689;
assign addr[17531] = -1839372356;
assign addr[17532] = -1829430172;
assign addr[17533] = -1819342925;
assign addr[17534] = -1809111415;
assign addr[17535] = -1798736454;
assign addr[17536] = -1788218865;
assign addr[17537] = -1777559480;
assign addr[17538] = -1766759146;
assign addr[17539] = -1755818718;
assign addr[17540] = -1744739065;
assign addr[17541] = -1733521064;
assign addr[17542] = -1722165606;
assign addr[17543] = -1710673591;
assign addr[17544] = -1699045930;
assign addr[17545] = -1687283545;
assign addr[17546] = -1675387369;
assign addr[17547] = -1663358344;
assign addr[17548] = -1651197426;
assign addr[17549] = -1638905577;
assign addr[17550] = -1626483774;
assign addr[17551] = -1613933000;
assign addr[17552] = -1601254251;
assign addr[17553] = -1588448533;
assign addr[17554] = -1575516860;
assign addr[17555] = -1562460258;
assign addr[17556] = -1549279763;
assign addr[17557] = -1535976419;
assign addr[17558] = -1522551282;
assign addr[17559] = -1509005416;
assign addr[17560] = -1495339895;
assign addr[17561] = -1481555802;
assign addr[17562] = -1467654232;
assign addr[17563] = -1453636285;
assign addr[17564] = -1439503074;
assign addr[17565] = -1425255719;
assign addr[17566] = -1410895350;
assign addr[17567] = -1396423105;
assign addr[17568] = -1381840133;
assign addr[17569] = -1367147589;
assign addr[17570] = -1352346639;
assign addr[17571] = -1337438456;
assign addr[17572] = -1322424222;
assign addr[17573] = -1307305128;
assign addr[17574] = -1292082373;
assign addr[17575] = -1276757164;
assign addr[17576] = -1261330715;
assign addr[17577] = -1245804251;
assign addr[17578] = -1230179002;
assign addr[17579] = -1214456207;
assign addr[17580] = -1198637114;
assign addr[17581] = -1182722976;
assign addr[17582] = -1166715055;
assign addr[17583] = -1150614620;
assign addr[17584] = -1134422949;
assign addr[17585] = -1118141326;
assign addr[17586] = -1101771040;
assign addr[17587] = -1085313391;
assign addr[17588] = -1068769683;
assign addr[17589] = -1052141228;
assign addr[17590] = -1035429345;
assign addr[17591] = -1018635358;
assign addr[17592] = -1001760600;
assign addr[17593] = -984806408;
assign addr[17594] = -967774128;
assign addr[17595] = -950665109;
assign addr[17596] = -933480707;
assign addr[17597] = -916222287;
assign addr[17598] = -898891215;
assign addr[17599] = -881488868;
assign addr[17600] = -864016623;
assign addr[17601] = -846475867;
assign addr[17602] = -828867991;
assign addr[17603] = -811194391;
assign addr[17604] = -793456467;
assign addr[17605] = -775655628;
assign addr[17606] = -757793284;
assign addr[17607] = -739870851;
assign addr[17608] = -721889752;
assign addr[17609] = -703851410;
assign addr[17610] = -685757258;
assign addr[17611] = -667608730;
assign addr[17612] = -649407264;
assign addr[17613] = -631154304;
assign addr[17614] = -612851297;
assign addr[17615] = -594499695;
assign addr[17616] = -576100953;
assign addr[17617] = -557656529;
assign addr[17618] = -539167887;
assign addr[17619] = -520636492;
assign addr[17620] = -502063814;
assign addr[17621] = -483451325;
assign addr[17622] = -464800501;
assign addr[17623] = -446112822;
assign addr[17624] = -427389768;
assign addr[17625] = -408632825;
assign addr[17626] = -389843480;
assign addr[17627] = -371023223;
assign addr[17628] = -352173546;
assign addr[17629] = -333295944;
assign addr[17630] = -314391913;
assign addr[17631] = -295462954;
assign addr[17632] = -276510565;
assign addr[17633] = -257536251;
assign addr[17634] = -238541516;
assign addr[17635] = -219527866;
assign addr[17636] = -200496809;
assign addr[17637] = -181449854;
assign addr[17638] = -162388511;
assign addr[17639] = -143314291;
assign addr[17640] = -124228708;
assign addr[17641] = -105133274;
assign addr[17642] = -86029503;
assign addr[17643] = -66918911;
assign addr[17644] = -47803013;
assign addr[17645] = -28683324;
assign addr[17646] = -9561361;
assign addr[17647] = 9561361;
assign addr[17648] = 28683324;
assign addr[17649] = 47803013;
assign addr[17650] = 66918911;
assign addr[17651] = 86029503;
assign addr[17652] = 105133274;
assign addr[17653] = 124228708;
assign addr[17654] = 143314291;
assign addr[17655] = 162388511;
assign addr[17656] = 181449854;
assign addr[17657] = 200496809;
assign addr[17658] = 219527866;
assign addr[17659] = 238541516;
assign addr[17660] = 257536251;
assign addr[17661] = 276510565;
assign addr[17662] = 295462954;
assign addr[17663] = 314391913;
assign addr[17664] = 333295944;
assign addr[17665] = 352173546;
assign addr[17666] = 371023223;
assign addr[17667] = 389843480;
assign addr[17668] = 408632825;
assign addr[17669] = 427389768;
assign addr[17670] = 446112822;
assign addr[17671] = 464800501;
assign addr[17672] = 483451325;
assign addr[17673] = 502063814;
assign addr[17674] = 520636492;
assign addr[17675] = 539167887;
assign addr[17676] = 557656529;
assign addr[17677] = 576100953;
assign addr[17678] = 594499695;
assign addr[17679] = 612851297;
assign addr[17680] = 631154304;
assign addr[17681] = 649407264;
assign addr[17682] = 667608730;
assign addr[17683] = 685757258;
assign addr[17684] = 703851410;
assign addr[17685] = 721889752;
assign addr[17686] = 739870851;
assign addr[17687] = 757793284;
assign addr[17688] = 775655628;
assign addr[17689] = 793456467;
assign addr[17690] = 811194391;
assign addr[17691] = 828867991;
assign addr[17692] = 846475867;
assign addr[17693] = 864016623;
assign addr[17694] = 881488868;
assign addr[17695] = 898891215;
assign addr[17696] = 916222287;
assign addr[17697] = 933480707;
assign addr[17698] = 950665109;
assign addr[17699] = 967774128;
assign addr[17700] = 984806408;
assign addr[17701] = 1001760600;
assign addr[17702] = 1018635358;
assign addr[17703] = 1035429345;
assign addr[17704] = 1052141228;
assign addr[17705] = 1068769683;
assign addr[17706] = 1085313391;
assign addr[17707] = 1101771040;
assign addr[17708] = 1118141326;
assign addr[17709] = 1134422949;
assign addr[17710] = 1150614620;
assign addr[17711] = 1166715055;
assign addr[17712] = 1182722976;
assign addr[17713] = 1198637114;
assign addr[17714] = 1214456207;
assign addr[17715] = 1230179002;
assign addr[17716] = 1245804251;
assign addr[17717] = 1261330715;
assign addr[17718] = 1276757164;
assign addr[17719] = 1292082373;
assign addr[17720] = 1307305128;
assign addr[17721] = 1322424222;
assign addr[17722] = 1337438456;
assign addr[17723] = 1352346639;
assign addr[17724] = 1367147589;
assign addr[17725] = 1381840133;
assign addr[17726] = 1396423105;
assign addr[17727] = 1410895350;
assign addr[17728] = 1425255719;
assign addr[17729] = 1439503074;
assign addr[17730] = 1453636285;
assign addr[17731] = 1467654232;
assign addr[17732] = 1481555802;
assign addr[17733] = 1495339895;
assign addr[17734] = 1509005416;
assign addr[17735] = 1522551282;
assign addr[17736] = 1535976419;
assign addr[17737] = 1549279763;
assign addr[17738] = 1562460258;
assign addr[17739] = 1575516860;
assign addr[17740] = 1588448533;
assign addr[17741] = 1601254251;
assign addr[17742] = 1613933000;
assign addr[17743] = 1626483774;
assign addr[17744] = 1638905577;
assign addr[17745] = 1651197426;
assign addr[17746] = 1663358344;
assign addr[17747] = 1675387369;
assign addr[17748] = 1687283545;
assign addr[17749] = 1699045930;
assign addr[17750] = 1710673591;
assign addr[17751] = 1722165606;
assign addr[17752] = 1733521064;
assign addr[17753] = 1744739065;
assign addr[17754] = 1755818718;
assign addr[17755] = 1766759146;
assign addr[17756] = 1777559480;
assign addr[17757] = 1788218865;
assign addr[17758] = 1798736454;
assign addr[17759] = 1809111415;
assign addr[17760] = 1819342925;
assign addr[17761] = 1829430172;
assign addr[17762] = 1839372356;
assign addr[17763] = 1849168689;
assign addr[17764] = 1858818395;
assign addr[17765] = 1868320707;
assign addr[17766] = 1877674873;
assign addr[17767] = 1886880151;
assign addr[17768] = 1895935811;
assign addr[17769] = 1904841135;
assign addr[17770] = 1913595416;
assign addr[17771] = 1922197961;
assign addr[17772] = 1930648088;
assign addr[17773] = 1938945125;
assign addr[17774] = 1947088417;
assign addr[17775] = 1955077316;
assign addr[17776] = 1962911189;
assign addr[17777] = 1970589416;
assign addr[17778] = 1978111387;
assign addr[17779] = 1985476506;
assign addr[17780] = 1992684188;
assign addr[17781] = 1999733863;
assign addr[17782] = 2006624971;
assign addr[17783] = 2013356967;
assign addr[17784] = 2019929315;
assign addr[17785] = 2026341495;
assign addr[17786] = 2032592999;
assign addr[17787] = 2038683330;
assign addr[17788] = 2044612007;
assign addr[17789] = 2050378558;
assign addr[17790] = 2055982526;
assign addr[17791] = 2061423468;
assign addr[17792] = 2066700952;
assign addr[17793] = 2071814558;
assign addr[17794] = 2076763883;
assign addr[17795] = 2081548533;
assign addr[17796] = 2086168128;
assign addr[17797] = 2090622304;
assign addr[17798] = 2094910706;
assign addr[17799] = 2099032994;
assign addr[17800] = 2102988841;
assign addr[17801] = 2106777935;
assign addr[17802] = 2110399974;
assign addr[17803] = 2113854671;
assign addr[17804] = 2117141752;
assign addr[17805] = 2120260957;
assign addr[17806] = 2123212038;
assign addr[17807] = 2125994762;
assign addr[17808] = 2128608907;
assign addr[17809] = 2131054266;
assign addr[17810] = 2133330646;
assign addr[17811] = 2135437865;
assign addr[17812] = 2137375758;
assign addr[17813] = 2139144169;
assign addr[17814] = 2140742960;
assign addr[17815] = 2142172003;
assign addr[17816] = 2143431184;
assign addr[17817] = 2144520405;
assign addr[17818] = 2145439578;
assign addr[17819] = 2146188631;
assign addr[17820] = 2146767505;
assign addr[17821] = 2147176152;
assign addr[17822] = 2147414542;
assign addr[17823] = 2147482655;
assign addr[17824] = 2147380486;
assign addr[17825] = 2147108043;
assign addr[17826] = 2146665347;
assign addr[17827] = 2146052433;
assign addr[17828] = 2145269351;
assign addr[17829] = 2144316162;
assign addr[17830] = 2143192942;
assign addr[17831] = 2141899780;
assign addr[17832] = 2140436778;
assign addr[17833] = 2138804053;
assign addr[17834] = 2137001733;
assign addr[17835] = 2135029962;
assign addr[17836] = 2132888897;
assign addr[17837] = 2130578706;
assign addr[17838] = 2128099574;
assign addr[17839] = 2125451696;
assign addr[17840] = 2122635283;
assign addr[17841] = 2119650558;
assign addr[17842] = 2116497758;
assign addr[17843] = 2113177132;
assign addr[17844] = 2109688944;
assign addr[17845] = 2106033471;
assign addr[17846] = 2102211002;
assign addr[17847] = 2098221841;
assign addr[17848] = 2094066304;
assign addr[17849] = 2089744719;
assign addr[17850] = 2085257431;
assign addr[17851] = 2080604795;
assign addr[17852] = 2075787180;
assign addr[17853] = 2070804967;
assign addr[17854] = 2065658552;
assign addr[17855] = 2060348343;
assign addr[17856] = 2054874761;
assign addr[17857] = 2049238240;
assign addr[17858] = 2043439226;
assign addr[17859] = 2037478181;
assign addr[17860] = 2031355576;
assign addr[17861] = 2025071897;
assign addr[17862] = 2018627642;
assign addr[17863] = 2012023322;
assign addr[17864] = 2005259462;
assign addr[17865] = 1998336596;
assign addr[17866] = 1991255274;
assign addr[17867] = 1984016058;
assign addr[17868] = 1976619522;
assign addr[17869] = 1969066252;
assign addr[17870] = 1961356847;
assign addr[17871] = 1953491918;
assign addr[17872] = 1945472089;
assign addr[17873] = 1937297997;
assign addr[17874] = 1928970288;
assign addr[17875] = 1920489624;
assign addr[17876] = 1911856677;
assign addr[17877] = 1903072131;
assign addr[17878] = 1894136683;
assign addr[17879] = 1885051042;
assign addr[17880] = 1875815927;
assign addr[17881] = 1866432072;
assign addr[17882] = 1856900221;
assign addr[17883] = 1847221128;
assign addr[17884] = 1837395562;
assign addr[17885] = 1827424302;
assign addr[17886] = 1817308138;
assign addr[17887] = 1807047873;
assign addr[17888] = 1796644320;
assign addr[17889] = 1786098304;
assign addr[17890] = 1775410662;
assign addr[17891] = 1764582240;
assign addr[17892] = 1753613897;
assign addr[17893] = 1742506504;
assign addr[17894] = 1731260941;
assign addr[17895] = 1719878099;
assign addr[17896] = 1708358881;
assign addr[17897] = 1696704201;
assign addr[17898] = 1684914983;
assign addr[17899] = 1672992161;
assign addr[17900] = 1660936681;
assign addr[17901] = 1648749499;
assign addr[17902] = 1636431582;
assign addr[17903] = 1623983905;
assign addr[17904] = 1611407456;
assign addr[17905] = 1598703233;
assign addr[17906] = 1585872242;
assign addr[17907] = 1572915501;
assign addr[17908] = 1559834037;
assign addr[17909] = 1546628888;
assign addr[17910] = 1533301101;
assign addr[17911] = 1519851733;
assign addr[17912] = 1506281850;
assign addr[17913] = 1492592527;
assign addr[17914] = 1478784851;
assign addr[17915] = 1464859917;
assign addr[17916] = 1450818828;
assign addr[17917] = 1436662698;
assign addr[17918] = 1422392650;
assign addr[17919] = 1408009814;
assign addr[17920] = 1393515332;
assign addr[17921] = 1378910353;
assign addr[17922] = 1364196034;
assign addr[17923] = 1349373543;
assign addr[17924] = 1334444055;
assign addr[17925] = 1319408754;
assign addr[17926] = 1304268832;
assign addr[17927] = 1289025489;
assign addr[17928] = 1273679934;
assign addr[17929] = 1258233384;
assign addr[17930] = 1242687064;
assign addr[17931] = 1227042207;
assign addr[17932] = 1211300053;
assign addr[17933] = 1195461849;
assign addr[17934] = 1179528853;
assign addr[17935] = 1163502328;
assign addr[17936] = 1147383544;
assign addr[17937] = 1131173780;
assign addr[17938] = 1114874320;
assign addr[17939] = 1098486458;
assign addr[17940] = 1082011492;
assign addr[17941] = 1065450729;
assign addr[17942] = 1048805483;
assign addr[17943] = 1032077073;
assign addr[17944] = 1015266825;
assign addr[17945] = 998376073;
assign addr[17946] = 981406156;
assign addr[17947] = 964358420;
assign addr[17948] = 947234215;
assign addr[17949] = 930034901;
assign addr[17950] = 912761841;
assign addr[17951] = 895416404;
assign addr[17952] = 877999966;
assign addr[17953] = 860513908;
assign addr[17954] = 842959617;
assign addr[17955] = 825338484;
assign addr[17956] = 807651907;
assign addr[17957] = 789901288;
assign addr[17958] = 772088034;
assign addr[17959] = 754213559;
assign addr[17960] = 736279279;
assign addr[17961] = 718286617;
assign addr[17962] = 700236999;
assign addr[17963] = 682131857;
assign addr[17964] = 663972625;
assign addr[17965] = 645760745;
assign addr[17966] = 627497660;
assign addr[17967] = 609184818;
assign addr[17968] = 590823671;
assign addr[17969] = 572415676;
assign addr[17970] = 553962291;
assign addr[17971] = 535464981;
assign addr[17972] = 516925212;
assign addr[17973] = 498344454;
assign addr[17974] = 479724180;
assign addr[17975] = 461065866;
assign addr[17976] = 442370993;
assign addr[17977] = 423641043;
assign addr[17978] = 404877501;
assign addr[17979] = 386081854;
assign addr[17980] = 367255594;
assign addr[17981] = 348400212;
assign addr[17982] = 329517204;
assign addr[17983] = 310608068;
assign addr[17984] = 291674302;
assign addr[17985] = 272717408;
assign addr[17986] = 253738890;
assign addr[17987] = 234740251;
assign addr[17988] = 215722999;
assign addr[17989] = 196688642;
assign addr[17990] = 177638688;
assign addr[17991] = 158574649;
assign addr[17992] = 139498035;
assign addr[17993] = 120410361;
assign addr[17994] = 101313138;
assign addr[17995] = 82207882;
assign addr[17996] = 63096108;
assign addr[17997] = 43979330;
assign addr[17998] = 24859065;
assign addr[17999] = 5736829;
assign addr[18000] = -13385863;
assign addr[18001] = -32507492;
assign addr[18002] = -51626544;
assign addr[18003] = -70741503;
assign addr[18004] = -89850852;
assign addr[18005] = -108953076;
assign addr[18006] = -128046661;
assign addr[18007] = -147130093;
assign addr[18008] = -166201858;
assign addr[18009] = -185260444;
assign addr[18010] = -204304341;
assign addr[18011] = -223332037;
assign addr[18012] = -242342025;
assign addr[18013] = -261332796;
assign addr[18014] = -280302845;
assign addr[18015] = -299250668;
assign addr[18016] = -318174762;
assign addr[18017] = -337073627;
assign addr[18018] = -355945764;
assign addr[18019] = -374789676;
assign addr[18020] = -393603870;
assign addr[18021] = -412386854;
assign addr[18022] = -431137138;
assign addr[18023] = -449853235;
assign addr[18024] = -468533662;
assign addr[18025] = -487176937;
assign addr[18026] = -505781581;
assign addr[18027] = -524346121;
assign addr[18028] = -542869083;
assign addr[18029] = -561348998;
assign addr[18030] = -579784402;
assign addr[18031] = -598173833;
assign addr[18032] = -616515832;
assign addr[18033] = -634808946;
assign addr[18034] = -653051723;
assign addr[18035] = -671242716;
assign addr[18036] = -689380485;
assign addr[18037] = -707463589;
assign addr[18038] = -725490597;
assign addr[18039] = -743460077;
assign addr[18040] = -761370605;
assign addr[18041] = -779220762;
assign addr[18042] = -797009130;
assign addr[18043] = -814734301;
assign addr[18044] = -832394869;
assign addr[18045] = -849989433;
assign addr[18046] = -867516597;
assign addr[18047] = -884974973;
assign addr[18048] = -902363176;
assign addr[18049] = -919679827;
assign addr[18050] = -936923553;
assign addr[18051] = -954092986;
assign addr[18052] = -971186766;
assign addr[18053] = -988203537;
assign addr[18054] = -1005141949;
assign addr[18055] = -1022000660;
assign addr[18056] = -1038778332;
assign addr[18057] = -1055473635;
assign addr[18058] = -1072085246;
assign addr[18059] = -1088611847;
assign addr[18060] = -1105052128;
assign addr[18061] = -1121404785;
assign addr[18062] = -1137668521;
assign addr[18063] = -1153842047;
assign addr[18064] = -1169924081;
assign addr[18065] = -1185913346;
assign addr[18066] = -1201808576;
assign addr[18067] = -1217608510;
assign addr[18068] = -1233311895;
assign addr[18069] = -1248917486;
assign addr[18070] = -1264424045;
assign addr[18071] = -1279830344;
assign addr[18072] = -1295135159;
assign addr[18073] = -1310337279;
assign addr[18074] = -1325435496;
assign addr[18075] = -1340428615;
assign addr[18076] = -1355315445;
assign addr[18077] = -1370094808;
assign addr[18078] = -1384765530;
assign addr[18079] = -1399326449;
assign addr[18080] = -1413776410;
assign addr[18081] = -1428114267;
assign addr[18082] = -1442338884;
assign addr[18083] = -1456449131;
assign addr[18084] = -1470443891;
assign addr[18085] = -1484322054;
assign addr[18086] = -1498082520;
assign addr[18087] = -1511724196;
assign addr[18088] = -1525246002;
assign addr[18089] = -1538646865;
assign addr[18090] = -1551925723;
assign addr[18091] = -1565081523;
assign addr[18092] = -1578113222;
assign addr[18093] = -1591019785;
assign addr[18094] = -1603800191;
assign addr[18095] = -1616453425;
assign addr[18096] = -1628978484;
assign addr[18097] = -1641374375;
assign addr[18098] = -1653640115;
assign addr[18099] = -1665774731;
assign addr[18100] = -1677777262;
assign addr[18101] = -1689646755;
assign addr[18102] = -1701382270;
assign addr[18103] = -1712982875;
assign addr[18104] = -1724447652;
assign addr[18105] = -1735775690;
assign addr[18106] = -1746966091;
assign addr[18107] = -1758017969;
assign addr[18108] = -1768930447;
assign addr[18109] = -1779702660;
assign addr[18110] = -1790333753;
assign addr[18111] = -1800822883;
assign addr[18112] = -1811169220;
assign addr[18113] = -1821371941;
assign addr[18114] = -1831430239;
assign addr[18115] = -1841343316;
assign addr[18116] = -1851110385;
assign addr[18117] = -1860730673;
assign addr[18118] = -1870203416;
assign addr[18119] = -1879527863;
assign addr[18120] = -1888703276;
assign addr[18121] = -1897728925;
assign addr[18122] = -1906604097;
assign addr[18123] = -1915328086;
assign addr[18124] = -1923900201;
assign addr[18125] = -1932319763;
assign addr[18126] = -1940586104;
assign addr[18127] = -1948698568;
assign addr[18128] = -1956656513;
assign addr[18129] = -1964459306;
assign addr[18130] = -1972106330;
assign addr[18131] = -1979596978;
assign addr[18132] = -1986930656;
assign addr[18133] = -1994106782;
assign addr[18134] = -2001124788;
assign addr[18135] = -2007984117;
assign addr[18136] = -2014684225;
assign addr[18137] = -2021224581;
assign addr[18138] = -2027604666;
assign addr[18139] = -2033823974;
assign addr[18140] = -2039882013;
assign addr[18141] = -2045778302;
assign addr[18142] = -2051512372;
assign addr[18143] = -2057083771;
assign addr[18144] = -2062492055;
assign addr[18145] = -2067736796;
assign addr[18146] = -2072817579;
assign addr[18147] = -2077733999;
assign addr[18148] = -2082485668;
assign addr[18149] = -2087072209;
assign addr[18150] = -2091493257;
assign addr[18151] = -2095748463;
assign addr[18152] = -2099837489;
assign addr[18153] = -2103760010;
assign addr[18154] = -2107515716;
assign addr[18155] = -2111104309;
assign addr[18156] = -2114525505;
assign addr[18157] = -2117779031;
assign addr[18158] = -2120864631;
assign addr[18159] = -2123782059;
assign addr[18160] = -2126531084;
assign addr[18161] = -2129111488;
assign addr[18162] = -2131523066;
assign addr[18163] = -2133765628;
assign addr[18164] = -2135838995;
assign addr[18165] = -2137743003;
assign addr[18166] = -2139477502;
assign addr[18167] = -2141042352;
assign addr[18168] = -2142437431;
assign addr[18169] = -2143662628;
assign addr[18170] = -2144717846;
assign addr[18171] = -2145603001;
assign addr[18172] = -2146318022;
assign addr[18173] = -2146862854;
assign addr[18174] = -2147237452;
assign addr[18175] = -2147441787;
assign addr[18176] = -2147475844;
assign addr[18177] = -2147339619;
assign addr[18178] = -2147033123;
assign addr[18179] = -2146556380;
assign addr[18180] = -2145909429;
assign addr[18181] = -2145092320;
assign addr[18182] = -2144105118;
assign addr[18183] = -2142947902;
assign addr[18184] = -2141620763;
assign addr[18185] = -2140123807;
assign addr[18186] = -2138457152;
assign addr[18187] = -2136620930;
assign addr[18188] = -2134615288;
assign addr[18189] = -2132440383;
assign addr[18190] = -2130096389;
assign addr[18191] = -2127583492;
assign addr[18192] = -2124901890;
assign addr[18193] = -2122051796;
assign addr[18194] = -2119033436;
assign addr[18195] = -2115847050;
assign addr[18196] = -2112492891;
assign addr[18197] = -2108971223;
assign addr[18198] = -2105282327;
assign addr[18199] = -2101426496;
assign addr[18200] = -2097404033;
assign addr[18201] = -2093215260;
assign addr[18202] = -2088860507;
assign addr[18203] = -2084340120;
assign addr[18204] = -2079654458;
assign addr[18205] = -2074803892;
assign addr[18206] = -2069788807;
assign addr[18207] = -2064609600;
assign addr[18208] = -2059266683;
assign addr[18209] = -2053760478;
assign addr[18210] = -2048091422;
assign addr[18211] = -2042259965;
assign addr[18212] = -2036266570;
assign addr[18213] = -2030111710;
assign addr[18214] = -2023795876;
assign addr[18215] = -2017319567;
assign addr[18216] = -2010683297;
assign addr[18217] = -2003887591;
assign addr[18218] = -1996932990;
assign addr[18219] = -1989820044;
assign addr[18220] = -1982549318;
assign addr[18221] = -1975121388;
assign addr[18222] = -1967536842;
assign addr[18223] = -1959796283;
assign addr[18224] = -1951900324;
assign addr[18225] = -1943849591;
assign addr[18226] = -1935644723;
assign addr[18227] = -1927286370;
assign addr[18228] = -1918775195;
assign addr[18229] = -1910111873;
assign addr[18230] = -1901297091;
assign addr[18231] = -1892331547;
assign addr[18232] = -1883215953;
assign addr[18233] = -1873951032;
assign addr[18234] = -1864537518;
assign addr[18235] = -1854976157;
assign addr[18236] = -1845267708;
assign addr[18237] = -1835412941;
assign addr[18238] = -1825412636;
assign addr[18239] = -1815267588;
assign addr[18240] = -1804978599;
assign addr[18241] = -1794546487;
assign addr[18242] = -1783972079;
assign addr[18243] = -1773256212;
assign addr[18244] = -1762399737;
assign addr[18245] = -1751403515;
assign addr[18246] = -1740268417;
assign addr[18247] = -1728995326;
assign addr[18248] = -1717585136;
assign addr[18249] = -1706038753;
assign addr[18250] = -1694357091;
assign addr[18251] = -1682541077;
assign addr[18252] = -1670591647;
assign addr[18253] = -1658509750;
assign addr[18254] = -1646296344;
assign addr[18255] = -1633952396;
assign addr[18256] = -1621478885;
assign addr[18257] = -1608876801;
assign addr[18258] = -1596147143;
assign addr[18259] = -1583290921;
assign addr[18260] = -1570309153;
assign addr[18261] = -1557202869;
assign addr[18262] = -1543973108;
assign addr[18263] = -1530620920;
assign addr[18264] = -1517147363;
assign addr[18265] = -1503553506;
assign addr[18266] = -1489840425;
assign addr[18267] = -1476009210;
assign addr[18268] = -1462060956;
assign addr[18269] = -1447996770;
assign addr[18270] = -1433817766;
assign addr[18271] = -1419525069;
assign addr[18272] = -1405119813;
assign addr[18273] = -1390603139;
assign addr[18274] = -1375976199;
assign addr[18275] = -1361240152;
assign addr[18276] = -1346396168;
assign addr[18277] = -1331445422;
assign addr[18278] = -1316389101;
assign addr[18279] = -1301228398;
assign addr[18280] = -1285964516;
assign addr[18281] = -1270598665;
assign addr[18282] = -1255132063;
assign addr[18283] = -1239565936;
assign addr[18284] = -1223901520;
assign addr[18285] = -1208140056;
assign addr[18286] = -1192282793;
assign addr[18287] = -1176330990;
assign addr[18288] = -1160285911;
assign addr[18289] = -1144148829;
assign addr[18290] = -1127921022;
assign addr[18291] = -1111603778;
assign addr[18292] = -1095198391;
assign addr[18293] = -1078706161;
assign addr[18294] = -1062128397;
assign addr[18295] = -1045466412;
assign addr[18296] = -1028721528;
assign addr[18297] = -1011895073;
assign addr[18298] = -994988380;
assign addr[18299] = -978002791;
assign addr[18300] = -960939653;
assign addr[18301] = -943800318;
assign addr[18302] = -926586145;
assign addr[18303] = -909298500;
assign addr[18304] = -891938752;
assign addr[18305] = -874508280;
assign addr[18306] = -857008464;
assign addr[18307] = -839440693;
assign addr[18308] = -821806359;
assign addr[18309] = -804106861;
assign addr[18310] = -786343603;
assign addr[18311] = -768517992;
assign addr[18312] = -750631442;
assign addr[18313] = -732685372;
assign addr[18314] = -714681204;
assign addr[18315] = -696620367;
assign addr[18316] = -678504291;
assign addr[18317] = -660334415;
assign addr[18318] = -642112178;
assign addr[18319] = -623839025;
assign addr[18320] = -605516406;
assign addr[18321] = -587145773;
assign addr[18322] = -568728583;
assign addr[18323] = -550266296;
assign addr[18324] = -531760377;
assign addr[18325] = -513212292;
assign addr[18326] = -494623513;
assign addr[18327] = -475995513;
assign addr[18328] = -457329769;
assign addr[18329] = -438627762;
assign addr[18330] = -419890975;
assign addr[18331] = -401120892;
assign addr[18332] = -382319004;
assign addr[18333] = -363486799;
assign addr[18334] = -344625773;
assign addr[18335] = -325737419;
assign addr[18336] = -306823237;
assign addr[18337] = -287884725;
assign addr[18338] = -268923386;
assign addr[18339] = -249940723;
assign addr[18340] = -230938242;
assign addr[18341] = -211917448;
assign addr[18342] = -192879850;
assign addr[18343] = -173826959;
assign addr[18344] = -154760284;
assign addr[18345] = -135681337;
assign addr[18346] = -116591632;
assign addr[18347] = -97492681;
assign addr[18348] = -78386000;
assign addr[18349] = -59273104;
assign addr[18350] = -40155507;
assign addr[18351] = -21034727;
assign addr[18352] = -1912278;
assign addr[18353] = 17210322;
assign addr[18354] = 36331557;
assign addr[18355] = 55449912;
assign addr[18356] = 74563870;
assign addr[18357] = 93671915;
assign addr[18358] = 112772533;
assign addr[18359] = 131864208;
assign addr[18360] = 150945428;
assign addr[18361] = 170014678;
assign addr[18362] = 189070447;
assign addr[18363] = 208111224;
assign addr[18364] = 227135500;
assign addr[18365] = 246141764;
assign addr[18366] = 265128512;
assign addr[18367] = 284094236;
assign addr[18368] = 303037433;
assign addr[18369] = 321956601;
assign addr[18370] = 340850240;
assign addr[18371] = 359716852;
assign addr[18372] = 378554940;
assign addr[18373] = 397363011;
assign addr[18374] = 416139574;
assign addr[18375] = 434883140;
assign addr[18376] = 453592221;
assign addr[18377] = 472265336;
assign addr[18378] = 490901003;
assign addr[18379] = 509497745;
assign addr[18380] = 528054086;
assign addr[18381] = 546568556;
assign addr[18382] = 565039687;
assign addr[18383] = 583466013;
assign addr[18384] = 601846074;
assign addr[18385] = 620178412;
assign addr[18386] = 638461574;
assign addr[18387] = 656694110;
assign addr[18388] = 674874574;
assign addr[18389] = 693001525;
assign addr[18390] = 711073524;
assign addr[18391] = 729089140;
assign addr[18392] = 747046944;
assign addr[18393] = 764945512;
assign addr[18394] = 782783424;
assign addr[18395] = 800559266;
assign addr[18396] = 818271628;
assign addr[18397] = 835919107;
assign addr[18398] = 853500302;
assign addr[18399] = 871013820;
assign addr[18400] = 888458272;
assign addr[18401] = 905832274;
assign addr[18402] = 923134450;
assign addr[18403] = 940363427;
assign addr[18404] = 957517838;
assign addr[18405] = 974596324;
assign addr[18406] = 991597531;
assign addr[18407] = 1008520110;
assign addr[18408] = 1025362720;
assign addr[18409] = 1042124025;
assign addr[18410] = 1058802695;
assign addr[18411] = 1075397409;
assign addr[18412] = 1091906851;
assign addr[18413] = 1108329711;
assign addr[18414] = 1124664687;
assign addr[18415] = 1140910484;
assign addr[18416] = 1157065814;
assign addr[18417] = 1173129396;
assign addr[18418] = 1189099956;
assign addr[18419] = 1204976227;
assign addr[18420] = 1220756951;
assign addr[18421] = 1236440877;
assign addr[18422] = 1252026760;
assign addr[18423] = 1267513365;
assign addr[18424] = 1282899464;
assign addr[18425] = 1298183838;
assign addr[18426] = 1313365273;
assign addr[18427] = 1328442566;
assign addr[18428] = 1343414522;
assign addr[18429] = 1358279953;
assign addr[18430] = 1373037681;
assign addr[18431] = 1387686535;
assign addr[18432] = 1402225355;
assign addr[18433] = 1416652986;
assign addr[18434] = 1430968286;
assign addr[18435] = 1445170118;
assign addr[18436] = 1459257358;
assign addr[18437] = 1473228887;
assign addr[18438] = 1487083598;
assign addr[18439] = 1500820393;
assign addr[18440] = 1514438181;
assign addr[18441] = 1527935884;
assign addr[18442] = 1541312431;
assign addr[18443] = 1554566762;
assign addr[18444] = 1567697824;
assign addr[18445] = 1580704578;
assign addr[18446] = 1593585992;
assign addr[18447] = 1606341043;
assign addr[18448] = 1618968722;
assign addr[18449] = 1631468027;
assign addr[18450] = 1643837966;
assign addr[18451] = 1656077559;
assign addr[18452] = 1668185835;
assign addr[18453] = 1680161834;
assign addr[18454] = 1692004606;
assign addr[18455] = 1703713213;
assign addr[18456] = 1715286726;
assign addr[18457] = 1726724227;
assign addr[18458] = 1738024810;
assign addr[18459] = 1749187577;
assign addr[18460] = 1760211645;
assign addr[18461] = 1771096139;
assign addr[18462] = 1781840195;
assign addr[18463] = 1792442963;
assign addr[18464] = 1802903601;
assign addr[18465] = 1813221279;
assign addr[18466] = 1823395180;
assign addr[18467] = 1833424497;
assign addr[18468] = 1843308435;
assign addr[18469] = 1853046210;
assign addr[18470] = 1862637049;
assign addr[18471] = 1872080193;
assign addr[18472] = 1881374892;
assign addr[18473] = 1890520410;
assign addr[18474] = 1899516021;
assign addr[18475] = 1908361011;
assign addr[18476] = 1917054681;
assign addr[18477] = 1925596340;
assign addr[18478] = 1933985310;
assign addr[18479] = 1942220928;
assign addr[18480] = 1950302539;
assign addr[18481] = 1958229503;
assign addr[18482] = 1966001192;
assign addr[18483] = 1973616989;
assign addr[18484] = 1981076290;
assign addr[18485] = 1988378503;
assign addr[18486] = 1995523051;
assign addr[18487] = 2002509365;
assign addr[18488] = 2009336893;
assign addr[18489] = 2016005093;
assign addr[18490] = 2022513436;
assign addr[18491] = 2028861406;
assign addr[18492] = 2035048499;
assign addr[18493] = 2041074226;
assign addr[18494] = 2046938108;
assign addr[18495] = 2052639680;
assign addr[18496] = 2058178491;
assign addr[18497] = 2063554100;
assign addr[18498] = 2068766083;
assign addr[18499] = 2073814024;
assign addr[18500] = 2078697525;
assign addr[18501] = 2083416198;
assign addr[18502] = 2087969669;
assign addr[18503] = 2092357577;
assign addr[18504] = 2096579573;
assign addr[18505] = 2100635323;
assign addr[18506] = 2104524506;
assign addr[18507] = 2108246813;
assign addr[18508] = 2111801949;
assign addr[18509] = 2115189632;
assign addr[18510] = 2118409593;
assign addr[18511] = 2121461578;
assign addr[18512] = 2124345343;
assign addr[18513] = 2127060661;
assign addr[18514] = 2129607316;
assign addr[18515] = 2131985106;
assign addr[18516] = 2134193842;
assign addr[18517] = 2136233350;
assign addr[18518] = 2138103468;
assign addr[18519] = 2139804048;
assign addr[18520] = 2141334954;
assign addr[18521] = 2142696065;
assign addr[18522] = 2143887273;
assign addr[18523] = 2144908484;
assign addr[18524] = 2145759618;
assign addr[18525] = 2146440605;
assign addr[18526] = 2146951393;
assign addr[18527] = 2147291941;
assign addr[18528] = 2147462221;
assign addr[18529] = 2147462221;
assign addr[18530] = 2147291941;
assign addr[18531] = 2146951393;
assign addr[18532] = 2146440605;
assign addr[18533] = 2145759618;
assign addr[18534] = 2144908484;
assign addr[18535] = 2143887273;
assign addr[18536] = 2142696065;
assign addr[18537] = 2141334954;
assign addr[18538] = 2139804048;
assign addr[18539] = 2138103468;
assign addr[18540] = 2136233350;
assign addr[18541] = 2134193842;
assign addr[18542] = 2131985106;
assign addr[18543] = 2129607316;
assign addr[18544] = 2127060661;
assign addr[18545] = 2124345343;
assign addr[18546] = 2121461578;
assign addr[18547] = 2118409593;
assign addr[18548] = 2115189632;
assign addr[18549] = 2111801949;
assign addr[18550] = 2108246813;
assign addr[18551] = 2104524506;
assign addr[18552] = 2100635323;
assign addr[18553] = 2096579573;
assign addr[18554] = 2092357577;
assign addr[18555] = 2087969669;
assign addr[18556] = 2083416198;
assign addr[18557] = 2078697525;
assign addr[18558] = 2073814024;
assign addr[18559] = 2068766083;
assign addr[18560] = 2063554100;
assign addr[18561] = 2058178491;
assign addr[18562] = 2052639680;
assign addr[18563] = 2046938108;
assign addr[18564] = 2041074226;
assign addr[18565] = 2035048499;
assign addr[18566] = 2028861406;
assign addr[18567] = 2022513436;
assign addr[18568] = 2016005093;
assign addr[18569] = 2009336893;
assign addr[18570] = 2002509365;
assign addr[18571] = 1995523051;
assign addr[18572] = 1988378503;
assign addr[18573] = 1981076290;
assign addr[18574] = 1973616989;
assign addr[18575] = 1966001192;
assign addr[18576] = 1958229503;
assign addr[18577] = 1950302539;
assign addr[18578] = 1942220928;
assign addr[18579] = 1933985310;
assign addr[18580] = 1925596340;
assign addr[18581] = 1917054681;
assign addr[18582] = 1908361011;
assign addr[18583] = 1899516021;
assign addr[18584] = 1890520410;
assign addr[18585] = 1881374892;
assign addr[18586] = 1872080193;
assign addr[18587] = 1862637049;
assign addr[18588] = 1853046210;
assign addr[18589] = 1843308435;
assign addr[18590] = 1833424497;
assign addr[18591] = 1823395180;
assign addr[18592] = 1813221279;
assign addr[18593] = 1802903601;
assign addr[18594] = 1792442963;
assign addr[18595] = 1781840195;
assign addr[18596] = 1771096139;
assign addr[18597] = 1760211645;
assign addr[18598] = 1749187577;
assign addr[18599] = 1738024810;
assign addr[18600] = 1726724227;
assign addr[18601] = 1715286726;
assign addr[18602] = 1703713213;
assign addr[18603] = 1692004606;
assign addr[18604] = 1680161834;
assign addr[18605] = 1668185835;
assign addr[18606] = 1656077559;
assign addr[18607] = 1643837966;
assign addr[18608] = 1631468027;
assign addr[18609] = 1618968722;
assign addr[18610] = 1606341043;
assign addr[18611] = 1593585992;
assign addr[18612] = 1580704578;
assign addr[18613] = 1567697824;
assign addr[18614] = 1554566762;
assign addr[18615] = 1541312431;
assign addr[18616] = 1527935884;
assign addr[18617] = 1514438181;
assign addr[18618] = 1500820393;
assign addr[18619] = 1487083598;
assign addr[18620] = 1473228887;
assign addr[18621] = 1459257358;
assign addr[18622] = 1445170118;
assign addr[18623] = 1430968286;
assign addr[18624] = 1416652986;
assign addr[18625] = 1402225355;
assign addr[18626] = 1387686535;
assign addr[18627] = 1373037681;
assign addr[18628] = 1358279953;
assign addr[18629] = 1343414522;
assign addr[18630] = 1328442566;
assign addr[18631] = 1313365273;
assign addr[18632] = 1298183838;
assign addr[18633] = 1282899464;
assign addr[18634] = 1267513365;
assign addr[18635] = 1252026760;
assign addr[18636] = 1236440877;
assign addr[18637] = 1220756951;
assign addr[18638] = 1204976227;
assign addr[18639] = 1189099956;
assign addr[18640] = 1173129396;
assign addr[18641] = 1157065814;
assign addr[18642] = 1140910484;
assign addr[18643] = 1124664687;
assign addr[18644] = 1108329711;
assign addr[18645] = 1091906851;
assign addr[18646] = 1075397409;
assign addr[18647] = 1058802695;
assign addr[18648] = 1042124025;
assign addr[18649] = 1025362720;
assign addr[18650] = 1008520110;
assign addr[18651] = 991597531;
assign addr[18652] = 974596324;
assign addr[18653] = 957517838;
assign addr[18654] = 940363427;
assign addr[18655] = 923134450;
assign addr[18656] = 905832274;
assign addr[18657] = 888458272;
assign addr[18658] = 871013820;
assign addr[18659] = 853500302;
assign addr[18660] = 835919107;
assign addr[18661] = 818271628;
assign addr[18662] = 800559266;
assign addr[18663] = 782783424;
assign addr[18664] = 764945512;
assign addr[18665] = 747046944;
assign addr[18666] = 729089140;
assign addr[18667] = 711073524;
assign addr[18668] = 693001525;
assign addr[18669] = 674874574;
assign addr[18670] = 656694110;
assign addr[18671] = 638461574;
assign addr[18672] = 620178412;
assign addr[18673] = 601846074;
assign addr[18674] = 583466013;
assign addr[18675] = 565039687;
assign addr[18676] = 546568556;
assign addr[18677] = 528054086;
assign addr[18678] = 509497745;
assign addr[18679] = 490901003;
assign addr[18680] = 472265336;
assign addr[18681] = 453592221;
assign addr[18682] = 434883140;
assign addr[18683] = 416139574;
assign addr[18684] = 397363011;
assign addr[18685] = 378554940;
assign addr[18686] = 359716852;
assign addr[18687] = 340850240;
assign addr[18688] = 321956601;
assign addr[18689] = 303037433;
assign addr[18690] = 284094236;
assign addr[18691] = 265128512;
assign addr[18692] = 246141764;
assign addr[18693] = 227135500;
assign addr[18694] = 208111224;
assign addr[18695] = 189070447;
assign addr[18696] = 170014678;
assign addr[18697] = 150945428;
assign addr[18698] = 131864208;
assign addr[18699] = 112772533;
assign addr[18700] = 93671915;
assign addr[18701] = 74563870;
assign addr[18702] = 55449912;
assign addr[18703] = 36331557;
assign addr[18704] = 17210322;
assign addr[18705] = -1912278;
assign addr[18706] = -21034727;
assign addr[18707] = -40155507;
assign addr[18708] = -59273104;
assign addr[18709] = -78386000;
assign addr[18710] = -97492681;
assign addr[18711] = -116591632;
assign addr[18712] = -135681337;
assign addr[18713] = -154760284;
assign addr[18714] = -173826959;
assign addr[18715] = -192879850;
assign addr[18716] = -211917448;
assign addr[18717] = -230938242;
assign addr[18718] = -249940723;
assign addr[18719] = -268923386;
assign addr[18720] = -287884725;
assign addr[18721] = -306823237;
assign addr[18722] = -325737419;
assign addr[18723] = -344625773;
assign addr[18724] = -363486799;
assign addr[18725] = -382319004;
assign addr[18726] = -401120892;
assign addr[18727] = -419890975;
assign addr[18728] = -438627762;
assign addr[18729] = -457329769;
assign addr[18730] = -475995513;
assign addr[18731] = -494623513;
assign addr[18732] = -513212292;
assign addr[18733] = -531760377;
assign addr[18734] = -550266296;
assign addr[18735] = -568728583;
assign addr[18736] = -587145773;
assign addr[18737] = -605516406;
assign addr[18738] = -623839025;
assign addr[18739] = -642112178;
assign addr[18740] = -660334415;
assign addr[18741] = -678504291;
assign addr[18742] = -696620367;
assign addr[18743] = -714681204;
assign addr[18744] = -732685372;
assign addr[18745] = -750631442;
assign addr[18746] = -768517992;
assign addr[18747] = -786343603;
assign addr[18748] = -804106861;
assign addr[18749] = -821806359;
assign addr[18750] = -839440693;
assign addr[18751] = -857008464;
assign addr[18752] = -874508280;
assign addr[18753] = -891938752;
assign addr[18754] = -909298500;
assign addr[18755] = -926586145;
assign addr[18756] = -943800318;
assign addr[18757] = -960939653;
assign addr[18758] = -978002791;
assign addr[18759] = -994988380;
assign addr[18760] = -1011895073;
assign addr[18761] = -1028721528;
assign addr[18762] = -1045466412;
assign addr[18763] = -1062128397;
assign addr[18764] = -1078706161;
assign addr[18765] = -1095198391;
assign addr[18766] = -1111603778;
assign addr[18767] = -1127921022;
assign addr[18768] = -1144148829;
assign addr[18769] = -1160285911;
assign addr[18770] = -1176330990;
assign addr[18771] = -1192282793;
assign addr[18772] = -1208140056;
assign addr[18773] = -1223901520;
assign addr[18774] = -1239565936;
assign addr[18775] = -1255132063;
assign addr[18776] = -1270598665;
assign addr[18777] = -1285964516;
assign addr[18778] = -1301228398;
assign addr[18779] = -1316389101;
assign addr[18780] = -1331445422;
assign addr[18781] = -1346396168;
assign addr[18782] = -1361240152;
assign addr[18783] = -1375976199;
assign addr[18784] = -1390603139;
assign addr[18785] = -1405119813;
assign addr[18786] = -1419525069;
assign addr[18787] = -1433817766;
assign addr[18788] = -1447996770;
assign addr[18789] = -1462060956;
assign addr[18790] = -1476009210;
assign addr[18791] = -1489840425;
assign addr[18792] = -1503553506;
assign addr[18793] = -1517147363;
assign addr[18794] = -1530620920;
assign addr[18795] = -1543973108;
assign addr[18796] = -1557202869;
assign addr[18797] = -1570309153;
assign addr[18798] = -1583290921;
assign addr[18799] = -1596147143;
assign addr[18800] = -1608876801;
assign addr[18801] = -1621478885;
assign addr[18802] = -1633952396;
assign addr[18803] = -1646296344;
assign addr[18804] = -1658509750;
assign addr[18805] = -1670591647;
assign addr[18806] = -1682541077;
assign addr[18807] = -1694357091;
assign addr[18808] = -1706038753;
assign addr[18809] = -1717585136;
assign addr[18810] = -1728995326;
assign addr[18811] = -1740268417;
assign addr[18812] = -1751403515;
assign addr[18813] = -1762399737;
assign addr[18814] = -1773256212;
assign addr[18815] = -1783972079;
assign addr[18816] = -1794546487;
assign addr[18817] = -1804978599;
assign addr[18818] = -1815267588;
assign addr[18819] = -1825412636;
assign addr[18820] = -1835412941;
assign addr[18821] = -1845267708;
assign addr[18822] = -1854976157;
assign addr[18823] = -1864537518;
assign addr[18824] = -1873951032;
assign addr[18825] = -1883215953;
assign addr[18826] = -1892331547;
assign addr[18827] = -1901297091;
assign addr[18828] = -1910111873;
assign addr[18829] = -1918775195;
assign addr[18830] = -1927286370;
assign addr[18831] = -1935644723;
assign addr[18832] = -1943849591;
assign addr[18833] = -1951900324;
assign addr[18834] = -1959796283;
assign addr[18835] = -1967536842;
assign addr[18836] = -1975121388;
assign addr[18837] = -1982549318;
assign addr[18838] = -1989820044;
assign addr[18839] = -1996932990;
assign addr[18840] = -2003887591;
assign addr[18841] = -2010683297;
assign addr[18842] = -2017319567;
assign addr[18843] = -2023795876;
assign addr[18844] = -2030111710;
assign addr[18845] = -2036266570;
assign addr[18846] = -2042259965;
assign addr[18847] = -2048091422;
assign addr[18848] = -2053760478;
assign addr[18849] = -2059266683;
assign addr[18850] = -2064609600;
assign addr[18851] = -2069788807;
assign addr[18852] = -2074803892;
assign addr[18853] = -2079654458;
assign addr[18854] = -2084340120;
assign addr[18855] = -2088860507;
assign addr[18856] = -2093215260;
assign addr[18857] = -2097404033;
assign addr[18858] = -2101426496;
assign addr[18859] = -2105282327;
assign addr[18860] = -2108971223;
assign addr[18861] = -2112492891;
assign addr[18862] = -2115847050;
assign addr[18863] = -2119033436;
assign addr[18864] = -2122051796;
assign addr[18865] = -2124901890;
assign addr[18866] = -2127583492;
assign addr[18867] = -2130096389;
assign addr[18868] = -2132440383;
assign addr[18869] = -2134615288;
assign addr[18870] = -2136620930;
assign addr[18871] = -2138457152;
assign addr[18872] = -2140123807;
assign addr[18873] = -2141620763;
assign addr[18874] = -2142947902;
assign addr[18875] = -2144105118;
assign addr[18876] = -2145092320;
assign addr[18877] = -2145909429;
assign addr[18878] = -2146556380;
assign addr[18879] = -2147033123;
assign addr[18880] = -2147339619;
assign addr[18881] = -2147475844;
assign addr[18882] = -2147441787;
assign addr[18883] = -2147237452;
assign addr[18884] = -2146862854;
assign addr[18885] = -2146318022;
assign addr[18886] = -2145603001;
assign addr[18887] = -2144717846;
assign addr[18888] = -2143662628;
assign addr[18889] = -2142437431;
assign addr[18890] = -2141042352;
assign addr[18891] = -2139477502;
assign addr[18892] = -2137743003;
assign addr[18893] = -2135838995;
assign addr[18894] = -2133765628;
assign addr[18895] = -2131523066;
assign addr[18896] = -2129111488;
assign addr[18897] = -2126531084;
assign addr[18898] = -2123782059;
assign addr[18899] = -2120864631;
assign addr[18900] = -2117779031;
assign addr[18901] = -2114525505;
assign addr[18902] = -2111104309;
assign addr[18903] = -2107515716;
assign addr[18904] = -2103760010;
assign addr[18905] = -2099837489;
assign addr[18906] = -2095748463;
assign addr[18907] = -2091493257;
assign addr[18908] = -2087072209;
assign addr[18909] = -2082485668;
assign addr[18910] = -2077733999;
assign addr[18911] = -2072817579;
assign addr[18912] = -2067736796;
assign addr[18913] = -2062492055;
assign addr[18914] = -2057083771;
assign addr[18915] = -2051512372;
assign addr[18916] = -2045778302;
assign addr[18917] = -2039882013;
assign addr[18918] = -2033823974;
assign addr[18919] = -2027604666;
assign addr[18920] = -2021224581;
assign addr[18921] = -2014684225;
assign addr[18922] = -2007984117;
assign addr[18923] = -2001124788;
assign addr[18924] = -1994106782;
assign addr[18925] = -1986930656;
assign addr[18926] = -1979596978;
assign addr[18927] = -1972106330;
assign addr[18928] = -1964459306;
assign addr[18929] = -1956656513;
assign addr[18930] = -1948698568;
assign addr[18931] = -1940586104;
assign addr[18932] = -1932319763;
assign addr[18933] = -1923900201;
assign addr[18934] = -1915328086;
assign addr[18935] = -1906604097;
assign addr[18936] = -1897728925;
assign addr[18937] = -1888703276;
assign addr[18938] = -1879527863;
assign addr[18939] = -1870203416;
assign addr[18940] = -1860730673;
assign addr[18941] = -1851110385;
assign addr[18942] = -1841343316;
assign addr[18943] = -1831430239;
assign addr[18944] = -1821371941;
assign addr[18945] = -1811169220;
assign addr[18946] = -1800822883;
assign addr[18947] = -1790333753;
assign addr[18948] = -1779702660;
assign addr[18949] = -1768930447;
assign addr[18950] = -1758017969;
assign addr[18951] = -1746966091;
assign addr[18952] = -1735775690;
assign addr[18953] = -1724447652;
assign addr[18954] = -1712982875;
assign addr[18955] = -1701382270;
assign addr[18956] = -1689646755;
assign addr[18957] = -1677777262;
assign addr[18958] = -1665774731;
assign addr[18959] = -1653640115;
assign addr[18960] = -1641374375;
assign addr[18961] = -1628978484;
assign addr[18962] = -1616453425;
assign addr[18963] = -1603800191;
assign addr[18964] = -1591019785;
assign addr[18965] = -1578113222;
assign addr[18966] = -1565081523;
assign addr[18967] = -1551925723;
assign addr[18968] = -1538646865;
assign addr[18969] = -1525246002;
assign addr[18970] = -1511724196;
assign addr[18971] = -1498082520;
assign addr[18972] = -1484322054;
assign addr[18973] = -1470443891;
assign addr[18974] = -1456449131;
assign addr[18975] = -1442338884;
assign addr[18976] = -1428114267;
assign addr[18977] = -1413776410;
assign addr[18978] = -1399326449;
assign addr[18979] = -1384765530;
assign addr[18980] = -1370094808;
assign addr[18981] = -1355315445;
assign addr[18982] = -1340428615;
assign addr[18983] = -1325435496;
assign addr[18984] = -1310337279;
assign addr[18985] = -1295135159;
assign addr[18986] = -1279830344;
assign addr[18987] = -1264424045;
assign addr[18988] = -1248917486;
assign addr[18989] = -1233311895;
assign addr[18990] = -1217608510;
assign addr[18991] = -1201808576;
assign addr[18992] = -1185913346;
assign addr[18993] = -1169924081;
assign addr[18994] = -1153842047;
assign addr[18995] = -1137668521;
assign addr[18996] = -1121404785;
assign addr[18997] = -1105052128;
assign addr[18998] = -1088611847;
assign addr[18999] = -1072085246;
assign addr[19000] = -1055473635;
assign addr[19001] = -1038778332;
assign addr[19002] = -1022000660;
assign addr[19003] = -1005141949;
assign addr[19004] = -988203537;
assign addr[19005] = -971186766;
assign addr[19006] = -954092986;
assign addr[19007] = -936923553;
assign addr[19008] = -919679827;
assign addr[19009] = -902363176;
assign addr[19010] = -884974973;
assign addr[19011] = -867516597;
assign addr[19012] = -849989433;
assign addr[19013] = -832394869;
assign addr[19014] = -814734301;
assign addr[19015] = -797009130;
assign addr[19016] = -779220762;
assign addr[19017] = -761370605;
assign addr[19018] = -743460077;
assign addr[19019] = -725490597;
assign addr[19020] = -707463589;
assign addr[19021] = -689380485;
assign addr[19022] = -671242716;
assign addr[19023] = -653051723;
assign addr[19024] = -634808946;
assign addr[19025] = -616515832;
assign addr[19026] = -598173833;
assign addr[19027] = -579784402;
assign addr[19028] = -561348998;
assign addr[19029] = -542869083;
assign addr[19030] = -524346121;
assign addr[19031] = -505781581;
assign addr[19032] = -487176937;
assign addr[19033] = -468533662;
assign addr[19034] = -449853235;
assign addr[19035] = -431137138;
assign addr[19036] = -412386854;
assign addr[19037] = -393603870;
assign addr[19038] = -374789676;
assign addr[19039] = -355945764;
assign addr[19040] = -337073627;
assign addr[19041] = -318174762;
assign addr[19042] = -299250668;
assign addr[19043] = -280302845;
assign addr[19044] = -261332796;
assign addr[19045] = -242342025;
assign addr[19046] = -223332037;
assign addr[19047] = -204304341;
assign addr[19048] = -185260444;
assign addr[19049] = -166201858;
assign addr[19050] = -147130093;
assign addr[19051] = -128046661;
assign addr[19052] = -108953076;
assign addr[19053] = -89850852;
assign addr[19054] = -70741503;
assign addr[19055] = -51626544;
assign addr[19056] = -32507492;
assign addr[19057] = -13385863;
assign addr[19058] = 5736829;
assign addr[19059] = 24859065;
assign addr[19060] = 43979330;
assign addr[19061] = 63096108;
assign addr[19062] = 82207882;
assign addr[19063] = 101313138;
assign addr[19064] = 120410361;
assign addr[19065] = 139498035;
assign addr[19066] = 158574649;
assign addr[19067] = 177638688;
assign addr[19068] = 196688642;
assign addr[19069] = 215722999;
assign addr[19070] = 234740251;
assign addr[19071] = 253738890;
assign addr[19072] = 272717408;
assign addr[19073] = 291674302;
assign addr[19074] = 310608068;
assign addr[19075] = 329517204;
assign addr[19076] = 348400212;
assign addr[19077] = 367255594;
assign addr[19078] = 386081854;
assign addr[19079] = 404877501;
assign addr[19080] = 423641043;
assign addr[19081] = 442370993;
assign addr[19082] = 461065866;
assign addr[19083] = 479724180;
assign addr[19084] = 498344454;
assign addr[19085] = 516925212;
assign addr[19086] = 535464981;
assign addr[19087] = 553962291;
assign addr[19088] = 572415676;
assign addr[19089] = 590823671;
assign addr[19090] = 609184818;
assign addr[19091] = 627497660;
assign addr[19092] = 645760745;
assign addr[19093] = 663972625;
assign addr[19094] = 682131857;
assign addr[19095] = 700236999;
assign addr[19096] = 718286617;
assign addr[19097] = 736279279;
assign addr[19098] = 754213559;
assign addr[19099] = 772088034;
assign addr[19100] = 789901288;
assign addr[19101] = 807651907;
assign addr[19102] = 825338484;
assign addr[19103] = 842959617;
assign addr[19104] = 860513908;
assign addr[19105] = 877999966;
assign addr[19106] = 895416404;
assign addr[19107] = 912761841;
assign addr[19108] = 930034901;
assign addr[19109] = 947234215;
assign addr[19110] = 964358420;
assign addr[19111] = 981406156;
assign addr[19112] = 998376073;
assign addr[19113] = 1015266825;
assign addr[19114] = 1032077073;
assign addr[19115] = 1048805483;
assign addr[19116] = 1065450729;
assign addr[19117] = 1082011492;
assign addr[19118] = 1098486458;
assign addr[19119] = 1114874320;
assign addr[19120] = 1131173780;
assign addr[19121] = 1147383544;
assign addr[19122] = 1163502328;
assign addr[19123] = 1179528853;
assign addr[19124] = 1195461849;
assign addr[19125] = 1211300053;
assign addr[19126] = 1227042207;
assign addr[19127] = 1242687064;
assign addr[19128] = 1258233384;
assign addr[19129] = 1273679934;
assign addr[19130] = 1289025489;
assign addr[19131] = 1304268832;
assign addr[19132] = 1319408754;
assign addr[19133] = 1334444055;
assign addr[19134] = 1349373543;
assign addr[19135] = 1364196034;
assign addr[19136] = 1378910353;
assign addr[19137] = 1393515332;
assign addr[19138] = 1408009814;
assign addr[19139] = 1422392650;
assign addr[19140] = 1436662698;
assign addr[19141] = 1450818828;
assign addr[19142] = 1464859917;
assign addr[19143] = 1478784851;
assign addr[19144] = 1492592527;
assign addr[19145] = 1506281850;
assign addr[19146] = 1519851733;
assign addr[19147] = 1533301101;
assign addr[19148] = 1546628888;
assign addr[19149] = 1559834037;
assign addr[19150] = 1572915501;
assign addr[19151] = 1585872242;
assign addr[19152] = 1598703233;
assign addr[19153] = 1611407456;
assign addr[19154] = 1623983905;
assign addr[19155] = 1636431582;
assign addr[19156] = 1648749499;
assign addr[19157] = 1660936681;
assign addr[19158] = 1672992161;
assign addr[19159] = 1684914983;
assign addr[19160] = 1696704201;
assign addr[19161] = 1708358881;
assign addr[19162] = 1719878099;
assign addr[19163] = 1731260941;
assign addr[19164] = 1742506504;
assign addr[19165] = 1753613897;
assign addr[19166] = 1764582240;
assign addr[19167] = 1775410662;
assign addr[19168] = 1786098304;
assign addr[19169] = 1796644320;
assign addr[19170] = 1807047873;
assign addr[19171] = 1817308138;
assign addr[19172] = 1827424302;
assign addr[19173] = 1837395562;
assign addr[19174] = 1847221128;
assign addr[19175] = 1856900221;
assign addr[19176] = 1866432072;
assign addr[19177] = 1875815927;
assign addr[19178] = 1885051042;
assign addr[19179] = 1894136683;
assign addr[19180] = 1903072131;
assign addr[19181] = 1911856677;
assign addr[19182] = 1920489624;
assign addr[19183] = 1928970288;
assign addr[19184] = 1937297997;
assign addr[19185] = 1945472089;
assign addr[19186] = 1953491918;
assign addr[19187] = 1961356847;
assign addr[19188] = 1969066252;
assign addr[19189] = 1976619522;
assign addr[19190] = 1984016058;
assign addr[19191] = 1991255274;
assign addr[19192] = 1998336596;
assign addr[19193] = 2005259462;
assign addr[19194] = 2012023322;
assign addr[19195] = 2018627642;
assign addr[19196] = 2025071897;
assign addr[19197] = 2031355576;
assign addr[19198] = 2037478181;
assign addr[19199] = 2043439226;
assign addr[19200] = 2049238240;
assign addr[19201] = 2054874761;
assign addr[19202] = 2060348343;
assign addr[19203] = 2065658552;
assign addr[19204] = 2070804967;
assign addr[19205] = 2075787180;
assign addr[19206] = 2080604795;
assign addr[19207] = 2085257431;
assign addr[19208] = 2089744719;
assign addr[19209] = 2094066304;
assign addr[19210] = 2098221841;
assign addr[19211] = 2102211002;
assign addr[19212] = 2106033471;
assign addr[19213] = 2109688944;
assign addr[19214] = 2113177132;
assign addr[19215] = 2116497758;
assign addr[19216] = 2119650558;
assign addr[19217] = 2122635283;
assign addr[19218] = 2125451696;
assign addr[19219] = 2128099574;
assign addr[19220] = 2130578706;
assign addr[19221] = 2132888897;
assign addr[19222] = 2135029962;
assign addr[19223] = 2137001733;
assign addr[19224] = 2138804053;
assign addr[19225] = 2140436778;
assign addr[19226] = 2141899780;
assign addr[19227] = 2143192942;
assign addr[19228] = 2144316162;
assign addr[19229] = 2145269351;
assign addr[19230] = 2146052433;
assign addr[19231] = 2146665347;
assign addr[19232] = 2147108043;
assign addr[19233] = 2147380486;
assign addr[19234] = 2147482655;
assign addr[19235] = 2147414542;
assign addr[19236] = 2147176152;
assign addr[19237] = 2146767505;
assign addr[19238] = 2146188631;
assign addr[19239] = 2145439578;
assign addr[19240] = 2144520405;
assign addr[19241] = 2143431184;
assign addr[19242] = 2142172003;
assign addr[19243] = 2140742960;
assign addr[19244] = 2139144169;
assign addr[19245] = 2137375758;
assign addr[19246] = 2135437865;
assign addr[19247] = 2133330646;
assign addr[19248] = 2131054266;
assign addr[19249] = 2128608907;
assign addr[19250] = 2125994762;
assign addr[19251] = 2123212038;
assign addr[19252] = 2120260957;
assign addr[19253] = 2117141752;
assign addr[19254] = 2113854671;
assign addr[19255] = 2110399974;
assign addr[19256] = 2106777935;
assign addr[19257] = 2102988841;
assign addr[19258] = 2099032994;
assign addr[19259] = 2094910706;
assign addr[19260] = 2090622304;
assign addr[19261] = 2086168128;
assign addr[19262] = 2081548533;
assign addr[19263] = 2076763883;
assign addr[19264] = 2071814558;
assign addr[19265] = 2066700952;
assign addr[19266] = 2061423468;
assign addr[19267] = 2055982526;
assign addr[19268] = 2050378558;
assign addr[19269] = 2044612007;
assign addr[19270] = 2038683330;
assign addr[19271] = 2032592999;
assign addr[19272] = 2026341495;
assign addr[19273] = 2019929315;
assign addr[19274] = 2013356967;
assign addr[19275] = 2006624971;
assign addr[19276] = 1999733863;
assign addr[19277] = 1992684188;
assign addr[19278] = 1985476506;
assign addr[19279] = 1978111387;
assign addr[19280] = 1970589416;
assign addr[19281] = 1962911189;
assign addr[19282] = 1955077316;
assign addr[19283] = 1947088417;
assign addr[19284] = 1938945125;
assign addr[19285] = 1930648088;
assign addr[19286] = 1922197961;
assign addr[19287] = 1913595416;
assign addr[19288] = 1904841135;
assign addr[19289] = 1895935811;
assign addr[19290] = 1886880151;
assign addr[19291] = 1877674873;
assign addr[19292] = 1868320707;
assign addr[19293] = 1858818395;
assign addr[19294] = 1849168689;
assign addr[19295] = 1839372356;
assign addr[19296] = 1829430172;
assign addr[19297] = 1819342925;
assign addr[19298] = 1809111415;
assign addr[19299] = 1798736454;
assign addr[19300] = 1788218865;
assign addr[19301] = 1777559480;
assign addr[19302] = 1766759146;
assign addr[19303] = 1755818718;
assign addr[19304] = 1744739065;
assign addr[19305] = 1733521064;
assign addr[19306] = 1722165606;
assign addr[19307] = 1710673591;
assign addr[19308] = 1699045930;
assign addr[19309] = 1687283545;
assign addr[19310] = 1675387369;
assign addr[19311] = 1663358344;
assign addr[19312] = 1651197426;
assign addr[19313] = 1638905577;
assign addr[19314] = 1626483774;
assign addr[19315] = 1613933000;
assign addr[19316] = 1601254251;
assign addr[19317] = 1588448533;
assign addr[19318] = 1575516860;
assign addr[19319] = 1562460258;
assign addr[19320] = 1549279763;
assign addr[19321] = 1535976419;
assign addr[19322] = 1522551282;
assign addr[19323] = 1509005416;
assign addr[19324] = 1495339895;
assign addr[19325] = 1481555802;
assign addr[19326] = 1467654232;
assign addr[19327] = 1453636285;
assign addr[19328] = 1439503074;
assign addr[19329] = 1425255719;
assign addr[19330] = 1410895350;
assign addr[19331] = 1396423105;
assign addr[19332] = 1381840133;
assign addr[19333] = 1367147589;
assign addr[19334] = 1352346639;
assign addr[19335] = 1337438456;
assign addr[19336] = 1322424222;
assign addr[19337] = 1307305128;
assign addr[19338] = 1292082373;
assign addr[19339] = 1276757164;
assign addr[19340] = 1261330715;
assign addr[19341] = 1245804251;
assign addr[19342] = 1230179002;
assign addr[19343] = 1214456207;
assign addr[19344] = 1198637114;
assign addr[19345] = 1182722976;
assign addr[19346] = 1166715055;
assign addr[19347] = 1150614620;
assign addr[19348] = 1134422949;
assign addr[19349] = 1118141326;
assign addr[19350] = 1101771040;
assign addr[19351] = 1085313391;
assign addr[19352] = 1068769683;
assign addr[19353] = 1052141228;
assign addr[19354] = 1035429345;
assign addr[19355] = 1018635358;
assign addr[19356] = 1001760600;
assign addr[19357] = 984806408;
assign addr[19358] = 967774128;
assign addr[19359] = 950665109;
assign addr[19360] = 933480707;
assign addr[19361] = 916222287;
assign addr[19362] = 898891215;
assign addr[19363] = 881488868;
assign addr[19364] = 864016623;
assign addr[19365] = 846475867;
assign addr[19366] = 828867991;
assign addr[19367] = 811194391;
assign addr[19368] = 793456467;
assign addr[19369] = 775655628;
assign addr[19370] = 757793284;
assign addr[19371] = 739870851;
assign addr[19372] = 721889752;
assign addr[19373] = 703851410;
assign addr[19374] = 685757258;
assign addr[19375] = 667608730;
assign addr[19376] = 649407264;
assign addr[19377] = 631154304;
assign addr[19378] = 612851297;
assign addr[19379] = 594499695;
assign addr[19380] = 576100953;
assign addr[19381] = 557656529;
assign addr[19382] = 539167887;
assign addr[19383] = 520636492;
assign addr[19384] = 502063814;
assign addr[19385] = 483451325;
assign addr[19386] = 464800501;
assign addr[19387] = 446112822;
assign addr[19388] = 427389768;
assign addr[19389] = 408632825;
assign addr[19390] = 389843480;
assign addr[19391] = 371023223;
assign addr[19392] = 352173546;
assign addr[19393] = 333295944;
assign addr[19394] = 314391913;
assign addr[19395] = 295462954;
assign addr[19396] = 276510565;
assign addr[19397] = 257536251;
assign addr[19398] = 238541516;
assign addr[19399] = 219527866;
assign addr[19400] = 200496809;
assign addr[19401] = 181449854;
assign addr[19402] = 162388511;
assign addr[19403] = 143314291;
assign addr[19404] = 124228708;
assign addr[19405] = 105133274;
assign addr[19406] = 86029503;
assign addr[19407] = 66918911;
assign addr[19408] = 47803013;
assign addr[19409] = 28683324;
assign addr[19410] = 9561361;
assign addr[19411] = -9561361;
assign addr[19412] = -28683324;
assign addr[19413] = -47803013;
assign addr[19414] = -66918911;
assign addr[19415] = -86029503;
assign addr[19416] = -105133274;
assign addr[19417] = -124228708;
assign addr[19418] = -143314291;
assign addr[19419] = -162388511;
assign addr[19420] = -181449854;
assign addr[19421] = -200496809;
assign addr[19422] = -219527866;
assign addr[19423] = -238541516;
assign addr[19424] = -257536251;
assign addr[19425] = -276510565;
assign addr[19426] = -295462953;
assign addr[19427] = -314391913;
assign addr[19428] = -333295944;
assign addr[19429] = -352173546;
assign addr[19430] = -371023223;
assign addr[19431] = -389843480;
assign addr[19432] = -408632825;
assign addr[19433] = -427389768;
assign addr[19434] = -446112822;
assign addr[19435] = -464800501;
assign addr[19436] = -483451325;
assign addr[19437] = -502063814;
assign addr[19438] = -520636492;
assign addr[19439] = -539167887;
assign addr[19440] = -557656529;
assign addr[19441] = -576100953;
assign addr[19442] = -594499695;
assign addr[19443] = -612851297;
assign addr[19444] = -631154304;
assign addr[19445] = -649407264;
assign addr[19446] = -667608730;
assign addr[19447] = -685757258;
assign addr[19448] = -703851410;
assign addr[19449] = -721889752;
assign addr[19450] = -739870851;
assign addr[19451] = -757793284;
assign addr[19452] = -775655628;
assign addr[19453] = -793456467;
assign addr[19454] = -811194391;
assign addr[19455] = -828867991;
assign addr[19456] = -846475867;
assign addr[19457] = -864016623;
assign addr[19458] = -881488868;
assign addr[19459] = -898891215;
assign addr[19460] = -916222287;
assign addr[19461] = -933480707;
assign addr[19462] = -950665109;
assign addr[19463] = -967774128;
assign addr[19464] = -984806408;
assign addr[19465] = -1001760600;
assign addr[19466] = -1018635358;
assign addr[19467] = -1035429345;
assign addr[19468] = -1052141228;
assign addr[19469] = -1068769683;
assign addr[19470] = -1085313391;
assign addr[19471] = -1101771040;
assign addr[19472] = -1118141326;
assign addr[19473] = -1134422949;
assign addr[19474] = -1150614620;
assign addr[19475] = -1166715055;
assign addr[19476] = -1182722976;
assign addr[19477] = -1198637114;
assign addr[19478] = -1214456207;
assign addr[19479] = -1230179002;
assign addr[19480] = -1245804251;
assign addr[19481] = -1261330715;
assign addr[19482] = -1276757164;
assign addr[19483] = -1292082373;
assign addr[19484] = -1307305128;
assign addr[19485] = -1322424222;
assign addr[19486] = -1337438456;
assign addr[19487] = -1352346639;
assign addr[19488] = -1367147589;
assign addr[19489] = -1381840133;
assign addr[19490] = -1396423105;
assign addr[19491] = -1410895350;
assign addr[19492] = -1425255719;
assign addr[19493] = -1439503074;
assign addr[19494] = -1453636285;
assign addr[19495] = -1467654232;
assign addr[19496] = -1481555802;
assign addr[19497] = -1495339895;
assign addr[19498] = -1509005416;
assign addr[19499] = -1522551282;
assign addr[19500] = -1535976419;
assign addr[19501] = -1549279763;
assign addr[19502] = -1562460258;
assign addr[19503] = -1575516860;
assign addr[19504] = -1588448533;
assign addr[19505] = -1601254251;
assign addr[19506] = -1613933000;
assign addr[19507] = -1626483774;
assign addr[19508] = -1638905577;
assign addr[19509] = -1651197426;
assign addr[19510] = -1663358344;
assign addr[19511] = -1675387369;
assign addr[19512] = -1687283545;
assign addr[19513] = -1699045930;
assign addr[19514] = -1710673591;
assign addr[19515] = -1722165606;
assign addr[19516] = -1733521064;
assign addr[19517] = -1744739065;
assign addr[19518] = -1755818718;
assign addr[19519] = -1766759146;
assign addr[19520] = -1777559480;
assign addr[19521] = -1788218865;
assign addr[19522] = -1798736454;
assign addr[19523] = -1809111415;
assign addr[19524] = -1819342925;
assign addr[19525] = -1829430172;
assign addr[19526] = -1839372356;
assign addr[19527] = -1849168689;
assign addr[19528] = -1858818395;
assign addr[19529] = -1868320707;
assign addr[19530] = -1877674873;
assign addr[19531] = -1886880151;
assign addr[19532] = -1895935811;
assign addr[19533] = -1904841135;
assign addr[19534] = -1913595416;
assign addr[19535] = -1922197961;
assign addr[19536] = -1930648088;
assign addr[19537] = -1938945125;
assign addr[19538] = -1947088417;
assign addr[19539] = -1955077316;
assign addr[19540] = -1962911189;
assign addr[19541] = -1970589416;
assign addr[19542] = -1978111387;
assign addr[19543] = -1985476506;
assign addr[19544] = -1992684188;
assign addr[19545] = -1999733863;
assign addr[19546] = -2006624971;
assign addr[19547] = -2013356967;
assign addr[19548] = -2019929315;
assign addr[19549] = -2026341495;
assign addr[19550] = -2032592999;
assign addr[19551] = -2038683330;
assign addr[19552] = -2044612007;
assign addr[19553] = -2050378558;
assign addr[19554] = -2055982526;
assign addr[19555] = -2061423468;
assign addr[19556] = -2066700952;
assign addr[19557] = -2071814558;
assign addr[19558] = -2076763883;
assign addr[19559] = -2081548533;
assign addr[19560] = -2086168128;
assign addr[19561] = -2090622304;
assign addr[19562] = -2094910706;
assign addr[19563] = -2099032994;
assign addr[19564] = -2102988841;
assign addr[19565] = -2106777935;
assign addr[19566] = -2110399974;
assign addr[19567] = -2113854671;
assign addr[19568] = -2117141752;
assign addr[19569] = -2120260957;
assign addr[19570] = -2123212038;
assign addr[19571] = -2125994762;
assign addr[19572] = -2128608907;
assign addr[19573] = -2131054266;
assign addr[19574] = -2133330646;
assign addr[19575] = -2135437865;
assign addr[19576] = -2137375758;
assign addr[19577] = -2139144169;
assign addr[19578] = -2140742960;
assign addr[19579] = -2142172003;
assign addr[19580] = -2143431184;
assign addr[19581] = -2144520405;
assign addr[19582] = -2145439578;
assign addr[19583] = -2146188631;
assign addr[19584] = -2146767505;
assign addr[19585] = -2147176152;
assign addr[19586] = -2147414542;
assign addr[19587] = -2147482655;
assign addr[19588] = -2147380486;
assign addr[19589] = -2147108043;
assign addr[19590] = -2146665347;
assign addr[19591] = -2146052433;
assign addr[19592] = -2145269351;
assign addr[19593] = -2144316162;
assign addr[19594] = -2143192942;
assign addr[19595] = -2141899780;
assign addr[19596] = -2140436778;
assign addr[19597] = -2138804053;
assign addr[19598] = -2137001733;
assign addr[19599] = -2135029962;
assign addr[19600] = -2132888897;
assign addr[19601] = -2130578706;
assign addr[19602] = -2128099574;
assign addr[19603] = -2125451696;
assign addr[19604] = -2122635283;
assign addr[19605] = -2119650558;
assign addr[19606] = -2116497758;
assign addr[19607] = -2113177132;
assign addr[19608] = -2109688944;
assign addr[19609] = -2106033471;
assign addr[19610] = -2102211002;
assign addr[19611] = -2098221841;
assign addr[19612] = -2094066304;
assign addr[19613] = -2089744719;
assign addr[19614] = -2085257431;
assign addr[19615] = -2080604795;
assign addr[19616] = -2075787180;
assign addr[19617] = -2070804967;
assign addr[19618] = -2065658552;
assign addr[19619] = -2060348343;
assign addr[19620] = -2054874761;
assign addr[19621] = -2049238240;
assign addr[19622] = -2043439226;
assign addr[19623] = -2037478181;
assign addr[19624] = -2031355576;
assign addr[19625] = -2025071897;
assign addr[19626] = -2018627642;
assign addr[19627] = -2012023322;
assign addr[19628] = -2005259462;
assign addr[19629] = -1998336596;
assign addr[19630] = -1991255274;
assign addr[19631] = -1984016058;
assign addr[19632] = -1976619522;
assign addr[19633] = -1969066252;
assign addr[19634] = -1961356847;
assign addr[19635] = -1953491918;
assign addr[19636] = -1945472089;
assign addr[19637] = -1937297997;
assign addr[19638] = -1928970288;
assign addr[19639] = -1920489624;
assign addr[19640] = -1911856677;
assign addr[19641] = -1903072131;
assign addr[19642] = -1894136683;
assign addr[19643] = -1885051042;
assign addr[19644] = -1875815927;
assign addr[19645] = -1866432072;
assign addr[19646] = -1856900221;
assign addr[19647] = -1847221128;
assign addr[19648] = -1837395562;
assign addr[19649] = -1827424302;
assign addr[19650] = -1817308138;
assign addr[19651] = -1807047873;
assign addr[19652] = -1796644320;
assign addr[19653] = -1786098304;
assign addr[19654] = -1775410662;
assign addr[19655] = -1764582240;
assign addr[19656] = -1753613897;
assign addr[19657] = -1742506504;
assign addr[19658] = -1731260941;
assign addr[19659] = -1719878099;
assign addr[19660] = -1708358881;
assign addr[19661] = -1696704201;
assign addr[19662] = -1684914983;
assign addr[19663] = -1672992161;
assign addr[19664] = -1660936681;
assign addr[19665] = -1648749499;
assign addr[19666] = -1636431582;
assign addr[19667] = -1623983905;
assign addr[19668] = -1611407456;
assign addr[19669] = -1598703233;
assign addr[19670] = -1585872242;
assign addr[19671] = -1572915501;
assign addr[19672] = -1559834037;
assign addr[19673] = -1546628888;
assign addr[19674] = -1533301101;
assign addr[19675] = -1519851733;
assign addr[19676] = -1506281850;
assign addr[19677] = -1492592527;
assign addr[19678] = -1478784851;
assign addr[19679] = -1464859917;
assign addr[19680] = -1450818828;
assign addr[19681] = -1436662698;
assign addr[19682] = -1422392650;
assign addr[19683] = -1408009814;
assign addr[19684] = -1393515332;
assign addr[19685] = -1378910353;
assign addr[19686] = -1364196034;
assign addr[19687] = -1349373543;
assign addr[19688] = -1334444055;
assign addr[19689] = -1319408754;
assign addr[19690] = -1304268832;
assign addr[19691] = -1289025489;
assign addr[19692] = -1273679934;
assign addr[19693] = -1258233384;
assign addr[19694] = -1242687064;
assign addr[19695] = -1227042207;
assign addr[19696] = -1211300053;
assign addr[19697] = -1195461849;
assign addr[19698] = -1179528853;
assign addr[19699] = -1163502328;
assign addr[19700] = -1147383544;
assign addr[19701] = -1131173780;
assign addr[19702] = -1114874320;
assign addr[19703] = -1098486458;
assign addr[19704] = -1082011492;
assign addr[19705] = -1065450729;
assign addr[19706] = -1048805483;
assign addr[19707] = -1032077073;
assign addr[19708] = -1015266825;
assign addr[19709] = -998376073;
assign addr[19710] = -981406156;
assign addr[19711] = -964358420;
assign addr[19712] = -947234215;
assign addr[19713] = -930034901;
assign addr[19714] = -912761841;
assign addr[19715] = -895416404;
assign addr[19716] = -877999966;
assign addr[19717] = -860513908;
assign addr[19718] = -842959617;
assign addr[19719] = -825338484;
assign addr[19720] = -807651907;
assign addr[19721] = -789901288;
assign addr[19722] = -772088034;
assign addr[19723] = -754213559;
assign addr[19724] = -736279279;
assign addr[19725] = -718286617;
assign addr[19726] = -700236999;
assign addr[19727] = -682131857;
assign addr[19728] = -663972625;
assign addr[19729] = -645760745;
assign addr[19730] = -627497660;
assign addr[19731] = -609184818;
assign addr[19732] = -590823671;
assign addr[19733] = -572415676;
assign addr[19734] = -553962291;
assign addr[19735] = -535464981;
assign addr[19736] = -516925212;
assign addr[19737] = -498344454;
assign addr[19738] = -479724180;
assign addr[19739] = -461065866;
assign addr[19740] = -442370993;
assign addr[19741] = -423641043;
assign addr[19742] = -404877501;
assign addr[19743] = -386081854;
assign addr[19744] = -367255594;
assign addr[19745] = -348400212;
assign addr[19746] = -329517204;
assign addr[19747] = -310608068;
assign addr[19748] = -291674302;
assign addr[19749] = -272717408;
assign addr[19750] = -253738890;
assign addr[19751] = -234740251;
assign addr[19752] = -215722999;
assign addr[19753] = -196688642;
assign addr[19754] = -177638688;
assign addr[19755] = -158574649;
assign addr[19756] = -139498035;
assign addr[19757] = -120410361;
assign addr[19758] = -101313138;
assign addr[19759] = -82207882;
assign addr[19760] = -63096108;
assign addr[19761] = -43979330;
assign addr[19762] = -24859065;
assign addr[19763] = -5736829;
assign addr[19764] = 13385863;
assign addr[19765] = 32507492;
assign addr[19766] = 51626544;
assign addr[19767] = 70741503;
assign addr[19768] = 89850852;
assign addr[19769] = 108953076;
assign addr[19770] = 128046661;
assign addr[19771] = 147130093;
assign addr[19772] = 166201858;
assign addr[19773] = 185260444;
assign addr[19774] = 204304341;
assign addr[19775] = 223332037;
assign addr[19776] = 242342025;
assign addr[19777] = 261332796;
assign addr[19778] = 280302845;
assign addr[19779] = 299250668;
assign addr[19780] = 318174762;
assign addr[19781] = 337073627;
assign addr[19782] = 355945764;
assign addr[19783] = 374789676;
assign addr[19784] = 393603870;
assign addr[19785] = 412386854;
assign addr[19786] = 431137138;
assign addr[19787] = 449853235;
assign addr[19788] = 468533662;
assign addr[19789] = 487176937;
assign addr[19790] = 505781581;
assign addr[19791] = 524346121;
assign addr[19792] = 542869083;
assign addr[19793] = 561348998;
assign addr[19794] = 579784402;
assign addr[19795] = 598173833;
assign addr[19796] = 616515832;
assign addr[19797] = 634808946;
assign addr[19798] = 653051723;
assign addr[19799] = 671242716;
assign addr[19800] = 689380485;
assign addr[19801] = 707463589;
assign addr[19802] = 725490597;
assign addr[19803] = 743460077;
assign addr[19804] = 761370605;
assign addr[19805] = 779220762;
assign addr[19806] = 797009130;
assign addr[19807] = 814734301;
assign addr[19808] = 832394869;
assign addr[19809] = 849989433;
assign addr[19810] = 867516597;
assign addr[19811] = 884974973;
assign addr[19812] = 902363176;
assign addr[19813] = 919679827;
assign addr[19814] = 936923553;
assign addr[19815] = 954092986;
assign addr[19816] = 971186766;
assign addr[19817] = 988203537;
assign addr[19818] = 1005141949;
assign addr[19819] = 1022000660;
assign addr[19820] = 1038778332;
assign addr[19821] = 1055473635;
assign addr[19822] = 1072085246;
assign addr[19823] = 1088611847;
assign addr[19824] = 1105052128;
assign addr[19825] = 1121404785;
assign addr[19826] = 1137668521;
assign addr[19827] = 1153842047;
assign addr[19828] = 1169924081;
assign addr[19829] = 1185913346;
assign addr[19830] = 1201808576;
assign addr[19831] = 1217608510;
assign addr[19832] = 1233311895;
assign addr[19833] = 1248917486;
assign addr[19834] = 1264424045;
assign addr[19835] = 1279830344;
assign addr[19836] = 1295135159;
assign addr[19837] = 1310337279;
assign addr[19838] = 1325435496;
assign addr[19839] = 1340428615;
assign addr[19840] = 1355315445;
assign addr[19841] = 1370094808;
assign addr[19842] = 1384765530;
assign addr[19843] = 1399326449;
assign addr[19844] = 1413776410;
assign addr[19845] = 1428114267;
assign addr[19846] = 1442338884;
assign addr[19847] = 1456449131;
assign addr[19848] = 1470443891;
assign addr[19849] = 1484322054;
assign addr[19850] = 1498082520;
assign addr[19851] = 1511724196;
assign addr[19852] = 1525246002;
assign addr[19853] = 1538646865;
assign addr[19854] = 1551925723;
assign addr[19855] = 1565081523;
assign addr[19856] = 1578113222;
assign addr[19857] = 1591019785;
assign addr[19858] = 1603800191;
assign addr[19859] = 1616453425;
assign addr[19860] = 1628978484;
assign addr[19861] = 1641374375;
assign addr[19862] = 1653640115;
assign addr[19863] = 1665774731;
assign addr[19864] = 1677777262;
assign addr[19865] = 1689646755;
assign addr[19866] = 1701382270;
assign addr[19867] = 1712982875;
assign addr[19868] = 1724447652;
assign addr[19869] = 1735775690;
assign addr[19870] = 1746966091;
assign addr[19871] = 1758017969;
assign addr[19872] = 1768930447;
assign addr[19873] = 1779702660;
assign addr[19874] = 1790333753;
assign addr[19875] = 1800822883;
assign addr[19876] = 1811169220;
assign addr[19877] = 1821371941;
assign addr[19878] = 1831430239;
assign addr[19879] = 1841343316;
assign addr[19880] = 1851110385;
assign addr[19881] = 1860730673;
assign addr[19882] = 1870203416;
assign addr[19883] = 1879527863;
assign addr[19884] = 1888703276;
assign addr[19885] = 1897728925;
assign addr[19886] = 1906604097;
assign addr[19887] = 1915328086;
assign addr[19888] = 1923900201;
assign addr[19889] = 1932319763;
assign addr[19890] = 1940586104;
assign addr[19891] = 1948698568;
assign addr[19892] = 1956656513;
assign addr[19893] = 1964459306;
assign addr[19894] = 1972106330;
assign addr[19895] = 1979596978;
assign addr[19896] = 1986930656;
assign addr[19897] = 1994106782;
assign addr[19898] = 2001124788;
assign addr[19899] = 2007984117;
assign addr[19900] = 2014684225;
assign addr[19901] = 2021224581;
assign addr[19902] = 2027604666;
assign addr[19903] = 2033823974;
assign addr[19904] = 2039882013;
assign addr[19905] = 2045778302;
assign addr[19906] = 2051512372;
assign addr[19907] = 2057083771;
assign addr[19908] = 2062492055;
assign addr[19909] = 2067736796;
assign addr[19910] = 2072817579;
assign addr[19911] = 2077733999;
assign addr[19912] = 2082485668;
assign addr[19913] = 2087072209;
assign addr[19914] = 2091493257;
assign addr[19915] = 2095748463;
assign addr[19916] = 2099837489;
assign addr[19917] = 2103760010;
assign addr[19918] = 2107515716;
assign addr[19919] = 2111104309;
assign addr[19920] = 2114525505;
assign addr[19921] = 2117779031;
assign addr[19922] = 2120864631;
assign addr[19923] = 2123782059;
assign addr[19924] = 2126531084;
assign addr[19925] = 2129111488;
assign addr[19926] = 2131523066;
assign addr[19927] = 2133765628;
assign addr[19928] = 2135838995;
assign addr[19929] = 2137743003;
assign addr[19930] = 2139477502;
assign addr[19931] = 2141042352;
assign addr[19932] = 2142437431;
assign addr[19933] = 2143662628;
assign addr[19934] = 2144717846;
assign addr[19935] = 2145603001;
assign addr[19936] = 2146318022;
assign addr[19937] = 2146862854;
assign addr[19938] = 2147237452;
assign addr[19939] = 2147441787;
assign addr[19940] = 2147475844;
assign addr[19941] = 2147339619;
assign addr[19942] = 2147033123;
assign addr[19943] = 2146556380;
assign addr[19944] = 2145909429;
assign addr[19945] = 2145092320;
assign addr[19946] = 2144105118;
assign addr[19947] = 2142947902;
assign addr[19948] = 2141620763;
assign addr[19949] = 2140123807;
assign addr[19950] = 2138457152;
assign addr[19951] = 2136620930;
assign addr[19952] = 2134615288;
assign addr[19953] = 2132440383;
assign addr[19954] = 2130096389;
assign addr[19955] = 2127583492;
assign addr[19956] = 2124901890;
assign addr[19957] = 2122051796;
assign addr[19958] = 2119033436;
assign addr[19959] = 2115847050;
assign addr[19960] = 2112492891;
assign addr[19961] = 2108971223;
assign addr[19962] = 2105282327;
assign addr[19963] = 2101426496;
assign addr[19964] = 2097404033;
assign addr[19965] = 2093215260;
assign addr[19966] = 2088860507;
assign addr[19967] = 2084340120;
assign addr[19968] = 2079654458;
assign addr[19969] = 2074803892;
assign addr[19970] = 2069788807;
assign addr[19971] = 2064609600;
assign addr[19972] = 2059266683;
assign addr[19973] = 2053760478;
assign addr[19974] = 2048091422;
assign addr[19975] = 2042259965;
assign addr[19976] = 2036266570;
assign addr[19977] = 2030111710;
assign addr[19978] = 2023795876;
assign addr[19979] = 2017319567;
assign addr[19980] = 2010683297;
assign addr[19981] = 2003887591;
assign addr[19982] = 1996932990;
assign addr[19983] = 1989820044;
assign addr[19984] = 1982549318;
assign addr[19985] = 1975121388;
assign addr[19986] = 1967536842;
assign addr[19987] = 1959796283;
assign addr[19988] = 1951900324;
assign addr[19989] = 1943849591;
assign addr[19990] = 1935644723;
assign addr[19991] = 1927286370;
assign addr[19992] = 1918775195;
assign addr[19993] = 1910111873;
assign addr[19994] = 1901297091;
assign addr[19995] = 1892331547;
assign addr[19996] = 1883215953;
assign addr[19997] = 1873951032;
assign addr[19998] = 1864537518;
assign addr[19999] = 1854976157;
assign addr[20000] = 1845267708;
assign addr[20001] = 1835412941;
assign addr[20002] = 1825412636;
assign addr[20003] = 1815267588;
assign addr[20004] = 1804978599;
assign addr[20005] = 1794546487;
assign addr[20006] = 1783972079;
assign addr[20007] = 1773256212;
assign addr[20008] = 1762399737;
assign addr[20009] = 1751403515;
assign addr[20010] = 1740268417;
assign addr[20011] = 1728995326;
assign addr[20012] = 1717585136;
assign addr[20013] = 1706038753;
assign addr[20014] = 1694357091;
assign addr[20015] = 1682541077;
assign addr[20016] = 1670591647;
assign addr[20017] = 1658509750;
assign addr[20018] = 1646296344;
assign addr[20019] = 1633952396;
assign addr[20020] = 1621478885;
assign addr[20021] = 1608876801;
assign addr[20022] = 1596147143;
assign addr[20023] = 1583290921;
assign addr[20024] = 1570309153;
assign addr[20025] = 1557202869;
assign addr[20026] = 1543973108;
assign addr[20027] = 1530620920;
assign addr[20028] = 1517147363;
assign addr[20029] = 1503553506;
assign addr[20030] = 1489840425;
assign addr[20031] = 1476009210;
assign addr[20032] = 1462060956;
assign addr[20033] = 1447996770;
assign addr[20034] = 1433817766;
assign addr[20035] = 1419525069;
assign addr[20036] = 1405119813;
assign addr[20037] = 1390603139;
assign addr[20038] = 1375976199;
assign addr[20039] = 1361240152;
assign addr[20040] = 1346396168;
assign addr[20041] = 1331445422;
assign addr[20042] = 1316389101;
assign addr[20043] = 1301228398;
assign addr[20044] = 1285964516;
assign addr[20045] = 1270598665;
assign addr[20046] = 1255132063;
assign addr[20047] = 1239565936;
assign addr[20048] = 1223901520;
assign addr[20049] = 1208140056;
assign addr[20050] = 1192282793;
assign addr[20051] = 1176330990;
assign addr[20052] = 1160285911;
assign addr[20053] = 1144148829;
assign addr[20054] = 1127921022;
assign addr[20055] = 1111603778;
assign addr[20056] = 1095198391;
assign addr[20057] = 1078706161;
assign addr[20058] = 1062128397;
assign addr[20059] = 1045466412;
assign addr[20060] = 1028721528;
assign addr[20061] = 1011895073;
assign addr[20062] = 994988380;
assign addr[20063] = 978002791;
assign addr[20064] = 960939653;
assign addr[20065] = 943800318;
assign addr[20066] = 926586145;
assign addr[20067] = 909298500;
assign addr[20068] = 891938752;
assign addr[20069] = 874508280;
assign addr[20070] = 857008464;
assign addr[20071] = 839440693;
assign addr[20072] = 821806359;
assign addr[20073] = 804106861;
assign addr[20074] = 786343603;
assign addr[20075] = 768517992;
assign addr[20076] = 750631442;
assign addr[20077] = 732685372;
assign addr[20078] = 714681204;
assign addr[20079] = 696620367;
assign addr[20080] = 678504291;
assign addr[20081] = 660334415;
assign addr[20082] = 642112178;
assign addr[20083] = 623839025;
assign addr[20084] = 605516406;
assign addr[20085] = 587145773;
assign addr[20086] = 568728583;
assign addr[20087] = 550266296;
assign addr[20088] = 531760377;
assign addr[20089] = 513212292;
assign addr[20090] = 494623513;
assign addr[20091] = 475995513;
assign addr[20092] = 457329769;
assign addr[20093] = 438627762;
assign addr[20094] = 419890975;
assign addr[20095] = 401120892;
assign addr[20096] = 382319004;
assign addr[20097] = 363486799;
assign addr[20098] = 344625773;
assign addr[20099] = 325737419;
assign addr[20100] = 306823237;
assign addr[20101] = 287884725;
assign addr[20102] = 268923386;
assign addr[20103] = 249940723;
assign addr[20104] = 230938242;
assign addr[20105] = 211917448;
assign addr[20106] = 192879850;
assign addr[20107] = 173826959;
assign addr[20108] = 154760284;
assign addr[20109] = 135681337;
assign addr[20110] = 116591632;
assign addr[20111] = 97492681;
assign addr[20112] = 78386000;
assign addr[20113] = 59273104;
assign addr[20114] = 40155507;
assign addr[20115] = 21034727;
assign addr[20116] = 1912278;
assign addr[20117] = -17210322;
assign addr[20118] = -36331557;
assign addr[20119] = -55449912;
assign addr[20120] = -74563870;
assign addr[20121] = -93671915;
assign addr[20122] = -112772533;
assign addr[20123] = -131864208;
assign addr[20124] = -150945428;
assign addr[20125] = -170014678;
assign addr[20126] = -189070447;
assign addr[20127] = -208111224;
assign addr[20128] = -227135500;
assign addr[20129] = -246141764;
assign addr[20130] = -265128512;
assign addr[20131] = -284094236;
assign addr[20132] = -303037433;
assign addr[20133] = -321956601;
assign addr[20134] = -340850240;
assign addr[20135] = -359716852;
assign addr[20136] = -378554940;
assign addr[20137] = -397363011;
assign addr[20138] = -416139574;
assign addr[20139] = -434883140;
assign addr[20140] = -453592221;
assign addr[20141] = -472265336;
assign addr[20142] = -490901003;
assign addr[20143] = -509497745;
assign addr[20144] = -528054086;
assign addr[20145] = -546568556;
assign addr[20146] = -565039687;
assign addr[20147] = -583466013;
assign addr[20148] = -601846074;
assign addr[20149] = -620178412;
assign addr[20150] = -638461574;
assign addr[20151] = -656694110;
assign addr[20152] = -674874574;
assign addr[20153] = -693001525;
assign addr[20154] = -711073524;
assign addr[20155] = -729089140;
assign addr[20156] = -747046944;
assign addr[20157] = -764945512;
assign addr[20158] = -782783424;
assign addr[20159] = -800559266;
assign addr[20160] = -818271628;
assign addr[20161] = -835919107;
assign addr[20162] = -853500302;
assign addr[20163] = -871013820;
assign addr[20164] = -888458272;
assign addr[20165] = -905832274;
assign addr[20166] = -923134450;
assign addr[20167] = -940363427;
assign addr[20168] = -957517838;
assign addr[20169] = -974596324;
assign addr[20170] = -991597531;
assign addr[20171] = -1008520110;
assign addr[20172] = -1025362720;
assign addr[20173] = -1042124025;
assign addr[20174] = -1058802695;
assign addr[20175] = -1075397409;
assign addr[20176] = -1091906851;
assign addr[20177] = -1108329711;
assign addr[20178] = -1124664687;
assign addr[20179] = -1140910484;
assign addr[20180] = -1157065814;
assign addr[20181] = -1173129396;
assign addr[20182] = -1189099956;
assign addr[20183] = -1204976227;
assign addr[20184] = -1220756951;
assign addr[20185] = -1236440877;
assign addr[20186] = -1252026760;
assign addr[20187] = -1267513365;
assign addr[20188] = -1282899464;
assign addr[20189] = -1298183838;
assign addr[20190] = -1313365273;
assign addr[20191] = -1328442566;
assign addr[20192] = -1343414522;
assign addr[20193] = -1358279953;
assign addr[20194] = -1373037681;
assign addr[20195] = -1387686535;
assign addr[20196] = -1402225355;
assign addr[20197] = -1416652986;
assign addr[20198] = -1430968286;
assign addr[20199] = -1445170118;
assign addr[20200] = -1459257358;
assign addr[20201] = -1473228887;
assign addr[20202] = -1487083598;
assign addr[20203] = -1500820393;
assign addr[20204] = -1514438181;
assign addr[20205] = -1527935884;
assign addr[20206] = -1541312431;
assign addr[20207] = -1554566762;
assign addr[20208] = -1567697824;
assign addr[20209] = -1580704578;
assign addr[20210] = -1593585992;
assign addr[20211] = -1606341043;
assign addr[20212] = -1618968722;
assign addr[20213] = -1631468027;
assign addr[20214] = -1643837966;
assign addr[20215] = -1656077559;
assign addr[20216] = -1668185835;
assign addr[20217] = -1680161834;
assign addr[20218] = -1692004606;
assign addr[20219] = -1703713213;
assign addr[20220] = -1715286726;
assign addr[20221] = -1726724227;
assign addr[20222] = -1738024810;
assign addr[20223] = -1749187577;
assign addr[20224] = -1760211645;
assign addr[20225] = -1771096139;
assign addr[20226] = -1781840195;
assign addr[20227] = -1792442963;
assign addr[20228] = -1802903601;
assign addr[20229] = -1813221279;
assign addr[20230] = -1823395180;
assign addr[20231] = -1833424497;
assign addr[20232] = -1843308435;
assign addr[20233] = -1853046210;
assign addr[20234] = -1862637049;
assign addr[20235] = -1872080193;
assign addr[20236] = -1881374892;
assign addr[20237] = -1890520410;
assign addr[20238] = -1899516021;
assign addr[20239] = -1908361011;
assign addr[20240] = -1917054681;
assign addr[20241] = -1925596340;
assign addr[20242] = -1933985310;
assign addr[20243] = -1942220928;
assign addr[20244] = -1950302539;
assign addr[20245] = -1958229503;
assign addr[20246] = -1966001192;
assign addr[20247] = -1973616989;
assign addr[20248] = -1981076290;
assign addr[20249] = -1988378503;
assign addr[20250] = -1995523051;
assign addr[20251] = -2002509365;
assign addr[20252] = -2009336893;
assign addr[20253] = -2016005093;
assign addr[20254] = -2022513436;
assign addr[20255] = -2028861406;
assign addr[20256] = -2035048499;
assign addr[20257] = -2041074226;
assign addr[20258] = -2046938108;
assign addr[20259] = -2052639680;
assign addr[20260] = -2058178491;
assign addr[20261] = -2063554100;
assign addr[20262] = -2068766083;
assign addr[20263] = -2073814024;
assign addr[20264] = -2078697525;
assign addr[20265] = -2083416198;
assign addr[20266] = -2087969669;
assign addr[20267] = -2092357577;
assign addr[20268] = -2096579573;
assign addr[20269] = -2100635323;
assign addr[20270] = -2104524506;
assign addr[20271] = -2108246813;
assign addr[20272] = -2111801949;
assign addr[20273] = -2115189632;
assign addr[20274] = -2118409593;
assign addr[20275] = -2121461578;
assign addr[20276] = -2124345343;
assign addr[20277] = -2127060661;
assign addr[20278] = -2129607316;
assign addr[20279] = -2131985106;
assign addr[20280] = -2134193842;
assign addr[20281] = -2136233350;
assign addr[20282] = -2138103468;
assign addr[20283] = -2139804048;
assign addr[20284] = -2141334954;
assign addr[20285] = -2142696065;
assign addr[20286] = -2143887273;
assign addr[20287] = -2144908484;
assign addr[20288] = -2145759618;
assign addr[20289] = -2146440605;
assign addr[20290] = -2146951393;
assign addr[20291] = -2147291941;
assign addr[20292] = -2147462221;
assign addr[20293] = -2147462221;
assign addr[20294] = -2147291941;
assign addr[20295] = -2146951393;
assign addr[20296] = -2146440605;
assign addr[20297] = -2145759618;
assign addr[20298] = -2144908484;
assign addr[20299] = -2143887273;
assign addr[20300] = -2142696065;
assign addr[20301] = -2141334954;
assign addr[20302] = -2139804048;
assign addr[20303] = -2138103468;
assign addr[20304] = -2136233350;
assign addr[20305] = -2134193842;
assign addr[20306] = -2131985106;
assign addr[20307] = -2129607316;
assign addr[20308] = -2127060661;
assign addr[20309] = -2124345343;
assign addr[20310] = -2121461578;
assign addr[20311] = -2118409593;
assign addr[20312] = -2115189632;
assign addr[20313] = -2111801949;
assign addr[20314] = -2108246813;
assign addr[20315] = -2104524506;
assign addr[20316] = -2100635323;
assign addr[20317] = -2096579573;
assign addr[20318] = -2092357577;
assign addr[20319] = -2087969669;
assign addr[20320] = -2083416198;
assign addr[20321] = -2078697525;
assign addr[20322] = -2073814024;
assign addr[20323] = -2068766083;
assign addr[20324] = -2063554100;
assign addr[20325] = -2058178491;
assign addr[20326] = -2052639680;
assign addr[20327] = -2046938108;
assign addr[20328] = -2041074226;
assign addr[20329] = -2035048499;
assign addr[20330] = -2028861406;
assign addr[20331] = -2022513436;
assign addr[20332] = -2016005093;
assign addr[20333] = -2009336893;
assign addr[20334] = -2002509365;
assign addr[20335] = -1995523051;
assign addr[20336] = -1988378503;
assign addr[20337] = -1981076290;
assign addr[20338] = -1973616989;
assign addr[20339] = -1966001192;
assign addr[20340] = -1958229503;
assign addr[20341] = -1950302539;
assign addr[20342] = -1942220928;
assign addr[20343] = -1933985310;
assign addr[20344] = -1925596340;
assign addr[20345] = -1917054681;
assign addr[20346] = -1908361011;
assign addr[20347] = -1899516021;
assign addr[20348] = -1890520410;
assign addr[20349] = -1881374892;
assign addr[20350] = -1872080193;
assign addr[20351] = -1862637049;
assign addr[20352] = -1853046210;
assign addr[20353] = -1843308435;
assign addr[20354] = -1833424497;
assign addr[20355] = -1823395180;
assign addr[20356] = -1813221279;
assign addr[20357] = -1802903601;
assign addr[20358] = -1792442963;
assign addr[20359] = -1781840195;
assign addr[20360] = -1771096139;
assign addr[20361] = -1760211645;
assign addr[20362] = -1749187577;
assign addr[20363] = -1738024810;
assign addr[20364] = -1726724227;
assign addr[20365] = -1715286726;
assign addr[20366] = -1703713213;
assign addr[20367] = -1692004606;
assign addr[20368] = -1680161834;
assign addr[20369] = -1668185835;
assign addr[20370] = -1656077559;
assign addr[20371] = -1643837966;
assign addr[20372] = -1631468027;
assign addr[20373] = -1618968722;
assign addr[20374] = -1606341043;
assign addr[20375] = -1593585992;
assign addr[20376] = -1580704578;
assign addr[20377] = -1567697824;
assign addr[20378] = -1554566762;
assign addr[20379] = -1541312431;
assign addr[20380] = -1527935884;
assign addr[20381] = -1514438181;
assign addr[20382] = -1500820393;
assign addr[20383] = -1487083598;
assign addr[20384] = -1473228887;
assign addr[20385] = -1459257358;
assign addr[20386] = -1445170118;
assign addr[20387] = -1430968286;
assign addr[20388] = -1416652986;
assign addr[20389] = -1402225355;
assign addr[20390] = -1387686535;
assign addr[20391] = -1373037681;
assign addr[20392] = -1358279953;
assign addr[20393] = -1343414522;
assign addr[20394] = -1328442566;
assign addr[20395] = -1313365273;
assign addr[20396] = -1298183838;
assign addr[20397] = -1282899464;
assign addr[20398] = -1267513365;
assign addr[20399] = -1252026760;
assign addr[20400] = -1236440877;
assign addr[20401] = -1220756951;
assign addr[20402] = -1204976227;
assign addr[20403] = -1189099956;
assign addr[20404] = -1173129396;
assign addr[20405] = -1157065814;
assign addr[20406] = -1140910484;
assign addr[20407] = -1124664687;
assign addr[20408] = -1108329711;
assign addr[20409] = -1091906851;
assign addr[20410] = -1075397409;
assign addr[20411] = -1058802695;
assign addr[20412] = -1042124025;
assign addr[20413] = -1025362720;
assign addr[20414] = -1008520110;
assign addr[20415] = -991597531;
assign addr[20416] = -974596324;
assign addr[20417] = -957517838;
assign addr[20418] = -940363427;
assign addr[20419] = -923134450;
assign addr[20420] = -905832274;
assign addr[20421] = -888458272;
assign addr[20422] = -871013820;
assign addr[20423] = -853500302;
assign addr[20424] = -835919107;
assign addr[20425] = -818271628;
assign addr[20426] = -800559266;
assign addr[20427] = -782783424;
assign addr[20428] = -764945512;
assign addr[20429] = -747046944;
assign addr[20430] = -729089140;
assign addr[20431] = -711073524;
assign addr[20432] = -693001525;
assign addr[20433] = -674874574;
assign addr[20434] = -656694110;
assign addr[20435] = -638461574;
assign addr[20436] = -620178412;
assign addr[20437] = -601846074;
assign addr[20438] = -583466013;
assign addr[20439] = -565039687;
assign addr[20440] = -546568556;
assign addr[20441] = -528054086;
assign addr[20442] = -509497745;
assign addr[20443] = -490901003;
assign addr[20444] = -472265336;
assign addr[20445] = -453592221;
assign addr[20446] = -434883140;
assign addr[20447] = -416139574;
assign addr[20448] = -397363011;
assign addr[20449] = -378554940;
assign addr[20450] = -359716852;
assign addr[20451] = -340850240;
assign addr[20452] = -321956601;
assign addr[20453] = -303037433;
assign addr[20454] = -284094236;
assign addr[20455] = -265128512;
assign addr[20456] = -246141764;
assign addr[20457] = -227135500;
assign addr[20458] = -208111224;
assign addr[20459] = -189070447;
assign addr[20460] = -170014678;
assign addr[20461] = -150945428;
assign addr[20462] = -131864208;
assign addr[20463] = -112772533;
assign addr[20464] = -93671915;
assign addr[20465] = -74563870;
assign addr[20466] = -55449912;
assign addr[20467] = -36331557;
assign addr[20468] = -17210322;
assign addr[20469] = 1912278;
assign addr[20470] = 21034727;
assign addr[20471] = 40155507;
assign addr[20472] = 59273104;
assign addr[20473] = 78386000;
assign addr[20474] = 97492681;
assign addr[20475] = 116591632;
assign addr[20476] = 135681337;
assign addr[20477] = 154760284;
assign addr[20478] = 173826959;
assign addr[20479] = 192879850;
assign addr[20480] = 211917448;
assign addr[20481] = 230938242;
assign addr[20482] = 249940723;
assign addr[20483] = 268923386;
assign addr[20484] = 287884725;
assign addr[20485] = 306823237;
assign addr[20486] = 325737419;
assign addr[20487] = 344625773;
assign addr[20488] = 363486799;
assign addr[20489] = 382319004;
assign addr[20490] = 401120892;
assign addr[20491] = 419890975;
assign addr[20492] = 438627762;
assign addr[20493] = 457329769;
assign addr[20494] = 475995513;
assign addr[20495] = 494623513;
assign addr[20496] = 513212292;
assign addr[20497] = 531760377;
assign addr[20498] = 550266296;
assign addr[20499] = 568728583;
assign addr[20500] = 587145773;
assign addr[20501] = 605516406;
assign addr[20502] = 623839025;
assign addr[20503] = 642112178;
assign addr[20504] = 660334415;
assign addr[20505] = 678504291;
assign addr[20506] = 696620367;
assign addr[20507] = 714681204;
assign addr[20508] = 732685372;
assign addr[20509] = 750631442;
assign addr[20510] = 768517992;
assign addr[20511] = 786343603;
assign addr[20512] = 804106861;
assign addr[20513] = 821806359;
assign addr[20514] = 839440693;
assign addr[20515] = 857008464;
assign addr[20516] = 874508280;
assign addr[20517] = 891938752;
assign addr[20518] = 909298500;
assign addr[20519] = 926586145;
assign addr[20520] = 943800318;
assign addr[20521] = 960939653;
assign addr[20522] = 978002791;
assign addr[20523] = 994988380;
assign addr[20524] = 1011895073;
assign addr[20525] = 1028721528;
assign addr[20526] = 1045466412;
assign addr[20527] = 1062128397;
assign addr[20528] = 1078706161;
assign addr[20529] = 1095198391;
assign addr[20530] = 1111603778;
assign addr[20531] = 1127921022;
assign addr[20532] = 1144148829;
assign addr[20533] = 1160285911;
assign addr[20534] = 1176330990;
assign addr[20535] = 1192282793;
assign addr[20536] = 1208140056;
assign addr[20537] = 1223901520;
assign addr[20538] = 1239565936;
assign addr[20539] = 1255132063;
assign addr[20540] = 1270598665;
assign addr[20541] = 1285964516;
assign addr[20542] = 1301228398;
assign addr[20543] = 1316389101;
assign addr[20544] = 1331445422;
assign addr[20545] = 1346396168;
assign addr[20546] = 1361240152;
assign addr[20547] = 1375976199;
assign addr[20548] = 1390603139;
assign addr[20549] = 1405119813;
assign addr[20550] = 1419525069;
assign addr[20551] = 1433817766;
assign addr[20552] = 1447996770;
assign addr[20553] = 1462060956;
assign addr[20554] = 1476009210;
assign addr[20555] = 1489840425;
assign addr[20556] = 1503553506;
assign addr[20557] = 1517147363;
assign addr[20558] = 1530620920;
assign addr[20559] = 1543973108;
assign addr[20560] = 1557202869;
assign addr[20561] = 1570309153;
assign addr[20562] = 1583290921;
assign addr[20563] = 1596147143;
assign addr[20564] = 1608876801;
assign addr[20565] = 1621478885;
assign addr[20566] = 1633952396;
assign addr[20567] = 1646296344;
assign addr[20568] = 1658509750;
assign addr[20569] = 1670591647;
assign addr[20570] = 1682541077;
assign addr[20571] = 1694357091;
assign addr[20572] = 1706038753;
assign addr[20573] = 1717585136;
assign addr[20574] = 1728995326;
assign addr[20575] = 1740268417;
assign addr[20576] = 1751403515;
assign addr[20577] = 1762399737;
assign addr[20578] = 1773256212;
assign addr[20579] = 1783972079;
assign addr[20580] = 1794546487;
assign addr[20581] = 1804978599;
assign addr[20582] = 1815267588;
assign addr[20583] = 1825412636;
assign addr[20584] = 1835412941;
assign addr[20585] = 1845267708;
assign addr[20586] = 1854976157;
assign addr[20587] = 1864537518;
assign addr[20588] = 1873951032;
assign addr[20589] = 1883215953;
assign addr[20590] = 1892331547;
assign addr[20591] = 1901297091;
assign addr[20592] = 1910111873;
assign addr[20593] = 1918775195;
assign addr[20594] = 1927286370;
assign addr[20595] = 1935644723;
assign addr[20596] = 1943849591;
assign addr[20597] = 1951900324;
assign addr[20598] = 1959796283;
assign addr[20599] = 1967536842;
assign addr[20600] = 1975121388;
assign addr[20601] = 1982549318;
assign addr[20602] = 1989820044;
assign addr[20603] = 1996932990;
assign addr[20604] = 2003887591;
assign addr[20605] = 2010683297;
assign addr[20606] = 2017319567;
assign addr[20607] = 2023795876;
assign addr[20608] = 2030111710;
assign addr[20609] = 2036266570;
assign addr[20610] = 2042259965;
assign addr[20611] = 2048091422;
assign addr[20612] = 2053760478;
assign addr[20613] = 2059266683;
assign addr[20614] = 2064609600;
assign addr[20615] = 2069788807;
assign addr[20616] = 2074803892;
assign addr[20617] = 2079654458;
assign addr[20618] = 2084340120;
assign addr[20619] = 2088860507;
assign addr[20620] = 2093215260;
assign addr[20621] = 2097404033;
assign addr[20622] = 2101426496;
assign addr[20623] = 2105282327;
assign addr[20624] = 2108971223;
assign addr[20625] = 2112492891;
assign addr[20626] = 2115847050;
assign addr[20627] = 2119033436;
assign addr[20628] = 2122051796;
assign addr[20629] = 2124901890;
assign addr[20630] = 2127583492;
assign addr[20631] = 2130096389;
assign addr[20632] = 2132440383;
assign addr[20633] = 2134615288;
assign addr[20634] = 2136620930;
assign addr[20635] = 2138457152;
assign addr[20636] = 2140123807;
assign addr[20637] = 2141620763;
assign addr[20638] = 2142947902;
assign addr[20639] = 2144105118;
assign addr[20640] = 2145092320;
assign addr[20641] = 2145909429;
assign addr[20642] = 2146556380;
assign addr[20643] = 2147033123;
assign addr[20644] = 2147339619;
assign addr[20645] = 2147475844;
assign addr[20646] = 2147441787;
assign addr[20647] = 2147237452;
assign addr[20648] = 2146862854;
assign addr[20649] = 2146318022;
assign addr[20650] = 2145603001;
assign addr[20651] = 2144717846;
assign addr[20652] = 2143662628;
assign addr[20653] = 2142437431;
assign addr[20654] = 2141042352;
assign addr[20655] = 2139477502;
assign addr[20656] = 2137743003;
assign addr[20657] = 2135838995;
assign addr[20658] = 2133765628;
assign addr[20659] = 2131523066;
assign addr[20660] = 2129111488;
assign addr[20661] = 2126531084;
assign addr[20662] = 2123782059;
assign addr[20663] = 2120864631;
assign addr[20664] = 2117779031;
assign addr[20665] = 2114525505;
assign addr[20666] = 2111104309;
assign addr[20667] = 2107515716;
assign addr[20668] = 2103760010;
assign addr[20669] = 2099837489;
assign addr[20670] = 2095748463;
assign addr[20671] = 2091493257;
assign addr[20672] = 2087072209;
assign addr[20673] = 2082485668;
assign addr[20674] = 2077733999;
assign addr[20675] = 2072817579;
assign addr[20676] = 2067736796;
assign addr[20677] = 2062492055;
assign addr[20678] = 2057083771;
assign addr[20679] = 2051512372;
assign addr[20680] = 2045778302;
assign addr[20681] = 2039882013;
assign addr[20682] = 2033823974;
assign addr[20683] = 2027604666;
assign addr[20684] = 2021224581;
assign addr[20685] = 2014684225;
assign addr[20686] = 2007984117;
assign addr[20687] = 2001124788;
assign addr[20688] = 1994106782;
assign addr[20689] = 1986930656;
assign addr[20690] = 1979596978;
assign addr[20691] = 1972106330;
assign addr[20692] = 1964459306;
assign addr[20693] = 1956656513;
assign addr[20694] = 1948698568;
assign addr[20695] = 1940586104;
assign addr[20696] = 1932319763;
assign addr[20697] = 1923900201;
assign addr[20698] = 1915328086;
assign addr[20699] = 1906604097;
assign addr[20700] = 1897728925;
assign addr[20701] = 1888703276;
assign addr[20702] = 1879527863;
assign addr[20703] = 1870203416;
assign addr[20704] = 1860730673;
assign addr[20705] = 1851110385;
assign addr[20706] = 1841343316;
assign addr[20707] = 1831430239;
assign addr[20708] = 1821371941;
assign addr[20709] = 1811169220;
assign addr[20710] = 1800822883;
assign addr[20711] = 1790333753;
assign addr[20712] = 1779702660;
assign addr[20713] = 1768930447;
assign addr[20714] = 1758017969;
assign addr[20715] = 1746966091;
assign addr[20716] = 1735775690;
assign addr[20717] = 1724447652;
assign addr[20718] = 1712982875;
assign addr[20719] = 1701382270;
assign addr[20720] = 1689646755;
assign addr[20721] = 1677777262;
assign addr[20722] = 1665774731;
assign addr[20723] = 1653640115;
assign addr[20724] = 1641374375;
assign addr[20725] = 1628978484;
assign addr[20726] = 1616453425;
assign addr[20727] = 1603800191;
assign addr[20728] = 1591019785;
assign addr[20729] = 1578113222;
assign addr[20730] = 1565081523;
assign addr[20731] = 1551925723;
assign addr[20732] = 1538646865;
assign addr[20733] = 1525246002;
assign addr[20734] = 1511724196;
assign addr[20735] = 1498082520;
assign addr[20736] = 1484322054;
assign addr[20737] = 1470443891;
assign addr[20738] = 1456449131;
assign addr[20739] = 1442338884;
assign addr[20740] = 1428114267;
assign addr[20741] = 1413776410;
assign addr[20742] = 1399326449;
assign addr[20743] = 1384765530;
assign addr[20744] = 1370094808;
assign addr[20745] = 1355315445;
assign addr[20746] = 1340428615;
assign addr[20747] = 1325435496;
assign addr[20748] = 1310337279;
assign addr[20749] = 1295135159;
assign addr[20750] = 1279830344;
assign addr[20751] = 1264424045;
assign addr[20752] = 1248917486;
assign addr[20753] = 1233311895;
assign addr[20754] = 1217608510;
assign addr[20755] = 1201808576;
assign addr[20756] = 1185913346;
assign addr[20757] = 1169924081;
assign addr[20758] = 1153842047;
assign addr[20759] = 1137668521;
assign addr[20760] = 1121404785;
assign addr[20761] = 1105052128;
assign addr[20762] = 1088611847;
assign addr[20763] = 1072085246;
assign addr[20764] = 1055473635;
assign addr[20765] = 1038778332;
assign addr[20766] = 1022000660;
assign addr[20767] = 1005141949;
assign addr[20768] = 988203537;
assign addr[20769] = 971186766;
assign addr[20770] = 954092986;
assign addr[20771] = 936923553;
assign addr[20772] = 919679827;
assign addr[20773] = 902363176;
assign addr[20774] = 884974973;
assign addr[20775] = 867516597;
assign addr[20776] = 849989433;
assign addr[20777] = 832394869;
assign addr[20778] = 814734301;
assign addr[20779] = 797009130;
assign addr[20780] = 779220762;
assign addr[20781] = 761370605;
assign addr[20782] = 743460077;
assign addr[20783] = 725490597;
assign addr[20784] = 707463589;
assign addr[20785] = 689380485;
assign addr[20786] = 671242716;
assign addr[20787] = 653051723;
assign addr[20788] = 634808946;
assign addr[20789] = 616515832;
assign addr[20790] = 598173833;
assign addr[20791] = 579784402;
assign addr[20792] = 561348998;
assign addr[20793] = 542869083;
assign addr[20794] = 524346121;
assign addr[20795] = 505781581;
assign addr[20796] = 487176937;
assign addr[20797] = 468533662;
assign addr[20798] = 449853235;
assign addr[20799] = 431137138;
assign addr[20800] = 412386854;
assign addr[20801] = 393603870;
assign addr[20802] = 374789676;
assign addr[20803] = 355945764;
assign addr[20804] = 337073627;
assign addr[20805] = 318174762;
assign addr[20806] = 299250668;
assign addr[20807] = 280302845;
assign addr[20808] = 261332796;
assign addr[20809] = 242342025;
assign addr[20810] = 223332037;
assign addr[20811] = 204304341;
assign addr[20812] = 185260444;
assign addr[20813] = 166201858;
assign addr[20814] = 147130093;
assign addr[20815] = 128046661;
assign addr[20816] = 108953076;
assign addr[20817] = 89850852;
assign addr[20818] = 70741503;
assign addr[20819] = 51626544;
assign addr[20820] = 32507492;
assign addr[20821] = 13385863;
assign addr[20822] = -5736829;
assign addr[20823] = -24859065;
assign addr[20824] = -43979330;
assign addr[20825] = -63096108;
assign addr[20826] = -82207882;
assign addr[20827] = -101313138;
assign addr[20828] = -120410361;
assign addr[20829] = -139498035;
assign addr[20830] = -158574649;
assign addr[20831] = -177638688;
assign addr[20832] = -196688642;
assign addr[20833] = -215722999;
assign addr[20834] = -234740251;
assign addr[20835] = -253738890;
assign addr[20836] = -272717408;
assign addr[20837] = -291674302;
assign addr[20838] = -310608068;
assign addr[20839] = -329517204;
assign addr[20840] = -348400212;
assign addr[20841] = -367255594;
assign addr[20842] = -386081854;
assign addr[20843] = -404877501;
assign addr[20844] = -423641043;
assign addr[20845] = -442370993;
assign addr[20846] = -461065866;
assign addr[20847] = -479724180;
assign addr[20848] = -498344454;
assign addr[20849] = -516925212;
assign addr[20850] = -535464981;
assign addr[20851] = -553962291;
assign addr[20852] = -572415676;
assign addr[20853] = -590823671;
assign addr[20854] = -609184818;
assign addr[20855] = -627497660;
assign addr[20856] = -645760745;
assign addr[20857] = -663972625;
assign addr[20858] = -682131857;
assign addr[20859] = -700236999;
assign addr[20860] = -718286617;
assign addr[20861] = -736279279;
assign addr[20862] = -754213559;
assign addr[20863] = -772088034;
assign addr[20864] = -789901288;
assign addr[20865] = -807651907;
assign addr[20866] = -825338484;
assign addr[20867] = -842959617;
assign addr[20868] = -860513908;
assign addr[20869] = -877999966;
assign addr[20870] = -895416404;
assign addr[20871] = -912761841;
assign addr[20872] = -930034901;
assign addr[20873] = -947234215;
assign addr[20874] = -964358420;
assign addr[20875] = -981406156;
assign addr[20876] = -998376073;
assign addr[20877] = -1015266825;
assign addr[20878] = -1032077073;
assign addr[20879] = -1048805483;
assign addr[20880] = -1065450729;
assign addr[20881] = -1082011492;
assign addr[20882] = -1098486458;
assign addr[20883] = -1114874320;
assign addr[20884] = -1131173780;
assign addr[20885] = -1147383544;
assign addr[20886] = -1163502328;
assign addr[20887] = -1179528853;
assign addr[20888] = -1195461849;
assign addr[20889] = -1211300053;
assign addr[20890] = -1227042207;
assign addr[20891] = -1242687064;
assign addr[20892] = -1258233384;
assign addr[20893] = -1273679934;
assign addr[20894] = -1289025489;
assign addr[20895] = -1304268832;
assign addr[20896] = -1319408754;
assign addr[20897] = -1334444055;
assign addr[20898] = -1349373543;
assign addr[20899] = -1364196034;
assign addr[20900] = -1378910353;
assign addr[20901] = -1393515332;
assign addr[20902] = -1408009814;
assign addr[20903] = -1422392650;
assign addr[20904] = -1436662698;
assign addr[20905] = -1450818828;
assign addr[20906] = -1464859917;
assign addr[20907] = -1478784851;
assign addr[20908] = -1492592527;
assign addr[20909] = -1506281850;
assign addr[20910] = -1519851733;
assign addr[20911] = -1533301101;
assign addr[20912] = -1546628888;
assign addr[20913] = -1559834037;
assign addr[20914] = -1572915501;
assign addr[20915] = -1585872242;
assign addr[20916] = -1598703233;
assign addr[20917] = -1611407456;
assign addr[20918] = -1623983905;
assign addr[20919] = -1636431582;
assign addr[20920] = -1648749499;
assign addr[20921] = -1660936681;
assign addr[20922] = -1672992161;
assign addr[20923] = -1684914983;
assign addr[20924] = -1696704201;
assign addr[20925] = -1708358881;
assign addr[20926] = -1719878099;
assign addr[20927] = -1731260941;
assign addr[20928] = -1742506504;
assign addr[20929] = -1753613897;
assign addr[20930] = -1764582240;
assign addr[20931] = -1775410662;
assign addr[20932] = -1786098304;
assign addr[20933] = -1796644320;
assign addr[20934] = -1807047873;
assign addr[20935] = -1817308138;
assign addr[20936] = -1827424302;
assign addr[20937] = -1837395562;
assign addr[20938] = -1847221128;
assign addr[20939] = -1856900221;
assign addr[20940] = -1866432072;
assign addr[20941] = -1875815927;
assign addr[20942] = -1885051042;
assign addr[20943] = -1894136683;
assign addr[20944] = -1903072131;
assign addr[20945] = -1911856677;
assign addr[20946] = -1920489624;
assign addr[20947] = -1928970288;
assign addr[20948] = -1937297997;
assign addr[20949] = -1945472089;
assign addr[20950] = -1953491918;
assign addr[20951] = -1961356847;
assign addr[20952] = -1969066252;
assign addr[20953] = -1976619522;
assign addr[20954] = -1984016058;
assign addr[20955] = -1991255274;
assign addr[20956] = -1998336596;
assign addr[20957] = -2005259462;
assign addr[20958] = -2012023322;
assign addr[20959] = -2018627642;
assign addr[20960] = -2025071897;
assign addr[20961] = -2031355576;
assign addr[20962] = -2037478181;
assign addr[20963] = -2043439226;
assign addr[20964] = -2049238240;
assign addr[20965] = -2054874761;
assign addr[20966] = -2060348343;
assign addr[20967] = -2065658552;
assign addr[20968] = -2070804967;
assign addr[20969] = -2075787180;
assign addr[20970] = -2080604795;
assign addr[20971] = -2085257431;
assign addr[20972] = -2089744719;
assign addr[20973] = -2094066304;
assign addr[20974] = -2098221841;
assign addr[20975] = -2102211002;
assign addr[20976] = -2106033471;
assign addr[20977] = -2109688944;
assign addr[20978] = -2113177132;
assign addr[20979] = -2116497758;
assign addr[20980] = -2119650558;
assign addr[20981] = -2122635283;
assign addr[20982] = -2125451696;
assign addr[20983] = -2128099574;
assign addr[20984] = -2130578706;
assign addr[20985] = -2132888897;
assign addr[20986] = -2135029962;
assign addr[20987] = -2137001733;
assign addr[20988] = -2138804053;
assign addr[20989] = -2140436778;
assign addr[20990] = -2141899780;
assign addr[20991] = -2143192942;
assign addr[20992] = -2144316162;
assign addr[20993] = -2145269351;
assign addr[20994] = -2146052433;
assign addr[20995] = -2146665347;
assign addr[20996] = -2147108043;
assign addr[20997] = -2147380486;
assign addr[20998] = -2147482655;
assign addr[20999] = -2147414542;
assign addr[21000] = -2147176152;
assign addr[21001] = -2146767505;
assign addr[21002] = -2146188631;
assign addr[21003] = -2145439578;
assign addr[21004] = -2144520405;
assign addr[21005] = -2143431184;
assign addr[21006] = -2142172003;
assign addr[21007] = -2140742960;
assign addr[21008] = -2139144169;
assign addr[21009] = -2137375758;
assign addr[21010] = -2135437865;
assign addr[21011] = -2133330646;
assign addr[21012] = -2131054266;
assign addr[21013] = -2128608907;
assign addr[21014] = -2125994762;
assign addr[21015] = -2123212038;
assign addr[21016] = -2120260957;
assign addr[21017] = -2117141752;
assign addr[21018] = -2113854671;
assign addr[21019] = -2110399974;
assign addr[21020] = -2106777935;
assign addr[21021] = -2102988841;
assign addr[21022] = -2099032994;
assign addr[21023] = -2094910706;
assign addr[21024] = -2090622304;
assign addr[21025] = -2086168128;
assign addr[21026] = -2081548533;
assign addr[21027] = -2076763883;
assign addr[21028] = -2071814558;
assign addr[21029] = -2066700952;
assign addr[21030] = -2061423468;
assign addr[21031] = -2055982526;
assign addr[21032] = -2050378558;
assign addr[21033] = -2044612007;
assign addr[21034] = -2038683330;
assign addr[21035] = -2032592999;
assign addr[21036] = -2026341495;
assign addr[21037] = -2019929315;
assign addr[21038] = -2013356967;
assign addr[21039] = -2006624971;
assign addr[21040] = -1999733863;
assign addr[21041] = -1992684188;
assign addr[21042] = -1985476506;
assign addr[21043] = -1978111387;
assign addr[21044] = -1970589416;
assign addr[21045] = -1962911189;
assign addr[21046] = -1955077316;
assign addr[21047] = -1947088417;
assign addr[21048] = -1938945125;
assign addr[21049] = -1930648088;
assign addr[21050] = -1922197961;
assign addr[21051] = -1913595416;
assign addr[21052] = -1904841135;
assign addr[21053] = -1895935811;
assign addr[21054] = -1886880151;
assign addr[21055] = -1877674873;
assign addr[21056] = -1868320707;
assign addr[21057] = -1858818395;
assign addr[21058] = -1849168689;
assign addr[21059] = -1839372356;
assign addr[21060] = -1829430172;
assign addr[21061] = -1819342925;
assign addr[21062] = -1809111415;
assign addr[21063] = -1798736454;
assign addr[21064] = -1788218865;
assign addr[21065] = -1777559480;
assign addr[21066] = -1766759146;
assign addr[21067] = -1755818718;
assign addr[21068] = -1744739065;
assign addr[21069] = -1733521064;
assign addr[21070] = -1722165606;
assign addr[21071] = -1710673591;
assign addr[21072] = -1699045930;
assign addr[21073] = -1687283545;
assign addr[21074] = -1675387369;
assign addr[21075] = -1663358344;
assign addr[21076] = -1651197426;
assign addr[21077] = -1638905577;
assign addr[21078] = -1626483774;
assign addr[21079] = -1613933000;
assign addr[21080] = -1601254251;
assign addr[21081] = -1588448533;
assign addr[21082] = -1575516860;
assign addr[21083] = -1562460258;
assign addr[21084] = -1549279763;
assign addr[21085] = -1535976419;
assign addr[21086] = -1522551282;
assign addr[21087] = -1509005416;
assign addr[21088] = -1495339895;
assign addr[21089] = -1481555802;
assign addr[21090] = -1467654232;
assign addr[21091] = -1453636285;
assign addr[21092] = -1439503074;
assign addr[21093] = -1425255719;
assign addr[21094] = -1410895350;
assign addr[21095] = -1396423105;
assign addr[21096] = -1381840133;
assign addr[21097] = -1367147589;
assign addr[21098] = -1352346639;
assign addr[21099] = -1337438456;
assign addr[21100] = -1322424222;
assign addr[21101] = -1307305128;
assign addr[21102] = -1292082373;
assign addr[21103] = -1276757164;
assign addr[21104] = -1261330715;
assign addr[21105] = -1245804251;
assign addr[21106] = -1230179002;
assign addr[21107] = -1214456207;
assign addr[21108] = -1198637114;
assign addr[21109] = -1182722976;
assign addr[21110] = -1166715055;
assign addr[21111] = -1150614620;
assign addr[21112] = -1134422949;
assign addr[21113] = -1118141326;
assign addr[21114] = -1101771040;
assign addr[21115] = -1085313391;
assign addr[21116] = -1068769683;
assign addr[21117] = -1052141228;
assign addr[21118] = -1035429345;
assign addr[21119] = -1018635358;
assign addr[21120] = -1001760600;
assign addr[21121] = -984806408;
assign addr[21122] = -967774128;
assign addr[21123] = -950665109;
assign addr[21124] = -933480707;
assign addr[21125] = -916222287;
assign addr[21126] = -898891215;
assign addr[21127] = -881488868;
assign addr[21128] = -864016623;
assign addr[21129] = -846475867;
assign addr[21130] = -828867991;
assign addr[21131] = -811194391;
assign addr[21132] = -793456467;
assign addr[21133] = -775655628;
assign addr[21134] = -757793284;
assign addr[21135] = -739870851;
assign addr[21136] = -721889752;
assign addr[21137] = -703851410;
assign addr[21138] = -685757258;
assign addr[21139] = -667608730;
assign addr[21140] = -649407264;
assign addr[21141] = -631154304;
assign addr[21142] = -612851297;
assign addr[21143] = -594499695;
assign addr[21144] = -576100953;
assign addr[21145] = -557656529;
assign addr[21146] = -539167887;
assign addr[21147] = -520636492;
assign addr[21148] = -502063814;
assign addr[21149] = -483451325;
assign addr[21150] = -464800501;
assign addr[21151] = -446112822;
assign addr[21152] = -427389768;
assign addr[21153] = -408632825;
assign addr[21154] = -389843480;
assign addr[21155] = -371023223;
assign addr[21156] = -352173546;
assign addr[21157] = -333295944;
assign addr[21158] = -314391913;
assign addr[21159] = -295462954;
assign addr[21160] = -276510565;
assign addr[21161] = -257536251;
assign addr[21162] = -238541516;
assign addr[21163] = -219527866;
assign addr[21164] = -200496809;
assign addr[21165] = -181449854;
assign addr[21166] = -162388511;
assign addr[21167] = -143314291;
assign addr[21168] = -124228708;
assign addr[21169] = -105133274;
assign addr[21170] = -86029503;
assign addr[21171] = -66918911;
assign addr[21172] = -47803013;
assign addr[21173] = -28683324;
assign addr[21174] = -9561361;
assign addr[21175] = 9561361;
assign addr[21176] = 28683324;
assign addr[21177] = 47803013;
assign addr[21178] = 66918911;
assign addr[21179] = 86029503;
assign addr[21180] = 105133274;
assign addr[21181] = 124228708;
assign addr[21182] = 143314291;
assign addr[21183] = 162388511;
assign addr[21184] = 181449854;
assign addr[21185] = 200496809;
assign addr[21186] = 219527866;
assign addr[21187] = 238541516;
assign addr[21188] = 257536251;
assign addr[21189] = 276510565;
assign addr[21190] = 295462954;
assign addr[21191] = 314391913;
assign addr[21192] = 333295944;
assign addr[21193] = 352173546;
assign addr[21194] = 371023223;
assign addr[21195] = 389843480;
assign addr[21196] = 408632825;
assign addr[21197] = 427389768;
assign addr[21198] = 446112822;
assign addr[21199] = 464800501;
assign addr[21200] = 483451325;
assign addr[21201] = 502063814;
assign addr[21202] = 520636492;
assign addr[21203] = 539167887;
assign addr[21204] = 557656529;
assign addr[21205] = 576100953;
assign addr[21206] = 594499695;
assign addr[21207] = 612851297;
assign addr[21208] = 631154304;
assign addr[21209] = 649407264;
assign addr[21210] = 667608730;
assign addr[21211] = 685757258;
assign addr[21212] = 703851410;
assign addr[21213] = 721889752;
assign addr[21214] = 739870851;
assign addr[21215] = 757793284;
assign addr[21216] = 775655628;
assign addr[21217] = 793456467;
assign addr[21218] = 811194391;
assign addr[21219] = 828867991;
assign addr[21220] = 846475867;
assign addr[21221] = 864016623;
assign addr[21222] = 881488868;
assign addr[21223] = 898891215;
assign addr[21224] = 916222287;
assign addr[21225] = 933480707;
assign addr[21226] = 950665109;
assign addr[21227] = 967774128;
assign addr[21228] = 984806408;
assign addr[21229] = 1001760600;
assign addr[21230] = 1018635358;
assign addr[21231] = 1035429345;
assign addr[21232] = 1052141228;
assign addr[21233] = 1068769683;
assign addr[21234] = 1085313391;
assign addr[21235] = 1101771040;
assign addr[21236] = 1118141326;
assign addr[21237] = 1134422949;
assign addr[21238] = 1150614620;
assign addr[21239] = 1166715055;
assign addr[21240] = 1182722976;
assign addr[21241] = 1198637114;
assign addr[21242] = 1214456207;
assign addr[21243] = 1230179002;
assign addr[21244] = 1245804251;
assign addr[21245] = 1261330715;
assign addr[21246] = 1276757164;
assign addr[21247] = 1292082373;
assign addr[21248] = 1307305128;
assign addr[21249] = 1322424222;
assign addr[21250] = 1337438456;
assign addr[21251] = 1352346639;
assign addr[21252] = 1367147589;
assign addr[21253] = 1381840133;
assign addr[21254] = 1396423105;
assign addr[21255] = 1410895350;
assign addr[21256] = 1425255719;
assign addr[21257] = 1439503074;
assign addr[21258] = 1453636285;
assign addr[21259] = 1467654232;
assign addr[21260] = 1481555802;
assign addr[21261] = 1495339895;
assign addr[21262] = 1509005416;
assign addr[21263] = 1522551282;
assign addr[21264] = 1535976419;
assign addr[21265] = 1549279763;
assign addr[21266] = 1562460258;
assign addr[21267] = 1575516860;
assign addr[21268] = 1588448533;
assign addr[21269] = 1601254251;
assign addr[21270] = 1613933000;
assign addr[21271] = 1626483774;
assign addr[21272] = 1638905577;
assign addr[21273] = 1651197426;
assign addr[21274] = 1663358344;
assign addr[21275] = 1675387369;
assign addr[21276] = 1687283545;
assign addr[21277] = 1699045930;
assign addr[21278] = 1710673591;
assign addr[21279] = 1722165606;
assign addr[21280] = 1733521064;
assign addr[21281] = 1744739065;
assign addr[21282] = 1755818718;
assign addr[21283] = 1766759146;
assign addr[21284] = 1777559480;
assign addr[21285] = 1788218865;
assign addr[21286] = 1798736454;
assign addr[21287] = 1809111415;
assign addr[21288] = 1819342925;
assign addr[21289] = 1829430172;
assign addr[21290] = 1839372356;
assign addr[21291] = 1849168689;
assign addr[21292] = 1858818395;
assign addr[21293] = 1868320707;
assign addr[21294] = 1877674873;
assign addr[21295] = 1886880151;
assign addr[21296] = 1895935811;
assign addr[21297] = 1904841135;
assign addr[21298] = 1913595416;
assign addr[21299] = 1922197961;
assign addr[21300] = 1930648088;
assign addr[21301] = 1938945125;
assign addr[21302] = 1947088417;
assign addr[21303] = 1955077316;
assign addr[21304] = 1962911189;
assign addr[21305] = 1970589416;
assign addr[21306] = 1978111387;
assign addr[21307] = 1985476506;
assign addr[21308] = 1992684188;
assign addr[21309] = 1999733863;
assign addr[21310] = 2006624971;
assign addr[21311] = 2013356967;
assign addr[21312] = 2019929315;
assign addr[21313] = 2026341495;
assign addr[21314] = 2032592999;
assign addr[21315] = 2038683330;
assign addr[21316] = 2044612007;
assign addr[21317] = 2050378558;
assign addr[21318] = 2055982526;
assign addr[21319] = 2061423468;
assign addr[21320] = 2066700952;
assign addr[21321] = 2071814558;
assign addr[21322] = 2076763883;
assign addr[21323] = 2081548533;
assign addr[21324] = 2086168128;
assign addr[21325] = 2090622304;
assign addr[21326] = 2094910706;
assign addr[21327] = 2099032994;
assign addr[21328] = 2102988841;
assign addr[21329] = 2106777935;
assign addr[21330] = 2110399974;
assign addr[21331] = 2113854671;
assign addr[21332] = 2117141752;
assign addr[21333] = 2120260957;
assign addr[21334] = 2123212038;
assign addr[21335] = 2125994762;
assign addr[21336] = 2128608907;
assign addr[21337] = 2131054266;
assign addr[21338] = 2133330646;
assign addr[21339] = 2135437865;
assign addr[21340] = 2137375758;
assign addr[21341] = 2139144169;
assign addr[21342] = 2140742960;
assign addr[21343] = 2142172003;
assign addr[21344] = 2143431184;
assign addr[21345] = 2144520405;
assign addr[21346] = 2145439578;
assign addr[21347] = 2146188631;
assign addr[21348] = 2146767505;
assign addr[21349] = 2147176152;
assign addr[21350] = 2147414542;
assign addr[21351] = 2147482655;
assign addr[21352] = 2147380486;
assign addr[21353] = 2147108043;
assign addr[21354] = 2146665347;
assign addr[21355] = 2146052433;
assign addr[21356] = 2145269351;
assign addr[21357] = 2144316162;
assign addr[21358] = 2143192942;
assign addr[21359] = 2141899780;
assign addr[21360] = 2140436778;
assign addr[21361] = 2138804053;
assign addr[21362] = 2137001733;
assign addr[21363] = 2135029962;
assign addr[21364] = 2132888897;
assign addr[21365] = 2130578706;
assign addr[21366] = 2128099574;
assign addr[21367] = 2125451696;
assign addr[21368] = 2122635283;
assign addr[21369] = 2119650558;
assign addr[21370] = 2116497758;
assign addr[21371] = 2113177132;
assign addr[21372] = 2109688944;
assign addr[21373] = 2106033471;
assign addr[21374] = 2102211002;
assign addr[21375] = 2098221841;
assign addr[21376] = 2094066304;
assign addr[21377] = 2089744719;
assign addr[21378] = 2085257431;
assign addr[21379] = 2080604795;
assign addr[21380] = 2075787180;
assign addr[21381] = 2070804967;
assign addr[21382] = 2065658552;
assign addr[21383] = 2060348343;
assign addr[21384] = 2054874761;
assign addr[21385] = 2049238240;
assign addr[21386] = 2043439226;
assign addr[21387] = 2037478181;
assign addr[21388] = 2031355576;
assign addr[21389] = 2025071897;
assign addr[21390] = 2018627642;
assign addr[21391] = 2012023322;
assign addr[21392] = 2005259462;
assign addr[21393] = 1998336596;
assign addr[21394] = 1991255274;
assign addr[21395] = 1984016058;
assign addr[21396] = 1976619522;
assign addr[21397] = 1969066252;
assign addr[21398] = 1961356847;
assign addr[21399] = 1953491918;
assign addr[21400] = 1945472089;
assign addr[21401] = 1937297997;
assign addr[21402] = 1928970288;
assign addr[21403] = 1920489624;
assign addr[21404] = 1911856677;
assign addr[21405] = 1903072131;
assign addr[21406] = 1894136683;
assign addr[21407] = 1885051042;
assign addr[21408] = 1875815927;
assign addr[21409] = 1866432072;
assign addr[21410] = 1856900221;
assign addr[21411] = 1847221128;
assign addr[21412] = 1837395562;
assign addr[21413] = 1827424302;
assign addr[21414] = 1817308138;
assign addr[21415] = 1807047873;
assign addr[21416] = 1796644320;
assign addr[21417] = 1786098304;
assign addr[21418] = 1775410662;
assign addr[21419] = 1764582240;
assign addr[21420] = 1753613897;
assign addr[21421] = 1742506504;
assign addr[21422] = 1731260941;
assign addr[21423] = 1719878099;
assign addr[21424] = 1708358881;
assign addr[21425] = 1696704201;
assign addr[21426] = 1684914983;
assign addr[21427] = 1672992161;
assign addr[21428] = 1660936681;
assign addr[21429] = 1648749499;
assign addr[21430] = 1636431582;
assign addr[21431] = 1623983905;
assign addr[21432] = 1611407456;
assign addr[21433] = 1598703233;
assign addr[21434] = 1585872242;
assign addr[21435] = 1572915501;
assign addr[21436] = 1559834037;
assign addr[21437] = 1546628888;
assign addr[21438] = 1533301101;
assign addr[21439] = 1519851733;
assign addr[21440] = 1506281850;
assign addr[21441] = 1492592527;
assign addr[21442] = 1478784851;
assign addr[21443] = 1464859917;
assign addr[21444] = 1450818828;
assign addr[21445] = 1436662698;
assign addr[21446] = 1422392650;
assign addr[21447] = 1408009814;
assign addr[21448] = 1393515332;
assign addr[21449] = 1378910353;
assign addr[21450] = 1364196034;
assign addr[21451] = 1349373543;
assign addr[21452] = 1334444055;
assign addr[21453] = 1319408754;
assign addr[21454] = 1304268832;
assign addr[21455] = 1289025489;
assign addr[21456] = 1273679934;
assign addr[21457] = 1258233384;
assign addr[21458] = 1242687064;
assign addr[21459] = 1227042207;
assign addr[21460] = 1211300053;
assign addr[21461] = 1195461849;
assign addr[21462] = 1179528853;
assign addr[21463] = 1163502328;
assign addr[21464] = 1147383544;
assign addr[21465] = 1131173780;
assign addr[21466] = 1114874320;
assign addr[21467] = 1098486458;
assign addr[21468] = 1082011492;
assign addr[21469] = 1065450729;
assign addr[21470] = 1048805483;
assign addr[21471] = 1032077073;
assign addr[21472] = 1015266825;
assign addr[21473] = 998376073;
assign addr[21474] = 981406156;
assign addr[21475] = 964358420;
assign addr[21476] = 947234215;
assign addr[21477] = 930034901;
assign addr[21478] = 912761841;
assign addr[21479] = 895416404;
assign addr[21480] = 877999966;
assign addr[21481] = 860513908;
assign addr[21482] = 842959617;
assign addr[21483] = 825338484;
assign addr[21484] = 807651907;
assign addr[21485] = 789901288;
assign addr[21486] = 772088034;
assign addr[21487] = 754213559;
assign addr[21488] = 736279279;
assign addr[21489] = 718286617;
assign addr[21490] = 700236999;
assign addr[21491] = 682131857;
assign addr[21492] = 663972625;
assign addr[21493] = 645760745;
assign addr[21494] = 627497660;
assign addr[21495] = 609184818;
assign addr[21496] = 590823671;
assign addr[21497] = 572415676;
assign addr[21498] = 553962291;
assign addr[21499] = 535464981;
assign addr[21500] = 516925212;
assign addr[21501] = 498344454;
assign addr[21502] = 479724180;
assign addr[21503] = 461065866;
assign addr[21504] = 442370993;
assign addr[21505] = 423641043;
assign addr[21506] = 404877501;
assign addr[21507] = 386081854;
assign addr[21508] = 367255594;
assign addr[21509] = 348400212;
assign addr[21510] = 329517204;
assign addr[21511] = 310608068;
assign addr[21512] = 291674302;
assign addr[21513] = 272717408;
assign addr[21514] = 253738890;
assign addr[21515] = 234740251;
assign addr[21516] = 215722999;
assign addr[21517] = 196688642;
assign addr[21518] = 177638688;
assign addr[21519] = 158574649;
assign addr[21520] = 139498035;
assign addr[21521] = 120410361;
assign addr[21522] = 101313138;
assign addr[21523] = 82207882;
assign addr[21524] = 63096108;
assign addr[21525] = 43979330;
assign addr[21526] = 24859065;
assign addr[21527] = 5736829;
assign addr[21528] = -13385863;
assign addr[21529] = -32507492;
assign addr[21530] = -51626544;
assign addr[21531] = -70741503;
assign addr[21532] = -89850852;
assign addr[21533] = -108953076;
assign addr[21534] = -128046661;
assign addr[21535] = -147130093;
assign addr[21536] = -166201858;
assign addr[21537] = -185260444;
assign addr[21538] = -204304341;
assign addr[21539] = -223332037;
assign addr[21540] = -242342025;
assign addr[21541] = -261332796;
assign addr[21542] = -280302845;
assign addr[21543] = -299250668;
assign addr[21544] = -318174762;
assign addr[21545] = -337073627;
assign addr[21546] = -355945764;
assign addr[21547] = -374789676;
assign addr[21548] = -393603870;
assign addr[21549] = -412386854;
assign addr[21550] = -431137138;
assign addr[21551] = -449853235;
assign addr[21552] = -468533662;
assign addr[21553] = -487176937;
assign addr[21554] = -505781581;
assign addr[21555] = -524346121;
assign addr[21556] = -542869083;
assign addr[21557] = -561348998;
assign addr[21558] = -579784402;
assign addr[21559] = -598173833;
assign addr[21560] = -616515832;
assign addr[21561] = -634808946;
assign addr[21562] = -653051723;
assign addr[21563] = -671242716;
assign addr[21564] = -689380485;
assign addr[21565] = -707463589;
assign addr[21566] = -725490597;
assign addr[21567] = -743460077;
assign addr[21568] = -761370605;
assign addr[21569] = -779220762;
assign addr[21570] = -797009130;
assign addr[21571] = -814734301;
assign addr[21572] = -832394869;
assign addr[21573] = -849989433;
assign addr[21574] = -867516597;
assign addr[21575] = -884974973;
assign addr[21576] = -902363176;
assign addr[21577] = -919679827;
assign addr[21578] = -936923553;
assign addr[21579] = -954092986;
assign addr[21580] = -971186766;
assign addr[21581] = -988203537;
assign addr[21582] = -1005141949;
assign addr[21583] = -1022000660;
assign addr[21584] = -1038778332;
assign addr[21585] = -1055473635;
assign addr[21586] = -1072085246;
assign addr[21587] = -1088611847;
assign addr[21588] = -1105052128;
assign addr[21589] = -1121404785;
assign addr[21590] = -1137668521;
assign addr[21591] = -1153842047;
assign addr[21592] = -1169924081;
assign addr[21593] = -1185913346;
assign addr[21594] = -1201808576;
assign addr[21595] = -1217608510;
assign addr[21596] = -1233311895;
assign addr[21597] = -1248917486;
assign addr[21598] = -1264424045;
assign addr[21599] = -1279830344;
assign addr[21600] = -1295135159;
assign addr[21601] = -1310337279;
assign addr[21602] = -1325435496;
assign addr[21603] = -1340428615;
assign addr[21604] = -1355315445;
assign addr[21605] = -1370094808;
assign addr[21606] = -1384765530;
assign addr[21607] = -1399326449;
assign addr[21608] = -1413776410;
assign addr[21609] = -1428114267;
assign addr[21610] = -1442338884;
assign addr[21611] = -1456449131;
assign addr[21612] = -1470443891;
assign addr[21613] = -1484322054;
assign addr[21614] = -1498082520;
assign addr[21615] = -1511724196;
assign addr[21616] = -1525246002;
assign addr[21617] = -1538646865;
assign addr[21618] = -1551925723;
assign addr[21619] = -1565081523;
assign addr[21620] = -1578113222;
assign addr[21621] = -1591019785;
assign addr[21622] = -1603800191;
assign addr[21623] = -1616453425;
assign addr[21624] = -1628978484;
assign addr[21625] = -1641374375;
assign addr[21626] = -1653640115;
assign addr[21627] = -1665774731;
assign addr[21628] = -1677777262;
assign addr[21629] = -1689646755;
assign addr[21630] = -1701382270;
assign addr[21631] = -1712982875;
assign addr[21632] = -1724447652;
assign addr[21633] = -1735775690;
assign addr[21634] = -1746966091;
assign addr[21635] = -1758017969;
assign addr[21636] = -1768930447;
assign addr[21637] = -1779702660;
assign addr[21638] = -1790333753;
assign addr[21639] = -1800822883;
assign addr[21640] = -1811169220;
assign addr[21641] = -1821371941;
assign addr[21642] = -1831430239;
assign addr[21643] = -1841343316;
assign addr[21644] = -1851110385;
assign addr[21645] = -1860730673;
assign addr[21646] = -1870203416;
assign addr[21647] = -1879527863;
assign addr[21648] = -1888703276;
assign addr[21649] = -1897728925;
assign addr[21650] = -1906604097;
assign addr[21651] = -1915328086;
assign addr[21652] = -1923900201;
assign addr[21653] = -1932319763;
assign addr[21654] = -1940586104;
assign addr[21655] = -1948698568;
assign addr[21656] = -1956656513;
assign addr[21657] = -1964459306;
assign addr[21658] = -1972106330;
assign addr[21659] = -1979596978;
assign addr[21660] = -1986930656;
assign addr[21661] = -1994106782;
assign addr[21662] = -2001124788;
assign addr[21663] = -2007984117;
assign addr[21664] = -2014684225;
assign addr[21665] = -2021224581;
assign addr[21666] = -2027604666;
assign addr[21667] = -2033823974;
assign addr[21668] = -2039882013;
assign addr[21669] = -2045778302;
assign addr[21670] = -2051512372;
assign addr[21671] = -2057083771;
assign addr[21672] = -2062492055;
assign addr[21673] = -2067736796;
assign addr[21674] = -2072817579;
assign addr[21675] = -2077733999;
assign addr[21676] = -2082485668;
assign addr[21677] = -2087072209;
assign addr[21678] = -2091493257;
assign addr[21679] = -2095748463;
assign addr[21680] = -2099837489;
assign addr[21681] = -2103760010;
assign addr[21682] = -2107515716;
assign addr[21683] = -2111104309;
assign addr[21684] = -2114525505;
assign addr[21685] = -2117779031;
assign addr[21686] = -2120864631;
assign addr[21687] = -2123782059;
assign addr[21688] = -2126531084;
assign addr[21689] = -2129111488;
assign addr[21690] = -2131523066;
assign addr[21691] = -2133765628;
assign addr[21692] = -2135838995;
assign addr[21693] = -2137743003;
assign addr[21694] = -2139477502;
assign addr[21695] = -2141042352;
assign addr[21696] = -2142437431;
assign addr[21697] = -2143662628;
assign addr[21698] = -2144717846;
assign addr[21699] = -2145603001;
assign addr[21700] = -2146318022;
assign addr[21701] = -2146862854;
assign addr[21702] = -2147237452;
assign addr[21703] = -2147441787;
assign addr[21704] = -2147475844;
assign addr[21705] = -2147339619;
assign addr[21706] = -2147033123;
assign addr[21707] = -2146556380;
assign addr[21708] = -2145909429;
assign addr[21709] = -2145092320;
assign addr[21710] = -2144105118;
assign addr[21711] = -2142947902;
assign addr[21712] = -2141620763;
assign addr[21713] = -2140123807;
assign addr[21714] = -2138457152;
assign addr[21715] = -2136620930;
assign addr[21716] = -2134615288;
assign addr[21717] = -2132440383;
assign addr[21718] = -2130096389;
assign addr[21719] = -2127583492;
assign addr[21720] = -2124901890;
assign addr[21721] = -2122051796;
assign addr[21722] = -2119033436;
assign addr[21723] = -2115847050;
assign addr[21724] = -2112492891;
assign addr[21725] = -2108971223;
assign addr[21726] = -2105282327;
assign addr[21727] = -2101426496;
assign addr[21728] = -2097404033;
assign addr[21729] = -2093215260;
assign addr[21730] = -2088860507;
assign addr[21731] = -2084340120;
assign addr[21732] = -2079654458;
assign addr[21733] = -2074803892;
assign addr[21734] = -2069788807;
assign addr[21735] = -2064609600;
assign addr[21736] = -2059266683;
assign addr[21737] = -2053760478;
assign addr[21738] = -2048091422;
assign addr[21739] = -2042259965;
assign addr[21740] = -2036266570;
assign addr[21741] = -2030111710;
assign addr[21742] = -2023795876;
assign addr[21743] = -2017319567;
assign addr[21744] = -2010683297;
assign addr[21745] = -2003887591;
assign addr[21746] = -1996932990;
assign addr[21747] = -1989820044;
assign addr[21748] = -1982549318;
assign addr[21749] = -1975121388;
assign addr[21750] = -1967536842;
assign addr[21751] = -1959796283;
assign addr[21752] = -1951900324;
assign addr[21753] = -1943849591;
assign addr[21754] = -1935644723;
assign addr[21755] = -1927286370;
assign addr[21756] = -1918775195;
assign addr[21757] = -1910111873;
assign addr[21758] = -1901297091;
assign addr[21759] = -1892331547;
assign addr[21760] = -1883215953;
assign addr[21761] = -1873951032;
assign addr[21762] = -1864537518;
assign addr[21763] = -1854976157;
assign addr[21764] = -1845267708;
assign addr[21765] = -1835412941;
assign addr[21766] = -1825412636;
assign addr[21767] = -1815267588;
assign addr[21768] = -1804978599;
assign addr[21769] = -1794546487;
assign addr[21770] = -1783972079;
assign addr[21771] = -1773256212;
assign addr[21772] = -1762399737;
assign addr[21773] = -1751403515;
assign addr[21774] = -1740268417;
assign addr[21775] = -1728995326;
assign addr[21776] = -1717585136;
assign addr[21777] = -1706038753;
assign addr[21778] = -1694357091;
assign addr[21779] = -1682541077;
assign addr[21780] = -1670591647;
assign addr[21781] = -1658509750;
assign addr[21782] = -1646296344;
assign addr[21783] = -1633952396;
assign addr[21784] = -1621478885;
assign addr[21785] = -1608876801;
assign addr[21786] = -1596147143;
assign addr[21787] = -1583290921;
assign addr[21788] = -1570309153;
assign addr[21789] = -1557202869;
assign addr[21790] = -1543973108;
assign addr[21791] = -1530620920;
assign addr[21792] = -1517147363;
assign addr[21793] = -1503553506;
assign addr[21794] = -1489840425;
assign addr[21795] = -1476009210;
assign addr[21796] = -1462060956;
assign addr[21797] = -1447996770;
assign addr[21798] = -1433817766;
assign addr[21799] = -1419525069;
assign addr[21800] = -1405119813;
assign addr[21801] = -1390603139;
assign addr[21802] = -1375976199;
assign addr[21803] = -1361240152;
assign addr[21804] = -1346396168;
assign addr[21805] = -1331445422;
assign addr[21806] = -1316389101;
assign addr[21807] = -1301228398;
assign addr[21808] = -1285964516;
assign addr[21809] = -1270598665;
assign addr[21810] = -1255132063;
assign addr[21811] = -1239565936;
assign addr[21812] = -1223901520;
assign addr[21813] = -1208140056;
assign addr[21814] = -1192282793;
assign addr[21815] = -1176330990;
assign addr[21816] = -1160285911;
assign addr[21817] = -1144148829;
assign addr[21818] = -1127921022;
assign addr[21819] = -1111603778;
assign addr[21820] = -1095198391;
assign addr[21821] = -1078706161;
assign addr[21822] = -1062128397;
assign addr[21823] = -1045466412;
assign addr[21824] = -1028721528;
assign addr[21825] = -1011895073;
assign addr[21826] = -994988380;
assign addr[21827] = -978002791;
assign addr[21828] = -960939653;
assign addr[21829] = -943800318;
assign addr[21830] = -926586145;
assign addr[21831] = -909298500;
assign addr[21832] = -891938752;
assign addr[21833] = -874508280;
assign addr[21834] = -857008464;
assign addr[21835] = -839440693;
assign addr[21836] = -821806359;
assign addr[21837] = -804106861;
assign addr[21838] = -786343603;
assign addr[21839] = -768517992;
assign addr[21840] = -750631442;
assign addr[21841] = -732685372;
assign addr[21842] = -714681204;
assign addr[21843] = -696620367;
assign addr[21844] = -678504291;
assign addr[21845] = -660334415;
assign addr[21846] = -642112178;
assign addr[21847] = -623839025;
assign addr[21848] = -605516406;
assign addr[21849] = -587145773;
assign addr[21850] = -568728583;
assign addr[21851] = -550266296;
assign addr[21852] = -531760377;
assign addr[21853] = -513212292;
assign addr[21854] = -494623513;
assign addr[21855] = -475995513;
assign addr[21856] = -457329769;
assign addr[21857] = -438627762;
assign addr[21858] = -419890975;
assign addr[21859] = -401120892;
assign addr[21860] = -382319004;
assign addr[21861] = -363486799;
assign addr[21862] = -344625773;
assign addr[21863] = -325737419;
assign addr[21864] = -306823237;
assign addr[21865] = -287884725;
assign addr[21866] = -268923386;
assign addr[21867] = -249940723;
assign addr[21868] = -230938242;
assign addr[21869] = -211917448;
assign addr[21870] = -192879850;
assign addr[21871] = -173826959;
assign addr[21872] = -154760284;
assign addr[21873] = -135681337;
assign addr[21874] = -116591632;
assign addr[21875] = -97492681;
assign addr[21876] = -78386000;
assign addr[21877] = -59273104;
assign addr[21878] = -40155507;
assign addr[21879] = -21034727;
assign addr[21880] = -1912278;
assign addr[21881] = 17210322;
assign addr[21882] = 36331557;
assign addr[21883] = 55449912;
assign addr[21884] = 74563870;
assign addr[21885] = 93671915;
assign addr[21886] = 112772533;
assign addr[21887] = 131864208;
assign addr[21888] = 150945428;
assign addr[21889] = 170014678;
assign addr[21890] = 189070447;
assign addr[21891] = 208111224;
assign addr[21892] = 227135500;
assign addr[21893] = 246141764;
assign addr[21894] = 265128512;
assign addr[21895] = 284094236;
assign addr[21896] = 303037433;
assign addr[21897] = 321956601;
assign addr[21898] = 340850240;
assign addr[21899] = 359716852;
assign addr[21900] = 378554940;
assign addr[21901] = 397363011;
assign addr[21902] = 416139574;
assign addr[21903] = 434883140;
assign addr[21904] = 453592221;
assign addr[21905] = 472265336;
assign addr[21906] = 490901003;
assign addr[21907] = 509497745;
assign addr[21908] = 528054086;
assign addr[21909] = 546568556;
assign addr[21910] = 565039687;
assign addr[21911] = 583466013;
assign addr[21912] = 601846074;
assign addr[21913] = 620178412;
assign addr[21914] = 638461574;
assign addr[21915] = 656694110;
assign addr[21916] = 674874574;
assign addr[21917] = 693001525;
assign addr[21918] = 711073524;
assign addr[21919] = 729089140;
assign addr[21920] = 747046944;
assign addr[21921] = 764945512;
assign addr[21922] = 782783424;
assign addr[21923] = 800559266;
assign addr[21924] = 818271628;
assign addr[21925] = 835919107;
assign addr[21926] = 853500302;
assign addr[21927] = 871013820;
assign addr[21928] = 888458272;
assign addr[21929] = 905832274;
assign addr[21930] = 923134450;
assign addr[21931] = 940363427;
assign addr[21932] = 957517838;
assign addr[21933] = 974596324;
assign addr[21934] = 991597531;
assign addr[21935] = 1008520110;
assign addr[21936] = 1025362720;
assign addr[21937] = 1042124025;
assign addr[21938] = 1058802695;
assign addr[21939] = 1075397409;
assign addr[21940] = 1091906851;
assign addr[21941] = 1108329711;
assign addr[21942] = 1124664687;
assign addr[21943] = 1140910484;
assign addr[21944] = 1157065814;
assign addr[21945] = 1173129396;
assign addr[21946] = 1189099956;
assign addr[21947] = 1204976227;
assign addr[21948] = 1220756951;
assign addr[21949] = 1236440877;
assign addr[21950] = 1252026760;
assign addr[21951] = 1267513365;
assign addr[21952] = 1282899464;
assign addr[21953] = 1298183838;
assign addr[21954] = 1313365273;
assign addr[21955] = 1328442566;
assign addr[21956] = 1343414522;
assign addr[21957] = 1358279953;
assign addr[21958] = 1373037681;
assign addr[21959] = 1387686535;
assign addr[21960] = 1402225355;
assign addr[21961] = 1416652986;
assign addr[21962] = 1430968286;
assign addr[21963] = 1445170118;
assign addr[21964] = 1459257358;
assign addr[21965] = 1473228887;
assign addr[21966] = 1487083598;
assign addr[21967] = 1500820393;
assign addr[21968] = 1514438181;
assign addr[21969] = 1527935884;
assign addr[21970] = 1541312431;
assign addr[21971] = 1554566762;
assign addr[21972] = 1567697824;
assign addr[21973] = 1580704578;
assign addr[21974] = 1593585992;
assign addr[21975] = 1606341043;
assign addr[21976] = 1618968722;
assign addr[21977] = 1631468027;
assign addr[21978] = 1643837966;
assign addr[21979] = 1656077559;
assign addr[21980] = 1668185835;
assign addr[21981] = 1680161834;
assign addr[21982] = 1692004606;
assign addr[21983] = 1703713213;
assign addr[21984] = 1715286726;
assign addr[21985] = 1726724227;
assign addr[21986] = 1738024810;
assign addr[21987] = 1749187577;
assign addr[21988] = 1760211645;
assign addr[21989] = 1771096139;
assign addr[21990] = 1781840195;
assign addr[21991] = 1792442963;
assign addr[21992] = 1802903601;
assign addr[21993] = 1813221279;
assign addr[21994] = 1823395180;
assign addr[21995] = 1833424497;
assign addr[21996] = 1843308435;
assign addr[21997] = 1853046210;
assign addr[21998] = 1862637049;
assign addr[21999] = 1872080193;
assign addr[22000] = 1881374892;
assign addr[22001] = 1890520410;
assign addr[22002] = 1899516021;
assign addr[22003] = 1908361011;
assign addr[22004] = 1917054681;
assign addr[22005] = 1925596340;
assign addr[22006] = 1933985310;
assign addr[22007] = 1942220928;
assign addr[22008] = 1950302539;
assign addr[22009] = 1958229503;
assign addr[22010] = 1966001192;
assign addr[22011] = 1973616989;
assign addr[22012] = 1981076290;
assign addr[22013] = 1988378503;
assign addr[22014] = 1995523051;
assign addr[22015] = 2002509365;
assign addr[22016] = 2009336893;
assign addr[22017] = 2016005093;
assign addr[22018] = 2022513436;
assign addr[22019] = 2028861406;
assign addr[22020] = 2035048499;
assign addr[22021] = 2041074226;
assign addr[22022] = 2046938108;
assign addr[22023] = 2052639680;
assign addr[22024] = 2058178491;
assign addr[22025] = 2063554100;
assign addr[22026] = 2068766083;
assign addr[22027] = 2073814024;
assign addr[22028] = 2078697525;
assign addr[22029] = 2083416198;
assign addr[22030] = 2087969669;
assign addr[22031] = 2092357577;
assign addr[22032] = 2096579573;
assign addr[22033] = 2100635323;
assign addr[22034] = 2104524506;
assign addr[22035] = 2108246813;
assign addr[22036] = 2111801949;
assign addr[22037] = 2115189632;
assign addr[22038] = 2118409593;
assign addr[22039] = 2121461578;
assign addr[22040] = 2124345343;
assign addr[22041] = 2127060661;
assign addr[22042] = 2129607316;
assign addr[22043] = 2131985106;
assign addr[22044] = 2134193842;
assign addr[22045] = 2136233350;
assign addr[22046] = 2138103468;
assign addr[22047] = 2139804048;
assign addr[22048] = 2141334954;
assign addr[22049] = 2142696065;
assign addr[22050] = 2143887273;
assign addr[22051] = 2144908484;
assign addr[22052] = 2145759618;
assign addr[22053] = 2146440605;
assign addr[22054] = 2146951393;
assign addr[22055] = 2147291941;
assign addr[22056] = 2147462221;
assign addr[22057] = 2147462221;
assign addr[22058] = 2147291941;
assign addr[22059] = 2146951393;
assign addr[22060] = 2146440605;
assign addr[22061] = 2145759618;
assign addr[22062] = 2144908484;
assign addr[22063] = 2143887273;
assign addr[22064] = 2142696065;
assign addr[22065] = 2141334954;
assign addr[22066] = 2139804048;
assign addr[22067] = 2138103468;
assign addr[22068] = 2136233350;
assign addr[22069] = 2134193842;
assign addr[22070] = 2131985106;
assign addr[22071] = 2129607316;
assign addr[22072] = 2127060661;
assign addr[22073] = 2124345343;
assign addr[22074] = 2121461578;
assign addr[22075] = 2118409593;
assign addr[22076] = 2115189632;
assign addr[22077] = 2111801949;
assign addr[22078] = 2108246813;
assign addr[22079] = 2104524506;
assign addr[22080] = 2100635323;
assign addr[22081] = 2096579573;
assign addr[22082] = 2092357577;
assign addr[22083] = 2087969669;
assign addr[22084] = 2083416198;
assign addr[22085] = 2078697525;
assign addr[22086] = 2073814024;
assign addr[22087] = 2068766083;
assign addr[22088] = 2063554100;
assign addr[22089] = 2058178491;
assign addr[22090] = 2052639680;
assign addr[22091] = 2046938108;
assign addr[22092] = 2041074226;
assign addr[22093] = 2035048499;
assign addr[22094] = 2028861406;
assign addr[22095] = 2022513436;
assign addr[22096] = 2016005093;
assign addr[22097] = 2009336893;
assign addr[22098] = 2002509365;
assign addr[22099] = 1995523051;
assign addr[22100] = 1988378503;
assign addr[22101] = 1981076290;
assign addr[22102] = 1973616989;
assign addr[22103] = 1966001192;
assign addr[22104] = 1958229503;
assign addr[22105] = 1950302539;
assign addr[22106] = 1942220928;
assign addr[22107] = 1933985310;
assign addr[22108] = 1925596340;
assign addr[22109] = 1917054681;
assign addr[22110] = 1908361011;
assign addr[22111] = 1899516021;
assign addr[22112] = 1890520410;
assign addr[22113] = 1881374892;
assign addr[22114] = 1872080193;
assign addr[22115] = 1862637049;
assign addr[22116] = 1853046210;
assign addr[22117] = 1843308435;
assign addr[22118] = 1833424497;
assign addr[22119] = 1823395180;
assign addr[22120] = 1813221279;
assign addr[22121] = 1802903601;
assign addr[22122] = 1792442963;
assign addr[22123] = 1781840195;
assign addr[22124] = 1771096139;
assign addr[22125] = 1760211645;
assign addr[22126] = 1749187577;
assign addr[22127] = 1738024810;
assign addr[22128] = 1726724227;
assign addr[22129] = 1715286726;
assign addr[22130] = 1703713213;
assign addr[22131] = 1692004606;
assign addr[22132] = 1680161834;
assign addr[22133] = 1668185835;
assign addr[22134] = 1656077559;
assign addr[22135] = 1643837966;
assign addr[22136] = 1631468027;
assign addr[22137] = 1618968722;
assign addr[22138] = 1606341043;
assign addr[22139] = 1593585992;
assign addr[22140] = 1580704578;
assign addr[22141] = 1567697824;
assign addr[22142] = 1554566762;
assign addr[22143] = 1541312431;
assign addr[22144] = 1527935884;
assign addr[22145] = 1514438181;
assign addr[22146] = 1500820393;
assign addr[22147] = 1487083598;
assign addr[22148] = 1473228887;
assign addr[22149] = 1459257358;
assign addr[22150] = 1445170118;
assign addr[22151] = 1430968286;
assign addr[22152] = 1416652986;
assign addr[22153] = 1402225355;
assign addr[22154] = 1387686535;
assign addr[22155] = 1373037681;
assign addr[22156] = 1358279953;
assign addr[22157] = 1343414522;
assign addr[22158] = 1328442566;
assign addr[22159] = 1313365273;
assign addr[22160] = 1298183838;
assign addr[22161] = 1282899464;
assign addr[22162] = 1267513365;
assign addr[22163] = 1252026760;
assign addr[22164] = 1236440877;
assign addr[22165] = 1220756951;
assign addr[22166] = 1204976227;
assign addr[22167] = 1189099956;
assign addr[22168] = 1173129396;
assign addr[22169] = 1157065814;
assign addr[22170] = 1140910484;
assign addr[22171] = 1124664687;
assign addr[22172] = 1108329711;
assign addr[22173] = 1091906851;
assign addr[22174] = 1075397409;
assign addr[22175] = 1058802695;
assign addr[22176] = 1042124025;
assign addr[22177] = 1025362720;
assign addr[22178] = 1008520110;
assign addr[22179] = 991597531;
assign addr[22180] = 974596324;
assign addr[22181] = 957517838;
assign addr[22182] = 940363427;
assign addr[22183] = 923134450;
assign addr[22184] = 905832274;
assign addr[22185] = 888458272;
assign addr[22186] = 871013820;
assign addr[22187] = 853500302;
assign addr[22188] = 835919107;
assign addr[22189] = 818271628;
assign addr[22190] = 800559266;
assign addr[22191] = 782783424;
assign addr[22192] = 764945512;
assign addr[22193] = 747046944;
assign addr[22194] = 729089140;
assign addr[22195] = 711073524;
assign addr[22196] = 693001525;
assign addr[22197] = 674874574;
assign addr[22198] = 656694110;
assign addr[22199] = 638461574;
assign addr[22200] = 620178412;
assign addr[22201] = 601846074;
assign addr[22202] = 583466013;
assign addr[22203] = 565039687;
assign addr[22204] = 546568556;
assign addr[22205] = 528054086;
assign addr[22206] = 509497745;
assign addr[22207] = 490901003;
assign addr[22208] = 472265336;
assign addr[22209] = 453592221;
assign addr[22210] = 434883140;
assign addr[22211] = 416139574;
assign addr[22212] = 397363011;
assign addr[22213] = 378554940;
assign addr[22214] = 359716852;
assign addr[22215] = 340850240;
assign addr[22216] = 321956601;
assign addr[22217] = 303037433;
assign addr[22218] = 284094236;
assign addr[22219] = 265128512;
assign addr[22220] = 246141764;
assign addr[22221] = 227135500;
assign addr[22222] = 208111224;
assign addr[22223] = 189070447;
assign addr[22224] = 170014678;
assign addr[22225] = 150945428;
assign addr[22226] = 131864208;
assign addr[22227] = 112772533;
assign addr[22228] = 93671915;
assign addr[22229] = 74563870;
assign addr[22230] = 55449912;
assign addr[22231] = 36331557;
assign addr[22232] = 17210322;
assign addr[22233] = -1912278;
assign addr[22234] = -21034727;
assign addr[22235] = -40155507;
assign addr[22236] = -59273104;
assign addr[22237] = -78386000;
assign addr[22238] = -97492681;
assign addr[22239] = -116591632;
assign addr[22240] = -135681337;
assign addr[22241] = -154760284;
assign addr[22242] = -173826959;
assign addr[22243] = -192879850;
assign addr[22244] = -211917448;
assign addr[22245] = -230938242;
assign addr[22246] = -249940723;
assign addr[22247] = -268923386;
assign addr[22248] = -287884725;
assign addr[22249] = -306823237;
assign addr[22250] = -325737419;
assign addr[22251] = -344625773;
assign addr[22252] = -363486799;
assign addr[22253] = -382319004;
assign addr[22254] = -401120892;
assign addr[22255] = -419890975;
assign addr[22256] = -438627762;
assign addr[22257] = -457329769;
assign addr[22258] = -475995513;
assign addr[22259] = -494623513;
assign addr[22260] = -513212292;
assign addr[22261] = -531760377;
assign addr[22262] = -550266296;
assign addr[22263] = -568728583;
assign addr[22264] = -587145773;
assign addr[22265] = -605516406;
assign addr[22266] = -623839025;
assign addr[22267] = -642112178;
assign addr[22268] = -660334415;
assign addr[22269] = -678504291;
assign addr[22270] = -696620367;
assign addr[22271] = -714681204;
assign addr[22272] = -732685372;
assign addr[22273] = -750631442;
assign addr[22274] = -768517992;
assign addr[22275] = -786343603;
assign addr[22276] = -804106861;
assign addr[22277] = -821806359;
assign addr[22278] = -839440693;
assign addr[22279] = -857008464;
assign addr[22280] = -874508280;
assign addr[22281] = -891938752;
assign addr[22282] = -909298500;
assign addr[22283] = -926586145;
assign addr[22284] = -943800318;
assign addr[22285] = -960939653;
assign addr[22286] = -978002791;
assign addr[22287] = -994988380;
assign addr[22288] = -1011895073;
assign addr[22289] = -1028721528;
assign addr[22290] = -1045466412;
assign addr[22291] = -1062128397;
assign addr[22292] = -1078706161;
assign addr[22293] = -1095198391;
assign addr[22294] = -1111603778;
assign addr[22295] = -1127921022;
assign addr[22296] = -1144148829;
assign addr[22297] = -1160285911;
assign addr[22298] = -1176330990;
assign addr[22299] = -1192282793;
assign addr[22300] = -1208140056;
assign addr[22301] = -1223901520;
assign addr[22302] = -1239565936;
assign addr[22303] = -1255132063;
assign addr[22304] = -1270598665;
assign addr[22305] = -1285964516;
assign addr[22306] = -1301228398;
assign addr[22307] = -1316389101;
assign addr[22308] = -1331445422;
assign addr[22309] = -1346396168;
assign addr[22310] = -1361240152;
assign addr[22311] = -1375976199;
assign addr[22312] = -1390603139;
assign addr[22313] = -1405119813;
assign addr[22314] = -1419525069;
assign addr[22315] = -1433817766;
assign addr[22316] = -1447996770;
assign addr[22317] = -1462060956;
assign addr[22318] = -1476009210;
assign addr[22319] = -1489840425;
assign addr[22320] = -1503553506;
assign addr[22321] = -1517147363;
assign addr[22322] = -1530620920;
assign addr[22323] = -1543973108;
assign addr[22324] = -1557202869;
assign addr[22325] = -1570309153;
assign addr[22326] = -1583290921;
assign addr[22327] = -1596147143;
assign addr[22328] = -1608876801;
assign addr[22329] = -1621478885;
assign addr[22330] = -1633952396;
assign addr[22331] = -1646296344;
assign addr[22332] = -1658509750;
assign addr[22333] = -1670591647;
assign addr[22334] = -1682541077;
assign addr[22335] = -1694357091;
assign addr[22336] = -1706038753;
assign addr[22337] = -1717585136;
assign addr[22338] = -1728995326;
assign addr[22339] = -1740268417;
assign addr[22340] = -1751403515;
assign addr[22341] = -1762399737;
assign addr[22342] = -1773256212;
assign addr[22343] = -1783972079;
assign addr[22344] = -1794546487;
assign addr[22345] = -1804978599;
assign addr[22346] = -1815267588;
assign addr[22347] = -1825412636;
assign addr[22348] = -1835412941;
assign addr[22349] = -1845267708;
assign addr[22350] = -1854976157;
assign addr[22351] = -1864537518;
assign addr[22352] = -1873951032;
assign addr[22353] = -1883215953;
assign addr[22354] = -1892331547;
assign addr[22355] = -1901297091;
assign addr[22356] = -1910111873;
assign addr[22357] = -1918775195;
assign addr[22358] = -1927286370;
assign addr[22359] = -1935644723;
assign addr[22360] = -1943849591;
assign addr[22361] = -1951900324;
assign addr[22362] = -1959796283;
assign addr[22363] = -1967536842;
assign addr[22364] = -1975121388;
assign addr[22365] = -1982549318;
assign addr[22366] = -1989820044;
assign addr[22367] = -1996932990;
assign addr[22368] = -2003887591;
assign addr[22369] = -2010683297;
assign addr[22370] = -2017319567;
assign addr[22371] = -2023795876;
assign addr[22372] = -2030111710;
assign addr[22373] = -2036266570;
assign addr[22374] = -2042259965;
assign addr[22375] = -2048091422;
assign addr[22376] = -2053760478;
assign addr[22377] = -2059266683;
assign addr[22378] = -2064609600;
assign addr[22379] = -2069788807;
assign addr[22380] = -2074803892;
assign addr[22381] = -2079654458;
assign addr[22382] = -2084340120;
assign addr[22383] = -2088860507;
assign addr[22384] = -2093215260;
assign addr[22385] = -2097404033;
assign addr[22386] = -2101426496;
assign addr[22387] = -2105282327;
assign addr[22388] = -2108971223;
assign addr[22389] = -2112492891;
assign addr[22390] = -2115847050;
assign addr[22391] = -2119033436;
assign addr[22392] = -2122051796;
assign addr[22393] = -2124901890;
assign addr[22394] = -2127583492;
assign addr[22395] = -2130096389;
assign addr[22396] = -2132440383;
assign addr[22397] = -2134615288;
assign addr[22398] = -2136620930;
assign addr[22399] = -2138457152;
assign addr[22400] = -2140123807;
assign addr[22401] = -2141620763;
assign addr[22402] = -2142947902;
assign addr[22403] = -2144105118;
assign addr[22404] = -2145092320;
assign addr[22405] = -2145909429;
assign addr[22406] = -2146556380;
assign addr[22407] = -2147033123;
assign addr[22408] = -2147339619;
assign addr[22409] = -2147475844;
assign addr[22410] = -2147441787;
assign addr[22411] = -2147237452;
assign addr[22412] = -2146862854;
assign addr[22413] = -2146318022;
assign addr[22414] = -2145603001;
assign addr[22415] = -2144717846;
assign addr[22416] = -2143662628;
assign addr[22417] = -2142437431;
assign addr[22418] = -2141042352;
assign addr[22419] = -2139477502;
assign addr[22420] = -2137743003;
assign addr[22421] = -2135838995;
assign addr[22422] = -2133765628;
assign addr[22423] = -2131523066;
assign addr[22424] = -2129111488;
assign addr[22425] = -2126531084;
assign addr[22426] = -2123782059;
assign addr[22427] = -2120864631;
assign addr[22428] = -2117779031;
assign addr[22429] = -2114525505;
assign addr[22430] = -2111104309;
assign addr[22431] = -2107515716;
assign addr[22432] = -2103760010;
assign addr[22433] = -2099837489;
assign addr[22434] = -2095748463;
assign addr[22435] = -2091493257;
assign addr[22436] = -2087072209;
assign addr[22437] = -2082485668;
assign addr[22438] = -2077733999;
assign addr[22439] = -2072817579;
assign addr[22440] = -2067736796;
assign addr[22441] = -2062492055;
assign addr[22442] = -2057083771;
assign addr[22443] = -2051512372;
assign addr[22444] = -2045778302;
assign addr[22445] = -2039882013;
assign addr[22446] = -2033823974;
assign addr[22447] = -2027604666;
assign addr[22448] = -2021224581;
assign addr[22449] = -2014684225;
assign addr[22450] = -2007984117;
assign addr[22451] = -2001124788;
assign addr[22452] = -1994106782;
assign addr[22453] = -1986930656;
assign addr[22454] = -1979596978;
assign addr[22455] = -1972106330;
assign addr[22456] = -1964459306;
assign addr[22457] = -1956656513;
assign addr[22458] = -1948698568;
assign addr[22459] = -1940586104;
assign addr[22460] = -1932319763;
assign addr[22461] = -1923900201;
assign addr[22462] = -1915328086;
assign addr[22463] = -1906604097;
assign addr[22464] = -1897728925;
assign addr[22465] = -1888703276;
assign addr[22466] = -1879527863;
assign addr[22467] = -1870203416;
assign addr[22468] = -1860730673;
assign addr[22469] = -1851110385;
assign addr[22470] = -1841343316;
assign addr[22471] = -1831430239;
assign addr[22472] = -1821371941;
assign addr[22473] = -1811169220;
assign addr[22474] = -1800822883;
assign addr[22475] = -1790333753;
assign addr[22476] = -1779702660;
assign addr[22477] = -1768930447;
assign addr[22478] = -1758017969;
assign addr[22479] = -1746966091;
assign addr[22480] = -1735775690;
assign addr[22481] = -1724447652;
assign addr[22482] = -1712982875;
assign addr[22483] = -1701382270;
assign addr[22484] = -1689646755;
assign addr[22485] = -1677777262;
assign addr[22486] = -1665774731;
assign addr[22487] = -1653640115;
assign addr[22488] = -1641374375;
assign addr[22489] = -1628978484;
assign addr[22490] = -1616453425;
assign addr[22491] = -1603800191;
assign addr[22492] = -1591019785;
assign addr[22493] = -1578113222;
assign addr[22494] = -1565081523;
assign addr[22495] = -1551925723;
assign addr[22496] = -1538646865;
assign addr[22497] = -1525246002;
assign addr[22498] = -1511724196;
assign addr[22499] = -1498082520;
assign addr[22500] = -1484322054;
assign addr[22501] = -1470443891;
assign addr[22502] = -1456449131;
assign addr[22503] = -1442338884;
assign addr[22504] = -1428114267;
assign addr[22505] = -1413776410;
assign addr[22506] = -1399326449;
assign addr[22507] = -1384765530;
assign addr[22508] = -1370094808;
assign addr[22509] = -1355315445;
assign addr[22510] = -1340428615;
assign addr[22511] = -1325435496;
assign addr[22512] = -1310337279;
assign addr[22513] = -1295135159;
assign addr[22514] = -1279830344;
assign addr[22515] = -1264424045;
assign addr[22516] = -1248917486;
assign addr[22517] = -1233311895;
assign addr[22518] = -1217608510;
assign addr[22519] = -1201808576;
assign addr[22520] = -1185913346;
assign addr[22521] = -1169924081;
assign addr[22522] = -1153842047;
assign addr[22523] = -1137668521;
assign addr[22524] = -1121404785;
assign addr[22525] = -1105052128;
assign addr[22526] = -1088611847;
assign addr[22527] = -1072085246;
assign addr[22528] = -1055473635;
assign addr[22529] = -1038778332;
assign addr[22530] = -1022000660;
assign addr[22531] = -1005141949;
assign addr[22532] = -988203537;
assign addr[22533] = -971186766;
assign addr[22534] = -954092986;
assign addr[22535] = -936923553;
assign addr[22536] = -919679827;
assign addr[22537] = -902363176;
assign addr[22538] = -884974973;
assign addr[22539] = -867516597;
assign addr[22540] = -849989433;
assign addr[22541] = -832394869;
assign addr[22542] = -814734301;
assign addr[22543] = -797009130;
assign addr[22544] = -779220762;
assign addr[22545] = -761370605;
assign addr[22546] = -743460077;
assign addr[22547] = -725490597;
assign addr[22548] = -707463589;
assign addr[22549] = -689380485;
assign addr[22550] = -671242716;
assign addr[22551] = -653051723;
assign addr[22552] = -634808946;
assign addr[22553] = -616515832;
assign addr[22554] = -598173833;
assign addr[22555] = -579784402;
assign addr[22556] = -561348998;
assign addr[22557] = -542869083;
assign addr[22558] = -524346121;
assign addr[22559] = -505781581;
assign addr[22560] = -487176937;
assign addr[22561] = -468533662;
assign addr[22562] = -449853235;
assign addr[22563] = -431137138;
assign addr[22564] = -412386854;
assign addr[22565] = -393603870;
assign addr[22566] = -374789676;
assign addr[22567] = -355945764;
assign addr[22568] = -337073627;
assign addr[22569] = -318174762;
assign addr[22570] = -299250668;
assign addr[22571] = -280302845;
assign addr[22572] = -261332796;
assign addr[22573] = -242342025;
assign addr[22574] = -223332037;
assign addr[22575] = -204304341;
assign addr[22576] = -185260444;
assign addr[22577] = -166201858;
assign addr[22578] = -147130093;
assign addr[22579] = -128046661;
assign addr[22580] = -108953076;
assign addr[22581] = -89850852;
assign addr[22582] = -70741503;
assign addr[22583] = -51626544;
assign addr[22584] = -32507492;
assign addr[22585] = -13385863;
assign addr[22586] = 5736829;
assign addr[22587] = 24859065;
assign addr[22588] = 43979330;
assign addr[22589] = 63096108;
assign addr[22590] = 82207882;
assign addr[22591] = 101313138;
assign addr[22592] = 120410361;
assign addr[22593] = 139498035;
assign addr[22594] = 158574649;
assign addr[22595] = 177638688;
assign addr[22596] = 196688642;
assign addr[22597] = 215722999;
assign addr[22598] = 234740251;
assign addr[22599] = 253738890;
assign addr[22600] = 272717408;
assign addr[22601] = 291674302;
assign addr[22602] = 310608068;
assign addr[22603] = 329517204;
assign addr[22604] = 348400212;
assign addr[22605] = 367255594;
assign addr[22606] = 386081854;
assign addr[22607] = 404877501;
assign addr[22608] = 423641043;
assign addr[22609] = 442370993;
assign addr[22610] = 461065866;
assign addr[22611] = 479724180;
assign addr[22612] = 498344454;
assign addr[22613] = 516925212;
assign addr[22614] = 535464981;
assign addr[22615] = 553962291;
assign addr[22616] = 572415676;
assign addr[22617] = 590823671;
assign addr[22618] = 609184818;
assign addr[22619] = 627497660;
assign addr[22620] = 645760745;
assign addr[22621] = 663972625;
assign addr[22622] = 682131857;
assign addr[22623] = 700236999;
assign addr[22624] = 718286617;
assign addr[22625] = 736279279;
assign addr[22626] = 754213559;
assign addr[22627] = 772088034;
assign addr[22628] = 789901288;
assign addr[22629] = 807651907;
assign addr[22630] = 825338484;
assign addr[22631] = 842959617;
assign addr[22632] = 860513908;
assign addr[22633] = 877999966;
assign addr[22634] = 895416404;
assign addr[22635] = 912761841;
assign addr[22636] = 930034901;
assign addr[22637] = 947234215;
assign addr[22638] = 964358420;
assign addr[22639] = 981406156;
assign addr[22640] = 998376073;
assign addr[22641] = 1015266825;
assign addr[22642] = 1032077073;
assign addr[22643] = 1048805483;
assign addr[22644] = 1065450729;
assign addr[22645] = 1082011492;
assign addr[22646] = 1098486458;
assign addr[22647] = 1114874320;
assign addr[22648] = 1131173780;
assign addr[22649] = 1147383544;
assign addr[22650] = 1163502328;
assign addr[22651] = 1179528853;
assign addr[22652] = 1195461849;
assign addr[22653] = 1211300053;
assign addr[22654] = 1227042207;
assign addr[22655] = 1242687064;
assign addr[22656] = 1258233384;
assign addr[22657] = 1273679934;
assign addr[22658] = 1289025489;
assign addr[22659] = 1304268832;
assign addr[22660] = 1319408754;
assign addr[22661] = 1334444055;
assign addr[22662] = 1349373543;
assign addr[22663] = 1364196034;
assign addr[22664] = 1378910353;
assign addr[22665] = 1393515332;
assign addr[22666] = 1408009814;
assign addr[22667] = 1422392650;
assign addr[22668] = 1436662698;
assign addr[22669] = 1450818828;
assign addr[22670] = 1464859917;
assign addr[22671] = 1478784851;
assign addr[22672] = 1492592527;
assign addr[22673] = 1506281850;
assign addr[22674] = 1519851733;
assign addr[22675] = 1533301101;
assign addr[22676] = 1546628888;
assign addr[22677] = 1559834037;
assign addr[22678] = 1572915501;
assign addr[22679] = 1585872242;
assign addr[22680] = 1598703233;
assign addr[22681] = 1611407456;
assign addr[22682] = 1623983905;
assign addr[22683] = 1636431582;
assign addr[22684] = 1648749499;
assign addr[22685] = 1660936681;
assign addr[22686] = 1672992161;
assign addr[22687] = 1684914983;
assign addr[22688] = 1696704201;
assign addr[22689] = 1708358881;
assign addr[22690] = 1719878099;
assign addr[22691] = 1731260941;
assign addr[22692] = 1742506504;
assign addr[22693] = 1753613897;
assign addr[22694] = 1764582240;
assign addr[22695] = 1775410662;
assign addr[22696] = 1786098304;
assign addr[22697] = 1796644320;
assign addr[22698] = 1807047873;
assign addr[22699] = 1817308138;
assign addr[22700] = 1827424302;
assign addr[22701] = 1837395562;
assign addr[22702] = 1847221128;
assign addr[22703] = 1856900221;
assign addr[22704] = 1866432072;
assign addr[22705] = 1875815927;
assign addr[22706] = 1885051042;
assign addr[22707] = 1894136683;
assign addr[22708] = 1903072131;
assign addr[22709] = 1911856677;
assign addr[22710] = 1920489624;
assign addr[22711] = 1928970288;
assign addr[22712] = 1937297997;
assign addr[22713] = 1945472089;
assign addr[22714] = 1953491918;
assign addr[22715] = 1961356847;
assign addr[22716] = 1969066252;
assign addr[22717] = 1976619522;
assign addr[22718] = 1984016058;
assign addr[22719] = 1991255274;
assign addr[22720] = 1998336596;
assign addr[22721] = 2005259462;
assign addr[22722] = 2012023322;
assign addr[22723] = 2018627642;
assign addr[22724] = 2025071897;
assign addr[22725] = 2031355576;
assign addr[22726] = 2037478181;
assign addr[22727] = 2043439226;
assign addr[22728] = 2049238240;
assign addr[22729] = 2054874761;
assign addr[22730] = 2060348343;
assign addr[22731] = 2065658552;
assign addr[22732] = 2070804967;
assign addr[22733] = 2075787180;
assign addr[22734] = 2080604795;
assign addr[22735] = 2085257431;
assign addr[22736] = 2089744719;
assign addr[22737] = 2094066304;
assign addr[22738] = 2098221841;
assign addr[22739] = 2102211002;
assign addr[22740] = 2106033471;
assign addr[22741] = 2109688944;
assign addr[22742] = 2113177132;
assign addr[22743] = 2116497758;
assign addr[22744] = 2119650558;
assign addr[22745] = 2122635283;
assign addr[22746] = 2125451696;
assign addr[22747] = 2128099574;
assign addr[22748] = 2130578706;
assign addr[22749] = 2132888897;
assign addr[22750] = 2135029962;
assign addr[22751] = 2137001733;
assign addr[22752] = 2138804053;
assign addr[22753] = 2140436778;
assign addr[22754] = 2141899780;
assign addr[22755] = 2143192942;
assign addr[22756] = 2144316162;
assign addr[22757] = 2145269351;
assign addr[22758] = 2146052433;
assign addr[22759] = 2146665347;
assign addr[22760] = 2147108043;
assign addr[22761] = 2147380486;
assign addr[22762] = 2147482655;
assign addr[22763] = 2147414542;
assign addr[22764] = 2147176152;
assign addr[22765] = 2146767505;
assign addr[22766] = 2146188631;
assign addr[22767] = 2145439578;
assign addr[22768] = 2144520405;
assign addr[22769] = 2143431184;
assign addr[22770] = 2142172003;
assign addr[22771] = 2140742960;
assign addr[22772] = 2139144169;
assign addr[22773] = 2137375758;
assign addr[22774] = 2135437865;
assign addr[22775] = 2133330646;
assign addr[22776] = 2131054266;
assign addr[22777] = 2128608907;
assign addr[22778] = 2125994762;
assign addr[22779] = 2123212038;
assign addr[22780] = 2120260957;
assign addr[22781] = 2117141752;
assign addr[22782] = 2113854671;
assign addr[22783] = 2110399974;
assign addr[22784] = 2106777935;
assign addr[22785] = 2102988841;
assign addr[22786] = 2099032994;
assign addr[22787] = 2094910706;
assign addr[22788] = 2090622304;
assign addr[22789] = 2086168128;
assign addr[22790] = 2081548533;
assign addr[22791] = 2076763883;
assign addr[22792] = 2071814558;
assign addr[22793] = 2066700952;
assign addr[22794] = 2061423468;
assign addr[22795] = 2055982526;
assign addr[22796] = 2050378558;
assign addr[22797] = 2044612007;
assign addr[22798] = 2038683330;
assign addr[22799] = 2032592999;
assign addr[22800] = 2026341495;
assign addr[22801] = 2019929315;
assign addr[22802] = 2013356967;
assign addr[22803] = 2006624971;
assign addr[22804] = 1999733863;
assign addr[22805] = 1992684188;
assign addr[22806] = 1985476506;
assign addr[22807] = 1978111387;
assign addr[22808] = 1970589416;
assign addr[22809] = 1962911189;
assign addr[22810] = 1955077316;
assign addr[22811] = 1947088417;
assign addr[22812] = 1938945125;
assign addr[22813] = 1930648088;
assign addr[22814] = 1922197961;
assign addr[22815] = 1913595416;
assign addr[22816] = 1904841135;
assign addr[22817] = 1895935811;
assign addr[22818] = 1886880151;
assign addr[22819] = 1877674873;
assign addr[22820] = 1868320707;
assign addr[22821] = 1858818395;
assign addr[22822] = 1849168689;
assign addr[22823] = 1839372356;
assign addr[22824] = 1829430172;
assign addr[22825] = 1819342925;
assign addr[22826] = 1809111415;
assign addr[22827] = 1798736454;
assign addr[22828] = 1788218865;
assign addr[22829] = 1777559480;
assign addr[22830] = 1766759146;
assign addr[22831] = 1755818718;
assign addr[22832] = 1744739065;
assign addr[22833] = 1733521064;
assign addr[22834] = 1722165606;
assign addr[22835] = 1710673591;
assign addr[22836] = 1699045930;
assign addr[22837] = 1687283545;
assign addr[22838] = 1675387369;
assign addr[22839] = 1663358344;
assign addr[22840] = 1651197426;
assign addr[22841] = 1638905577;
assign addr[22842] = 1626483774;
assign addr[22843] = 1613933000;
assign addr[22844] = 1601254251;
assign addr[22845] = 1588448533;
assign addr[22846] = 1575516860;
assign addr[22847] = 1562460258;
assign addr[22848] = 1549279763;
assign addr[22849] = 1535976419;
assign addr[22850] = 1522551282;
assign addr[22851] = 1509005416;
assign addr[22852] = 1495339895;
assign addr[22853] = 1481555802;
assign addr[22854] = 1467654232;
assign addr[22855] = 1453636285;
assign addr[22856] = 1439503074;
assign addr[22857] = 1425255719;
assign addr[22858] = 1410895350;
assign addr[22859] = 1396423105;
assign addr[22860] = 1381840133;
assign addr[22861] = 1367147589;
assign addr[22862] = 1352346639;
assign addr[22863] = 1337438456;
assign addr[22864] = 1322424222;
assign addr[22865] = 1307305128;
assign addr[22866] = 1292082373;
assign addr[22867] = 1276757164;
assign addr[22868] = 1261330715;
assign addr[22869] = 1245804251;
assign addr[22870] = 1230179002;
assign addr[22871] = 1214456207;
assign addr[22872] = 1198637114;
assign addr[22873] = 1182722976;
assign addr[22874] = 1166715055;
assign addr[22875] = 1150614620;
assign addr[22876] = 1134422949;
assign addr[22877] = 1118141326;
assign addr[22878] = 1101771040;
assign addr[22879] = 1085313391;
assign addr[22880] = 1068769683;
assign addr[22881] = 1052141228;
assign addr[22882] = 1035429345;
assign addr[22883] = 1018635358;
assign addr[22884] = 1001760600;
assign addr[22885] = 984806408;
assign addr[22886] = 967774128;
assign addr[22887] = 950665109;
assign addr[22888] = 933480707;
assign addr[22889] = 916222287;
assign addr[22890] = 898891215;
assign addr[22891] = 881488868;
assign addr[22892] = 864016623;
assign addr[22893] = 846475867;
assign addr[22894] = 828867991;
assign addr[22895] = 811194391;
assign addr[22896] = 793456467;
assign addr[22897] = 775655628;
assign addr[22898] = 757793284;
assign addr[22899] = 739870851;
assign addr[22900] = 721889752;
assign addr[22901] = 703851410;
assign addr[22902] = 685757258;
assign addr[22903] = 667608730;
assign addr[22904] = 649407264;
assign addr[22905] = 631154304;
assign addr[22906] = 612851297;
assign addr[22907] = 594499695;
assign addr[22908] = 576100953;
assign addr[22909] = 557656529;
assign addr[22910] = 539167887;
assign addr[22911] = 520636492;
assign addr[22912] = 502063814;
assign addr[22913] = 483451325;
assign addr[22914] = 464800501;
assign addr[22915] = 446112822;
assign addr[22916] = 427389768;
assign addr[22917] = 408632825;
assign addr[22918] = 389843480;
assign addr[22919] = 371023223;
assign addr[22920] = 352173546;
assign addr[22921] = 333295944;
assign addr[22922] = 314391913;
assign addr[22923] = 295462954;
assign addr[22924] = 276510565;
assign addr[22925] = 257536251;
assign addr[22926] = 238541516;
assign addr[22927] = 219527866;
assign addr[22928] = 200496809;
assign addr[22929] = 181449854;
assign addr[22930] = 162388511;
assign addr[22931] = 143314291;
assign addr[22932] = 124228708;
assign addr[22933] = 105133274;
assign addr[22934] = 86029503;
assign addr[22935] = 66918911;
assign addr[22936] = 47803013;
assign addr[22937] = 28683324;
assign addr[22938] = 9561361;
assign addr[22939] = -9561361;
assign addr[22940] = -28683324;
assign addr[22941] = -47803013;
assign addr[22942] = -66918911;
assign addr[22943] = -86029503;
assign addr[22944] = -105133274;
assign addr[22945] = -124228708;
assign addr[22946] = -143314291;
assign addr[22947] = -162388511;
assign addr[22948] = -181449854;
assign addr[22949] = -200496809;
assign addr[22950] = -219527866;
assign addr[22951] = -238541516;
assign addr[22952] = -257536251;
assign addr[22953] = -276510565;
assign addr[22954] = -295462953;
assign addr[22955] = -314391913;
assign addr[22956] = -333295944;
assign addr[22957] = -352173546;
assign addr[22958] = -371023223;
assign addr[22959] = -389843480;
assign addr[22960] = -408632825;
assign addr[22961] = -427389768;
assign addr[22962] = -446112822;
assign addr[22963] = -464800501;
assign addr[22964] = -483451325;
assign addr[22965] = -502063814;
assign addr[22966] = -520636492;
assign addr[22967] = -539167887;
assign addr[22968] = -557656529;
assign addr[22969] = -576100953;
assign addr[22970] = -594499695;
assign addr[22971] = -612851297;
assign addr[22972] = -631154304;
assign addr[22973] = -649407264;
assign addr[22974] = -667608730;
assign addr[22975] = -685757258;
assign addr[22976] = -703851410;
assign addr[22977] = -721889752;
assign addr[22978] = -739870851;
assign addr[22979] = -757793284;
assign addr[22980] = -775655628;
assign addr[22981] = -793456467;
assign addr[22982] = -811194391;
assign addr[22983] = -828867991;
assign addr[22984] = -846475867;
assign addr[22985] = -864016623;
assign addr[22986] = -881488868;
assign addr[22987] = -898891215;
assign addr[22988] = -916222287;
assign addr[22989] = -933480707;
assign addr[22990] = -950665109;
assign addr[22991] = -967774128;
assign addr[22992] = -984806408;
assign addr[22993] = -1001760600;
assign addr[22994] = -1018635358;
assign addr[22995] = -1035429345;
assign addr[22996] = -1052141228;
assign addr[22997] = -1068769683;
assign addr[22998] = -1085313391;
assign addr[22999] = -1101771040;
assign addr[23000] = -1118141326;
assign addr[23001] = -1134422949;
assign addr[23002] = -1150614620;
assign addr[23003] = -1166715055;
assign addr[23004] = -1182722976;
assign addr[23005] = -1198637114;
assign addr[23006] = -1214456207;
assign addr[23007] = -1230179002;
assign addr[23008] = -1245804251;
assign addr[23009] = -1261330715;
assign addr[23010] = -1276757164;
assign addr[23011] = -1292082373;
assign addr[23012] = -1307305128;
assign addr[23013] = -1322424222;
assign addr[23014] = -1337438456;
assign addr[23015] = -1352346639;
assign addr[23016] = -1367147589;
assign addr[23017] = -1381840133;
assign addr[23018] = -1396423105;
assign addr[23019] = -1410895350;
assign addr[23020] = -1425255719;
assign addr[23021] = -1439503074;
assign addr[23022] = -1453636285;
assign addr[23023] = -1467654232;
assign addr[23024] = -1481555802;
assign addr[23025] = -1495339895;
assign addr[23026] = -1509005416;
assign addr[23027] = -1522551282;
assign addr[23028] = -1535976419;
assign addr[23029] = -1549279763;
assign addr[23030] = -1562460258;
assign addr[23031] = -1575516860;
assign addr[23032] = -1588448533;
assign addr[23033] = -1601254251;
assign addr[23034] = -1613933000;
assign addr[23035] = -1626483774;
assign addr[23036] = -1638905577;
assign addr[23037] = -1651197426;
assign addr[23038] = -1663358344;
assign addr[23039] = -1675387369;
assign addr[23040] = -1687283545;
assign addr[23041] = -1699045930;
assign addr[23042] = -1710673591;
assign addr[23043] = -1722165606;
assign addr[23044] = -1733521064;
assign addr[23045] = -1744739065;
assign addr[23046] = -1755818718;
assign addr[23047] = -1766759146;
assign addr[23048] = -1777559480;
assign addr[23049] = -1788218865;
assign addr[23050] = -1798736454;
assign addr[23051] = -1809111415;
assign addr[23052] = -1819342925;
assign addr[23053] = -1829430172;
assign addr[23054] = -1839372356;
assign addr[23055] = -1849168689;
assign addr[23056] = -1858818395;
assign addr[23057] = -1868320707;
assign addr[23058] = -1877674873;
assign addr[23059] = -1886880151;
assign addr[23060] = -1895935811;
assign addr[23061] = -1904841135;
assign addr[23062] = -1913595416;
assign addr[23063] = -1922197961;
assign addr[23064] = -1930648088;
assign addr[23065] = -1938945125;
assign addr[23066] = -1947088417;
assign addr[23067] = -1955077316;
assign addr[23068] = -1962911189;
assign addr[23069] = -1970589416;
assign addr[23070] = -1978111387;
assign addr[23071] = -1985476506;
assign addr[23072] = -1992684188;
assign addr[23073] = -1999733863;
assign addr[23074] = -2006624971;
assign addr[23075] = -2013356967;
assign addr[23076] = -2019929315;
assign addr[23077] = -2026341495;
assign addr[23078] = -2032592999;
assign addr[23079] = -2038683330;
assign addr[23080] = -2044612007;
assign addr[23081] = -2050378558;
assign addr[23082] = -2055982526;
assign addr[23083] = -2061423468;
assign addr[23084] = -2066700952;
assign addr[23085] = -2071814558;
assign addr[23086] = -2076763883;
assign addr[23087] = -2081548533;
assign addr[23088] = -2086168128;
assign addr[23089] = -2090622304;
assign addr[23090] = -2094910706;
assign addr[23091] = -2099032994;
assign addr[23092] = -2102988841;
assign addr[23093] = -2106777935;
assign addr[23094] = -2110399974;
assign addr[23095] = -2113854671;
assign addr[23096] = -2117141752;
assign addr[23097] = -2120260957;
assign addr[23098] = -2123212038;
assign addr[23099] = -2125994762;
assign addr[23100] = -2128608907;
assign addr[23101] = -2131054266;
assign addr[23102] = -2133330646;
assign addr[23103] = -2135437865;
assign addr[23104] = -2137375758;
assign addr[23105] = -2139144169;
assign addr[23106] = -2140742960;
assign addr[23107] = -2142172003;
assign addr[23108] = -2143431184;
assign addr[23109] = -2144520405;
assign addr[23110] = -2145439578;
assign addr[23111] = -2146188631;
assign addr[23112] = -2146767505;
assign addr[23113] = -2147176152;
assign addr[23114] = -2147414542;
assign addr[23115] = -2147482655;
assign addr[23116] = -2147380486;
assign addr[23117] = -2147108043;
assign addr[23118] = -2146665347;
assign addr[23119] = -2146052433;
assign addr[23120] = -2145269351;
assign addr[23121] = -2144316162;
assign addr[23122] = -2143192942;
assign addr[23123] = -2141899780;
assign addr[23124] = -2140436778;
assign addr[23125] = -2138804053;
assign addr[23126] = -2137001733;
assign addr[23127] = -2135029962;
assign addr[23128] = -2132888897;
assign addr[23129] = -2130578706;
assign addr[23130] = -2128099574;
assign addr[23131] = -2125451696;
assign addr[23132] = -2122635283;
assign addr[23133] = -2119650558;
assign addr[23134] = -2116497758;
assign addr[23135] = -2113177132;
assign addr[23136] = -2109688944;
assign addr[23137] = -2106033471;
assign addr[23138] = -2102211002;
assign addr[23139] = -2098221841;
assign addr[23140] = -2094066304;
assign addr[23141] = -2089744719;
assign addr[23142] = -2085257431;
assign addr[23143] = -2080604795;
assign addr[23144] = -2075787180;
assign addr[23145] = -2070804967;
assign addr[23146] = -2065658552;
assign addr[23147] = -2060348343;
assign addr[23148] = -2054874761;
assign addr[23149] = -2049238240;
assign addr[23150] = -2043439226;
assign addr[23151] = -2037478181;
assign addr[23152] = -2031355576;
assign addr[23153] = -2025071897;
assign addr[23154] = -2018627642;
assign addr[23155] = -2012023322;
assign addr[23156] = -2005259462;
assign addr[23157] = -1998336596;
assign addr[23158] = -1991255274;
assign addr[23159] = -1984016058;
assign addr[23160] = -1976619522;
assign addr[23161] = -1969066252;
assign addr[23162] = -1961356847;
assign addr[23163] = -1953491918;
assign addr[23164] = -1945472089;
assign addr[23165] = -1937297997;
assign addr[23166] = -1928970288;
assign addr[23167] = -1920489624;
assign addr[23168] = -1911856677;
assign addr[23169] = -1903072131;
assign addr[23170] = -1894136683;
assign addr[23171] = -1885051042;
assign addr[23172] = -1875815927;
assign addr[23173] = -1866432072;
assign addr[23174] = -1856900221;
assign addr[23175] = -1847221128;
assign addr[23176] = -1837395562;
assign addr[23177] = -1827424302;
assign addr[23178] = -1817308138;
assign addr[23179] = -1807047873;
assign addr[23180] = -1796644320;
assign addr[23181] = -1786098304;
assign addr[23182] = -1775410662;
assign addr[23183] = -1764582240;
assign addr[23184] = -1753613897;
assign addr[23185] = -1742506504;
assign addr[23186] = -1731260941;
assign addr[23187] = -1719878099;
assign addr[23188] = -1708358881;
assign addr[23189] = -1696704201;
assign addr[23190] = -1684914983;
assign addr[23191] = -1672992161;
assign addr[23192] = -1660936681;
assign addr[23193] = -1648749499;
assign addr[23194] = -1636431582;
assign addr[23195] = -1623983905;
assign addr[23196] = -1611407456;
assign addr[23197] = -1598703233;
assign addr[23198] = -1585872242;
assign addr[23199] = -1572915501;
assign addr[23200] = -1559834037;
assign addr[23201] = -1546628888;
assign addr[23202] = -1533301101;
assign addr[23203] = -1519851733;
assign addr[23204] = -1506281850;
assign addr[23205] = -1492592527;
assign addr[23206] = -1478784851;
assign addr[23207] = -1464859917;
assign addr[23208] = -1450818828;
assign addr[23209] = -1436662698;
assign addr[23210] = -1422392650;
assign addr[23211] = -1408009814;
assign addr[23212] = -1393515332;
assign addr[23213] = -1378910353;
assign addr[23214] = -1364196034;
assign addr[23215] = -1349373543;
assign addr[23216] = -1334444055;
assign addr[23217] = -1319408754;
assign addr[23218] = -1304268832;
assign addr[23219] = -1289025489;
assign addr[23220] = -1273679934;
assign addr[23221] = -1258233384;
assign addr[23222] = -1242687064;
assign addr[23223] = -1227042207;
assign addr[23224] = -1211300053;
assign addr[23225] = -1195461849;
assign addr[23226] = -1179528853;
assign addr[23227] = -1163502328;
assign addr[23228] = -1147383544;
assign addr[23229] = -1131173780;
assign addr[23230] = -1114874320;
assign addr[23231] = -1098486458;
assign addr[23232] = -1082011492;
assign addr[23233] = -1065450729;
assign addr[23234] = -1048805483;
assign addr[23235] = -1032077073;
assign addr[23236] = -1015266825;
assign addr[23237] = -998376073;
assign addr[23238] = -981406156;
assign addr[23239] = -964358420;
assign addr[23240] = -947234215;
assign addr[23241] = -930034901;
assign addr[23242] = -912761841;
assign addr[23243] = -895416404;
assign addr[23244] = -877999966;
assign addr[23245] = -860513908;
assign addr[23246] = -842959617;
assign addr[23247] = -825338484;
assign addr[23248] = -807651907;
assign addr[23249] = -789901288;
assign addr[23250] = -772088034;
assign addr[23251] = -754213559;
assign addr[23252] = -736279279;
assign addr[23253] = -718286617;
assign addr[23254] = -700236999;
assign addr[23255] = -682131857;
assign addr[23256] = -663972625;
assign addr[23257] = -645760745;
assign addr[23258] = -627497660;
assign addr[23259] = -609184818;
assign addr[23260] = -590823671;
assign addr[23261] = -572415676;
assign addr[23262] = -553962291;
assign addr[23263] = -535464981;
assign addr[23264] = -516925212;
assign addr[23265] = -498344454;
assign addr[23266] = -479724180;
assign addr[23267] = -461065866;
assign addr[23268] = -442370993;
assign addr[23269] = -423641043;
assign addr[23270] = -404877501;
assign addr[23271] = -386081854;
assign addr[23272] = -367255594;
assign addr[23273] = -348400212;
assign addr[23274] = -329517204;
assign addr[23275] = -310608068;
assign addr[23276] = -291674302;
assign addr[23277] = -272717408;
assign addr[23278] = -253738890;
assign addr[23279] = -234740251;
assign addr[23280] = -215722999;
assign addr[23281] = -196688642;
assign addr[23282] = -177638688;
assign addr[23283] = -158574649;
assign addr[23284] = -139498035;
assign addr[23285] = -120410361;
assign addr[23286] = -101313138;
assign addr[23287] = -82207882;
assign addr[23288] = -63096108;
assign addr[23289] = -43979330;
assign addr[23290] = -24859065;
assign addr[23291] = -5736829;
assign addr[23292] = 13385863;
assign addr[23293] = 32507492;
assign addr[23294] = 51626544;
assign addr[23295] = 70741503;
assign addr[23296] = 89850852;
assign addr[23297] = 108953076;
assign addr[23298] = 128046661;
assign addr[23299] = 147130093;
assign addr[23300] = 166201858;
assign addr[23301] = 185260444;
assign addr[23302] = 204304341;
assign addr[23303] = 223332037;
assign addr[23304] = 242342025;
assign addr[23305] = 261332796;
assign addr[23306] = 280302845;
assign addr[23307] = 299250668;
assign addr[23308] = 318174762;
assign addr[23309] = 337073627;
assign addr[23310] = 355945764;
assign addr[23311] = 374789676;
assign addr[23312] = 393603870;
assign addr[23313] = 412386854;
assign addr[23314] = 431137138;
assign addr[23315] = 449853235;
assign addr[23316] = 468533662;
assign addr[23317] = 487176937;
assign addr[23318] = 505781581;
assign addr[23319] = 524346121;
assign addr[23320] = 542869083;
assign addr[23321] = 561348998;
assign addr[23322] = 579784402;
assign addr[23323] = 598173833;
assign addr[23324] = 616515832;
assign addr[23325] = 634808946;
assign addr[23326] = 653051723;
assign addr[23327] = 671242716;
assign addr[23328] = 689380485;
assign addr[23329] = 707463589;
assign addr[23330] = 725490597;
assign addr[23331] = 743460077;
assign addr[23332] = 761370605;
assign addr[23333] = 779220762;
assign addr[23334] = 797009130;
assign addr[23335] = 814734301;
assign addr[23336] = 832394869;
assign addr[23337] = 849989433;
assign addr[23338] = 867516597;
assign addr[23339] = 884974973;
assign addr[23340] = 902363176;
assign addr[23341] = 919679827;
assign addr[23342] = 936923553;
assign addr[23343] = 954092986;
assign addr[23344] = 971186766;
assign addr[23345] = 988203537;
assign addr[23346] = 1005141949;
assign addr[23347] = 1022000660;
assign addr[23348] = 1038778332;
assign addr[23349] = 1055473635;
assign addr[23350] = 1072085246;
assign addr[23351] = 1088611847;
assign addr[23352] = 1105052128;
assign addr[23353] = 1121404785;
assign addr[23354] = 1137668521;
assign addr[23355] = 1153842047;
assign addr[23356] = 1169924081;
assign addr[23357] = 1185913346;
assign addr[23358] = 1201808576;
assign addr[23359] = 1217608510;
assign addr[23360] = 1233311895;
assign addr[23361] = 1248917486;
assign addr[23362] = 1264424045;
assign addr[23363] = 1279830344;
assign addr[23364] = 1295135159;
assign addr[23365] = 1310337279;
assign addr[23366] = 1325435496;
assign addr[23367] = 1340428615;
assign addr[23368] = 1355315445;
assign addr[23369] = 1370094808;
assign addr[23370] = 1384765530;
assign addr[23371] = 1399326449;
assign addr[23372] = 1413776410;
assign addr[23373] = 1428114267;
assign addr[23374] = 1442338884;
assign addr[23375] = 1456449131;
assign addr[23376] = 1470443891;
assign addr[23377] = 1484322054;
assign addr[23378] = 1498082520;
assign addr[23379] = 1511724196;
assign addr[23380] = 1525246002;
assign addr[23381] = 1538646865;
assign addr[23382] = 1551925723;
assign addr[23383] = 1565081523;
assign addr[23384] = 1578113222;
assign addr[23385] = 1591019785;
assign addr[23386] = 1603800191;
assign addr[23387] = 1616453425;
assign addr[23388] = 1628978484;
assign addr[23389] = 1641374375;
assign addr[23390] = 1653640115;
assign addr[23391] = 1665774731;
assign addr[23392] = 1677777262;
assign addr[23393] = 1689646755;
assign addr[23394] = 1701382270;
assign addr[23395] = 1712982875;
assign addr[23396] = 1724447652;
assign addr[23397] = 1735775690;
assign addr[23398] = 1746966091;
assign addr[23399] = 1758017969;
assign addr[23400] = 1768930447;
assign addr[23401] = 1779702660;
assign addr[23402] = 1790333753;
assign addr[23403] = 1800822883;
assign addr[23404] = 1811169220;
assign addr[23405] = 1821371941;
assign addr[23406] = 1831430239;
assign addr[23407] = 1841343316;
assign addr[23408] = 1851110385;
assign addr[23409] = 1860730673;
assign addr[23410] = 1870203416;
assign addr[23411] = 1879527863;
assign addr[23412] = 1888703276;
assign addr[23413] = 1897728925;
assign addr[23414] = 1906604097;
assign addr[23415] = 1915328086;
assign addr[23416] = 1923900201;
assign addr[23417] = 1932319763;
assign addr[23418] = 1940586104;
assign addr[23419] = 1948698568;
assign addr[23420] = 1956656513;
assign addr[23421] = 1964459306;
assign addr[23422] = 1972106330;
assign addr[23423] = 1979596978;
assign addr[23424] = 1986930656;
assign addr[23425] = 1994106782;
assign addr[23426] = 2001124788;
assign addr[23427] = 2007984117;
assign addr[23428] = 2014684225;
assign addr[23429] = 2021224581;
assign addr[23430] = 2027604666;
assign addr[23431] = 2033823974;
assign addr[23432] = 2039882013;
assign addr[23433] = 2045778302;
assign addr[23434] = 2051512372;
assign addr[23435] = 2057083771;
assign addr[23436] = 2062492055;
assign addr[23437] = 2067736796;
assign addr[23438] = 2072817579;
assign addr[23439] = 2077733999;
assign addr[23440] = 2082485668;
assign addr[23441] = 2087072209;
assign addr[23442] = 2091493257;
assign addr[23443] = 2095748463;
assign addr[23444] = 2099837489;
assign addr[23445] = 2103760010;
assign addr[23446] = 2107515716;
assign addr[23447] = 2111104309;
assign addr[23448] = 2114525505;
assign addr[23449] = 2117779031;
assign addr[23450] = 2120864631;
assign addr[23451] = 2123782059;
assign addr[23452] = 2126531084;
assign addr[23453] = 2129111488;
assign addr[23454] = 2131523066;
assign addr[23455] = 2133765628;
assign addr[23456] = 2135838995;
assign addr[23457] = 2137743003;
assign addr[23458] = 2139477502;
assign addr[23459] = 2141042352;
assign addr[23460] = 2142437431;
assign addr[23461] = 2143662628;
assign addr[23462] = 2144717846;
assign addr[23463] = 2145603001;
assign addr[23464] = 2146318022;
assign addr[23465] = 2146862854;
assign addr[23466] = 2147237452;
assign addr[23467] = 2147441787;
assign addr[23468] = 2147475844;
assign addr[23469] = 2147339619;
assign addr[23470] = 2147033123;
assign addr[23471] = 2146556380;
assign addr[23472] = 2145909429;
assign addr[23473] = 2145092320;
assign addr[23474] = 2144105118;
assign addr[23475] = 2142947902;
assign addr[23476] = 2141620763;
assign addr[23477] = 2140123807;
assign addr[23478] = 2138457152;
assign addr[23479] = 2136620930;
assign addr[23480] = 2134615288;
assign addr[23481] = 2132440383;
assign addr[23482] = 2130096389;
assign addr[23483] = 2127583492;
assign addr[23484] = 2124901890;
assign addr[23485] = 2122051796;
assign addr[23486] = 2119033436;
assign addr[23487] = 2115847050;
assign addr[23488] = 2112492891;
assign addr[23489] = 2108971223;
assign addr[23490] = 2105282327;
assign addr[23491] = 2101426496;
assign addr[23492] = 2097404033;
assign addr[23493] = 2093215260;
assign addr[23494] = 2088860507;
assign addr[23495] = 2084340120;
assign addr[23496] = 2079654458;
assign addr[23497] = 2074803892;
assign addr[23498] = 2069788807;
assign addr[23499] = 2064609600;
assign addr[23500] = 2059266683;
assign addr[23501] = 2053760478;
assign addr[23502] = 2048091422;
assign addr[23503] = 2042259965;
assign addr[23504] = 2036266570;
assign addr[23505] = 2030111710;
assign addr[23506] = 2023795876;
assign addr[23507] = 2017319567;
assign addr[23508] = 2010683297;
assign addr[23509] = 2003887591;
assign addr[23510] = 1996932990;
assign addr[23511] = 1989820044;
assign addr[23512] = 1982549318;
assign addr[23513] = 1975121388;
assign addr[23514] = 1967536842;
assign addr[23515] = 1959796283;
assign addr[23516] = 1951900324;
assign addr[23517] = 1943849591;
assign addr[23518] = 1935644723;
assign addr[23519] = 1927286370;
assign addr[23520] = 1918775195;
assign addr[23521] = 1910111873;
assign addr[23522] = 1901297091;
assign addr[23523] = 1892331547;
assign addr[23524] = 1883215953;
assign addr[23525] = 1873951032;
assign addr[23526] = 1864537518;
assign addr[23527] = 1854976157;
assign addr[23528] = 1845267708;
assign addr[23529] = 1835412941;
assign addr[23530] = 1825412636;
assign addr[23531] = 1815267588;
assign addr[23532] = 1804978599;
assign addr[23533] = 1794546487;
assign addr[23534] = 1783972079;
assign addr[23535] = 1773256212;
assign addr[23536] = 1762399737;
assign addr[23537] = 1751403515;
assign addr[23538] = 1740268417;
assign addr[23539] = 1728995326;
assign addr[23540] = 1717585136;
assign addr[23541] = 1706038753;
assign addr[23542] = 1694357091;
assign addr[23543] = 1682541077;
assign addr[23544] = 1670591647;
assign addr[23545] = 1658509750;
assign addr[23546] = 1646296344;
assign addr[23547] = 1633952396;
assign addr[23548] = 1621478885;
assign addr[23549] = 1608876801;
assign addr[23550] = 1596147143;
assign addr[23551] = 1583290921;
assign addr[23552] = 1570309153;
assign addr[23553] = 1557202869;
assign addr[23554] = 1543973108;
assign addr[23555] = 1530620920;
assign addr[23556] = 1517147363;
assign addr[23557] = 1503553506;
assign addr[23558] = 1489840425;
assign addr[23559] = 1476009210;
assign addr[23560] = 1462060956;
assign addr[23561] = 1447996770;
assign addr[23562] = 1433817766;
assign addr[23563] = 1419525069;
assign addr[23564] = 1405119813;
assign addr[23565] = 1390603139;
assign addr[23566] = 1375976199;
assign addr[23567] = 1361240152;
assign addr[23568] = 1346396168;
assign addr[23569] = 1331445422;
assign addr[23570] = 1316389101;
assign addr[23571] = 1301228398;
assign addr[23572] = 1285964516;
assign addr[23573] = 1270598665;
assign addr[23574] = 1255132063;
assign addr[23575] = 1239565936;
assign addr[23576] = 1223901520;
assign addr[23577] = 1208140056;
assign addr[23578] = 1192282793;
assign addr[23579] = 1176330990;
assign addr[23580] = 1160285911;
assign addr[23581] = 1144148829;
assign addr[23582] = 1127921022;
assign addr[23583] = 1111603778;
assign addr[23584] = 1095198391;
assign addr[23585] = 1078706161;
assign addr[23586] = 1062128397;
assign addr[23587] = 1045466412;
assign addr[23588] = 1028721528;
assign addr[23589] = 1011895073;
assign addr[23590] = 994988380;
assign addr[23591] = 978002791;
assign addr[23592] = 960939653;
assign addr[23593] = 943800318;
assign addr[23594] = 926586145;
assign addr[23595] = 909298500;
assign addr[23596] = 891938752;
assign addr[23597] = 874508280;
assign addr[23598] = 857008464;
assign addr[23599] = 839440693;
assign addr[23600] = 821806359;
assign addr[23601] = 804106861;
assign addr[23602] = 786343603;
assign addr[23603] = 768517992;
assign addr[23604] = 750631442;
assign addr[23605] = 732685372;
assign addr[23606] = 714681204;
assign addr[23607] = 696620367;
assign addr[23608] = 678504291;
assign addr[23609] = 660334415;
assign addr[23610] = 642112178;
assign addr[23611] = 623839025;
assign addr[23612] = 605516406;
assign addr[23613] = 587145773;
assign addr[23614] = 568728583;
assign addr[23615] = 550266296;
assign addr[23616] = 531760377;
assign addr[23617] = 513212292;
assign addr[23618] = 494623513;
assign addr[23619] = 475995513;
assign addr[23620] = 457329769;
assign addr[23621] = 438627762;
assign addr[23622] = 419890975;
assign addr[23623] = 401120892;
assign addr[23624] = 382319004;
assign addr[23625] = 363486799;
assign addr[23626] = 344625773;
assign addr[23627] = 325737419;
assign addr[23628] = 306823237;
assign addr[23629] = 287884725;
assign addr[23630] = 268923386;
assign addr[23631] = 249940723;
assign addr[23632] = 230938242;
assign addr[23633] = 211917448;
assign addr[23634] = 192879850;
assign addr[23635] = 173826959;
assign addr[23636] = 154760284;
assign addr[23637] = 135681337;
assign addr[23638] = 116591632;
assign addr[23639] = 97492681;
assign addr[23640] = 78386000;
assign addr[23641] = 59273104;
assign addr[23642] = 40155507;
assign addr[23643] = 21034727;
assign addr[23644] = 1912278;
assign addr[23645] = -17210322;
assign addr[23646] = -36331557;
assign addr[23647] = -55449912;
assign addr[23648] = -74563870;
assign addr[23649] = -93671915;
assign addr[23650] = -112772533;
assign addr[23651] = -131864208;
assign addr[23652] = -150945428;
assign addr[23653] = -170014678;
assign addr[23654] = -189070447;
assign addr[23655] = -208111224;
assign addr[23656] = -227135500;
assign addr[23657] = -246141764;
assign addr[23658] = -265128512;
assign addr[23659] = -284094236;
assign addr[23660] = -303037433;
assign addr[23661] = -321956601;
assign addr[23662] = -340850240;
assign addr[23663] = -359716852;
assign addr[23664] = -378554940;
assign addr[23665] = -397363011;
assign addr[23666] = -416139574;
assign addr[23667] = -434883140;
assign addr[23668] = -453592221;
assign addr[23669] = -472265336;
assign addr[23670] = -490901003;
assign addr[23671] = -509497745;
assign addr[23672] = -528054086;
assign addr[23673] = -546568556;
assign addr[23674] = -565039687;
assign addr[23675] = -583466013;
assign addr[23676] = -601846074;
assign addr[23677] = -620178412;
assign addr[23678] = -638461574;
assign addr[23679] = -656694110;
assign addr[23680] = -674874574;
assign addr[23681] = -693001525;
assign addr[23682] = -711073524;
assign addr[23683] = -729089140;
assign addr[23684] = -747046944;
assign addr[23685] = -764945512;
assign addr[23686] = -782783424;
assign addr[23687] = -800559266;
assign addr[23688] = -818271628;
assign addr[23689] = -835919107;
assign addr[23690] = -853500302;
assign addr[23691] = -871013820;
assign addr[23692] = -888458272;
assign addr[23693] = -905832274;
assign addr[23694] = -923134450;
assign addr[23695] = -940363427;
assign addr[23696] = -957517838;
assign addr[23697] = -974596324;
assign addr[23698] = -991597531;
assign addr[23699] = -1008520110;
assign addr[23700] = -1025362720;
assign addr[23701] = -1042124025;
assign addr[23702] = -1058802695;
assign addr[23703] = -1075397409;
assign addr[23704] = -1091906851;
assign addr[23705] = -1108329711;
assign addr[23706] = -1124664687;
assign addr[23707] = -1140910484;
assign addr[23708] = -1157065814;
assign addr[23709] = -1173129396;
assign addr[23710] = -1189099956;
assign addr[23711] = -1204976227;
assign addr[23712] = -1220756951;
assign addr[23713] = -1236440877;
assign addr[23714] = -1252026760;
assign addr[23715] = -1267513365;
assign addr[23716] = -1282899464;
assign addr[23717] = -1298183838;
assign addr[23718] = -1313365273;
assign addr[23719] = -1328442566;
assign addr[23720] = -1343414522;
assign addr[23721] = -1358279953;
assign addr[23722] = -1373037681;
assign addr[23723] = -1387686535;
assign addr[23724] = -1402225355;
assign addr[23725] = -1416652986;
assign addr[23726] = -1430968286;
assign addr[23727] = -1445170118;
assign addr[23728] = -1459257358;
assign addr[23729] = -1473228887;
assign addr[23730] = -1487083598;
assign addr[23731] = -1500820393;
assign addr[23732] = -1514438181;
assign addr[23733] = -1527935884;
assign addr[23734] = -1541312431;
assign addr[23735] = -1554566762;
assign addr[23736] = -1567697824;
assign addr[23737] = -1580704578;
assign addr[23738] = -1593585992;
assign addr[23739] = -1606341043;
assign addr[23740] = -1618968722;
assign addr[23741] = -1631468027;
assign addr[23742] = -1643837966;
assign addr[23743] = -1656077559;
assign addr[23744] = -1668185835;
assign addr[23745] = -1680161834;
assign addr[23746] = -1692004606;
assign addr[23747] = -1703713213;
assign addr[23748] = -1715286726;
assign addr[23749] = -1726724227;
assign addr[23750] = -1738024810;
assign addr[23751] = -1749187577;
assign addr[23752] = -1760211645;
assign addr[23753] = -1771096139;
assign addr[23754] = -1781840195;
assign addr[23755] = -1792442963;
assign addr[23756] = -1802903601;
assign addr[23757] = -1813221279;
assign addr[23758] = -1823395180;
assign addr[23759] = -1833424497;
assign addr[23760] = -1843308435;
assign addr[23761] = -1853046210;
assign addr[23762] = -1862637049;
assign addr[23763] = -1872080193;
assign addr[23764] = -1881374892;
assign addr[23765] = -1890520410;
assign addr[23766] = -1899516021;
assign addr[23767] = -1908361011;
assign addr[23768] = -1917054681;
assign addr[23769] = -1925596340;
assign addr[23770] = -1933985310;
assign addr[23771] = -1942220928;
assign addr[23772] = -1950302539;
assign addr[23773] = -1958229503;
assign addr[23774] = -1966001192;
assign addr[23775] = -1973616989;
assign addr[23776] = -1981076290;
assign addr[23777] = -1988378503;
assign addr[23778] = -1995523051;
assign addr[23779] = -2002509365;
assign addr[23780] = -2009336893;
assign addr[23781] = -2016005093;
assign addr[23782] = -2022513436;
assign addr[23783] = -2028861406;
assign addr[23784] = -2035048499;
assign addr[23785] = -2041074226;
assign addr[23786] = -2046938108;
assign addr[23787] = -2052639680;
assign addr[23788] = -2058178491;
assign addr[23789] = -2063554100;
assign addr[23790] = -2068766083;
assign addr[23791] = -2073814024;
assign addr[23792] = -2078697525;
assign addr[23793] = -2083416198;
assign addr[23794] = -2087969669;
assign addr[23795] = -2092357577;
assign addr[23796] = -2096579573;
assign addr[23797] = -2100635323;
assign addr[23798] = -2104524506;
assign addr[23799] = -2108246813;
assign addr[23800] = -2111801949;
assign addr[23801] = -2115189632;
assign addr[23802] = -2118409593;
assign addr[23803] = -2121461578;
assign addr[23804] = -2124345343;
assign addr[23805] = -2127060661;
assign addr[23806] = -2129607316;
assign addr[23807] = -2131985106;
assign addr[23808] = -2134193842;
assign addr[23809] = -2136233350;
assign addr[23810] = -2138103468;
assign addr[23811] = -2139804048;
assign addr[23812] = -2141334954;
assign addr[23813] = -2142696065;
assign addr[23814] = -2143887273;
assign addr[23815] = -2144908484;
assign addr[23816] = -2145759618;
assign addr[23817] = -2146440605;
assign addr[23818] = -2146951393;
assign addr[23819] = -2147291941;
assign addr[23820] = -2147462221;
assign addr[23821] = -2147462221;
assign addr[23822] = -2147291941;
assign addr[23823] = -2146951393;
assign addr[23824] = -2146440605;
assign addr[23825] = -2145759618;
assign addr[23826] = -2144908484;
assign addr[23827] = -2143887273;
assign addr[23828] = -2142696065;
assign addr[23829] = -2141334954;
assign addr[23830] = -2139804048;
assign addr[23831] = -2138103468;
assign addr[23832] = -2136233350;
assign addr[23833] = -2134193842;
assign addr[23834] = -2131985106;
assign addr[23835] = -2129607316;
assign addr[23836] = -2127060661;
assign addr[23837] = -2124345343;
assign addr[23838] = -2121461578;
assign addr[23839] = -2118409593;
assign addr[23840] = -2115189632;
assign addr[23841] = -2111801949;
assign addr[23842] = -2108246813;
assign addr[23843] = -2104524506;
assign addr[23844] = -2100635323;
assign addr[23845] = -2096579573;
assign addr[23846] = -2092357577;
assign addr[23847] = -2087969669;
assign addr[23848] = -2083416198;
assign addr[23849] = -2078697525;
assign addr[23850] = -2073814024;
assign addr[23851] = -2068766083;
assign addr[23852] = -2063554100;
assign addr[23853] = -2058178491;
assign addr[23854] = -2052639680;
assign addr[23855] = -2046938108;
assign addr[23856] = -2041074226;
assign addr[23857] = -2035048499;
assign addr[23858] = -2028861406;
assign addr[23859] = -2022513436;
assign addr[23860] = -2016005093;
assign addr[23861] = -2009336893;
assign addr[23862] = -2002509365;
assign addr[23863] = -1995523051;
assign addr[23864] = -1988378503;
assign addr[23865] = -1981076290;
assign addr[23866] = -1973616989;
assign addr[23867] = -1966001192;
assign addr[23868] = -1958229503;
assign addr[23869] = -1950302539;
assign addr[23870] = -1942220928;
assign addr[23871] = -1933985310;
assign addr[23872] = -1925596340;
assign addr[23873] = -1917054681;
assign addr[23874] = -1908361011;
assign addr[23875] = -1899516021;
assign addr[23876] = -1890520410;
assign addr[23877] = -1881374892;
assign addr[23878] = -1872080193;
assign addr[23879] = -1862637049;
assign addr[23880] = -1853046210;
assign addr[23881] = -1843308435;
assign addr[23882] = -1833424497;
assign addr[23883] = -1823395180;
assign addr[23884] = -1813221279;
assign addr[23885] = -1802903601;
assign addr[23886] = -1792442963;
assign addr[23887] = -1781840195;
assign addr[23888] = -1771096139;
assign addr[23889] = -1760211645;
assign addr[23890] = -1749187577;
assign addr[23891] = -1738024810;
assign addr[23892] = -1726724227;
assign addr[23893] = -1715286726;
assign addr[23894] = -1703713213;
assign addr[23895] = -1692004606;
assign addr[23896] = -1680161834;
assign addr[23897] = -1668185835;
assign addr[23898] = -1656077559;
assign addr[23899] = -1643837966;
assign addr[23900] = -1631468027;
assign addr[23901] = -1618968722;
assign addr[23902] = -1606341043;
assign addr[23903] = -1593585992;
assign addr[23904] = -1580704578;
assign addr[23905] = -1567697824;
assign addr[23906] = -1554566762;
assign addr[23907] = -1541312431;
assign addr[23908] = -1527935884;
assign addr[23909] = -1514438181;
assign addr[23910] = -1500820393;
assign addr[23911] = -1487083598;
assign addr[23912] = -1473228887;
assign addr[23913] = -1459257358;
assign addr[23914] = -1445170118;
assign addr[23915] = -1430968286;
assign addr[23916] = -1416652986;
assign addr[23917] = -1402225355;
assign addr[23918] = -1387686535;
assign addr[23919] = -1373037681;
assign addr[23920] = -1358279953;
assign addr[23921] = -1343414522;
assign addr[23922] = -1328442566;
assign addr[23923] = -1313365273;
assign addr[23924] = -1298183838;
assign addr[23925] = -1282899464;
assign addr[23926] = -1267513365;
assign addr[23927] = -1252026760;
assign addr[23928] = -1236440877;
assign addr[23929] = -1220756951;
assign addr[23930] = -1204976227;
assign addr[23931] = -1189099956;
assign addr[23932] = -1173129396;
assign addr[23933] = -1157065814;
assign addr[23934] = -1140910484;
assign addr[23935] = -1124664687;
assign addr[23936] = -1108329711;
assign addr[23937] = -1091906851;
assign addr[23938] = -1075397409;
assign addr[23939] = -1058802695;
assign addr[23940] = -1042124025;
assign addr[23941] = -1025362720;
assign addr[23942] = -1008520110;
assign addr[23943] = -991597531;
assign addr[23944] = -974596324;
assign addr[23945] = -957517838;
assign addr[23946] = -940363427;
assign addr[23947] = -923134450;
assign addr[23948] = -905832274;
assign addr[23949] = -888458272;
assign addr[23950] = -871013820;
assign addr[23951] = -853500302;
assign addr[23952] = -835919107;
assign addr[23953] = -818271628;
assign addr[23954] = -800559266;
assign addr[23955] = -782783424;
assign addr[23956] = -764945512;
assign addr[23957] = -747046944;
assign addr[23958] = -729089140;
assign addr[23959] = -711073524;
assign addr[23960] = -693001525;
assign addr[23961] = -674874574;
assign addr[23962] = -656694110;
assign addr[23963] = -638461574;
assign addr[23964] = -620178412;
assign addr[23965] = -601846074;
assign addr[23966] = -583466013;
assign addr[23967] = -565039687;
assign addr[23968] = -546568556;
assign addr[23969] = -528054086;
assign addr[23970] = -509497745;
assign addr[23971] = -490901003;
assign addr[23972] = -472265336;
assign addr[23973] = -453592221;
assign addr[23974] = -434883140;
assign addr[23975] = -416139574;
assign addr[23976] = -397363011;
assign addr[23977] = -378554940;
assign addr[23978] = -359716852;
assign addr[23979] = -340850240;
assign addr[23980] = -321956601;
assign addr[23981] = -303037433;
assign addr[23982] = -284094236;
assign addr[23983] = -265128512;
assign addr[23984] = -246141764;
assign addr[23985] = -227135500;
assign addr[23986] = -208111224;
assign addr[23987] = -189070447;
assign addr[23988] = -170014678;
assign addr[23989] = -150945428;
assign addr[23990] = -131864208;
assign addr[23991] = -112772533;
assign addr[23992] = -93671915;
assign addr[23993] = -74563870;
assign addr[23994] = -55449912;
assign addr[23995] = -36331557;
assign addr[23996] = -17210322;
assign addr[23997] = 1912278;
assign addr[23998] = 21034727;
assign addr[23999] = 40155507;
assign addr[24000] = 59273104;
assign addr[24001] = 78386000;
assign addr[24002] = 97492681;
assign addr[24003] = 116591632;
assign addr[24004] = 135681337;
assign addr[24005] = 154760284;
assign addr[24006] = 173826959;
assign addr[24007] = 192879850;
assign addr[24008] = 211917448;
assign addr[24009] = 230938242;
assign addr[24010] = 249940723;
assign addr[24011] = 268923386;
assign addr[24012] = 287884725;
assign addr[24013] = 306823237;
assign addr[24014] = 325737419;
assign addr[24015] = 344625773;
assign addr[24016] = 363486799;
assign addr[24017] = 382319004;
assign addr[24018] = 401120892;
assign addr[24019] = 419890975;
assign addr[24020] = 438627762;
assign addr[24021] = 457329769;
assign addr[24022] = 475995513;
assign addr[24023] = 494623513;
assign addr[24024] = 513212292;
assign addr[24025] = 531760377;
assign addr[24026] = 550266296;
assign addr[24027] = 568728583;
assign addr[24028] = 587145773;
assign addr[24029] = 605516406;
assign addr[24030] = 623839025;
assign addr[24031] = 642112178;
assign addr[24032] = 660334415;
assign addr[24033] = 678504291;
assign addr[24034] = 696620367;
assign addr[24035] = 714681204;
assign addr[24036] = 732685372;
assign addr[24037] = 750631442;
assign addr[24038] = 768517992;
assign addr[24039] = 786343603;
assign addr[24040] = 804106861;
assign addr[24041] = 821806359;
assign addr[24042] = 839440693;
assign addr[24043] = 857008464;
assign addr[24044] = 874508280;
assign addr[24045] = 891938752;
assign addr[24046] = 909298500;
assign addr[24047] = 926586145;
assign addr[24048] = 943800318;
assign addr[24049] = 960939653;
assign addr[24050] = 978002791;
assign addr[24051] = 994988380;
assign addr[24052] = 1011895073;
assign addr[24053] = 1028721528;
assign addr[24054] = 1045466412;
assign addr[24055] = 1062128397;
assign addr[24056] = 1078706161;
assign addr[24057] = 1095198391;
assign addr[24058] = 1111603778;
assign addr[24059] = 1127921022;
assign addr[24060] = 1144148829;
assign addr[24061] = 1160285911;
assign addr[24062] = 1176330990;
assign addr[24063] = 1192282793;
assign addr[24064] = 1208140056;
assign addr[24065] = 1223901520;
assign addr[24066] = 1239565936;
assign addr[24067] = 1255132063;
assign addr[24068] = 1270598665;
assign addr[24069] = 1285964516;
assign addr[24070] = 1301228398;
assign addr[24071] = 1316389101;
assign addr[24072] = 1331445422;
assign addr[24073] = 1346396168;
assign addr[24074] = 1361240152;
assign addr[24075] = 1375976199;
assign addr[24076] = 1390603139;
assign addr[24077] = 1405119813;
assign addr[24078] = 1419525069;
assign addr[24079] = 1433817766;
assign addr[24080] = 1447996770;
assign addr[24081] = 1462060956;
assign addr[24082] = 1476009210;
assign addr[24083] = 1489840425;
assign addr[24084] = 1503553506;
assign addr[24085] = 1517147363;
assign addr[24086] = 1530620920;
assign addr[24087] = 1543973108;
assign addr[24088] = 1557202869;
assign addr[24089] = 1570309153;
assign addr[24090] = 1583290921;
assign addr[24091] = 1596147143;
assign addr[24092] = 1608876801;
assign addr[24093] = 1621478885;
assign addr[24094] = 1633952396;
assign addr[24095] = 1646296344;
assign addr[24096] = 1658509750;
assign addr[24097] = 1670591647;
assign addr[24098] = 1682541077;
assign addr[24099] = 1694357091;
assign addr[24100] = 1706038753;
assign addr[24101] = 1717585136;
assign addr[24102] = 1728995326;
assign addr[24103] = 1740268417;
assign addr[24104] = 1751403515;
assign addr[24105] = 1762399737;
assign addr[24106] = 1773256212;
assign addr[24107] = 1783972079;
assign addr[24108] = 1794546487;
assign addr[24109] = 1804978599;
assign addr[24110] = 1815267588;
assign addr[24111] = 1825412636;
assign addr[24112] = 1835412941;
assign addr[24113] = 1845267708;
assign addr[24114] = 1854976157;
assign addr[24115] = 1864537518;
assign addr[24116] = 1873951032;
assign addr[24117] = 1883215953;
assign addr[24118] = 1892331547;
assign addr[24119] = 1901297091;
assign addr[24120] = 1910111873;
assign addr[24121] = 1918775195;
assign addr[24122] = 1927286370;
assign addr[24123] = 1935644723;
assign addr[24124] = 1943849591;
assign addr[24125] = 1951900324;
assign addr[24126] = 1959796283;
assign addr[24127] = 1967536842;
assign addr[24128] = 1975121388;
assign addr[24129] = 1982549318;
assign addr[24130] = 1989820044;
assign addr[24131] = 1996932990;
assign addr[24132] = 2003887591;
assign addr[24133] = 2010683297;
assign addr[24134] = 2017319567;
assign addr[24135] = 2023795876;
assign addr[24136] = 2030111710;
assign addr[24137] = 2036266570;
assign addr[24138] = 2042259965;
assign addr[24139] = 2048091422;
assign addr[24140] = 2053760478;
assign addr[24141] = 2059266683;
assign addr[24142] = 2064609600;
assign addr[24143] = 2069788807;
assign addr[24144] = 2074803892;
assign addr[24145] = 2079654458;
assign addr[24146] = 2084340120;
assign addr[24147] = 2088860507;
assign addr[24148] = 2093215260;
assign addr[24149] = 2097404033;
assign addr[24150] = 2101426496;
assign addr[24151] = 2105282327;
assign addr[24152] = 2108971223;
assign addr[24153] = 2112492891;
assign addr[24154] = 2115847050;
assign addr[24155] = 2119033436;
assign addr[24156] = 2122051796;
assign addr[24157] = 2124901890;
assign addr[24158] = 2127583492;
assign addr[24159] = 2130096389;
assign addr[24160] = 2132440383;
assign addr[24161] = 2134615288;
assign addr[24162] = 2136620930;
assign addr[24163] = 2138457152;
assign addr[24164] = 2140123807;
assign addr[24165] = 2141620763;
assign addr[24166] = 2142947902;
assign addr[24167] = 2144105118;
assign addr[24168] = 2145092320;
assign addr[24169] = 2145909429;
assign addr[24170] = 2146556380;
assign addr[24171] = 2147033123;
assign addr[24172] = 2147339619;
assign addr[24173] = 2147475844;
assign addr[24174] = 2147441787;
assign addr[24175] = 2147237452;
assign addr[24176] = 2146862854;
assign addr[24177] = 2146318022;
assign addr[24178] = 2145603001;
assign addr[24179] = 2144717846;
assign addr[24180] = 2143662628;
assign addr[24181] = 2142437431;
assign addr[24182] = 2141042352;
assign addr[24183] = 2139477502;
assign addr[24184] = 2137743003;
assign addr[24185] = 2135838995;
assign addr[24186] = 2133765628;
assign addr[24187] = 2131523066;
assign addr[24188] = 2129111488;
assign addr[24189] = 2126531084;
assign addr[24190] = 2123782059;
assign addr[24191] = 2120864631;
assign addr[24192] = 2117779031;
assign addr[24193] = 2114525505;
assign addr[24194] = 2111104309;
assign addr[24195] = 2107515716;
assign addr[24196] = 2103760010;
assign addr[24197] = 2099837489;
assign addr[24198] = 2095748463;
assign addr[24199] = 2091493257;
assign addr[24200] = 2087072209;
assign addr[24201] = 2082485668;
assign addr[24202] = 2077733999;
assign addr[24203] = 2072817579;
assign addr[24204] = 2067736796;
assign addr[24205] = 2062492055;
assign addr[24206] = 2057083771;
assign addr[24207] = 2051512372;
assign addr[24208] = 2045778302;
assign addr[24209] = 2039882013;
assign addr[24210] = 2033823974;
assign addr[24211] = 2027604666;
assign addr[24212] = 2021224581;
assign addr[24213] = 2014684225;
assign addr[24214] = 2007984117;
assign addr[24215] = 2001124788;
assign addr[24216] = 1994106782;
assign addr[24217] = 1986930656;
assign addr[24218] = 1979596978;
assign addr[24219] = 1972106330;
assign addr[24220] = 1964459306;
assign addr[24221] = 1956656513;
assign addr[24222] = 1948698568;
assign addr[24223] = 1940586104;
assign addr[24224] = 1932319763;
assign addr[24225] = 1923900201;
assign addr[24226] = 1915328086;
assign addr[24227] = 1906604097;
assign addr[24228] = 1897728925;
assign addr[24229] = 1888703276;
assign addr[24230] = 1879527863;
assign addr[24231] = 1870203416;
assign addr[24232] = 1860730673;
assign addr[24233] = 1851110385;
assign addr[24234] = 1841343316;
assign addr[24235] = 1831430239;
assign addr[24236] = 1821371941;
assign addr[24237] = 1811169220;
assign addr[24238] = 1800822883;
assign addr[24239] = 1790333753;
assign addr[24240] = 1779702660;
assign addr[24241] = 1768930447;
assign addr[24242] = 1758017969;
assign addr[24243] = 1746966091;
assign addr[24244] = 1735775690;
assign addr[24245] = 1724447652;
assign addr[24246] = 1712982875;
assign addr[24247] = 1701382270;
assign addr[24248] = 1689646755;
assign addr[24249] = 1677777262;
assign addr[24250] = 1665774731;
assign addr[24251] = 1653640115;
assign addr[24252] = 1641374375;
assign addr[24253] = 1628978484;
assign addr[24254] = 1616453425;
assign addr[24255] = 1603800191;
assign addr[24256] = 1591019785;
assign addr[24257] = 1578113222;
assign addr[24258] = 1565081523;
assign addr[24259] = 1551925723;
assign addr[24260] = 1538646865;
assign addr[24261] = 1525246002;
assign addr[24262] = 1511724196;
assign addr[24263] = 1498082520;
assign addr[24264] = 1484322054;
assign addr[24265] = 1470443891;
assign addr[24266] = 1456449131;
assign addr[24267] = 1442338884;
assign addr[24268] = 1428114267;
assign addr[24269] = 1413776410;
assign addr[24270] = 1399326449;
assign addr[24271] = 1384765530;
assign addr[24272] = 1370094808;
assign addr[24273] = 1355315445;
assign addr[24274] = 1340428615;
assign addr[24275] = 1325435496;
assign addr[24276] = 1310337279;
assign addr[24277] = 1295135159;
assign addr[24278] = 1279830344;
assign addr[24279] = 1264424045;
assign addr[24280] = 1248917486;
assign addr[24281] = 1233311895;
assign addr[24282] = 1217608510;
assign addr[24283] = 1201808576;
assign addr[24284] = 1185913346;
assign addr[24285] = 1169924081;
assign addr[24286] = 1153842047;
assign addr[24287] = 1137668521;
assign addr[24288] = 1121404785;
assign addr[24289] = 1105052128;
assign addr[24290] = 1088611847;
assign addr[24291] = 1072085246;
assign addr[24292] = 1055473635;
assign addr[24293] = 1038778332;
assign addr[24294] = 1022000660;
assign addr[24295] = 1005141949;
assign addr[24296] = 988203537;
assign addr[24297] = 971186766;
assign addr[24298] = 954092986;
assign addr[24299] = 936923553;
assign addr[24300] = 919679827;
assign addr[24301] = 902363176;
assign addr[24302] = 884974973;
assign addr[24303] = 867516597;
assign addr[24304] = 849989433;
assign addr[24305] = 832394869;
assign addr[24306] = 814734301;
assign addr[24307] = 797009130;
assign addr[24308] = 779220762;
assign addr[24309] = 761370605;
assign addr[24310] = 743460077;
assign addr[24311] = 725490597;
assign addr[24312] = 707463589;
assign addr[24313] = 689380485;
assign addr[24314] = 671242716;
assign addr[24315] = 653051723;
assign addr[24316] = 634808946;
assign addr[24317] = 616515832;
assign addr[24318] = 598173833;
assign addr[24319] = 579784402;
assign addr[24320] = 561348998;
assign addr[24321] = 542869083;
assign addr[24322] = 524346121;
assign addr[24323] = 505781581;
assign addr[24324] = 487176937;
assign addr[24325] = 468533662;
assign addr[24326] = 449853235;
assign addr[24327] = 431137138;
assign addr[24328] = 412386854;
assign addr[24329] = 393603870;
assign addr[24330] = 374789676;
assign addr[24331] = 355945764;
assign addr[24332] = 337073627;
assign addr[24333] = 318174762;
assign addr[24334] = 299250668;
assign addr[24335] = 280302845;
assign addr[24336] = 261332796;
assign addr[24337] = 242342025;
assign addr[24338] = 223332037;
assign addr[24339] = 204304341;
assign addr[24340] = 185260444;
assign addr[24341] = 166201858;
assign addr[24342] = 147130093;
assign addr[24343] = 128046661;
assign addr[24344] = 108953076;
assign addr[24345] = 89850852;
assign addr[24346] = 70741503;
assign addr[24347] = 51626544;
assign addr[24348] = 32507492;
assign addr[24349] = 13385863;
assign addr[24350] = -5736829;
assign addr[24351] = -24859065;
assign addr[24352] = -43979330;
assign addr[24353] = -63096108;
assign addr[24354] = -82207882;
assign addr[24355] = -101313138;
assign addr[24356] = -120410361;
assign addr[24357] = -139498035;
assign addr[24358] = -158574649;
assign addr[24359] = -177638688;
assign addr[24360] = -196688642;
assign addr[24361] = -215722999;
assign addr[24362] = -234740251;
assign addr[24363] = -253738890;
assign addr[24364] = -272717408;
assign addr[24365] = -291674302;
assign addr[24366] = -310608068;
assign addr[24367] = -329517204;
assign addr[24368] = -348400212;
assign addr[24369] = -367255594;
assign addr[24370] = -386081854;
assign addr[24371] = -404877501;
assign addr[24372] = -423641043;
assign addr[24373] = -442370993;
assign addr[24374] = -461065866;
assign addr[24375] = -479724180;
assign addr[24376] = -498344454;
assign addr[24377] = -516925212;
assign addr[24378] = -535464981;
assign addr[24379] = -553962291;
assign addr[24380] = -572415676;
assign addr[24381] = -590823671;
assign addr[24382] = -609184818;
assign addr[24383] = -627497660;
assign addr[24384] = -645760745;
assign addr[24385] = -663972625;
assign addr[24386] = -682131857;
assign addr[24387] = -700236999;
assign addr[24388] = -718286617;
assign addr[24389] = -736279279;
assign addr[24390] = -754213559;
assign addr[24391] = -772088034;
assign addr[24392] = -789901288;
assign addr[24393] = -807651907;
assign addr[24394] = -825338484;
assign addr[24395] = -842959617;
assign addr[24396] = -860513908;
assign addr[24397] = -877999966;
assign addr[24398] = -895416404;
assign addr[24399] = -912761841;
assign addr[24400] = -930034901;
assign addr[24401] = -947234215;
assign addr[24402] = -964358420;
assign addr[24403] = -981406156;
assign addr[24404] = -998376073;
assign addr[24405] = -1015266825;
assign addr[24406] = -1032077073;
assign addr[24407] = -1048805483;
assign addr[24408] = -1065450729;
assign addr[24409] = -1082011492;
assign addr[24410] = -1098486458;
assign addr[24411] = -1114874320;
assign addr[24412] = -1131173780;
assign addr[24413] = -1147383544;
assign addr[24414] = -1163502328;
assign addr[24415] = -1179528853;
assign addr[24416] = -1195461849;
assign addr[24417] = -1211300053;
assign addr[24418] = -1227042207;
assign addr[24419] = -1242687064;
assign addr[24420] = -1258233384;
assign addr[24421] = -1273679934;
assign addr[24422] = -1289025489;
assign addr[24423] = -1304268832;
assign addr[24424] = -1319408754;
assign addr[24425] = -1334444055;
assign addr[24426] = -1349373543;
assign addr[24427] = -1364196034;
assign addr[24428] = -1378910353;
assign addr[24429] = -1393515332;
assign addr[24430] = -1408009814;
assign addr[24431] = -1422392650;
assign addr[24432] = -1436662698;
assign addr[24433] = -1450818828;
assign addr[24434] = -1464859917;
assign addr[24435] = -1478784851;
assign addr[24436] = -1492592527;
assign addr[24437] = -1506281850;
assign addr[24438] = -1519851733;
assign addr[24439] = -1533301101;
assign addr[24440] = -1546628888;
assign addr[24441] = -1559834037;
assign addr[24442] = -1572915501;
assign addr[24443] = -1585872242;
assign addr[24444] = -1598703233;
assign addr[24445] = -1611407456;
assign addr[24446] = -1623983905;
assign addr[24447] = -1636431582;
assign addr[24448] = -1648749499;
assign addr[24449] = -1660936681;
assign addr[24450] = -1672992161;
assign addr[24451] = -1684914983;
assign addr[24452] = -1696704201;
assign addr[24453] = -1708358881;
assign addr[24454] = -1719878099;
assign addr[24455] = -1731260941;
assign addr[24456] = -1742506504;
assign addr[24457] = -1753613897;
assign addr[24458] = -1764582240;
assign addr[24459] = -1775410662;
assign addr[24460] = -1786098304;
assign addr[24461] = -1796644320;
assign addr[24462] = -1807047873;
assign addr[24463] = -1817308138;
assign addr[24464] = -1827424302;
assign addr[24465] = -1837395562;
assign addr[24466] = -1847221128;
assign addr[24467] = -1856900221;
assign addr[24468] = -1866432072;
assign addr[24469] = -1875815927;
assign addr[24470] = -1885051042;
assign addr[24471] = -1894136683;
assign addr[24472] = -1903072131;
assign addr[24473] = -1911856677;
assign addr[24474] = -1920489624;
assign addr[24475] = -1928970288;
assign addr[24476] = -1937297997;
assign addr[24477] = -1945472089;
assign addr[24478] = -1953491918;
assign addr[24479] = -1961356847;
assign addr[24480] = -1969066252;
assign addr[24481] = -1976619522;
assign addr[24482] = -1984016058;
assign addr[24483] = -1991255274;
assign addr[24484] = -1998336596;
assign addr[24485] = -2005259462;
assign addr[24486] = -2012023322;
assign addr[24487] = -2018627642;
assign addr[24488] = -2025071897;
assign addr[24489] = -2031355576;
assign addr[24490] = -2037478181;
assign addr[24491] = -2043439226;
assign addr[24492] = -2049238240;
assign addr[24493] = -2054874761;
assign addr[24494] = -2060348343;
assign addr[24495] = -2065658552;
assign addr[24496] = -2070804967;
assign addr[24497] = -2075787180;
assign addr[24498] = -2080604795;
assign addr[24499] = -2085257431;
assign addr[24500] = -2089744719;
assign addr[24501] = -2094066304;
assign addr[24502] = -2098221841;
assign addr[24503] = -2102211002;
assign addr[24504] = -2106033471;
assign addr[24505] = -2109688944;
assign addr[24506] = -2113177132;
assign addr[24507] = -2116497758;
assign addr[24508] = -2119650558;
assign addr[24509] = -2122635283;
assign addr[24510] = -2125451696;
assign addr[24511] = -2128099574;
assign addr[24512] = -2130578706;
assign addr[24513] = -2132888897;
assign addr[24514] = -2135029962;
assign addr[24515] = -2137001733;
assign addr[24516] = -2138804053;
assign addr[24517] = -2140436778;
assign addr[24518] = -2141899780;
assign addr[24519] = -2143192942;
assign addr[24520] = -2144316162;
assign addr[24521] = -2145269351;
assign addr[24522] = -2146052433;
assign addr[24523] = -2146665347;
assign addr[24524] = -2147108043;
assign addr[24525] = -2147380486;
assign addr[24526] = -2147482655;
assign addr[24527] = -2147414542;
assign addr[24528] = -2147176152;
assign addr[24529] = -2146767505;
assign addr[24530] = -2146188631;
assign addr[24531] = -2145439578;
assign addr[24532] = -2144520405;
assign addr[24533] = -2143431184;
assign addr[24534] = -2142172003;
assign addr[24535] = -2140742960;
assign addr[24536] = -2139144169;
assign addr[24537] = -2137375758;
assign addr[24538] = -2135437865;
assign addr[24539] = -2133330646;
assign addr[24540] = -2131054266;
assign addr[24541] = -2128608907;
assign addr[24542] = -2125994762;
assign addr[24543] = -2123212038;
assign addr[24544] = -2120260957;
assign addr[24545] = -2117141752;
assign addr[24546] = -2113854671;
assign addr[24547] = -2110399974;
assign addr[24548] = -2106777935;
assign addr[24549] = -2102988841;
assign addr[24550] = -2099032994;
assign addr[24551] = -2094910706;
assign addr[24552] = -2090622304;
assign addr[24553] = -2086168128;
assign addr[24554] = -2081548533;
assign addr[24555] = -2076763883;
assign addr[24556] = -2071814558;
assign addr[24557] = -2066700952;
assign addr[24558] = -2061423468;
assign addr[24559] = -2055982526;
assign addr[24560] = -2050378558;
assign addr[24561] = -2044612007;
assign addr[24562] = -2038683330;
assign addr[24563] = -2032592999;
assign addr[24564] = -2026341495;
assign addr[24565] = -2019929315;
assign addr[24566] = -2013356967;
assign addr[24567] = -2006624971;
assign addr[24568] = -1999733863;
assign addr[24569] = -1992684188;
assign addr[24570] = -1985476506;
assign addr[24571] = -1978111387;
assign addr[24572] = -1970589416;
assign addr[24573] = -1962911189;
assign addr[24574] = -1955077316;
assign addr[24575] = -1947088417;
assign addr[24576] = -1938945125;
assign addr[24577] = -1930648088;
assign addr[24578] = -1922197961;
assign addr[24579] = -1913595416;
assign addr[24580] = -1904841135;
assign addr[24581] = -1895935811;
assign addr[24582] = -1886880151;
assign addr[24583] = -1877674873;
assign addr[24584] = -1868320707;
assign addr[24585] = -1858818395;
assign addr[24586] = -1849168689;
assign addr[24587] = -1839372356;
assign addr[24588] = -1829430172;
assign addr[24589] = -1819342925;
assign addr[24590] = -1809111415;
assign addr[24591] = -1798736454;
assign addr[24592] = -1788218865;
assign addr[24593] = -1777559480;
assign addr[24594] = -1766759146;
assign addr[24595] = -1755818718;
assign addr[24596] = -1744739065;
assign addr[24597] = -1733521064;
assign addr[24598] = -1722165606;
assign addr[24599] = -1710673591;
assign addr[24600] = -1699045930;
assign addr[24601] = -1687283545;
assign addr[24602] = -1675387369;
assign addr[24603] = -1663358344;
assign addr[24604] = -1651197426;
assign addr[24605] = -1638905577;
assign addr[24606] = -1626483774;
assign addr[24607] = -1613933000;
assign addr[24608] = -1601254251;
assign addr[24609] = -1588448533;
assign addr[24610] = -1575516860;
assign addr[24611] = -1562460258;
assign addr[24612] = -1549279763;
assign addr[24613] = -1535976419;
assign addr[24614] = -1522551282;
assign addr[24615] = -1509005416;
assign addr[24616] = -1495339895;
assign addr[24617] = -1481555802;
assign addr[24618] = -1467654232;
assign addr[24619] = -1453636285;
assign addr[24620] = -1439503074;
assign addr[24621] = -1425255719;
assign addr[24622] = -1410895350;
assign addr[24623] = -1396423105;
assign addr[24624] = -1381840133;
assign addr[24625] = -1367147589;
assign addr[24626] = -1352346639;
assign addr[24627] = -1337438456;
assign addr[24628] = -1322424222;
assign addr[24629] = -1307305128;
assign addr[24630] = -1292082373;
assign addr[24631] = -1276757164;
assign addr[24632] = -1261330715;
assign addr[24633] = -1245804251;
assign addr[24634] = -1230179002;
assign addr[24635] = -1214456207;
assign addr[24636] = -1198637114;
assign addr[24637] = -1182722976;
assign addr[24638] = -1166715055;
assign addr[24639] = -1150614620;
assign addr[24640] = -1134422949;
assign addr[24641] = -1118141326;
assign addr[24642] = -1101771040;
assign addr[24643] = -1085313391;
assign addr[24644] = -1068769683;
assign addr[24645] = -1052141228;
assign addr[24646] = -1035429345;
assign addr[24647] = -1018635358;
assign addr[24648] = -1001760600;
assign addr[24649] = -984806408;
assign addr[24650] = -967774128;
assign addr[24651] = -950665109;
assign addr[24652] = -933480707;
assign addr[24653] = -916222287;
assign addr[24654] = -898891215;
assign addr[24655] = -881488868;
assign addr[24656] = -864016623;
assign addr[24657] = -846475867;
assign addr[24658] = -828867991;
assign addr[24659] = -811194391;
assign addr[24660] = -793456467;
assign addr[24661] = -775655628;
assign addr[24662] = -757793284;
assign addr[24663] = -739870851;
assign addr[24664] = -721889752;
assign addr[24665] = -703851410;
assign addr[24666] = -685757258;
assign addr[24667] = -667608730;
assign addr[24668] = -649407264;
assign addr[24669] = -631154304;
assign addr[24670] = -612851297;
assign addr[24671] = -594499695;
assign addr[24672] = -576100953;
assign addr[24673] = -557656529;
assign addr[24674] = -539167887;
assign addr[24675] = -520636492;
assign addr[24676] = -502063814;
assign addr[24677] = -483451325;
assign addr[24678] = -464800501;
assign addr[24679] = -446112822;
assign addr[24680] = -427389768;
assign addr[24681] = -408632825;
assign addr[24682] = -389843480;
assign addr[24683] = -371023223;
assign addr[24684] = -352173546;
assign addr[24685] = -333295944;
assign addr[24686] = -314391913;
assign addr[24687] = -295462954;
assign addr[24688] = -276510565;
assign addr[24689] = -257536251;
assign addr[24690] = -238541516;
assign addr[24691] = -219527866;
assign addr[24692] = -200496809;
assign addr[24693] = -181449854;
assign addr[24694] = -162388511;
assign addr[24695] = -143314291;
assign addr[24696] = -124228708;
assign addr[24697] = -105133274;
assign addr[24698] = -86029503;
assign addr[24699] = -66918911;
assign addr[24700] = -47803013;
assign addr[24701] = -28683324;
assign addr[24702] = -9561361;
assign addr[24703] = 9561361;
assign addr[24704] = 28683324;
assign addr[24705] = 47803013;
assign addr[24706] = 66918911;
assign addr[24707] = 86029503;
assign addr[24708] = 105133274;
assign addr[24709] = 124228708;
assign addr[24710] = 143314291;
assign addr[24711] = 162388511;
assign addr[24712] = 181449854;
assign addr[24713] = 200496809;
assign addr[24714] = 219527866;
assign addr[24715] = 238541516;
assign addr[24716] = 257536251;
assign addr[24717] = 276510565;
assign addr[24718] = 295462954;
assign addr[24719] = 314391913;
assign addr[24720] = 333295944;
assign addr[24721] = 352173546;
assign addr[24722] = 371023223;
assign addr[24723] = 389843480;
assign addr[24724] = 408632825;
assign addr[24725] = 427389768;
assign addr[24726] = 446112822;
assign addr[24727] = 464800501;
assign addr[24728] = 483451325;
assign addr[24729] = 502063814;
assign addr[24730] = 520636492;
assign addr[24731] = 539167887;
assign addr[24732] = 557656529;
assign addr[24733] = 576100953;
assign addr[24734] = 594499695;
assign addr[24735] = 612851297;
assign addr[24736] = 631154304;
assign addr[24737] = 649407264;
assign addr[24738] = 667608730;
assign addr[24739] = 685757258;
assign addr[24740] = 703851410;
assign addr[24741] = 721889752;
assign addr[24742] = 739870851;
assign addr[24743] = 757793284;
assign addr[24744] = 775655628;
assign addr[24745] = 793456467;
assign addr[24746] = 811194391;
assign addr[24747] = 828867991;
assign addr[24748] = 846475867;
assign addr[24749] = 864016623;
assign addr[24750] = 881488868;
assign addr[24751] = 898891215;
assign addr[24752] = 916222287;
assign addr[24753] = 933480707;
assign addr[24754] = 950665109;
assign addr[24755] = 967774128;
assign addr[24756] = 984806408;
assign addr[24757] = 1001760600;
assign addr[24758] = 1018635358;
assign addr[24759] = 1035429345;
assign addr[24760] = 1052141228;
assign addr[24761] = 1068769683;
assign addr[24762] = 1085313391;
assign addr[24763] = 1101771040;
assign addr[24764] = 1118141326;
assign addr[24765] = 1134422949;
assign addr[24766] = 1150614620;
assign addr[24767] = 1166715055;
assign addr[24768] = 1182722976;
assign addr[24769] = 1198637114;
assign addr[24770] = 1214456207;
assign addr[24771] = 1230179002;
assign addr[24772] = 1245804251;
assign addr[24773] = 1261330715;
assign addr[24774] = 1276757164;
assign addr[24775] = 1292082373;
assign addr[24776] = 1307305128;
assign addr[24777] = 1322424222;
assign addr[24778] = 1337438456;
assign addr[24779] = 1352346639;
assign addr[24780] = 1367147589;
assign addr[24781] = 1381840133;
assign addr[24782] = 1396423105;
assign addr[24783] = 1410895350;
assign addr[24784] = 1425255719;
assign addr[24785] = 1439503074;
assign addr[24786] = 1453636285;
assign addr[24787] = 1467654232;
assign addr[24788] = 1481555802;
assign addr[24789] = 1495339895;
assign addr[24790] = 1509005416;
assign addr[24791] = 1522551282;
assign addr[24792] = 1535976419;
assign addr[24793] = 1549279763;
assign addr[24794] = 1562460258;
assign addr[24795] = 1575516860;
assign addr[24796] = 1588448533;
assign addr[24797] = 1601254251;
assign addr[24798] = 1613933000;
assign addr[24799] = 1626483774;
assign addr[24800] = 1638905577;
assign addr[24801] = 1651197426;
assign addr[24802] = 1663358344;
assign addr[24803] = 1675387369;
assign addr[24804] = 1687283545;
assign addr[24805] = 1699045930;
assign addr[24806] = 1710673591;
assign addr[24807] = 1722165606;
assign addr[24808] = 1733521064;
assign addr[24809] = 1744739065;
assign addr[24810] = 1755818718;
assign addr[24811] = 1766759146;
assign addr[24812] = 1777559480;
assign addr[24813] = 1788218865;
assign addr[24814] = 1798736454;
assign addr[24815] = 1809111415;
assign addr[24816] = 1819342925;
assign addr[24817] = 1829430172;
assign addr[24818] = 1839372356;
assign addr[24819] = 1849168689;
assign addr[24820] = 1858818395;
assign addr[24821] = 1868320707;
assign addr[24822] = 1877674873;
assign addr[24823] = 1886880151;
assign addr[24824] = 1895935811;
assign addr[24825] = 1904841135;
assign addr[24826] = 1913595416;
assign addr[24827] = 1922197961;
assign addr[24828] = 1930648088;
assign addr[24829] = 1938945125;
assign addr[24830] = 1947088417;
assign addr[24831] = 1955077316;
assign addr[24832] = 1962911189;
assign addr[24833] = 1970589416;
assign addr[24834] = 1978111387;
assign addr[24835] = 1985476506;
assign addr[24836] = 1992684188;
assign addr[24837] = 1999733863;
assign addr[24838] = 2006624971;
assign addr[24839] = 2013356967;
assign addr[24840] = 2019929315;
assign addr[24841] = 2026341495;
assign addr[24842] = 2032592999;
assign addr[24843] = 2038683330;
assign addr[24844] = 2044612007;
assign addr[24845] = 2050378558;
assign addr[24846] = 2055982526;
assign addr[24847] = 2061423468;
assign addr[24848] = 2066700952;
assign addr[24849] = 2071814558;
assign addr[24850] = 2076763883;
assign addr[24851] = 2081548533;
assign addr[24852] = 2086168128;
assign addr[24853] = 2090622304;
assign addr[24854] = 2094910706;
assign addr[24855] = 2099032994;
assign addr[24856] = 2102988841;
assign addr[24857] = 2106777935;
assign addr[24858] = 2110399974;
assign addr[24859] = 2113854671;
assign addr[24860] = 2117141752;
assign addr[24861] = 2120260957;
assign addr[24862] = 2123212038;
assign addr[24863] = 2125994762;
assign addr[24864] = 2128608907;
assign addr[24865] = 2131054266;
assign addr[24866] = 2133330646;
assign addr[24867] = 2135437865;
assign addr[24868] = 2137375758;
assign addr[24869] = 2139144169;
assign addr[24870] = 2140742960;
assign addr[24871] = 2142172003;
assign addr[24872] = 2143431184;
assign addr[24873] = 2144520405;
assign addr[24874] = 2145439578;
assign addr[24875] = 2146188631;
assign addr[24876] = 2146767505;
assign addr[24877] = 2147176152;
assign addr[24878] = 2147414542;
assign addr[24879] = 2147482655;
assign addr[24880] = 2147380486;
assign addr[24881] = 2147108043;
assign addr[24882] = 2146665347;
assign addr[24883] = 2146052433;
assign addr[24884] = 2145269351;
assign addr[24885] = 2144316162;
assign addr[24886] = 2143192942;
assign addr[24887] = 2141899780;
assign addr[24888] = 2140436778;
assign addr[24889] = 2138804053;
assign addr[24890] = 2137001733;
assign addr[24891] = 2135029962;
assign addr[24892] = 2132888897;
assign addr[24893] = 2130578706;
assign addr[24894] = 2128099574;
assign addr[24895] = 2125451696;
assign addr[24896] = 2122635283;
assign addr[24897] = 2119650558;
assign addr[24898] = 2116497758;
assign addr[24899] = 2113177132;
assign addr[24900] = 2109688944;
assign addr[24901] = 2106033471;
assign addr[24902] = 2102211002;
assign addr[24903] = 2098221841;
assign addr[24904] = 2094066304;
assign addr[24905] = 2089744719;
assign addr[24906] = 2085257431;
assign addr[24907] = 2080604795;
assign addr[24908] = 2075787180;
assign addr[24909] = 2070804967;
assign addr[24910] = 2065658552;
assign addr[24911] = 2060348343;
assign addr[24912] = 2054874761;
assign addr[24913] = 2049238240;
assign addr[24914] = 2043439226;
assign addr[24915] = 2037478181;
assign addr[24916] = 2031355576;
assign addr[24917] = 2025071897;
assign addr[24918] = 2018627642;
assign addr[24919] = 2012023322;
assign addr[24920] = 2005259462;
assign addr[24921] = 1998336596;
assign addr[24922] = 1991255274;
assign addr[24923] = 1984016058;
assign addr[24924] = 1976619522;
assign addr[24925] = 1969066252;
assign addr[24926] = 1961356847;
assign addr[24927] = 1953491918;
assign addr[24928] = 1945472089;
assign addr[24929] = 1937297997;
assign addr[24930] = 1928970288;
assign addr[24931] = 1920489624;
assign addr[24932] = 1911856677;
assign addr[24933] = 1903072131;
assign addr[24934] = 1894136683;
assign addr[24935] = 1885051042;
assign addr[24936] = 1875815927;
assign addr[24937] = 1866432072;
assign addr[24938] = 1856900221;
assign addr[24939] = 1847221128;
assign addr[24940] = 1837395562;
assign addr[24941] = 1827424302;
assign addr[24942] = 1817308138;
assign addr[24943] = 1807047873;
assign addr[24944] = 1796644320;
assign addr[24945] = 1786098304;
assign addr[24946] = 1775410662;
assign addr[24947] = 1764582240;
assign addr[24948] = 1753613897;
assign addr[24949] = 1742506504;
assign addr[24950] = 1731260941;
assign addr[24951] = 1719878099;
assign addr[24952] = 1708358881;
assign addr[24953] = 1696704201;
assign addr[24954] = 1684914983;
assign addr[24955] = 1672992161;
assign addr[24956] = 1660936681;
assign addr[24957] = 1648749499;
assign addr[24958] = 1636431582;
assign addr[24959] = 1623983905;
assign addr[24960] = 1611407456;
assign addr[24961] = 1598703233;
assign addr[24962] = 1585872242;
assign addr[24963] = 1572915501;
assign addr[24964] = 1559834037;
assign addr[24965] = 1546628888;
assign addr[24966] = 1533301101;
assign addr[24967] = 1519851733;
assign addr[24968] = 1506281850;
assign addr[24969] = 1492592527;
assign addr[24970] = 1478784851;
assign addr[24971] = 1464859917;
assign addr[24972] = 1450818828;
assign addr[24973] = 1436662698;
assign addr[24974] = 1422392650;
assign addr[24975] = 1408009814;
assign addr[24976] = 1393515332;
assign addr[24977] = 1378910353;
assign addr[24978] = 1364196034;
assign addr[24979] = 1349373543;
assign addr[24980] = 1334444055;
assign addr[24981] = 1319408754;
assign addr[24982] = 1304268832;
assign addr[24983] = 1289025489;
assign addr[24984] = 1273679934;
assign addr[24985] = 1258233384;
assign addr[24986] = 1242687064;
assign addr[24987] = 1227042207;
assign addr[24988] = 1211300053;
assign addr[24989] = 1195461849;
assign addr[24990] = 1179528853;
assign addr[24991] = 1163502328;
assign addr[24992] = 1147383544;
assign addr[24993] = 1131173780;
assign addr[24994] = 1114874320;
assign addr[24995] = 1098486458;
assign addr[24996] = 1082011492;
assign addr[24997] = 1065450729;
assign addr[24998] = 1048805483;
assign addr[24999] = 1032077073;
assign addr[25000] = 1015266825;
assign addr[25001] = 998376073;
assign addr[25002] = 981406156;
assign addr[25003] = 964358420;
assign addr[25004] = 947234215;
assign addr[25005] = 930034901;
assign addr[25006] = 912761841;
assign addr[25007] = 895416404;
assign addr[25008] = 877999966;
assign addr[25009] = 860513908;
assign addr[25010] = 842959617;
assign addr[25011] = 825338484;
assign addr[25012] = 807651907;
assign addr[25013] = 789901288;
assign addr[25014] = 772088034;
assign addr[25015] = 754213559;
assign addr[25016] = 736279279;
assign addr[25017] = 718286617;
assign addr[25018] = 700236999;
assign addr[25019] = 682131857;
assign addr[25020] = 663972625;
assign addr[25021] = 645760745;
assign addr[25022] = 627497660;
assign addr[25023] = 609184818;
assign addr[25024] = 590823671;
assign addr[25025] = 572415676;
assign addr[25026] = 553962291;
assign addr[25027] = 535464981;
assign addr[25028] = 516925212;
assign addr[25029] = 498344454;
assign addr[25030] = 479724180;
assign addr[25031] = 461065866;
assign addr[25032] = 442370993;
assign addr[25033] = 423641043;
assign addr[25034] = 404877501;
assign addr[25035] = 386081854;
assign addr[25036] = 367255594;
assign addr[25037] = 348400212;
assign addr[25038] = 329517204;
assign addr[25039] = 310608068;
assign addr[25040] = 291674302;
assign addr[25041] = 272717408;
assign addr[25042] = 253738890;
assign addr[25043] = 234740251;
assign addr[25044] = 215722999;
assign addr[25045] = 196688642;
assign addr[25046] = 177638688;
assign addr[25047] = 158574649;
assign addr[25048] = 139498035;
assign addr[25049] = 120410361;
assign addr[25050] = 101313138;
assign addr[25051] = 82207882;
assign addr[25052] = 63096108;
assign addr[25053] = 43979330;
assign addr[25054] = 24859065;
assign addr[25055] = 5736829;
assign addr[25056] = -13385863;
assign addr[25057] = -32507492;
assign addr[25058] = -51626544;
assign addr[25059] = -70741503;
assign addr[25060] = -89850852;
assign addr[25061] = -108953076;
assign addr[25062] = -128046661;
assign addr[25063] = -147130093;
assign addr[25064] = -166201858;
assign addr[25065] = -185260444;
assign addr[25066] = -204304341;
assign addr[25067] = -223332037;
assign addr[25068] = -242342025;
assign addr[25069] = -261332796;
assign addr[25070] = -280302845;
assign addr[25071] = -299250668;
assign addr[25072] = -318174762;
assign addr[25073] = -337073627;
assign addr[25074] = -355945764;
assign addr[25075] = -374789676;
assign addr[25076] = -393603870;
assign addr[25077] = -412386854;
assign addr[25078] = -431137138;
assign addr[25079] = -449853235;
assign addr[25080] = -468533662;
assign addr[25081] = -487176937;
assign addr[25082] = -505781581;
assign addr[25083] = -524346121;
assign addr[25084] = -542869083;
assign addr[25085] = -561348998;
assign addr[25086] = -579784402;
assign addr[25087] = -598173833;
assign addr[25088] = -616515832;
assign addr[25089] = -634808946;
assign addr[25090] = -653051723;
assign addr[25091] = -671242716;
assign addr[25092] = -689380485;
assign addr[25093] = -707463589;
assign addr[25094] = -725490597;
assign addr[25095] = -743460077;
assign addr[25096] = -761370605;
assign addr[25097] = -779220762;
assign addr[25098] = -797009130;
assign addr[25099] = -814734301;
assign addr[25100] = -832394869;
assign addr[25101] = -849989433;
assign addr[25102] = -867516597;
assign addr[25103] = -884974973;
assign addr[25104] = -902363176;
assign addr[25105] = -919679827;
assign addr[25106] = -936923553;
assign addr[25107] = -954092986;
assign addr[25108] = -971186766;
assign addr[25109] = -988203537;
assign addr[25110] = -1005141949;
assign addr[25111] = -1022000660;
assign addr[25112] = -1038778332;
assign addr[25113] = -1055473635;
assign addr[25114] = -1072085246;
assign addr[25115] = -1088611847;
assign addr[25116] = -1105052128;
assign addr[25117] = -1121404785;
assign addr[25118] = -1137668521;
assign addr[25119] = -1153842047;
assign addr[25120] = -1169924081;
assign addr[25121] = -1185913346;
assign addr[25122] = -1201808576;
assign addr[25123] = -1217608510;
assign addr[25124] = -1233311895;
assign addr[25125] = -1248917486;
assign addr[25126] = -1264424045;
assign addr[25127] = -1279830344;
assign addr[25128] = -1295135159;
assign addr[25129] = -1310337279;
assign addr[25130] = -1325435496;
assign addr[25131] = -1340428615;
assign addr[25132] = -1355315445;
assign addr[25133] = -1370094808;
assign addr[25134] = -1384765530;
assign addr[25135] = -1399326449;
assign addr[25136] = -1413776410;
assign addr[25137] = -1428114267;
assign addr[25138] = -1442338884;
assign addr[25139] = -1456449131;
assign addr[25140] = -1470443891;
assign addr[25141] = -1484322054;
assign addr[25142] = -1498082520;
assign addr[25143] = -1511724196;
assign addr[25144] = -1525246002;
assign addr[25145] = -1538646865;
assign addr[25146] = -1551925723;
assign addr[25147] = -1565081523;
assign addr[25148] = -1578113222;
assign addr[25149] = -1591019785;
assign addr[25150] = -1603800191;
assign addr[25151] = -1616453425;
assign addr[25152] = -1628978484;
assign addr[25153] = -1641374375;
assign addr[25154] = -1653640115;
assign addr[25155] = -1665774731;
assign addr[25156] = -1677777262;
assign addr[25157] = -1689646755;
assign addr[25158] = -1701382270;
assign addr[25159] = -1712982875;
assign addr[25160] = -1724447652;
assign addr[25161] = -1735775690;
assign addr[25162] = -1746966091;
assign addr[25163] = -1758017969;
assign addr[25164] = -1768930447;
assign addr[25165] = -1779702660;
assign addr[25166] = -1790333753;
assign addr[25167] = -1800822883;
assign addr[25168] = -1811169220;
assign addr[25169] = -1821371941;
assign addr[25170] = -1831430239;
assign addr[25171] = -1841343316;
assign addr[25172] = -1851110385;
assign addr[25173] = -1860730673;
assign addr[25174] = -1870203416;
assign addr[25175] = -1879527863;
assign addr[25176] = -1888703276;
assign addr[25177] = -1897728925;
assign addr[25178] = -1906604097;
assign addr[25179] = -1915328086;
assign addr[25180] = -1923900201;
assign addr[25181] = -1932319763;
assign addr[25182] = -1940586104;
assign addr[25183] = -1948698568;
assign addr[25184] = -1956656513;
assign addr[25185] = -1964459306;
assign addr[25186] = -1972106330;
assign addr[25187] = -1979596978;
assign addr[25188] = -1986930656;
assign addr[25189] = -1994106782;
assign addr[25190] = -2001124788;
assign addr[25191] = -2007984117;
assign addr[25192] = -2014684225;
assign addr[25193] = -2021224581;
assign addr[25194] = -2027604666;
assign addr[25195] = -2033823974;
assign addr[25196] = -2039882013;
assign addr[25197] = -2045778302;
assign addr[25198] = -2051512372;
assign addr[25199] = -2057083771;
assign addr[25200] = -2062492055;
assign addr[25201] = -2067736796;
assign addr[25202] = -2072817579;
assign addr[25203] = -2077733999;
assign addr[25204] = -2082485668;
assign addr[25205] = -2087072209;
assign addr[25206] = -2091493257;
assign addr[25207] = -2095748463;
assign addr[25208] = -2099837489;
assign addr[25209] = -2103760010;
assign addr[25210] = -2107515716;
assign addr[25211] = -2111104309;
assign addr[25212] = -2114525505;
assign addr[25213] = -2117779031;
assign addr[25214] = -2120864631;
assign addr[25215] = -2123782059;
assign addr[25216] = -2126531084;
assign addr[25217] = -2129111488;
assign addr[25218] = -2131523066;
assign addr[25219] = -2133765628;
assign addr[25220] = -2135838995;
assign addr[25221] = -2137743003;
assign addr[25222] = -2139477502;
assign addr[25223] = -2141042352;
assign addr[25224] = -2142437431;
assign addr[25225] = -2143662628;
assign addr[25226] = -2144717846;
assign addr[25227] = -2145603001;
assign addr[25228] = -2146318022;
assign addr[25229] = -2146862854;
assign addr[25230] = -2147237452;
assign addr[25231] = -2147441787;
assign addr[25232] = -2147475844;
assign addr[25233] = -2147339619;
assign addr[25234] = -2147033123;
assign addr[25235] = -2146556380;
assign addr[25236] = -2145909429;
assign addr[25237] = -2145092320;
assign addr[25238] = -2144105118;
assign addr[25239] = -2142947902;
assign addr[25240] = -2141620763;
assign addr[25241] = -2140123807;
assign addr[25242] = -2138457152;
assign addr[25243] = -2136620930;
assign addr[25244] = -2134615288;
assign addr[25245] = -2132440383;
assign addr[25246] = -2130096389;
assign addr[25247] = -2127583492;
assign addr[25248] = -2124901890;
assign addr[25249] = -2122051796;
assign addr[25250] = -2119033436;
assign addr[25251] = -2115847050;
assign addr[25252] = -2112492891;
assign addr[25253] = -2108971223;
assign addr[25254] = -2105282327;
assign addr[25255] = -2101426496;
assign addr[25256] = -2097404033;
assign addr[25257] = -2093215260;
assign addr[25258] = -2088860507;
assign addr[25259] = -2084340120;
assign addr[25260] = -2079654458;
assign addr[25261] = -2074803892;
assign addr[25262] = -2069788807;
assign addr[25263] = -2064609600;
assign addr[25264] = -2059266683;
assign addr[25265] = -2053760478;
assign addr[25266] = -2048091422;
assign addr[25267] = -2042259965;
assign addr[25268] = -2036266570;
assign addr[25269] = -2030111710;
assign addr[25270] = -2023795876;
assign addr[25271] = -2017319567;
assign addr[25272] = -2010683297;
assign addr[25273] = -2003887591;
assign addr[25274] = -1996932990;
assign addr[25275] = -1989820044;
assign addr[25276] = -1982549318;
assign addr[25277] = -1975121388;
assign addr[25278] = -1967536842;
assign addr[25279] = -1959796283;
assign addr[25280] = -1951900324;
assign addr[25281] = -1943849591;
assign addr[25282] = -1935644723;
assign addr[25283] = -1927286370;
assign addr[25284] = -1918775195;
assign addr[25285] = -1910111873;
assign addr[25286] = -1901297091;
assign addr[25287] = -1892331547;
assign addr[25288] = -1883215953;
assign addr[25289] = -1873951032;
assign addr[25290] = -1864537518;
assign addr[25291] = -1854976157;
assign addr[25292] = -1845267708;
assign addr[25293] = -1835412941;
assign addr[25294] = -1825412636;
assign addr[25295] = -1815267588;
assign addr[25296] = -1804978599;
assign addr[25297] = -1794546487;
assign addr[25298] = -1783972079;
assign addr[25299] = -1773256212;
assign addr[25300] = -1762399737;
assign addr[25301] = -1751403515;
assign addr[25302] = -1740268417;
assign addr[25303] = -1728995326;
assign addr[25304] = -1717585136;
assign addr[25305] = -1706038753;
assign addr[25306] = -1694357091;
assign addr[25307] = -1682541077;
assign addr[25308] = -1670591647;
assign addr[25309] = -1658509750;
assign addr[25310] = -1646296344;
assign addr[25311] = -1633952396;
assign addr[25312] = -1621478885;
assign addr[25313] = -1608876801;
assign addr[25314] = -1596147143;
assign addr[25315] = -1583290921;
assign addr[25316] = -1570309153;
assign addr[25317] = -1557202869;
assign addr[25318] = -1543973108;
assign addr[25319] = -1530620920;
assign addr[25320] = -1517147363;
assign addr[25321] = -1503553506;
assign addr[25322] = -1489840425;
assign addr[25323] = -1476009210;
assign addr[25324] = -1462060956;
assign addr[25325] = -1447996770;
assign addr[25326] = -1433817766;
assign addr[25327] = -1419525069;
assign addr[25328] = -1405119813;
assign addr[25329] = -1390603139;
assign addr[25330] = -1375976199;
assign addr[25331] = -1361240152;
assign addr[25332] = -1346396168;
assign addr[25333] = -1331445422;
assign addr[25334] = -1316389101;
assign addr[25335] = -1301228398;
assign addr[25336] = -1285964516;
assign addr[25337] = -1270598665;
assign addr[25338] = -1255132063;
assign addr[25339] = -1239565936;
assign addr[25340] = -1223901520;
assign addr[25341] = -1208140056;
assign addr[25342] = -1192282793;
assign addr[25343] = -1176330990;
assign addr[25344] = -1160285911;
assign addr[25345] = -1144148829;
assign addr[25346] = -1127921022;
assign addr[25347] = -1111603778;
assign addr[25348] = -1095198391;
assign addr[25349] = -1078706161;
assign addr[25350] = -1062128397;
assign addr[25351] = -1045466412;
assign addr[25352] = -1028721528;
assign addr[25353] = -1011895073;
assign addr[25354] = -994988380;
assign addr[25355] = -978002791;
assign addr[25356] = -960939653;
assign addr[25357] = -943800318;
assign addr[25358] = -926586145;
assign addr[25359] = -909298500;
assign addr[25360] = -891938752;
assign addr[25361] = -874508280;
assign addr[25362] = -857008464;
assign addr[25363] = -839440693;
assign addr[25364] = -821806359;
assign addr[25365] = -804106861;
assign addr[25366] = -786343603;
assign addr[25367] = -768517992;
assign addr[25368] = -750631442;
assign addr[25369] = -732685372;
assign addr[25370] = -714681204;
assign addr[25371] = -696620367;
assign addr[25372] = -678504291;
assign addr[25373] = -660334415;
assign addr[25374] = -642112178;
assign addr[25375] = -623839025;
assign addr[25376] = -605516406;
assign addr[25377] = -587145773;
assign addr[25378] = -568728583;
assign addr[25379] = -550266296;
assign addr[25380] = -531760377;
assign addr[25381] = -513212292;
assign addr[25382] = -494623513;
assign addr[25383] = -475995513;
assign addr[25384] = -457329769;
assign addr[25385] = -438627762;
assign addr[25386] = -419890975;
assign addr[25387] = -401120892;
assign addr[25388] = -382319004;
assign addr[25389] = -363486799;
assign addr[25390] = -344625773;
assign addr[25391] = -325737419;
assign addr[25392] = -306823237;
assign addr[25393] = -287884725;
assign addr[25394] = -268923386;
assign addr[25395] = -249940723;
assign addr[25396] = -230938242;
assign addr[25397] = -211917448;
assign addr[25398] = -192879850;
assign addr[25399] = -173826959;
assign addr[25400] = -154760284;
assign addr[25401] = -135681337;
assign addr[25402] = -116591632;
assign addr[25403] = -97492681;
assign addr[25404] = -78386000;
assign addr[25405] = -59273104;
assign addr[25406] = -40155507;
assign addr[25407] = -21034727;
assign addr[25408] = -1912278;
assign addr[25409] = 17210322;
assign addr[25410] = 36331557;
assign addr[25411] = 55449912;
assign addr[25412] = 74563870;
assign addr[25413] = 93671915;
assign addr[25414] = 112772533;
assign addr[25415] = 131864208;
assign addr[25416] = 150945428;
assign addr[25417] = 170014678;
assign addr[25418] = 189070447;
assign addr[25419] = 208111224;
assign addr[25420] = 227135500;
assign addr[25421] = 246141764;
assign addr[25422] = 265128512;
assign addr[25423] = 284094236;
assign addr[25424] = 303037433;
assign addr[25425] = 321956601;
assign addr[25426] = 340850240;
assign addr[25427] = 359716852;
assign addr[25428] = 378554940;
assign addr[25429] = 397363011;
assign addr[25430] = 416139574;
assign addr[25431] = 434883140;
assign addr[25432] = 453592221;
assign addr[25433] = 472265336;
assign addr[25434] = 490901003;
assign addr[25435] = 509497745;
assign addr[25436] = 528054086;
assign addr[25437] = 546568556;
assign addr[25438] = 565039687;
assign addr[25439] = 583466013;
assign addr[25440] = 601846074;
assign addr[25441] = 620178412;
assign addr[25442] = 638461574;
assign addr[25443] = 656694110;
assign addr[25444] = 674874574;
assign addr[25445] = 693001525;
assign addr[25446] = 711073524;
assign addr[25447] = 729089140;
assign addr[25448] = 747046944;
assign addr[25449] = 764945512;
assign addr[25450] = 782783424;
assign addr[25451] = 800559266;
assign addr[25452] = 818271628;
assign addr[25453] = 835919107;
assign addr[25454] = 853500302;
assign addr[25455] = 871013820;
assign addr[25456] = 888458272;
assign addr[25457] = 905832274;
assign addr[25458] = 923134450;
assign addr[25459] = 940363427;
assign addr[25460] = 957517838;
assign addr[25461] = 974596324;
assign addr[25462] = 991597531;
assign addr[25463] = 1008520110;
assign addr[25464] = 1025362720;
assign addr[25465] = 1042124025;
assign addr[25466] = 1058802695;
assign addr[25467] = 1075397409;
assign addr[25468] = 1091906851;
assign addr[25469] = 1108329711;
assign addr[25470] = 1124664687;
assign addr[25471] = 1140910484;
assign addr[25472] = 1157065814;
assign addr[25473] = 1173129396;
assign addr[25474] = 1189099956;
assign addr[25475] = 1204976227;
assign addr[25476] = 1220756951;
assign addr[25477] = 1236440877;
assign addr[25478] = 1252026760;
assign addr[25479] = 1267513365;
assign addr[25480] = 1282899464;
assign addr[25481] = 1298183838;
assign addr[25482] = 1313365273;
assign addr[25483] = 1328442566;
assign addr[25484] = 1343414522;
assign addr[25485] = 1358279953;
assign addr[25486] = 1373037681;
assign addr[25487] = 1387686535;
assign addr[25488] = 1402225355;
assign addr[25489] = 1416652986;
assign addr[25490] = 1430968286;
assign addr[25491] = 1445170118;
assign addr[25492] = 1459257358;
assign addr[25493] = 1473228887;
assign addr[25494] = 1487083598;
assign addr[25495] = 1500820393;
assign addr[25496] = 1514438181;
assign addr[25497] = 1527935884;
assign addr[25498] = 1541312431;
assign addr[25499] = 1554566762;
assign addr[25500] = 1567697824;
assign addr[25501] = 1580704578;
assign addr[25502] = 1593585992;
assign addr[25503] = 1606341043;
assign addr[25504] = 1618968722;
assign addr[25505] = 1631468027;
assign addr[25506] = 1643837966;
assign addr[25507] = 1656077559;
assign addr[25508] = 1668185835;
assign addr[25509] = 1680161834;
assign addr[25510] = 1692004606;
assign addr[25511] = 1703713213;
assign addr[25512] = 1715286726;
assign addr[25513] = 1726724227;
assign addr[25514] = 1738024810;
assign addr[25515] = 1749187577;
assign addr[25516] = 1760211645;
assign addr[25517] = 1771096139;
assign addr[25518] = 1781840195;
assign addr[25519] = 1792442963;
assign addr[25520] = 1802903601;
assign addr[25521] = 1813221279;
assign addr[25522] = 1823395180;
assign addr[25523] = 1833424497;
assign addr[25524] = 1843308435;
assign addr[25525] = 1853046210;
assign addr[25526] = 1862637049;
assign addr[25527] = 1872080193;
assign addr[25528] = 1881374892;
assign addr[25529] = 1890520410;
assign addr[25530] = 1899516021;
assign addr[25531] = 1908361011;
assign addr[25532] = 1917054681;
assign addr[25533] = 1925596340;
assign addr[25534] = 1933985310;
assign addr[25535] = 1942220928;
assign addr[25536] = 1950302539;
assign addr[25537] = 1958229503;
assign addr[25538] = 1966001192;
assign addr[25539] = 1973616989;
assign addr[25540] = 1981076290;
assign addr[25541] = 1988378503;
assign addr[25542] = 1995523051;
assign addr[25543] = 2002509365;
assign addr[25544] = 2009336893;
assign addr[25545] = 2016005093;
assign addr[25546] = 2022513436;
assign addr[25547] = 2028861406;
assign addr[25548] = 2035048499;
assign addr[25549] = 2041074226;
assign addr[25550] = 2046938108;
assign addr[25551] = 2052639680;
assign addr[25552] = 2058178491;
assign addr[25553] = 2063554100;
assign addr[25554] = 2068766083;
assign addr[25555] = 2073814024;
assign addr[25556] = 2078697525;
assign addr[25557] = 2083416198;
assign addr[25558] = 2087969669;
assign addr[25559] = 2092357577;
assign addr[25560] = 2096579573;
assign addr[25561] = 2100635323;
assign addr[25562] = 2104524506;
assign addr[25563] = 2108246813;
assign addr[25564] = 2111801949;
assign addr[25565] = 2115189632;
assign addr[25566] = 2118409593;
assign addr[25567] = 2121461578;
assign addr[25568] = 2124345343;
assign addr[25569] = 2127060661;
assign addr[25570] = 2129607316;
assign addr[25571] = 2131985106;
assign addr[25572] = 2134193842;
assign addr[25573] = 2136233350;
assign addr[25574] = 2138103468;
assign addr[25575] = 2139804048;
assign addr[25576] = 2141334954;
assign addr[25577] = 2142696065;
assign addr[25578] = 2143887273;
assign addr[25579] = 2144908484;
assign addr[25580] = 2145759618;
assign addr[25581] = 2146440605;
assign addr[25582] = 2146951393;
assign addr[25583] = 2147291941;
assign addr[25584] = 2147462221;
assign addr[25585] = 2147462221;
assign addr[25586] = 2147291941;
assign addr[25587] = 2146951393;
assign addr[25588] = 2146440605;
assign addr[25589] = 2145759618;
assign addr[25590] = 2144908484;
assign addr[25591] = 2143887273;
assign addr[25592] = 2142696065;
assign addr[25593] = 2141334954;
assign addr[25594] = 2139804048;
assign addr[25595] = 2138103468;
assign addr[25596] = 2136233350;
assign addr[25597] = 2134193842;
assign addr[25598] = 2131985106;
assign addr[25599] = 2129607316;
assign addr[25600] = 2127060661;
assign addr[25601] = 2124345343;
assign addr[25602] = 2121461578;
assign addr[25603] = 2118409593;
assign addr[25604] = 2115189632;
assign addr[25605] = 2111801949;
assign addr[25606] = 2108246813;
assign addr[25607] = 2104524506;
assign addr[25608] = 2100635323;
assign addr[25609] = 2096579573;
assign addr[25610] = 2092357577;
assign addr[25611] = 2087969669;
assign addr[25612] = 2083416198;
assign addr[25613] = 2078697525;
assign addr[25614] = 2073814024;
assign addr[25615] = 2068766083;
assign addr[25616] = 2063554100;
assign addr[25617] = 2058178491;
assign addr[25618] = 2052639680;
assign addr[25619] = 2046938108;
assign addr[25620] = 2041074226;
assign addr[25621] = 2035048499;
assign addr[25622] = 2028861406;
assign addr[25623] = 2022513436;
assign addr[25624] = 2016005093;
assign addr[25625] = 2009336893;
assign addr[25626] = 2002509365;
assign addr[25627] = 1995523051;
assign addr[25628] = 1988378503;
assign addr[25629] = 1981076290;
assign addr[25630] = 1973616989;
assign addr[25631] = 1966001192;
assign addr[25632] = 1958229503;
assign addr[25633] = 1950302539;
assign addr[25634] = 1942220928;
assign addr[25635] = 1933985310;
assign addr[25636] = 1925596340;
assign addr[25637] = 1917054681;
assign addr[25638] = 1908361011;
assign addr[25639] = 1899516021;
assign addr[25640] = 1890520410;
assign addr[25641] = 1881374892;
assign addr[25642] = 1872080193;
assign addr[25643] = 1862637049;
assign addr[25644] = 1853046210;
assign addr[25645] = 1843308435;
assign addr[25646] = 1833424497;
assign addr[25647] = 1823395180;
assign addr[25648] = 1813221279;
assign addr[25649] = 1802903601;
assign addr[25650] = 1792442963;
assign addr[25651] = 1781840195;
assign addr[25652] = 1771096139;
assign addr[25653] = 1760211645;
assign addr[25654] = 1749187577;
assign addr[25655] = 1738024810;
assign addr[25656] = 1726724227;
assign addr[25657] = 1715286726;
assign addr[25658] = 1703713213;
assign addr[25659] = 1692004606;
assign addr[25660] = 1680161834;
assign addr[25661] = 1668185835;
assign addr[25662] = 1656077559;
assign addr[25663] = 1643837966;
assign addr[25664] = 1631468027;
assign addr[25665] = 1618968722;
assign addr[25666] = 1606341043;
assign addr[25667] = 1593585992;
assign addr[25668] = 1580704578;
assign addr[25669] = 1567697824;
assign addr[25670] = 1554566762;
assign addr[25671] = 1541312431;
assign addr[25672] = 1527935884;
assign addr[25673] = 1514438181;
assign addr[25674] = 1500820393;
assign addr[25675] = 1487083598;
assign addr[25676] = 1473228887;
assign addr[25677] = 1459257358;
assign addr[25678] = 1445170118;
assign addr[25679] = 1430968286;
assign addr[25680] = 1416652986;
assign addr[25681] = 1402225355;
assign addr[25682] = 1387686535;
assign addr[25683] = 1373037681;
assign addr[25684] = 1358279953;
assign addr[25685] = 1343414522;
assign addr[25686] = 1328442566;
assign addr[25687] = 1313365273;
assign addr[25688] = 1298183838;
assign addr[25689] = 1282899464;
assign addr[25690] = 1267513365;
assign addr[25691] = 1252026760;
assign addr[25692] = 1236440877;
assign addr[25693] = 1220756951;
assign addr[25694] = 1204976227;
assign addr[25695] = 1189099956;
assign addr[25696] = 1173129396;
assign addr[25697] = 1157065814;
assign addr[25698] = 1140910484;
assign addr[25699] = 1124664687;
assign addr[25700] = 1108329711;
assign addr[25701] = 1091906851;
assign addr[25702] = 1075397409;
assign addr[25703] = 1058802695;
assign addr[25704] = 1042124025;
assign addr[25705] = 1025362720;
assign addr[25706] = 1008520110;
assign addr[25707] = 991597531;
assign addr[25708] = 974596324;
assign addr[25709] = 957517838;
assign addr[25710] = 940363427;
assign addr[25711] = 923134450;
assign addr[25712] = 905832274;
assign addr[25713] = 888458272;
assign addr[25714] = 871013820;
assign addr[25715] = 853500302;
assign addr[25716] = 835919107;
assign addr[25717] = 818271628;
assign addr[25718] = 800559266;
assign addr[25719] = 782783424;
assign addr[25720] = 764945512;
assign addr[25721] = 747046944;
assign addr[25722] = 729089140;
assign addr[25723] = 711073524;
assign addr[25724] = 693001525;
assign addr[25725] = 674874574;
assign addr[25726] = 656694110;
assign addr[25727] = 638461574;
assign addr[25728] = 620178412;
assign addr[25729] = 601846074;
assign addr[25730] = 583466013;
assign addr[25731] = 565039687;
assign addr[25732] = 546568556;
assign addr[25733] = 528054086;
assign addr[25734] = 509497745;
assign addr[25735] = 490901003;
assign addr[25736] = 472265336;
assign addr[25737] = 453592221;
assign addr[25738] = 434883140;
assign addr[25739] = 416139574;
assign addr[25740] = 397363011;
assign addr[25741] = 378554940;
assign addr[25742] = 359716852;
assign addr[25743] = 340850240;
assign addr[25744] = 321956601;
assign addr[25745] = 303037433;
assign addr[25746] = 284094236;
assign addr[25747] = 265128512;
assign addr[25748] = 246141764;
assign addr[25749] = 227135500;
assign addr[25750] = 208111224;
assign addr[25751] = 189070447;
assign addr[25752] = 170014678;
assign addr[25753] = 150945428;
assign addr[25754] = 131864208;
assign addr[25755] = 112772533;
assign addr[25756] = 93671915;
assign addr[25757] = 74563870;
assign addr[25758] = 55449912;
assign addr[25759] = 36331557;
assign addr[25760] = 17210322;
assign addr[25761] = -1912278;
assign addr[25762] = -21034727;
assign addr[25763] = -40155507;
assign addr[25764] = -59273104;
assign addr[25765] = -78386000;
assign addr[25766] = -97492681;
assign addr[25767] = -116591632;
assign addr[25768] = -135681337;
assign addr[25769] = -154760284;
assign addr[25770] = -173826959;
assign addr[25771] = -192879850;
assign addr[25772] = -211917448;
assign addr[25773] = -230938242;
assign addr[25774] = -249940723;
assign addr[25775] = -268923386;
assign addr[25776] = -287884725;
assign addr[25777] = -306823237;
assign addr[25778] = -325737419;
assign addr[25779] = -344625773;
assign addr[25780] = -363486799;
assign addr[25781] = -382319004;
assign addr[25782] = -401120892;
assign addr[25783] = -419890975;
assign addr[25784] = -438627762;
assign addr[25785] = -457329769;
assign addr[25786] = -475995513;
assign addr[25787] = -494623513;
assign addr[25788] = -513212292;
assign addr[25789] = -531760377;
assign addr[25790] = -550266296;
assign addr[25791] = -568728583;
assign addr[25792] = -587145773;
assign addr[25793] = -605516406;
assign addr[25794] = -623839025;
assign addr[25795] = -642112178;
assign addr[25796] = -660334415;
assign addr[25797] = -678504291;
assign addr[25798] = -696620367;
assign addr[25799] = -714681204;
assign addr[25800] = -732685372;
assign addr[25801] = -750631442;
assign addr[25802] = -768517992;
assign addr[25803] = -786343603;
assign addr[25804] = -804106861;
assign addr[25805] = -821806359;
assign addr[25806] = -839440693;
assign addr[25807] = -857008464;
assign addr[25808] = -874508280;
assign addr[25809] = -891938752;
assign addr[25810] = -909298500;
assign addr[25811] = -926586145;
assign addr[25812] = -943800318;
assign addr[25813] = -960939653;
assign addr[25814] = -978002791;
assign addr[25815] = -994988380;
assign addr[25816] = -1011895073;
assign addr[25817] = -1028721528;
assign addr[25818] = -1045466412;
assign addr[25819] = -1062128397;
assign addr[25820] = -1078706161;
assign addr[25821] = -1095198391;
assign addr[25822] = -1111603778;
assign addr[25823] = -1127921022;
assign addr[25824] = -1144148829;
assign addr[25825] = -1160285911;
assign addr[25826] = -1176330990;
assign addr[25827] = -1192282793;
assign addr[25828] = -1208140056;
assign addr[25829] = -1223901520;
assign addr[25830] = -1239565936;
assign addr[25831] = -1255132063;
assign addr[25832] = -1270598665;
assign addr[25833] = -1285964516;
assign addr[25834] = -1301228398;
assign addr[25835] = -1316389101;
assign addr[25836] = -1331445422;
assign addr[25837] = -1346396168;
assign addr[25838] = -1361240152;
assign addr[25839] = -1375976199;
assign addr[25840] = -1390603139;
assign addr[25841] = -1405119813;
assign addr[25842] = -1419525069;
assign addr[25843] = -1433817766;
assign addr[25844] = -1447996770;
assign addr[25845] = -1462060956;
assign addr[25846] = -1476009210;
assign addr[25847] = -1489840425;
assign addr[25848] = -1503553506;
assign addr[25849] = -1517147363;
assign addr[25850] = -1530620920;
assign addr[25851] = -1543973108;
assign addr[25852] = -1557202869;
assign addr[25853] = -1570309153;
assign addr[25854] = -1583290921;
assign addr[25855] = -1596147143;
assign addr[25856] = -1608876801;
assign addr[25857] = -1621478885;
assign addr[25858] = -1633952396;
assign addr[25859] = -1646296344;
assign addr[25860] = -1658509750;
assign addr[25861] = -1670591647;
assign addr[25862] = -1682541077;
assign addr[25863] = -1694357091;
assign addr[25864] = -1706038753;
assign addr[25865] = -1717585136;
assign addr[25866] = -1728995326;
assign addr[25867] = -1740268417;
assign addr[25868] = -1751403515;
assign addr[25869] = -1762399737;
assign addr[25870] = -1773256212;
assign addr[25871] = -1783972079;
assign addr[25872] = -1794546487;
assign addr[25873] = -1804978599;
assign addr[25874] = -1815267588;
assign addr[25875] = -1825412636;
assign addr[25876] = -1835412941;
assign addr[25877] = -1845267708;
assign addr[25878] = -1854976157;
assign addr[25879] = -1864537518;
assign addr[25880] = -1873951032;
assign addr[25881] = -1883215953;
assign addr[25882] = -1892331547;
assign addr[25883] = -1901297091;
assign addr[25884] = -1910111873;
assign addr[25885] = -1918775195;
assign addr[25886] = -1927286370;
assign addr[25887] = -1935644723;
assign addr[25888] = -1943849591;
assign addr[25889] = -1951900324;
assign addr[25890] = -1959796283;
assign addr[25891] = -1967536842;
assign addr[25892] = -1975121388;
assign addr[25893] = -1982549318;
assign addr[25894] = -1989820044;
assign addr[25895] = -1996932990;
assign addr[25896] = -2003887591;
assign addr[25897] = -2010683297;
assign addr[25898] = -2017319567;
assign addr[25899] = -2023795876;
assign addr[25900] = -2030111710;
assign addr[25901] = -2036266570;
assign addr[25902] = -2042259965;
assign addr[25903] = -2048091422;
assign addr[25904] = -2053760478;
assign addr[25905] = -2059266683;
assign addr[25906] = -2064609600;
assign addr[25907] = -2069788807;
assign addr[25908] = -2074803892;
assign addr[25909] = -2079654458;
assign addr[25910] = -2084340120;
assign addr[25911] = -2088860507;
assign addr[25912] = -2093215260;
assign addr[25913] = -2097404033;
assign addr[25914] = -2101426496;
assign addr[25915] = -2105282327;
assign addr[25916] = -2108971223;
assign addr[25917] = -2112492891;
assign addr[25918] = -2115847050;
assign addr[25919] = -2119033436;
assign addr[25920] = -2122051796;
assign addr[25921] = -2124901890;
assign addr[25922] = -2127583492;
assign addr[25923] = -2130096389;
assign addr[25924] = -2132440383;
assign addr[25925] = -2134615288;
assign addr[25926] = -2136620930;
assign addr[25927] = -2138457152;
assign addr[25928] = -2140123807;
assign addr[25929] = -2141620763;
assign addr[25930] = -2142947902;
assign addr[25931] = -2144105118;
assign addr[25932] = -2145092320;
assign addr[25933] = -2145909429;
assign addr[25934] = -2146556380;
assign addr[25935] = -2147033123;
assign addr[25936] = -2147339619;
assign addr[25937] = -2147475844;
assign addr[25938] = -2147441787;
assign addr[25939] = -2147237452;
assign addr[25940] = -2146862854;
assign addr[25941] = -2146318022;
assign addr[25942] = -2145603001;
assign addr[25943] = -2144717846;
assign addr[25944] = -2143662628;
assign addr[25945] = -2142437431;
assign addr[25946] = -2141042352;
assign addr[25947] = -2139477502;
assign addr[25948] = -2137743003;
assign addr[25949] = -2135838995;
assign addr[25950] = -2133765628;
assign addr[25951] = -2131523066;
assign addr[25952] = -2129111488;
assign addr[25953] = -2126531084;
assign addr[25954] = -2123782059;
assign addr[25955] = -2120864631;
assign addr[25956] = -2117779031;
assign addr[25957] = -2114525505;
assign addr[25958] = -2111104309;
assign addr[25959] = -2107515716;
assign addr[25960] = -2103760010;
assign addr[25961] = -2099837489;
assign addr[25962] = -2095748463;
assign addr[25963] = -2091493257;
assign addr[25964] = -2087072209;
assign addr[25965] = -2082485668;
assign addr[25966] = -2077733999;
assign addr[25967] = -2072817579;
assign addr[25968] = -2067736796;
assign addr[25969] = -2062492055;
assign addr[25970] = -2057083771;
assign addr[25971] = -2051512372;
assign addr[25972] = -2045778302;
assign addr[25973] = -2039882013;
assign addr[25974] = -2033823974;
assign addr[25975] = -2027604666;
assign addr[25976] = -2021224581;
assign addr[25977] = -2014684225;
assign addr[25978] = -2007984117;
assign addr[25979] = -2001124788;
assign addr[25980] = -1994106782;
assign addr[25981] = -1986930656;
assign addr[25982] = -1979596978;
assign addr[25983] = -1972106330;
assign addr[25984] = -1964459306;
assign addr[25985] = -1956656513;
assign addr[25986] = -1948698568;
assign addr[25987] = -1940586104;
assign addr[25988] = -1932319763;
assign addr[25989] = -1923900201;
assign addr[25990] = -1915328086;
assign addr[25991] = -1906604097;
assign addr[25992] = -1897728925;
assign addr[25993] = -1888703276;
assign addr[25994] = -1879527863;
assign addr[25995] = -1870203416;
assign addr[25996] = -1860730673;
assign addr[25997] = -1851110385;
assign addr[25998] = -1841343316;
assign addr[25999] = -1831430239;
assign addr[26000] = -1821371941;
assign addr[26001] = -1811169220;
assign addr[26002] = -1800822883;
assign addr[26003] = -1790333753;
assign addr[26004] = -1779702660;
assign addr[26005] = -1768930447;
assign addr[26006] = -1758017969;
assign addr[26007] = -1746966091;
assign addr[26008] = -1735775690;
assign addr[26009] = -1724447652;
assign addr[26010] = -1712982875;
assign addr[26011] = -1701382270;
assign addr[26012] = -1689646755;
assign addr[26013] = -1677777262;
assign addr[26014] = -1665774731;
assign addr[26015] = -1653640115;
assign addr[26016] = -1641374375;
assign addr[26017] = -1628978484;
assign addr[26018] = -1616453425;
assign addr[26019] = -1603800191;
assign addr[26020] = -1591019785;
assign addr[26021] = -1578113222;
assign addr[26022] = -1565081523;
assign addr[26023] = -1551925723;
assign addr[26024] = -1538646865;
assign addr[26025] = -1525246002;
assign addr[26026] = -1511724196;
assign addr[26027] = -1498082520;
assign addr[26028] = -1484322054;
assign addr[26029] = -1470443891;
assign addr[26030] = -1456449131;
assign addr[26031] = -1442338884;
assign addr[26032] = -1428114267;
assign addr[26033] = -1413776410;
assign addr[26034] = -1399326449;
assign addr[26035] = -1384765530;
assign addr[26036] = -1370094808;
assign addr[26037] = -1355315445;
assign addr[26038] = -1340428615;
assign addr[26039] = -1325435496;
assign addr[26040] = -1310337279;
assign addr[26041] = -1295135159;
assign addr[26042] = -1279830344;
assign addr[26043] = -1264424045;
assign addr[26044] = -1248917486;
assign addr[26045] = -1233311895;
assign addr[26046] = -1217608510;
assign addr[26047] = -1201808576;
assign addr[26048] = -1185913346;
assign addr[26049] = -1169924081;
assign addr[26050] = -1153842047;
assign addr[26051] = -1137668521;
assign addr[26052] = -1121404785;
assign addr[26053] = -1105052128;
assign addr[26054] = -1088611847;
assign addr[26055] = -1072085246;
assign addr[26056] = -1055473635;
assign addr[26057] = -1038778332;
assign addr[26058] = -1022000660;
assign addr[26059] = -1005141949;
assign addr[26060] = -988203537;
assign addr[26061] = -971186766;
assign addr[26062] = -954092986;
assign addr[26063] = -936923553;
assign addr[26064] = -919679827;
assign addr[26065] = -902363176;
assign addr[26066] = -884974973;
assign addr[26067] = -867516597;
assign addr[26068] = -849989433;
assign addr[26069] = -832394869;
assign addr[26070] = -814734301;
assign addr[26071] = -797009130;
assign addr[26072] = -779220762;
assign addr[26073] = -761370605;
assign addr[26074] = -743460077;
assign addr[26075] = -725490597;
assign addr[26076] = -707463589;
assign addr[26077] = -689380485;
assign addr[26078] = -671242716;
assign addr[26079] = -653051723;
assign addr[26080] = -634808946;
assign addr[26081] = -616515832;
assign addr[26082] = -598173833;
assign addr[26083] = -579784402;
assign addr[26084] = -561348998;
assign addr[26085] = -542869083;
assign addr[26086] = -524346121;
assign addr[26087] = -505781581;
assign addr[26088] = -487176937;
assign addr[26089] = -468533662;
assign addr[26090] = -449853235;
assign addr[26091] = -431137138;
assign addr[26092] = -412386854;
assign addr[26093] = -393603870;
assign addr[26094] = -374789676;
assign addr[26095] = -355945764;
assign addr[26096] = -337073627;
assign addr[26097] = -318174762;
assign addr[26098] = -299250668;
assign addr[26099] = -280302845;
assign addr[26100] = -261332796;
assign addr[26101] = -242342025;
assign addr[26102] = -223332037;
assign addr[26103] = -204304341;
assign addr[26104] = -185260444;
assign addr[26105] = -166201858;
assign addr[26106] = -147130093;
assign addr[26107] = -128046661;
assign addr[26108] = -108953076;
assign addr[26109] = -89850852;
assign addr[26110] = -70741503;
assign addr[26111] = -51626544;
assign addr[26112] = -32507492;
assign addr[26113] = -13385863;
assign addr[26114] = 5736829;
assign addr[26115] = 24859065;
assign addr[26116] = 43979330;
assign addr[26117] = 63096108;
assign addr[26118] = 82207882;
assign addr[26119] = 101313138;
assign addr[26120] = 120410361;
assign addr[26121] = 139498035;
assign addr[26122] = 158574649;
assign addr[26123] = 177638688;
assign addr[26124] = 196688642;
assign addr[26125] = 215722999;
assign addr[26126] = 234740251;
assign addr[26127] = 253738890;
assign addr[26128] = 272717408;
assign addr[26129] = 291674302;
assign addr[26130] = 310608068;
assign addr[26131] = 329517204;
assign addr[26132] = 348400212;
assign addr[26133] = 367255594;
assign addr[26134] = 386081854;
assign addr[26135] = 404877501;
assign addr[26136] = 423641043;
assign addr[26137] = 442370993;
assign addr[26138] = 461065866;
assign addr[26139] = 479724180;
assign addr[26140] = 498344454;
assign addr[26141] = 516925212;
assign addr[26142] = 535464981;
assign addr[26143] = 553962291;
assign addr[26144] = 572415676;
assign addr[26145] = 590823671;
assign addr[26146] = 609184818;
assign addr[26147] = 627497660;
assign addr[26148] = 645760745;
assign addr[26149] = 663972625;
assign addr[26150] = 682131857;
assign addr[26151] = 700236999;
assign addr[26152] = 718286617;
assign addr[26153] = 736279279;
assign addr[26154] = 754213559;
assign addr[26155] = 772088034;
assign addr[26156] = 789901288;
assign addr[26157] = 807651907;
assign addr[26158] = 825338484;
assign addr[26159] = 842959617;
assign addr[26160] = 860513908;
assign addr[26161] = 877999966;
assign addr[26162] = 895416404;
assign addr[26163] = 912761841;
assign addr[26164] = 930034901;
assign addr[26165] = 947234215;
assign addr[26166] = 964358420;
assign addr[26167] = 981406156;
assign addr[26168] = 998376073;
assign addr[26169] = 1015266825;
assign addr[26170] = 1032077073;
assign addr[26171] = 1048805483;
assign addr[26172] = 1065450729;
assign addr[26173] = 1082011492;
assign addr[26174] = 1098486458;
assign addr[26175] = 1114874320;
assign addr[26176] = 1131173780;
assign addr[26177] = 1147383544;
assign addr[26178] = 1163502328;
assign addr[26179] = 1179528853;
assign addr[26180] = 1195461849;
assign addr[26181] = 1211300053;
assign addr[26182] = 1227042207;
assign addr[26183] = 1242687064;
assign addr[26184] = 1258233384;
assign addr[26185] = 1273679934;
assign addr[26186] = 1289025489;
assign addr[26187] = 1304268832;
assign addr[26188] = 1319408754;
assign addr[26189] = 1334444055;
assign addr[26190] = 1349373543;
assign addr[26191] = 1364196034;
assign addr[26192] = 1378910353;
assign addr[26193] = 1393515332;
assign addr[26194] = 1408009814;
assign addr[26195] = 1422392650;
assign addr[26196] = 1436662698;
assign addr[26197] = 1450818828;
assign addr[26198] = 1464859917;
assign addr[26199] = 1478784851;
assign addr[26200] = 1492592527;
assign addr[26201] = 1506281850;
assign addr[26202] = 1519851733;
assign addr[26203] = 1533301101;
assign addr[26204] = 1546628888;
assign addr[26205] = 1559834037;
assign addr[26206] = 1572915501;
assign addr[26207] = 1585872242;
assign addr[26208] = 1598703233;
assign addr[26209] = 1611407456;
assign addr[26210] = 1623983905;
assign addr[26211] = 1636431582;
assign addr[26212] = 1648749499;
assign addr[26213] = 1660936681;
assign addr[26214] = 1672992161;
assign addr[26215] = 1684914983;
assign addr[26216] = 1696704201;
assign addr[26217] = 1708358881;
assign addr[26218] = 1719878099;
assign addr[26219] = 1731260941;
assign addr[26220] = 1742506504;
assign addr[26221] = 1753613897;
assign addr[26222] = 1764582240;
assign addr[26223] = 1775410662;
assign addr[26224] = 1786098304;
assign addr[26225] = 1796644320;
assign addr[26226] = 1807047873;
assign addr[26227] = 1817308138;
assign addr[26228] = 1827424302;
assign addr[26229] = 1837395562;
assign addr[26230] = 1847221128;
assign addr[26231] = 1856900221;
assign addr[26232] = 1866432072;
assign addr[26233] = 1875815927;
assign addr[26234] = 1885051042;
assign addr[26235] = 1894136683;
assign addr[26236] = 1903072131;
assign addr[26237] = 1911856677;
assign addr[26238] = 1920489624;
assign addr[26239] = 1928970288;
assign addr[26240] = 1937297997;
assign addr[26241] = 1945472089;
assign addr[26242] = 1953491918;
assign addr[26243] = 1961356847;
assign addr[26244] = 1969066252;
assign addr[26245] = 1976619522;
assign addr[26246] = 1984016058;
assign addr[26247] = 1991255274;
assign addr[26248] = 1998336596;
assign addr[26249] = 2005259462;
assign addr[26250] = 2012023322;
assign addr[26251] = 2018627642;
assign addr[26252] = 2025071897;
assign addr[26253] = 2031355576;
assign addr[26254] = 2037478181;
assign addr[26255] = 2043439226;
assign addr[26256] = 2049238240;
assign addr[26257] = 2054874761;
assign addr[26258] = 2060348343;
assign addr[26259] = 2065658552;
assign addr[26260] = 2070804967;
assign addr[26261] = 2075787180;
assign addr[26262] = 2080604795;
assign addr[26263] = 2085257431;
assign addr[26264] = 2089744719;
assign addr[26265] = 2094066304;
assign addr[26266] = 2098221841;
assign addr[26267] = 2102211002;
assign addr[26268] = 2106033471;
assign addr[26269] = 2109688944;
assign addr[26270] = 2113177132;
assign addr[26271] = 2116497758;
assign addr[26272] = 2119650558;
assign addr[26273] = 2122635283;
assign addr[26274] = 2125451696;
assign addr[26275] = 2128099574;
assign addr[26276] = 2130578706;
assign addr[26277] = 2132888897;
assign addr[26278] = 2135029962;
assign addr[26279] = 2137001733;
assign addr[26280] = 2138804053;
assign addr[26281] = 2140436778;
assign addr[26282] = 2141899780;
assign addr[26283] = 2143192942;
assign addr[26284] = 2144316162;
assign addr[26285] = 2145269351;
assign addr[26286] = 2146052433;
assign addr[26287] = 2146665347;
assign addr[26288] = 2147108043;
assign addr[26289] = 2147380486;
assign addr[26290] = 2147482655;
assign addr[26291] = 2147414542;
assign addr[26292] = 2147176152;
assign addr[26293] = 2146767505;
assign addr[26294] = 2146188631;
assign addr[26295] = 2145439578;
assign addr[26296] = 2144520405;
assign addr[26297] = 2143431184;
assign addr[26298] = 2142172003;
assign addr[26299] = 2140742960;
assign addr[26300] = 2139144169;
assign addr[26301] = 2137375758;
assign addr[26302] = 2135437865;
assign addr[26303] = 2133330646;
assign addr[26304] = 2131054266;
assign addr[26305] = 2128608907;
assign addr[26306] = 2125994762;
assign addr[26307] = 2123212038;
assign addr[26308] = 2120260957;
assign addr[26309] = 2117141752;
assign addr[26310] = 2113854671;
assign addr[26311] = 2110399974;
assign addr[26312] = 2106777935;
assign addr[26313] = 2102988841;
assign addr[26314] = 2099032994;
assign addr[26315] = 2094910706;
assign addr[26316] = 2090622304;
assign addr[26317] = 2086168128;
assign addr[26318] = 2081548533;
assign addr[26319] = 2076763883;
assign addr[26320] = 2071814558;
assign addr[26321] = 2066700952;
assign addr[26322] = 2061423468;
assign addr[26323] = 2055982526;
assign addr[26324] = 2050378558;
assign addr[26325] = 2044612007;
assign addr[26326] = 2038683330;
assign addr[26327] = 2032592999;
assign addr[26328] = 2026341495;
assign addr[26329] = 2019929315;
assign addr[26330] = 2013356967;
assign addr[26331] = 2006624971;
assign addr[26332] = 1999733863;
assign addr[26333] = 1992684188;
assign addr[26334] = 1985476506;
assign addr[26335] = 1978111387;
assign addr[26336] = 1970589416;
assign addr[26337] = 1962911189;
assign addr[26338] = 1955077316;
assign addr[26339] = 1947088417;
assign addr[26340] = 1938945125;
assign addr[26341] = 1930648088;
assign addr[26342] = 1922197961;
assign addr[26343] = 1913595416;
assign addr[26344] = 1904841135;
assign addr[26345] = 1895935811;
assign addr[26346] = 1886880151;
assign addr[26347] = 1877674873;
assign addr[26348] = 1868320707;
assign addr[26349] = 1858818395;
assign addr[26350] = 1849168689;
assign addr[26351] = 1839372356;
assign addr[26352] = 1829430172;
assign addr[26353] = 1819342925;
assign addr[26354] = 1809111415;
assign addr[26355] = 1798736454;
assign addr[26356] = 1788218865;
assign addr[26357] = 1777559480;
assign addr[26358] = 1766759146;
assign addr[26359] = 1755818718;
assign addr[26360] = 1744739065;
assign addr[26361] = 1733521064;
assign addr[26362] = 1722165606;
assign addr[26363] = 1710673591;
assign addr[26364] = 1699045930;
assign addr[26365] = 1687283545;
assign addr[26366] = 1675387369;
assign addr[26367] = 1663358344;
assign addr[26368] = 1651197426;
assign addr[26369] = 1638905577;
assign addr[26370] = 1626483774;
assign addr[26371] = 1613933000;
assign addr[26372] = 1601254251;
assign addr[26373] = 1588448533;
assign addr[26374] = 1575516860;
assign addr[26375] = 1562460258;
assign addr[26376] = 1549279763;
assign addr[26377] = 1535976419;
assign addr[26378] = 1522551282;
assign addr[26379] = 1509005416;
assign addr[26380] = 1495339895;
assign addr[26381] = 1481555802;
assign addr[26382] = 1467654232;
assign addr[26383] = 1453636285;
assign addr[26384] = 1439503074;
assign addr[26385] = 1425255719;
assign addr[26386] = 1410895350;
assign addr[26387] = 1396423105;
assign addr[26388] = 1381840133;
assign addr[26389] = 1367147589;
assign addr[26390] = 1352346639;
assign addr[26391] = 1337438456;
assign addr[26392] = 1322424222;
assign addr[26393] = 1307305128;
assign addr[26394] = 1292082373;
assign addr[26395] = 1276757164;
assign addr[26396] = 1261330715;
assign addr[26397] = 1245804251;
assign addr[26398] = 1230179002;
assign addr[26399] = 1214456207;
assign addr[26400] = 1198637114;
assign addr[26401] = 1182722976;
assign addr[26402] = 1166715055;
assign addr[26403] = 1150614620;
assign addr[26404] = 1134422949;
assign addr[26405] = 1118141326;
assign addr[26406] = 1101771040;
assign addr[26407] = 1085313391;
assign addr[26408] = 1068769683;
assign addr[26409] = 1052141228;
assign addr[26410] = 1035429345;
assign addr[26411] = 1018635358;
assign addr[26412] = 1001760600;
assign addr[26413] = 984806408;
assign addr[26414] = 967774128;
assign addr[26415] = 950665109;
assign addr[26416] = 933480707;
assign addr[26417] = 916222287;
assign addr[26418] = 898891215;
assign addr[26419] = 881488868;
assign addr[26420] = 864016623;
assign addr[26421] = 846475867;
assign addr[26422] = 828867991;
assign addr[26423] = 811194391;
assign addr[26424] = 793456467;
assign addr[26425] = 775655628;
assign addr[26426] = 757793284;
assign addr[26427] = 739870851;
assign addr[26428] = 721889752;
assign addr[26429] = 703851410;
assign addr[26430] = 685757258;
assign addr[26431] = 667608730;
assign addr[26432] = 649407264;
assign addr[26433] = 631154304;
assign addr[26434] = 612851297;
assign addr[26435] = 594499695;
assign addr[26436] = 576100953;
assign addr[26437] = 557656529;
assign addr[26438] = 539167887;
assign addr[26439] = 520636492;
assign addr[26440] = 502063814;
assign addr[26441] = 483451325;
assign addr[26442] = 464800501;
assign addr[26443] = 446112822;
assign addr[26444] = 427389768;
assign addr[26445] = 408632825;
assign addr[26446] = 389843480;
assign addr[26447] = 371023223;
assign addr[26448] = 352173546;
assign addr[26449] = 333295944;
assign addr[26450] = 314391913;
assign addr[26451] = 295462954;
assign addr[26452] = 276510565;
assign addr[26453] = 257536251;
assign addr[26454] = 238541516;
assign addr[26455] = 219527866;
assign addr[26456] = 200496809;
assign addr[26457] = 181449854;
assign addr[26458] = 162388511;
assign addr[26459] = 143314291;
assign addr[26460] = 124228708;
assign addr[26461] = 105133274;
assign addr[26462] = 86029503;
assign addr[26463] = 66918911;
assign addr[26464] = 47803013;
assign addr[26465] = 28683324;
assign addr[26466] = 9561361;
assign addr[26467] = -9561361;
assign addr[26468] = -28683324;
assign addr[26469] = -47803013;
assign addr[26470] = -66918911;
assign addr[26471] = -86029503;
assign addr[26472] = -105133274;
assign addr[26473] = -124228708;
assign addr[26474] = -143314291;
assign addr[26475] = -162388511;
assign addr[26476] = -181449854;
assign addr[26477] = -200496809;
assign addr[26478] = -219527866;
assign addr[26479] = -238541516;
assign addr[26480] = -257536251;
assign addr[26481] = -276510565;
assign addr[26482] = -295462953;
assign addr[26483] = -314391913;
assign addr[26484] = -333295944;
assign addr[26485] = -352173546;
assign addr[26486] = -371023223;
assign addr[26487] = -389843480;
assign addr[26488] = -408632825;
assign addr[26489] = -427389768;
assign addr[26490] = -446112822;
assign addr[26491] = -464800501;
assign addr[26492] = -483451325;
assign addr[26493] = -502063814;
assign addr[26494] = -520636492;
assign addr[26495] = -539167887;
assign addr[26496] = -557656529;
assign addr[26497] = -576100953;
assign addr[26498] = -594499695;
assign addr[26499] = -612851297;
assign addr[26500] = -631154304;
assign addr[26501] = -649407264;
assign addr[26502] = -667608730;
assign addr[26503] = -685757258;
assign addr[26504] = -703851410;
assign addr[26505] = -721889752;
assign addr[26506] = -739870851;
assign addr[26507] = -757793284;
assign addr[26508] = -775655628;
assign addr[26509] = -793456467;
assign addr[26510] = -811194391;
assign addr[26511] = -828867991;
assign addr[26512] = -846475867;
assign addr[26513] = -864016623;
assign addr[26514] = -881488868;
assign addr[26515] = -898891215;
assign addr[26516] = -916222287;
assign addr[26517] = -933480707;
assign addr[26518] = -950665109;
assign addr[26519] = -967774128;
assign addr[26520] = -984806408;
assign addr[26521] = -1001760600;
assign addr[26522] = -1018635358;
assign addr[26523] = -1035429345;
assign addr[26524] = -1052141228;
assign addr[26525] = -1068769683;
assign addr[26526] = -1085313391;
assign addr[26527] = -1101771040;
assign addr[26528] = -1118141326;
assign addr[26529] = -1134422949;
assign addr[26530] = -1150614620;
assign addr[26531] = -1166715055;
assign addr[26532] = -1182722976;
assign addr[26533] = -1198637114;
assign addr[26534] = -1214456207;
assign addr[26535] = -1230179002;
assign addr[26536] = -1245804251;
assign addr[26537] = -1261330715;
assign addr[26538] = -1276757164;
assign addr[26539] = -1292082373;
assign addr[26540] = -1307305128;
assign addr[26541] = -1322424222;
assign addr[26542] = -1337438456;
assign addr[26543] = -1352346639;
assign addr[26544] = -1367147589;
assign addr[26545] = -1381840133;
assign addr[26546] = -1396423105;
assign addr[26547] = -1410895350;
assign addr[26548] = -1425255719;
assign addr[26549] = -1439503074;
assign addr[26550] = -1453636285;
assign addr[26551] = -1467654232;
assign addr[26552] = -1481555802;
assign addr[26553] = -1495339895;
assign addr[26554] = -1509005416;
assign addr[26555] = -1522551282;
assign addr[26556] = -1535976419;
assign addr[26557] = -1549279763;
assign addr[26558] = -1562460258;
assign addr[26559] = -1575516860;
assign addr[26560] = -1588448533;
assign addr[26561] = -1601254251;
assign addr[26562] = -1613933000;
assign addr[26563] = -1626483774;
assign addr[26564] = -1638905577;
assign addr[26565] = -1651197426;
assign addr[26566] = -1663358344;
assign addr[26567] = -1675387369;
assign addr[26568] = -1687283545;
assign addr[26569] = -1699045930;
assign addr[26570] = -1710673591;
assign addr[26571] = -1722165606;
assign addr[26572] = -1733521064;
assign addr[26573] = -1744739065;
assign addr[26574] = -1755818718;
assign addr[26575] = -1766759146;
assign addr[26576] = -1777559480;
assign addr[26577] = -1788218865;
assign addr[26578] = -1798736454;
assign addr[26579] = -1809111415;
assign addr[26580] = -1819342925;
assign addr[26581] = -1829430172;
assign addr[26582] = -1839372356;
assign addr[26583] = -1849168689;
assign addr[26584] = -1858818395;
assign addr[26585] = -1868320707;
assign addr[26586] = -1877674873;
assign addr[26587] = -1886880151;
assign addr[26588] = -1895935811;
assign addr[26589] = -1904841135;
assign addr[26590] = -1913595416;
assign addr[26591] = -1922197961;
assign addr[26592] = -1930648088;
assign addr[26593] = -1938945125;
assign addr[26594] = -1947088417;
assign addr[26595] = -1955077316;
assign addr[26596] = -1962911189;
assign addr[26597] = -1970589416;
assign addr[26598] = -1978111387;
assign addr[26599] = -1985476506;
assign addr[26600] = -1992684188;
assign addr[26601] = -1999733863;
assign addr[26602] = -2006624971;
assign addr[26603] = -2013356967;
assign addr[26604] = -2019929315;
assign addr[26605] = -2026341495;
assign addr[26606] = -2032592999;
assign addr[26607] = -2038683330;
assign addr[26608] = -2044612007;
assign addr[26609] = -2050378558;
assign addr[26610] = -2055982526;
assign addr[26611] = -2061423468;
assign addr[26612] = -2066700952;
assign addr[26613] = -2071814558;
assign addr[26614] = -2076763883;
assign addr[26615] = -2081548533;
assign addr[26616] = -2086168128;
assign addr[26617] = -2090622304;
assign addr[26618] = -2094910706;
assign addr[26619] = -2099032994;
assign addr[26620] = -2102988841;
assign addr[26621] = -2106777935;
assign addr[26622] = -2110399974;
assign addr[26623] = -2113854671;
assign addr[26624] = -2117141752;
assign addr[26625] = -2120260957;
assign addr[26626] = -2123212038;
assign addr[26627] = -2125994762;
assign addr[26628] = -2128608907;
assign addr[26629] = -2131054266;
assign addr[26630] = -2133330646;
assign addr[26631] = -2135437865;
assign addr[26632] = -2137375758;
assign addr[26633] = -2139144169;
assign addr[26634] = -2140742960;
assign addr[26635] = -2142172003;
assign addr[26636] = -2143431184;
assign addr[26637] = -2144520405;
assign addr[26638] = -2145439578;
assign addr[26639] = -2146188631;
assign addr[26640] = -2146767505;
assign addr[26641] = -2147176152;
assign addr[26642] = -2147414542;
assign addr[26643] = -2147482655;
assign addr[26644] = -2147380486;
assign addr[26645] = -2147108043;
assign addr[26646] = -2146665347;
assign addr[26647] = -2146052433;
assign addr[26648] = -2145269351;
assign addr[26649] = -2144316162;
assign addr[26650] = -2143192942;
assign addr[26651] = -2141899780;
assign addr[26652] = -2140436778;
assign addr[26653] = -2138804053;
assign addr[26654] = -2137001733;
assign addr[26655] = -2135029962;
assign addr[26656] = -2132888897;
assign addr[26657] = -2130578706;
assign addr[26658] = -2128099574;
assign addr[26659] = -2125451696;
assign addr[26660] = -2122635283;
assign addr[26661] = -2119650558;
assign addr[26662] = -2116497758;
assign addr[26663] = -2113177132;
assign addr[26664] = -2109688944;
assign addr[26665] = -2106033471;
assign addr[26666] = -2102211002;
assign addr[26667] = -2098221841;
assign addr[26668] = -2094066304;
assign addr[26669] = -2089744719;
assign addr[26670] = -2085257431;
assign addr[26671] = -2080604795;
assign addr[26672] = -2075787180;
assign addr[26673] = -2070804967;
assign addr[26674] = -2065658552;
assign addr[26675] = -2060348343;
assign addr[26676] = -2054874761;
assign addr[26677] = -2049238240;
assign addr[26678] = -2043439226;
assign addr[26679] = -2037478181;
assign addr[26680] = -2031355576;
assign addr[26681] = -2025071897;
assign addr[26682] = -2018627642;
assign addr[26683] = -2012023322;
assign addr[26684] = -2005259462;
assign addr[26685] = -1998336596;
assign addr[26686] = -1991255274;
assign addr[26687] = -1984016058;
assign addr[26688] = -1976619522;
assign addr[26689] = -1969066252;
assign addr[26690] = -1961356847;
assign addr[26691] = -1953491918;
assign addr[26692] = -1945472089;
assign addr[26693] = -1937297997;
assign addr[26694] = -1928970288;
assign addr[26695] = -1920489624;
assign addr[26696] = -1911856677;
assign addr[26697] = -1903072131;
assign addr[26698] = -1894136683;
assign addr[26699] = -1885051042;
assign addr[26700] = -1875815927;
assign addr[26701] = -1866432072;
assign addr[26702] = -1856900221;
assign addr[26703] = -1847221128;
assign addr[26704] = -1837395562;
assign addr[26705] = -1827424302;
assign addr[26706] = -1817308138;
assign addr[26707] = -1807047873;
assign addr[26708] = -1796644320;
assign addr[26709] = -1786098304;
assign addr[26710] = -1775410662;
assign addr[26711] = -1764582240;
assign addr[26712] = -1753613897;
assign addr[26713] = -1742506504;
assign addr[26714] = -1731260941;
assign addr[26715] = -1719878099;
assign addr[26716] = -1708358881;
assign addr[26717] = -1696704201;
assign addr[26718] = -1684914983;
assign addr[26719] = -1672992161;
assign addr[26720] = -1660936681;
assign addr[26721] = -1648749499;
assign addr[26722] = -1636431582;
assign addr[26723] = -1623983905;
assign addr[26724] = -1611407456;
assign addr[26725] = -1598703233;
assign addr[26726] = -1585872242;
assign addr[26727] = -1572915501;
assign addr[26728] = -1559834037;
assign addr[26729] = -1546628888;
assign addr[26730] = -1533301101;
assign addr[26731] = -1519851733;
assign addr[26732] = -1506281850;
assign addr[26733] = -1492592527;
assign addr[26734] = -1478784851;
assign addr[26735] = -1464859917;
assign addr[26736] = -1450818828;
assign addr[26737] = -1436662698;
assign addr[26738] = -1422392650;
assign addr[26739] = -1408009814;
assign addr[26740] = -1393515332;
assign addr[26741] = -1378910353;
assign addr[26742] = -1364196034;
assign addr[26743] = -1349373543;
assign addr[26744] = -1334444055;
assign addr[26745] = -1319408754;
assign addr[26746] = -1304268832;
assign addr[26747] = -1289025489;
assign addr[26748] = -1273679934;
assign addr[26749] = -1258233384;
assign addr[26750] = -1242687064;
assign addr[26751] = -1227042207;
assign addr[26752] = -1211300053;
assign addr[26753] = -1195461849;
assign addr[26754] = -1179528853;
assign addr[26755] = -1163502328;
assign addr[26756] = -1147383544;
assign addr[26757] = -1131173780;
assign addr[26758] = -1114874320;
assign addr[26759] = -1098486458;
assign addr[26760] = -1082011492;
assign addr[26761] = -1065450729;
assign addr[26762] = -1048805483;
assign addr[26763] = -1032077073;
assign addr[26764] = -1015266825;
assign addr[26765] = -998376073;
assign addr[26766] = -981406156;
assign addr[26767] = -964358420;
assign addr[26768] = -947234215;
assign addr[26769] = -930034901;
assign addr[26770] = -912761841;
assign addr[26771] = -895416404;
assign addr[26772] = -877999966;
assign addr[26773] = -860513908;
assign addr[26774] = -842959617;
assign addr[26775] = -825338484;
assign addr[26776] = -807651907;
assign addr[26777] = -789901288;
assign addr[26778] = -772088034;
assign addr[26779] = -754213559;
assign addr[26780] = -736279279;
assign addr[26781] = -718286617;
assign addr[26782] = -700236999;
assign addr[26783] = -682131857;
assign addr[26784] = -663972625;
assign addr[26785] = -645760745;
assign addr[26786] = -627497660;
assign addr[26787] = -609184818;
assign addr[26788] = -590823671;
assign addr[26789] = -572415676;
assign addr[26790] = -553962291;
assign addr[26791] = -535464981;
assign addr[26792] = -516925212;
assign addr[26793] = -498344454;
assign addr[26794] = -479724180;
assign addr[26795] = -461065866;
assign addr[26796] = -442370993;
assign addr[26797] = -423641043;
assign addr[26798] = -404877501;
assign addr[26799] = -386081854;
assign addr[26800] = -367255594;
assign addr[26801] = -348400212;
assign addr[26802] = -329517204;
assign addr[26803] = -310608068;
assign addr[26804] = -291674302;
assign addr[26805] = -272717408;
assign addr[26806] = -253738890;
assign addr[26807] = -234740251;
assign addr[26808] = -215722999;
assign addr[26809] = -196688642;
assign addr[26810] = -177638688;
assign addr[26811] = -158574649;
assign addr[26812] = -139498035;
assign addr[26813] = -120410361;
assign addr[26814] = -101313138;
assign addr[26815] = -82207882;
assign addr[26816] = -63096108;
assign addr[26817] = -43979330;
assign addr[26818] = -24859065;
assign addr[26819] = -5736829;
assign addr[26820] = 13385863;
assign addr[26821] = 32507492;
assign addr[26822] = 51626544;
assign addr[26823] = 70741503;
assign addr[26824] = 89850852;
assign addr[26825] = 108953076;
assign addr[26826] = 128046661;
assign addr[26827] = 147130093;
assign addr[26828] = 166201858;
assign addr[26829] = 185260444;
assign addr[26830] = 204304341;
assign addr[26831] = 223332037;
assign addr[26832] = 242342025;
assign addr[26833] = 261332796;
assign addr[26834] = 280302845;
assign addr[26835] = 299250668;
assign addr[26836] = 318174762;
assign addr[26837] = 337073627;
assign addr[26838] = 355945764;
assign addr[26839] = 374789676;
assign addr[26840] = 393603870;
assign addr[26841] = 412386854;
assign addr[26842] = 431137138;
assign addr[26843] = 449853235;
assign addr[26844] = 468533662;
assign addr[26845] = 487176937;
assign addr[26846] = 505781581;
assign addr[26847] = 524346121;
assign addr[26848] = 542869083;
assign addr[26849] = 561348998;
assign addr[26850] = 579784402;
assign addr[26851] = 598173833;
assign addr[26852] = 616515832;
assign addr[26853] = 634808946;
assign addr[26854] = 653051723;
assign addr[26855] = 671242716;
assign addr[26856] = 689380485;
assign addr[26857] = 707463589;
assign addr[26858] = 725490597;
assign addr[26859] = 743460077;
assign addr[26860] = 761370605;
assign addr[26861] = 779220762;
assign addr[26862] = 797009130;
assign addr[26863] = 814734301;
assign addr[26864] = 832394869;
assign addr[26865] = 849989433;
assign addr[26866] = 867516597;
assign addr[26867] = 884974973;
assign addr[26868] = 902363176;
assign addr[26869] = 919679827;
assign addr[26870] = 936923553;
assign addr[26871] = 954092986;
assign addr[26872] = 971186766;
assign addr[26873] = 988203537;
assign addr[26874] = 1005141949;
assign addr[26875] = 1022000660;
assign addr[26876] = 1038778332;
assign addr[26877] = 1055473635;
assign addr[26878] = 1072085246;
assign addr[26879] = 1088611847;
assign addr[26880] = 1105052128;
assign addr[26881] = 1121404785;
assign addr[26882] = 1137668521;
assign addr[26883] = 1153842047;
assign addr[26884] = 1169924081;
assign addr[26885] = 1185913346;
assign addr[26886] = 1201808576;
assign addr[26887] = 1217608510;
assign addr[26888] = 1233311895;
assign addr[26889] = 1248917486;
assign addr[26890] = 1264424045;
assign addr[26891] = 1279830344;
assign addr[26892] = 1295135159;
assign addr[26893] = 1310337279;
assign addr[26894] = 1325435496;
assign addr[26895] = 1340428615;
assign addr[26896] = 1355315445;
assign addr[26897] = 1370094808;
assign addr[26898] = 1384765530;
assign addr[26899] = 1399326449;
assign addr[26900] = 1413776410;
assign addr[26901] = 1428114267;
assign addr[26902] = 1442338884;
assign addr[26903] = 1456449131;
assign addr[26904] = 1470443891;
assign addr[26905] = 1484322054;
assign addr[26906] = 1498082520;
assign addr[26907] = 1511724196;
assign addr[26908] = 1525246002;
assign addr[26909] = 1538646865;
assign addr[26910] = 1551925723;
assign addr[26911] = 1565081523;
assign addr[26912] = 1578113222;
assign addr[26913] = 1591019785;
assign addr[26914] = 1603800191;
assign addr[26915] = 1616453425;
assign addr[26916] = 1628978484;
assign addr[26917] = 1641374375;
assign addr[26918] = 1653640115;
assign addr[26919] = 1665774731;
assign addr[26920] = 1677777262;
assign addr[26921] = 1689646755;
assign addr[26922] = 1701382270;
assign addr[26923] = 1712982875;
assign addr[26924] = 1724447652;
assign addr[26925] = 1735775690;
assign addr[26926] = 1746966091;
assign addr[26927] = 1758017969;
assign addr[26928] = 1768930447;
assign addr[26929] = 1779702660;
assign addr[26930] = 1790333753;
assign addr[26931] = 1800822883;
assign addr[26932] = 1811169220;
assign addr[26933] = 1821371941;
assign addr[26934] = 1831430239;
assign addr[26935] = 1841343316;
assign addr[26936] = 1851110385;
assign addr[26937] = 1860730673;
assign addr[26938] = 1870203416;
assign addr[26939] = 1879527863;
assign addr[26940] = 1888703276;
assign addr[26941] = 1897728925;
assign addr[26942] = 1906604097;
assign addr[26943] = 1915328086;
assign addr[26944] = 1923900201;
assign addr[26945] = 1932319763;
assign addr[26946] = 1940586104;
assign addr[26947] = 1948698568;
assign addr[26948] = 1956656513;
assign addr[26949] = 1964459306;
assign addr[26950] = 1972106330;
assign addr[26951] = 1979596978;
assign addr[26952] = 1986930656;
assign addr[26953] = 1994106782;
assign addr[26954] = 2001124788;
assign addr[26955] = 2007984117;
assign addr[26956] = 2014684225;
assign addr[26957] = 2021224581;
assign addr[26958] = 2027604666;
assign addr[26959] = 2033823974;
assign addr[26960] = 2039882013;
assign addr[26961] = 2045778302;
assign addr[26962] = 2051512372;
assign addr[26963] = 2057083771;
assign addr[26964] = 2062492055;
assign addr[26965] = 2067736796;
assign addr[26966] = 2072817579;
assign addr[26967] = 2077733999;
assign addr[26968] = 2082485668;
assign addr[26969] = 2087072209;
assign addr[26970] = 2091493257;
assign addr[26971] = 2095748463;
assign addr[26972] = 2099837489;
assign addr[26973] = 2103760010;
assign addr[26974] = 2107515716;
assign addr[26975] = 2111104309;
assign addr[26976] = 2114525505;
assign addr[26977] = 2117779031;
assign addr[26978] = 2120864631;
assign addr[26979] = 2123782059;
assign addr[26980] = 2126531084;
assign addr[26981] = 2129111488;
assign addr[26982] = 2131523066;
assign addr[26983] = 2133765628;
assign addr[26984] = 2135838995;
assign addr[26985] = 2137743003;
assign addr[26986] = 2139477502;
assign addr[26987] = 2141042352;
assign addr[26988] = 2142437431;
assign addr[26989] = 2143662628;
assign addr[26990] = 2144717846;
assign addr[26991] = 2145603001;
assign addr[26992] = 2146318022;
assign addr[26993] = 2146862854;
assign addr[26994] = 2147237452;
assign addr[26995] = 2147441787;
assign addr[26996] = 2147475844;
assign addr[26997] = 2147339619;
assign addr[26998] = 2147033123;
assign addr[26999] = 2146556380;
assign addr[27000] = 2145909429;
assign addr[27001] = 2145092320;
assign addr[27002] = 2144105118;
assign addr[27003] = 2142947902;
assign addr[27004] = 2141620763;
assign addr[27005] = 2140123807;
assign addr[27006] = 2138457152;
assign addr[27007] = 2136620930;
assign addr[27008] = 2134615288;
assign addr[27009] = 2132440383;
assign addr[27010] = 2130096389;
assign addr[27011] = 2127583492;
assign addr[27012] = 2124901890;
assign addr[27013] = 2122051796;
assign addr[27014] = 2119033436;
assign addr[27015] = 2115847050;
assign addr[27016] = 2112492891;
assign addr[27017] = 2108971223;
assign addr[27018] = 2105282327;
assign addr[27019] = 2101426496;
assign addr[27020] = 2097404033;
assign addr[27021] = 2093215260;
assign addr[27022] = 2088860507;
assign addr[27023] = 2084340120;
assign addr[27024] = 2079654458;
assign addr[27025] = 2074803892;
assign addr[27026] = 2069788807;
assign addr[27027] = 2064609600;
assign addr[27028] = 2059266683;
assign addr[27029] = 2053760478;
assign addr[27030] = 2048091422;
assign addr[27031] = 2042259965;
assign addr[27032] = 2036266570;
assign addr[27033] = 2030111710;
assign addr[27034] = 2023795876;
assign addr[27035] = 2017319567;
assign addr[27036] = 2010683297;
assign addr[27037] = 2003887591;
assign addr[27038] = 1996932990;
assign addr[27039] = 1989820044;
assign addr[27040] = 1982549318;
assign addr[27041] = 1975121388;
assign addr[27042] = 1967536842;
assign addr[27043] = 1959796283;
assign addr[27044] = 1951900324;
assign addr[27045] = 1943849591;
assign addr[27046] = 1935644723;
assign addr[27047] = 1927286370;
assign addr[27048] = 1918775195;
assign addr[27049] = 1910111873;
assign addr[27050] = 1901297091;
assign addr[27051] = 1892331547;
assign addr[27052] = 1883215953;
assign addr[27053] = 1873951032;
assign addr[27054] = 1864537518;
assign addr[27055] = 1854976157;
assign addr[27056] = 1845267708;
assign addr[27057] = 1835412941;
assign addr[27058] = 1825412636;
assign addr[27059] = 1815267588;
assign addr[27060] = 1804978599;
assign addr[27061] = 1794546487;
assign addr[27062] = 1783972079;
assign addr[27063] = 1773256212;
assign addr[27064] = 1762399737;
assign addr[27065] = 1751403515;
assign addr[27066] = 1740268417;
assign addr[27067] = 1728995326;
assign addr[27068] = 1717585136;
assign addr[27069] = 1706038753;
assign addr[27070] = 1694357091;
assign addr[27071] = 1682541077;
assign addr[27072] = 1670591647;
assign addr[27073] = 1658509750;
assign addr[27074] = 1646296344;
assign addr[27075] = 1633952396;
assign addr[27076] = 1621478885;
assign addr[27077] = 1608876801;
assign addr[27078] = 1596147143;
assign addr[27079] = 1583290921;
assign addr[27080] = 1570309153;
assign addr[27081] = 1557202869;
assign addr[27082] = 1543973108;
assign addr[27083] = 1530620920;
assign addr[27084] = 1517147363;
assign addr[27085] = 1503553506;
assign addr[27086] = 1489840425;
assign addr[27087] = 1476009210;
assign addr[27088] = 1462060956;
assign addr[27089] = 1447996770;
assign addr[27090] = 1433817766;
assign addr[27091] = 1419525069;
assign addr[27092] = 1405119813;
assign addr[27093] = 1390603139;
assign addr[27094] = 1375976199;
assign addr[27095] = 1361240152;
assign addr[27096] = 1346396168;
assign addr[27097] = 1331445422;
assign addr[27098] = 1316389101;
assign addr[27099] = 1301228398;
assign addr[27100] = 1285964516;
assign addr[27101] = 1270598665;
assign addr[27102] = 1255132063;
assign addr[27103] = 1239565936;
assign addr[27104] = 1223901520;
assign addr[27105] = 1208140056;
assign addr[27106] = 1192282793;
assign addr[27107] = 1176330990;
assign addr[27108] = 1160285911;
assign addr[27109] = 1144148829;
assign addr[27110] = 1127921022;
assign addr[27111] = 1111603778;
assign addr[27112] = 1095198391;
assign addr[27113] = 1078706161;
assign addr[27114] = 1062128397;
assign addr[27115] = 1045466412;
assign addr[27116] = 1028721528;
assign addr[27117] = 1011895073;
assign addr[27118] = 994988380;
assign addr[27119] = 978002791;
assign addr[27120] = 960939653;
assign addr[27121] = 943800318;
assign addr[27122] = 926586145;
assign addr[27123] = 909298500;
assign addr[27124] = 891938752;
assign addr[27125] = 874508280;
assign addr[27126] = 857008464;
assign addr[27127] = 839440693;
assign addr[27128] = 821806359;
assign addr[27129] = 804106861;
assign addr[27130] = 786343603;
assign addr[27131] = 768517992;
assign addr[27132] = 750631442;
assign addr[27133] = 732685372;
assign addr[27134] = 714681204;
assign addr[27135] = 696620367;
assign addr[27136] = 678504291;
assign addr[27137] = 660334415;
assign addr[27138] = 642112178;
assign addr[27139] = 623839025;
assign addr[27140] = 605516406;
assign addr[27141] = 587145773;
assign addr[27142] = 568728583;
assign addr[27143] = 550266296;
assign addr[27144] = 531760377;
assign addr[27145] = 513212292;
assign addr[27146] = 494623513;
assign addr[27147] = 475995513;
assign addr[27148] = 457329769;
assign addr[27149] = 438627762;
assign addr[27150] = 419890975;
assign addr[27151] = 401120892;
assign addr[27152] = 382319004;
assign addr[27153] = 363486799;
assign addr[27154] = 344625773;
assign addr[27155] = 325737419;
assign addr[27156] = 306823237;
assign addr[27157] = 287884725;
assign addr[27158] = 268923386;
assign addr[27159] = 249940723;
assign addr[27160] = 230938242;
assign addr[27161] = 211917448;
assign addr[27162] = 192879850;
assign addr[27163] = 173826959;
assign addr[27164] = 154760284;
assign addr[27165] = 135681337;
assign addr[27166] = 116591632;
assign addr[27167] = 97492681;
assign addr[27168] = 78386000;
assign addr[27169] = 59273104;
assign addr[27170] = 40155507;
assign addr[27171] = 21034727;
assign addr[27172] = 1912278;
assign addr[27173] = -17210322;
assign addr[27174] = -36331557;
assign addr[27175] = -55449912;
assign addr[27176] = -74563870;
assign addr[27177] = -93671915;
assign addr[27178] = -112772533;
assign addr[27179] = -131864208;
assign addr[27180] = -150945428;
assign addr[27181] = -170014678;
assign addr[27182] = -189070447;
assign addr[27183] = -208111224;
assign addr[27184] = -227135500;
assign addr[27185] = -246141764;
assign addr[27186] = -265128512;
assign addr[27187] = -284094236;
assign addr[27188] = -303037433;
assign addr[27189] = -321956601;
assign addr[27190] = -340850240;
assign addr[27191] = -359716852;
assign addr[27192] = -378554940;
assign addr[27193] = -397363011;
assign addr[27194] = -416139574;
assign addr[27195] = -434883140;
assign addr[27196] = -453592221;
assign addr[27197] = -472265336;
assign addr[27198] = -490901003;
assign addr[27199] = -509497745;
assign addr[27200] = -528054086;
assign addr[27201] = -546568556;
assign addr[27202] = -565039687;
assign addr[27203] = -583466013;
assign addr[27204] = -601846074;
assign addr[27205] = -620178412;
assign addr[27206] = -638461574;
assign addr[27207] = -656694110;
assign addr[27208] = -674874574;
assign addr[27209] = -693001525;
assign addr[27210] = -711073524;
assign addr[27211] = -729089140;
assign addr[27212] = -747046944;
assign addr[27213] = -764945512;
assign addr[27214] = -782783424;
assign addr[27215] = -800559266;
assign addr[27216] = -818271628;
assign addr[27217] = -835919107;
assign addr[27218] = -853500302;
assign addr[27219] = -871013820;
assign addr[27220] = -888458272;
assign addr[27221] = -905832274;
assign addr[27222] = -923134450;
assign addr[27223] = -940363427;
assign addr[27224] = -957517838;
assign addr[27225] = -974596324;
assign addr[27226] = -991597531;
assign addr[27227] = -1008520110;
assign addr[27228] = -1025362720;
assign addr[27229] = -1042124025;
assign addr[27230] = -1058802695;
assign addr[27231] = -1075397409;
assign addr[27232] = -1091906851;
assign addr[27233] = -1108329711;
assign addr[27234] = -1124664687;
assign addr[27235] = -1140910484;
assign addr[27236] = -1157065814;
assign addr[27237] = -1173129396;
assign addr[27238] = -1189099956;
assign addr[27239] = -1204976227;
assign addr[27240] = -1220756951;
assign addr[27241] = -1236440877;
assign addr[27242] = -1252026760;
assign addr[27243] = -1267513365;
assign addr[27244] = -1282899464;
assign addr[27245] = -1298183838;
assign addr[27246] = -1313365273;
assign addr[27247] = -1328442566;
assign addr[27248] = -1343414522;
assign addr[27249] = -1358279953;
assign addr[27250] = -1373037681;
assign addr[27251] = -1387686535;
assign addr[27252] = -1402225355;
assign addr[27253] = -1416652986;
assign addr[27254] = -1430968286;
assign addr[27255] = -1445170118;
assign addr[27256] = -1459257358;
assign addr[27257] = -1473228887;
assign addr[27258] = -1487083598;
assign addr[27259] = -1500820393;
assign addr[27260] = -1514438181;
assign addr[27261] = -1527935884;
assign addr[27262] = -1541312431;
assign addr[27263] = -1554566762;
assign addr[27264] = -1567697824;
assign addr[27265] = -1580704578;
assign addr[27266] = -1593585992;
assign addr[27267] = -1606341043;
assign addr[27268] = -1618968722;
assign addr[27269] = -1631468027;
assign addr[27270] = -1643837966;
assign addr[27271] = -1656077559;
assign addr[27272] = -1668185835;
assign addr[27273] = -1680161834;
assign addr[27274] = -1692004606;
assign addr[27275] = -1703713213;
assign addr[27276] = -1715286726;
assign addr[27277] = -1726724227;
assign addr[27278] = -1738024810;
assign addr[27279] = -1749187577;
assign addr[27280] = -1760211645;
assign addr[27281] = -1771096139;
assign addr[27282] = -1781840195;
assign addr[27283] = -1792442963;
assign addr[27284] = -1802903601;
assign addr[27285] = -1813221279;
assign addr[27286] = -1823395180;
assign addr[27287] = -1833424497;
assign addr[27288] = -1843308435;
assign addr[27289] = -1853046210;
assign addr[27290] = -1862637049;
assign addr[27291] = -1872080193;
assign addr[27292] = -1881374892;
assign addr[27293] = -1890520410;
assign addr[27294] = -1899516021;
assign addr[27295] = -1908361011;
assign addr[27296] = -1917054681;
assign addr[27297] = -1925596340;
assign addr[27298] = -1933985310;
assign addr[27299] = -1942220928;
assign addr[27300] = -1950302539;
assign addr[27301] = -1958229503;
assign addr[27302] = -1966001192;
assign addr[27303] = -1973616989;
assign addr[27304] = -1981076290;
assign addr[27305] = -1988378503;
assign addr[27306] = -1995523051;
assign addr[27307] = -2002509365;
assign addr[27308] = -2009336893;
assign addr[27309] = -2016005093;
assign addr[27310] = -2022513436;
assign addr[27311] = -2028861406;
assign addr[27312] = -2035048499;
assign addr[27313] = -2041074226;
assign addr[27314] = -2046938108;
assign addr[27315] = -2052639680;
assign addr[27316] = -2058178491;
assign addr[27317] = -2063554100;
assign addr[27318] = -2068766083;
assign addr[27319] = -2073814024;
assign addr[27320] = -2078697525;
assign addr[27321] = -2083416198;
assign addr[27322] = -2087969669;
assign addr[27323] = -2092357577;
assign addr[27324] = -2096579573;
assign addr[27325] = -2100635323;
assign addr[27326] = -2104524506;
assign addr[27327] = -2108246813;
assign addr[27328] = -2111801949;
assign addr[27329] = -2115189632;
assign addr[27330] = -2118409593;
assign addr[27331] = -2121461578;
assign addr[27332] = -2124345343;
assign addr[27333] = -2127060661;
assign addr[27334] = -2129607316;
assign addr[27335] = -2131985106;
assign addr[27336] = -2134193842;
assign addr[27337] = -2136233350;
assign addr[27338] = -2138103468;
assign addr[27339] = -2139804048;
assign addr[27340] = -2141334954;
assign addr[27341] = -2142696065;
assign addr[27342] = -2143887273;
assign addr[27343] = -2144908484;
assign addr[27344] = -2145759618;
assign addr[27345] = -2146440605;
assign addr[27346] = -2146951393;
assign addr[27347] = -2147291941;
assign addr[27348] = -2147462221;
assign addr[27349] = -2147462221;
assign addr[27350] = -2147291941;
assign addr[27351] = -2146951393;
assign addr[27352] = -2146440605;
assign addr[27353] = -2145759618;
assign addr[27354] = -2144908484;
assign addr[27355] = -2143887273;
assign addr[27356] = -2142696065;
assign addr[27357] = -2141334954;
assign addr[27358] = -2139804048;
assign addr[27359] = -2138103468;
assign addr[27360] = -2136233350;
assign addr[27361] = -2134193842;
assign addr[27362] = -2131985106;
assign addr[27363] = -2129607316;
assign addr[27364] = -2127060661;
assign addr[27365] = -2124345343;
assign addr[27366] = -2121461578;
assign addr[27367] = -2118409593;
assign addr[27368] = -2115189632;
assign addr[27369] = -2111801949;
assign addr[27370] = -2108246813;
assign addr[27371] = -2104524506;
assign addr[27372] = -2100635323;
assign addr[27373] = -2096579573;
assign addr[27374] = -2092357577;
assign addr[27375] = -2087969669;
assign addr[27376] = -2083416198;
assign addr[27377] = -2078697525;
assign addr[27378] = -2073814024;
assign addr[27379] = -2068766083;
assign addr[27380] = -2063554100;
assign addr[27381] = -2058178491;
assign addr[27382] = -2052639680;
assign addr[27383] = -2046938108;
assign addr[27384] = -2041074226;
assign addr[27385] = -2035048499;
assign addr[27386] = -2028861406;
assign addr[27387] = -2022513436;
assign addr[27388] = -2016005093;
assign addr[27389] = -2009336893;
assign addr[27390] = -2002509365;
assign addr[27391] = -1995523051;
assign addr[27392] = -1988378503;
assign addr[27393] = -1981076290;
assign addr[27394] = -1973616989;
assign addr[27395] = -1966001192;
assign addr[27396] = -1958229503;
assign addr[27397] = -1950302539;
assign addr[27398] = -1942220928;
assign addr[27399] = -1933985310;
assign addr[27400] = -1925596340;
assign addr[27401] = -1917054681;
assign addr[27402] = -1908361011;
assign addr[27403] = -1899516021;
assign addr[27404] = -1890520410;
assign addr[27405] = -1881374892;
assign addr[27406] = -1872080193;
assign addr[27407] = -1862637049;
assign addr[27408] = -1853046210;
assign addr[27409] = -1843308435;
assign addr[27410] = -1833424497;
assign addr[27411] = -1823395180;
assign addr[27412] = -1813221279;
assign addr[27413] = -1802903601;
assign addr[27414] = -1792442963;
assign addr[27415] = -1781840195;
assign addr[27416] = -1771096139;
assign addr[27417] = -1760211645;
assign addr[27418] = -1749187577;
assign addr[27419] = -1738024810;
assign addr[27420] = -1726724227;
assign addr[27421] = -1715286726;
assign addr[27422] = -1703713213;
assign addr[27423] = -1692004606;
assign addr[27424] = -1680161834;
assign addr[27425] = -1668185835;
assign addr[27426] = -1656077559;
assign addr[27427] = -1643837966;
assign addr[27428] = -1631468027;
assign addr[27429] = -1618968722;
assign addr[27430] = -1606341043;
assign addr[27431] = -1593585992;
assign addr[27432] = -1580704578;
assign addr[27433] = -1567697824;
assign addr[27434] = -1554566762;
assign addr[27435] = -1541312431;
assign addr[27436] = -1527935884;
assign addr[27437] = -1514438181;
assign addr[27438] = -1500820393;
assign addr[27439] = -1487083598;
assign addr[27440] = -1473228887;
assign addr[27441] = -1459257358;
assign addr[27442] = -1445170118;
assign addr[27443] = -1430968286;
assign addr[27444] = -1416652986;
assign addr[27445] = -1402225355;
assign addr[27446] = -1387686535;
assign addr[27447] = -1373037681;
assign addr[27448] = -1358279953;
assign addr[27449] = -1343414522;
assign addr[27450] = -1328442566;
assign addr[27451] = -1313365273;
assign addr[27452] = -1298183838;
assign addr[27453] = -1282899464;
assign addr[27454] = -1267513365;
assign addr[27455] = -1252026760;
assign addr[27456] = -1236440877;
assign addr[27457] = -1220756951;
assign addr[27458] = -1204976227;
assign addr[27459] = -1189099956;
assign addr[27460] = -1173129396;
assign addr[27461] = -1157065814;
assign addr[27462] = -1140910484;
assign addr[27463] = -1124664687;
assign addr[27464] = -1108329711;
assign addr[27465] = -1091906851;
assign addr[27466] = -1075397409;
assign addr[27467] = -1058802695;
assign addr[27468] = -1042124025;
assign addr[27469] = -1025362720;
assign addr[27470] = -1008520110;
assign addr[27471] = -991597531;
assign addr[27472] = -974596324;
assign addr[27473] = -957517838;
assign addr[27474] = -940363427;
assign addr[27475] = -923134450;
assign addr[27476] = -905832274;
assign addr[27477] = -888458272;
assign addr[27478] = -871013820;
assign addr[27479] = -853500302;
assign addr[27480] = -835919107;
assign addr[27481] = -818271628;
assign addr[27482] = -800559266;
assign addr[27483] = -782783424;
assign addr[27484] = -764945512;
assign addr[27485] = -747046944;
assign addr[27486] = -729089140;
assign addr[27487] = -711073524;
assign addr[27488] = -693001525;
assign addr[27489] = -674874574;
assign addr[27490] = -656694110;
assign addr[27491] = -638461574;
assign addr[27492] = -620178412;
assign addr[27493] = -601846074;
assign addr[27494] = -583466013;
assign addr[27495] = -565039687;
assign addr[27496] = -546568556;
assign addr[27497] = -528054086;
assign addr[27498] = -509497745;
assign addr[27499] = -490901003;
assign addr[27500] = -472265336;
assign addr[27501] = -453592221;
assign addr[27502] = -434883140;
assign addr[27503] = -416139574;
assign addr[27504] = -397363011;
assign addr[27505] = -378554940;
assign addr[27506] = -359716852;
assign addr[27507] = -340850240;
assign addr[27508] = -321956601;
assign addr[27509] = -303037433;
assign addr[27510] = -284094236;
assign addr[27511] = -265128512;
assign addr[27512] = -246141764;
assign addr[27513] = -227135500;
assign addr[27514] = -208111224;
assign addr[27515] = -189070447;
assign addr[27516] = -170014678;
assign addr[27517] = -150945428;
assign addr[27518] = -131864208;
assign addr[27519] = -112772533;
assign addr[27520] = -93671915;
assign addr[27521] = -74563870;
assign addr[27522] = -55449912;
assign addr[27523] = -36331557;
assign addr[27524] = -17210322;
assign addr[27525] = 1912278;
assign addr[27526] = 21034727;
assign addr[27527] = 40155507;
assign addr[27528] = 59273104;
assign addr[27529] = 78386000;
assign addr[27530] = 97492681;
assign addr[27531] = 116591632;
assign addr[27532] = 135681337;
assign addr[27533] = 154760284;
assign addr[27534] = 173826959;
assign addr[27535] = 192879850;
assign addr[27536] = 211917448;
assign addr[27537] = 230938242;
assign addr[27538] = 249940723;
assign addr[27539] = 268923386;
assign addr[27540] = 287884725;
assign addr[27541] = 306823237;
assign addr[27542] = 325737419;
assign addr[27543] = 344625773;
assign addr[27544] = 363486799;
assign addr[27545] = 382319004;
assign addr[27546] = 401120892;
assign addr[27547] = 419890975;
assign addr[27548] = 438627762;
assign addr[27549] = 457329769;
assign addr[27550] = 475995513;
assign addr[27551] = 494623513;
assign addr[27552] = 513212292;
assign addr[27553] = 531760377;
assign addr[27554] = 550266296;
assign addr[27555] = 568728583;
assign addr[27556] = 587145773;
assign addr[27557] = 605516406;
assign addr[27558] = 623839025;
assign addr[27559] = 642112178;
assign addr[27560] = 660334415;
assign addr[27561] = 678504291;
assign addr[27562] = 696620367;
assign addr[27563] = 714681204;
assign addr[27564] = 732685372;
assign addr[27565] = 750631442;
assign addr[27566] = 768517992;
assign addr[27567] = 786343603;
assign addr[27568] = 804106861;
assign addr[27569] = 821806359;
assign addr[27570] = 839440693;
assign addr[27571] = 857008464;
assign addr[27572] = 874508280;
assign addr[27573] = 891938752;
assign addr[27574] = 909298500;
assign addr[27575] = 926586145;
assign addr[27576] = 943800318;
assign addr[27577] = 960939653;
assign addr[27578] = 978002791;
assign addr[27579] = 994988380;
assign addr[27580] = 1011895073;
assign addr[27581] = 1028721528;
assign addr[27582] = 1045466412;
assign addr[27583] = 1062128397;
assign addr[27584] = 1078706161;
assign addr[27585] = 1095198391;
assign addr[27586] = 1111603778;
assign addr[27587] = 1127921022;
assign addr[27588] = 1144148829;
assign addr[27589] = 1160285911;
assign addr[27590] = 1176330990;
assign addr[27591] = 1192282793;
assign addr[27592] = 1208140056;
assign addr[27593] = 1223901520;
assign addr[27594] = 1239565936;
assign addr[27595] = 1255132063;
assign addr[27596] = 1270598665;
assign addr[27597] = 1285964516;
assign addr[27598] = 1301228398;
assign addr[27599] = 1316389101;
assign addr[27600] = 1331445422;
assign addr[27601] = 1346396168;
assign addr[27602] = 1361240152;
assign addr[27603] = 1375976199;
assign addr[27604] = 1390603139;
assign addr[27605] = 1405119813;
assign addr[27606] = 1419525069;
assign addr[27607] = 1433817766;
assign addr[27608] = 1447996770;
assign addr[27609] = 1462060956;
assign addr[27610] = 1476009210;
assign addr[27611] = 1489840425;
assign addr[27612] = 1503553506;
assign addr[27613] = 1517147363;
assign addr[27614] = 1530620920;
assign addr[27615] = 1543973108;
assign addr[27616] = 1557202869;
assign addr[27617] = 1570309153;
assign addr[27618] = 1583290921;
assign addr[27619] = 1596147143;
assign addr[27620] = 1608876801;
assign addr[27621] = 1621478885;
assign addr[27622] = 1633952396;
assign addr[27623] = 1646296344;
assign addr[27624] = 1658509750;
assign addr[27625] = 1670591647;
assign addr[27626] = 1682541077;
assign addr[27627] = 1694357091;
assign addr[27628] = 1706038753;
assign addr[27629] = 1717585136;
assign addr[27630] = 1728995326;
assign addr[27631] = 1740268417;
assign addr[27632] = 1751403515;
assign addr[27633] = 1762399737;
assign addr[27634] = 1773256212;
assign addr[27635] = 1783972079;
assign addr[27636] = 1794546487;
assign addr[27637] = 1804978599;
assign addr[27638] = 1815267588;
assign addr[27639] = 1825412636;
assign addr[27640] = 1835412941;
assign addr[27641] = 1845267708;
assign addr[27642] = 1854976157;
assign addr[27643] = 1864537518;
assign addr[27644] = 1873951032;
assign addr[27645] = 1883215953;
assign addr[27646] = 1892331547;
assign addr[27647] = 1901297091;
assign addr[27648] = 1910111873;
assign addr[27649] = 1918775195;
assign addr[27650] = 1927286370;
assign addr[27651] = 1935644723;
assign addr[27652] = 1943849591;
assign addr[27653] = 1951900324;
assign addr[27654] = 1959796283;
assign addr[27655] = 1967536842;
assign addr[27656] = 1975121388;
assign addr[27657] = 1982549318;
assign addr[27658] = 1989820044;
assign addr[27659] = 1996932990;
assign addr[27660] = 2003887591;
assign addr[27661] = 2010683297;
assign addr[27662] = 2017319567;
assign addr[27663] = 2023795876;
assign addr[27664] = 2030111710;
assign addr[27665] = 2036266570;
assign addr[27666] = 2042259965;
assign addr[27667] = 2048091422;
assign addr[27668] = 2053760478;
assign addr[27669] = 2059266683;
assign addr[27670] = 2064609600;
assign addr[27671] = 2069788807;
assign addr[27672] = 2074803892;
assign addr[27673] = 2079654458;
assign addr[27674] = 2084340120;
assign addr[27675] = 2088860507;
assign addr[27676] = 2093215260;
assign addr[27677] = 2097404033;
assign addr[27678] = 2101426496;
assign addr[27679] = 2105282327;
assign addr[27680] = 2108971223;
assign addr[27681] = 2112492891;
assign addr[27682] = 2115847050;
assign addr[27683] = 2119033436;
assign addr[27684] = 2122051796;
assign addr[27685] = 2124901890;
assign addr[27686] = 2127583492;
assign addr[27687] = 2130096389;
assign addr[27688] = 2132440383;
assign addr[27689] = 2134615288;
assign addr[27690] = 2136620930;
assign addr[27691] = 2138457152;
assign addr[27692] = 2140123807;
assign addr[27693] = 2141620763;
assign addr[27694] = 2142947902;
assign addr[27695] = 2144105118;
assign addr[27696] = 2145092320;
assign addr[27697] = 2145909429;
assign addr[27698] = 2146556380;
assign addr[27699] = 2147033123;
assign addr[27700] = 2147339619;
assign addr[27701] = 2147475844;
assign addr[27702] = 2147441787;
assign addr[27703] = 2147237452;
assign addr[27704] = 2146862854;
assign addr[27705] = 2146318022;
assign addr[27706] = 2145603001;
assign addr[27707] = 2144717846;
assign addr[27708] = 2143662628;
assign addr[27709] = 2142437431;
assign addr[27710] = 2141042352;
assign addr[27711] = 2139477502;
assign addr[27712] = 2137743003;
assign addr[27713] = 2135838995;
assign addr[27714] = 2133765628;
assign addr[27715] = 2131523066;
assign addr[27716] = 2129111488;
assign addr[27717] = 2126531084;
assign addr[27718] = 2123782059;
assign addr[27719] = 2120864631;
assign addr[27720] = 2117779031;
assign addr[27721] = 2114525505;
assign addr[27722] = 2111104309;
assign addr[27723] = 2107515716;
assign addr[27724] = 2103760010;
assign addr[27725] = 2099837489;
assign addr[27726] = 2095748463;
assign addr[27727] = 2091493257;
assign addr[27728] = 2087072209;
assign addr[27729] = 2082485668;
assign addr[27730] = 2077733999;
assign addr[27731] = 2072817579;
assign addr[27732] = 2067736796;
assign addr[27733] = 2062492055;
assign addr[27734] = 2057083771;
assign addr[27735] = 2051512372;
assign addr[27736] = 2045778302;
assign addr[27737] = 2039882013;
assign addr[27738] = 2033823974;
assign addr[27739] = 2027604666;
assign addr[27740] = 2021224581;
assign addr[27741] = 2014684225;
assign addr[27742] = 2007984117;
assign addr[27743] = 2001124788;
assign addr[27744] = 1994106782;
assign addr[27745] = 1986930656;
assign addr[27746] = 1979596978;
assign addr[27747] = 1972106330;
assign addr[27748] = 1964459306;
assign addr[27749] = 1956656513;
assign addr[27750] = 1948698568;
assign addr[27751] = 1940586104;
assign addr[27752] = 1932319763;
assign addr[27753] = 1923900201;
assign addr[27754] = 1915328086;
assign addr[27755] = 1906604097;
assign addr[27756] = 1897728925;
assign addr[27757] = 1888703276;
assign addr[27758] = 1879527863;
assign addr[27759] = 1870203416;
assign addr[27760] = 1860730673;
assign addr[27761] = 1851110385;
assign addr[27762] = 1841343316;
assign addr[27763] = 1831430239;
assign addr[27764] = 1821371941;
assign addr[27765] = 1811169220;
assign addr[27766] = 1800822883;
assign addr[27767] = 1790333753;
assign addr[27768] = 1779702660;
assign addr[27769] = 1768930447;
assign addr[27770] = 1758017969;
assign addr[27771] = 1746966091;
assign addr[27772] = 1735775690;
assign addr[27773] = 1724447652;
assign addr[27774] = 1712982875;
assign addr[27775] = 1701382270;
assign addr[27776] = 1689646755;
assign addr[27777] = 1677777262;
assign addr[27778] = 1665774731;
assign addr[27779] = 1653640115;
assign addr[27780] = 1641374375;
assign addr[27781] = 1628978484;
assign addr[27782] = 1616453425;
assign addr[27783] = 1603800191;
assign addr[27784] = 1591019785;
assign addr[27785] = 1578113222;
assign addr[27786] = 1565081523;
assign addr[27787] = 1551925723;
assign addr[27788] = 1538646865;
assign addr[27789] = 1525246002;
assign addr[27790] = 1511724196;
assign addr[27791] = 1498082520;
assign addr[27792] = 1484322054;
assign addr[27793] = 1470443891;
assign addr[27794] = 1456449131;
assign addr[27795] = 1442338884;
assign addr[27796] = 1428114267;
assign addr[27797] = 1413776410;
assign addr[27798] = 1399326449;
assign addr[27799] = 1384765530;
assign addr[27800] = 1370094808;
assign addr[27801] = 1355315445;
assign addr[27802] = 1340428615;
assign addr[27803] = 1325435496;
assign addr[27804] = 1310337279;
assign addr[27805] = 1295135159;
assign addr[27806] = 1279830344;
assign addr[27807] = 1264424045;
assign addr[27808] = 1248917486;
assign addr[27809] = 1233311895;
assign addr[27810] = 1217608510;
assign addr[27811] = 1201808576;
assign addr[27812] = 1185913346;
assign addr[27813] = 1169924081;
assign addr[27814] = 1153842047;
assign addr[27815] = 1137668521;
assign addr[27816] = 1121404785;
assign addr[27817] = 1105052128;
assign addr[27818] = 1088611847;
assign addr[27819] = 1072085246;
assign addr[27820] = 1055473635;
assign addr[27821] = 1038778332;
assign addr[27822] = 1022000660;
assign addr[27823] = 1005141949;
assign addr[27824] = 988203537;
assign addr[27825] = 971186766;
assign addr[27826] = 954092986;
assign addr[27827] = 936923553;
assign addr[27828] = 919679827;
assign addr[27829] = 902363176;
assign addr[27830] = 884974973;
assign addr[27831] = 867516597;
assign addr[27832] = 849989433;
assign addr[27833] = 832394869;
assign addr[27834] = 814734301;
assign addr[27835] = 797009130;
assign addr[27836] = 779220762;
assign addr[27837] = 761370605;
assign addr[27838] = 743460077;
assign addr[27839] = 725490597;
assign addr[27840] = 707463589;
assign addr[27841] = 689380485;
assign addr[27842] = 671242716;
assign addr[27843] = 653051723;
assign addr[27844] = 634808946;
assign addr[27845] = 616515832;
assign addr[27846] = 598173833;
assign addr[27847] = 579784402;
assign addr[27848] = 561348998;
assign addr[27849] = 542869083;
assign addr[27850] = 524346121;
assign addr[27851] = 505781581;
assign addr[27852] = 487176937;
assign addr[27853] = 468533662;
assign addr[27854] = 449853235;
assign addr[27855] = 431137138;
assign addr[27856] = 412386854;
assign addr[27857] = 393603870;
assign addr[27858] = 374789676;
assign addr[27859] = 355945764;
assign addr[27860] = 337073627;
assign addr[27861] = 318174762;
assign addr[27862] = 299250668;
assign addr[27863] = 280302845;
assign addr[27864] = 261332796;
assign addr[27865] = 242342025;
assign addr[27866] = 223332037;
assign addr[27867] = 204304341;
assign addr[27868] = 185260444;
assign addr[27869] = 166201858;
assign addr[27870] = 147130093;
assign addr[27871] = 128046661;
assign addr[27872] = 108953076;
assign addr[27873] = 89850852;
assign addr[27874] = 70741503;
assign addr[27875] = 51626544;
assign addr[27876] = 32507492;
assign addr[27877] = 13385863;
assign addr[27878] = -5736829;
assign addr[27879] = -24859065;
assign addr[27880] = -43979330;
assign addr[27881] = -63096108;
assign addr[27882] = -82207882;
assign addr[27883] = -101313138;
assign addr[27884] = -120410361;
assign addr[27885] = -139498035;
assign addr[27886] = -158574649;
assign addr[27887] = -177638688;
assign addr[27888] = -196688642;
assign addr[27889] = -215722999;
assign addr[27890] = -234740251;
assign addr[27891] = -253738890;
assign addr[27892] = -272717408;
assign addr[27893] = -291674302;
assign addr[27894] = -310608068;
assign addr[27895] = -329517204;
assign addr[27896] = -348400212;
assign addr[27897] = -367255594;
assign addr[27898] = -386081854;
assign addr[27899] = -404877501;
assign addr[27900] = -423641043;
assign addr[27901] = -442370993;
assign addr[27902] = -461065866;
assign addr[27903] = -479724180;
assign addr[27904] = -498344454;
assign addr[27905] = -516925212;
assign addr[27906] = -535464981;
assign addr[27907] = -553962291;
assign addr[27908] = -572415676;
assign addr[27909] = -590823671;
assign addr[27910] = -609184818;
assign addr[27911] = -627497660;
assign addr[27912] = -645760745;
assign addr[27913] = -663972625;
assign addr[27914] = -682131857;
assign addr[27915] = -700236999;
assign addr[27916] = -718286617;
assign addr[27917] = -736279279;
assign addr[27918] = -754213559;
assign addr[27919] = -772088034;
assign addr[27920] = -789901288;
assign addr[27921] = -807651907;
assign addr[27922] = -825338484;
assign addr[27923] = -842959617;
assign addr[27924] = -860513908;
assign addr[27925] = -877999966;
assign addr[27926] = -895416404;
assign addr[27927] = -912761841;
assign addr[27928] = -930034901;
assign addr[27929] = -947234215;
assign addr[27930] = -964358420;
assign addr[27931] = -981406156;
assign addr[27932] = -998376073;
assign addr[27933] = -1015266825;
assign addr[27934] = -1032077073;
assign addr[27935] = -1048805483;
assign addr[27936] = -1065450729;
assign addr[27937] = -1082011492;
assign addr[27938] = -1098486458;
assign addr[27939] = -1114874320;
assign addr[27940] = -1131173780;
assign addr[27941] = -1147383544;
assign addr[27942] = -1163502328;
assign addr[27943] = -1179528853;
assign addr[27944] = -1195461849;
assign addr[27945] = -1211300053;
assign addr[27946] = -1227042207;
assign addr[27947] = -1242687064;
assign addr[27948] = -1258233384;
assign addr[27949] = -1273679934;
assign addr[27950] = -1289025489;
assign addr[27951] = -1304268832;
assign addr[27952] = -1319408754;
assign addr[27953] = -1334444055;
assign addr[27954] = -1349373543;
assign addr[27955] = -1364196034;
assign addr[27956] = -1378910353;
assign addr[27957] = -1393515332;
assign addr[27958] = -1408009814;
assign addr[27959] = -1422392650;
assign addr[27960] = -1436662698;
assign addr[27961] = -1450818828;
assign addr[27962] = -1464859917;
assign addr[27963] = -1478784851;
assign addr[27964] = -1492592527;
assign addr[27965] = -1506281850;
assign addr[27966] = -1519851733;
assign addr[27967] = -1533301101;
assign addr[27968] = -1546628888;
assign addr[27969] = -1559834037;
assign addr[27970] = -1572915501;
assign addr[27971] = -1585872242;
assign addr[27972] = -1598703233;
assign addr[27973] = -1611407456;
assign addr[27974] = -1623983905;
assign addr[27975] = -1636431582;
assign addr[27976] = -1648749499;
assign addr[27977] = -1660936681;
assign addr[27978] = -1672992161;
assign addr[27979] = -1684914983;
assign addr[27980] = -1696704201;
assign addr[27981] = -1708358881;
assign addr[27982] = -1719878099;
assign addr[27983] = -1731260941;
assign addr[27984] = -1742506504;
assign addr[27985] = -1753613897;
assign addr[27986] = -1764582240;
assign addr[27987] = -1775410662;
assign addr[27988] = -1786098304;
assign addr[27989] = -1796644320;
assign addr[27990] = -1807047873;
assign addr[27991] = -1817308138;
assign addr[27992] = -1827424302;
assign addr[27993] = -1837395562;
assign addr[27994] = -1847221128;
assign addr[27995] = -1856900221;
assign addr[27996] = -1866432072;
assign addr[27997] = -1875815927;
assign addr[27998] = -1885051042;
assign addr[27999] = -1894136683;
assign addr[28000] = -1903072131;
assign addr[28001] = -1911856677;
assign addr[28002] = -1920489624;
assign addr[28003] = -1928970288;
assign addr[28004] = -1937297997;
assign addr[28005] = -1945472089;
assign addr[28006] = -1953491918;
assign addr[28007] = -1961356847;
assign addr[28008] = -1969066252;
assign addr[28009] = -1976619522;
assign addr[28010] = -1984016058;
assign addr[28011] = -1991255274;
assign addr[28012] = -1998336596;
assign addr[28013] = -2005259462;
assign addr[28014] = -2012023322;
assign addr[28015] = -2018627642;
assign addr[28016] = -2025071897;
assign addr[28017] = -2031355576;
assign addr[28018] = -2037478181;
assign addr[28019] = -2043439226;
assign addr[28020] = -2049238240;
assign addr[28021] = -2054874761;
assign addr[28022] = -2060348343;
assign addr[28023] = -2065658552;
assign addr[28024] = -2070804967;
assign addr[28025] = -2075787180;
assign addr[28026] = -2080604795;
assign addr[28027] = -2085257431;
assign addr[28028] = -2089744719;
assign addr[28029] = -2094066304;
assign addr[28030] = -2098221841;
assign addr[28031] = -2102211002;
assign addr[28032] = -2106033471;
assign addr[28033] = -2109688944;
assign addr[28034] = -2113177132;
assign addr[28035] = -2116497758;
assign addr[28036] = -2119650558;
assign addr[28037] = -2122635283;
assign addr[28038] = -2125451696;
assign addr[28039] = -2128099574;
assign addr[28040] = -2130578706;
assign addr[28041] = -2132888897;
assign addr[28042] = -2135029962;
assign addr[28043] = -2137001733;
assign addr[28044] = -2138804053;
assign addr[28045] = -2140436778;
assign addr[28046] = -2141899780;
assign addr[28047] = -2143192942;
assign addr[28048] = -2144316162;
assign addr[28049] = -2145269351;
assign addr[28050] = -2146052433;
assign addr[28051] = -2146665347;
assign addr[28052] = -2147108043;
assign addr[28053] = -2147380486;
assign addr[28054] = -2147482655;
assign addr[28055] = -2147414542;
assign addr[28056] = -2147176152;
assign addr[28057] = -2146767505;
assign addr[28058] = -2146188631;
assign addr[28059] = -2145439578;
assign addr[28060] = -2144520405;
assign addr[28061] = -2143431184;
assign addr[28062] = -2142172003;
assign addr[28063] = -2140742960;
assign addr[28064] = -2139144169;
assign addr[28065] = -2137375758;
assign addr[28066] = -2135437865;
assign addr[28067] = -2133330646;
assign addr[28068] = -2131054266;
assign addr[28069] = -2128608907;
assign addr[28070] = -2125994762;
assign addr[28071] = -2123212038;
assign addr[28072] = -2120260957;
assign addr[28073] = -2117141752;
assign addr[28074] = -2113854671;
assign addr[28075] = -2110399974;
assign addr[28076] = -2106777935;
assign addr[28077] = -2102988841;
assign addr[28078] = -2099032994;
assign addr[28079] = -2094910706;
assign addr[28080] = -2090622304;
assign addr[28081] = -2086168128;
assign addr[28082] = -2081548533;
assign addr[28083] = -2076763883;
assign addr[28084] = -2071814558;
assign addr[28085] = -2066700952;
assign addr[28086] = -2061423468;
assign addr[28087] = -2055982526;
assign addr[28088] = -2050378558;
assign addr[28089] = -2044612007;
assign addr[28090] = -2038683330;
assign addr[28091] = -2032592999;
assign addr[28092] = -2026341495;
assign addr[28093] = -2019929315;
assign addr[28094] = -2013356967;
assign addr[28095] = -2006624971;
assign addr[28096] = -1999733863;
assign addr[28097] = -1992684188;
assign addr[28098] = -1985476506;
assign addr[28099] = -1978111387;
assign addr[28100] = -1970589416;
assign addr[28101] = -1962911189;
assign addr[28102] = -1955077316;
assign addr[28103] = -1947088417;
assign addr[28104] = -1938945125;
assign addr[28105] = -1930648088;
assign addr[28106] = -1922197961;
assign addr[28107] = -1913595416;
assign addr[28108] = -1904841135;
assign addr[28109] = -1895935811;
assign addr[28110] = -1886880151;
assign addr[28111] = -1877674873;
assign addr[28112] = -1868320707;
assign addr[28113] = -1858818395;
assign addr[28114] = -1849168689;
assign addr[28115] = -1839372356;
assign addr[28116] = -1829430172;
assign addr[28117] = -1819342925;
assign addr[28118] = -1809111415;
assign addr[28119] = -1798736454;
assign addr[28120] = -1788218865;
assign addr[28121] = -1777559480;
assign addr[28122] = -1766759146;
assign addr[28123] = -1755818718;
assign addr[28124] = -1744739065;
assign addr[28125] = -1733521064;
assign addr[28126] = -1722165606;
assign addr[28127] = -1710673591;
assign addr[28128] = -1699045930;
assign addr[28129] = -1687283545;
assign addr[28130] = -1675387369;
assign addr[28131] = -1663358344;
assign addr[28132] = -1651197426;
assign addr[28133] = -1638905577;
assign addr[28134] = -1626483774;
assign addr[28135] = -1613933000;
assign addr[28136] = -1601254251;
assign addr[28137] = -1588448533;
assign addr[28138] = -1575516860;
assign addr[28139] = -1562460258;
assign addr[28140] = -1549279763;
assign addr[28141] = -1535976419;
assign addr[28142] = -1522551282;
assign addr[28143] = -1509005416;
assign addr[28144] = -1495339895;
assign addr[28145] = -1481555802;
assign addr[28146] = -1467654232;
assign addr[28147] = -1453636285;
assign addr[28148] = -1439503074;
assign addr[28149] = -1425255719;
assign addr[28150] = -1410895350;
assign addr[28151] = -1396423105;
assign addr[28152] = -1381840133;
assign addr[28153] = -1367147589;
assign addr[28154] = -1352346639;
assign addr[28155] = -1337438456;
assign addr[28156] = -1322424222;
assign addr[28157] = -1307305128;
assign addr[28158] = -1292082373;
assign addr[28159] = -1276757164;
assign addr[28160] = -1261330715;
assign addr[28161] = -1245804251;
assign addr[28162] = -1230179002;
assign addr[28163] = -1214456207;
assign addr[28164] = -1198637114;
assign addr[28165] = -1182722976;
assign addr[28166] = -1166715055;
assign addr[28167] = -1150614620;
assign addr[28168] = -1134422949;
assign addr[28169] = -1118141326;
assign addr[28170] = -1101771040;
assign addr[28171] = -1085313391;
assign addr[28172] = -1068769683;
assign addr[28173] = -1052141228;
assign addr[28174] = -1035429345;
assign addr[28175] = -1018635358;
assign addr[28176] = -1001760600;
assign addr[28177] = -984806408;
assign addr[28178] = -967774128;
assign addr[28179] = -950665109;
assign addr[28180] = -933480707;
assign addr[28181] = -916222287;
assign addr[28182] = -898891215;
assign addr[28183] = -881488868;
assign addr[28184] = -864016623;
assign addr[28185] = -846475867;
assign addr[28186] = -828867991;
assign addr[28187] = -811194391;
assign addr[28188] = -793456467;
assign addr[28189] = -775655628;
assign addr[28190] = -757793284;
assign addr[28191] = -739870851;
assign addr[28192] = -721889752;
assign addr[28193] = -703851410;
assign addr[28194] = -685757258;
assign addr[28195] = -667608730;
assign addr[28196] = -649407264;
assign addr[28197] = -631154304;
assign addr[28198] = -612851297;
assign addr[28199] = -594499695;
assign addr[28200] = -576100953;
assign addr[28201] = -557656529;
assign addr[28202] = -539167887;
assign addr[28203] = -520636492;
assign addr[28204] = -502063814;
assign addr[28205] = -483451325;
assign addr[28206] = -464800501;
assign addr[28207] = -446112822;
assign addr[28208] = -427389768;
assign addr[28209] = -408632825;
assign addr[28210] = -389843480;
assign addr[28211] = -371023223;
assign addr[28212] = -352173546;
assign addr[28213] = -333295944;
assign addr[28214] = -314391913;
assign addr[28215] = -295462954;
assign addr[28216] = -276510565;
assign addr[28217] = -257536251;
assign addr[28218] = -238541516;
assign addr[28219] = -219527866;
assign addr[28220] = -200496809;
assign addr[28221] = -181449854;
assign addr[28222] = -162388511;
assign addr[28223] = -143314291;
assign addr[28224] = -124228708;
assign addr[28225] = -105133274;
assign addr[28226] = -86029503;
assign addr[28227] = -66918911;
assign addr[28228] = -47803013;
assign addr[28229] = -28683324;
assign addr[28230] = -9561361;
assign addr[28231] = 9561361;
assign addr[28232] = 28683324;
assign addr[28233] = 47803013;
assign addr[28234] = 66918911;
assign addr[28235] = 86029503;
assign addr[28236] = 105133274;
assign addr[28237] = 124228708;
assign addr[28238] = 143314291;
assign addr[28239] = 162388511;
assign addr[28240] = 181449854;
assign addr[28241] = 200496809;
assign addr[28242] = 219527866;
assign addr[28243] = 238541516;
assign addr[28244] = 257536251;
assign addr[28245] = 276510565;
assign addr[28246] = 295462953;
assign addr[28247] = 314391913;
assign addr[28248] = 333295944;
assign addr[28249] = 352173546;
assign addr[28250] = 371023223;
assign addr[28251] = 389843480;
assign addr[28252] = 408632825;
assign addr[28253] = 427389768;
assign addr[28254] = 446112822;
assign addr[28255] = 464800501;
assign addr[28256] = 483451325;
assign addr[28257] = 502063814;
assign addr[28258] = 520636492;
assign addr[28259] = 539167887;
assign addr[28260] = 557656529;
assign addr[28261] = 576100953;
assign addr[28262] = 594499695;
assign addr[28263] = 612851297;
assign addr[28264] = 631154304;
assign addr[28265] = 649407264;
assign addr[28266] = 667608730;
assign addr[28267] = 685757258;
assign addr[28268] = 703851410;
assign addr[28269] = 721889752;
assign addr[28270] = 739870851;
assign addr[28271] = 757793284;
assign addr[28272] = 775655628;
assign addr[28273] = 793456467;
assign addr[28274] = 811194391;
assign addr[28275] = 828867991;
assign addr[28276] = 846475867;
assign addr[28277] = 864016623;
assign addr[28278] = 881488868;
assign addr[28279] = 898891215;
assign addr[28280] = 916222287;
assign addr[28281] = 933480707;
assign addr[28282] = 950665109;
assign addr[28283] = 967774128;
assign addr[28284] = 984806408;
assign addr[28285] = 1001760600;
assign addr[28286] = 1018635358;
assign addr[28287] = 1035429345;
assign addr[28288] = 1052141228;
assign addr[28289] = 1068769683;
assign addr[28290] = 1085313391;
assign addr[28291] = 1101771040;
assign addr[28292] = 1118141326;
assign addr[28293] = 1134422949;
assign addr[28294] = 1150614620;
assign addr[28295] = 1166715055;
assign addr[28296] = 1182722976;
assign addr[28297] = 1198637114;
assign addr[28298] = 1214456207;
assign addr[28299] = 1230179002;
assign addr[28300] = 1245804251;
assign addr[28301] = 1261330715;
assign addr[28302] = 1276757164;
assign addr[28303] = 1292082373;
assign addr[28304] = 1307305128;
assign addr[28305] = 1322424222;
assign addr[28306] = 1337438456;
assign addr[28307] = 1352346639;
assign addr[28308] = 1367147589;
assign addr[28309] = 1381840133;
assign addr[28310] = 1396423105;
assign addr[28311] = 1410895350;
assign addr[28312] = 1425255719;
assign addr[28313] = 1439503074;
assign addr[28314] = 1453636285;
assign addr[28315] = 1467654232;
assign addr[28316] = 1481555802;
assign addr[28317] = 1495339895;
assign addr[28318] = 1509005416;
assign addr[28319] = 1522551282;
assign addr[28320] = 1535976419;
assign addr[28321] = 1549279763;
assign addr[28322] = 1562460258;
assign addr[28323] = 1575516860;
assign addr[28324] = 1588448533;
assign addr[28325] = 1601254251;
assign addr[28326] = 1613933000;
assign addr[28327] = 1626483774;
assign addr[28328] = 1638905577;
assign addr[28329] = 1651197426;
assign addr[28330] = 1663358344;
assign addr[28331] = 1675387369;
assign addr[28332] = 1687283545;
assign addr[28333] = 1699045930;
assign addr[28334] = 1710673591;
assign addr[28335] = 1722165606;
assign addr[28336] = 1733521064;
assign addr[28337] = 1744739065;
assign addr[28338] = 1755818718;
assign addr[28339] = 1766759146;
assign addr[28340] = 1777559480;
assign addr[28341] = 1788218865;
assign addr[28342] = 1798736454;
assign addr[28343] = 1809111415;
assign addr[28344] = 1819342925;
assign addr[28345] = 1829430172;
assign addr[28346] = 1839372356;
assign addr[28347] = 1849168689;
assign addr[28348] = 1858818395;
assign addr[28349] = 1868320707;
assign addr[28350] = 1877674873;
assign addr[28351] = 1886880151;
assign addr[28352] = 1895935811;
assign addr[28353] = 1904841135;
assign addr[28354] = 1913595416;
assign addr[28355] = 1922197961;
assign addr[28356] = 1930648088;
assign addr[28357] = 1938945125;
assign addr[28358] = 1947088417;
assign addr[28359] = 1955077316;
assign addr[28360] = 1962911189;
assign addr[28361] = 1970589416;
assign addr[28362] = 1978111387;
assign addr[28363] = 1985476506;
assign addr[28364] = 1992684188;
assign addr[28365] = 1999733863;
assign addr[28366] = 2006624971;
assign addr[28367] = 2013356967;
assign addr[28368] = 2019929315;
assign addr[28369] = 2026341495;
assign addr[28370] = 2032592999;
assign addr[28371] = 2038683330;
assign addr[28372] = 2044612007;
assign addr[28373] = 2050378558;
assign addr[28374] = 2055982526;
assign addr[28375] = 2061423468;
assign addr[28376] = 2066700952;
assign addr[28377] = 2071814558;
assign addr[28378] = 2076763883;
assign addr[28379] = 2081548533;
assign addr[28380] = 2086168128;
assign addr[28381] = 2090622304;
assign addr[28382] = 2094910706;
assign addr[28383] = 2099032994;
assign addr[28384] = 2102988841;
assign addr[28385] = 2106777935;
assign addr[28386] = 2110399974;
assign addr[28387] = 2113854671;
assign addr[28388] = 2117141752;
assign addr[28389] = 2120260957;
assign addr[28390] = 2123212038;
assign addr[28391] = 2125994762;
assign addr[28392] = 2128608907;
assign addr[28393] = 2131054266;
assign addr[28394] = 2133330646;
assign addr[28395] = 2135437865;
assign addr[28396] = 2137375758;
assign addr[28397] = 2139144169;
assign addr[28398] = 2140742960;
assign addr[28399] = 2142172003;
assign addr[28400] = 2143431184;
assign addr[28401] = 2144520405;
assign addr[28402] = 2145439578;
assign addr[28403] = 2146188631;
assign addr[28404] = 2146767505;
assign addr[28405] = 2147176152;
assign addr[28406] = 2147414542;
assign addr[28407] = 2147482655;
assign addr[28408] = 2147380486;
assign addr[28409] = 2147108043;
assign addr[28410] = 2146665347;
assign addr[28411] = 2146052433;
assign addr[28412] = 2145269351;
assign addr[28413] = 2144316162;
assign addr[28414] = 2143192942;
assign addr[28415] = 2141899780;
assign addr[28416] = 2140436778;
assign addr[28417] = 2138804053;
assign addr[28418] = 2137001733;
assign addr[28419] = 2135029962;
assign addr[28420] = 2132888897;
assign addr[28421] = 2130578706;
assign addr[28422] = 2128099574;
assign addr[28423] = 2125451696;
assign addr[28424] = 2122635283;
assign addr[28425] = 2119650558;
assign addr[28426] = 2116497758;
assign addr[28427] = 2113177132;
assign addr[28428] = 2109688944;
assign addr[28429] = 2106033471;
assign addr[28430] = 2102211002;
assign addr[28431] = 2098221841;
assign addr[28432] = 2094066304;
assign addr[28433] = 2089744719;
assign addr[28434] = 2085257431;
assign addr[28435] = 2080604795;
assign addr[28436] = 2075787180;
assign addr[28437] = 2070804967;
assign addr[28438] = 2065658552;
assign addr[28439] = 2060348343;
assign addr[28440] = 2054874761;
assign addr[28441] = 2049238240;
assign addr[28442] = 2043439226;
assign addr[28443] = 2037478181;
assign addr[28444] = 2031355576;
assign addr[28445] = 2025071897;
assign addr[28446] = 2018627642;
assign addr[28447] = 2012023322;
assign addr[28448] = 2005259462;
assign addr[28449] = 1998336596;
assign addr[28450] = 1991255274;
assign addr[28451] = 1984016058;
assign addr[28452] = 1976619522;
assign addr[28453] = 1969066252;
assign addr[28454] = 1961356847;
assign addr[28455] = 1953491918;
assign addr[28456] = 1945472089;
assign addr[28457] = 1937297997;
assign addr[28458] = 1928970288;
assign addr[28459] = 1920489624;
assign addr[28460] = 1911856677;
assign addr[28461] = 1903072131;
assign addr[28462] = 1894136683;
assign addr[28463] = 1885051042;
assign addr[28464] = 1875815927;
assign addr[28465] = 1866432072;
assign addr[28466] = 1856900221;
assign addr[28467] = 1847221128;
assign addr[28468] = 1837395562;
assign addr[28469] = 1827424302;
assign addr[28470] = 1817308138;
assign addr[28471] = 1807047873;
assign addr[28472] = 1796644320;
assign addr[28473] = 1786098304;
assign addr[28474] = 1775410662;
assign addr[28475] = 1764582240;
assign addr[28476] = 1753613897;
assign addr[28477] = 1742506504;
assign addr[28478] = 1731260941;
assign addr[28479] = 1719878099;
assign addr[28480] = 1708358881;
assign addr[28481] = 1696704201;
assign addr[28482] = 1684914983;
assign addr[28483] = 1672992161;
assign addr[28484] = 1660936681;
assign addr[28485] = 1648749499;
assign addr[28486] = 1636431582;
assign addr[28487] = 1623983905;
assign addr[28488] = 1611407456;
assign addr[28489] = 1598703233;
assign addr[28490] = 1585872242;
assign addr[28491] = 1572915501;
assign addr[28492] = 1559834037;
assign addr[28493] = 1546628888;
assign addr[28494] = 1533301101;
assign addr[28495] = 1519851733;
assign addr[28496] = 1506281850;
assign addr[28497] = 1492592527;
assign addr[28498] = 1478784851;
assign addr[28499] = 1464859917;
assign addr[28500] = 1450818828;
assign addr[28501] = 1436662698;
assign addr[28502] = 1422392650;
assign addr[28503] = 1408009814;
assign addr[28504] = 1393515332;
assign addr[28505] = 1378910353;
assign addr[28506] = 1364196034;
assign addr[28507] = 1349373543;
assign addr[28508] = 1334444055;
assign addr[28509] = 1319408754;
assign addr[28510] = 1304268832;
assign addr[28511] = 1289025489;
assign addr[28512] = 1273679934;
assign addr[28513] = 1258233384;
assign addr[28514] = 1242687064;
assign addr[28515] = 1227042207;
assign addr[28516] = 1211300053;
assign addr[28517] = 1195461849;
assign addr[28518] = 1179528853;
assign addr[28519] = 1163502328;
assign addr[28520] = 1147383544;
assign addr[28521] = 1131173780;
assign addr[28522] = 1114874320;
assign addr[28523] = 1098486458;
assign addr[28524] = 1082011492;
assign addr[28525] = 1065450729;
assign addr[28526] = 1048805483;
assign addr[28527] = 1032077073;
assign addr[28528] = 1015266825;
assign addr[28529] = 998376073;
assign addr[28530] = 981406156;
assign addr[28531] = 964358420;
assign addr[28532] = 947234215;
assign addr[28533] = 930034901;
assign addr[28534] = 912761841;
assign addr[28535] = 895416404;
assign addr[28536] = 877999966;
assign addr[28537] = 860513908;
assign addr[28538] = 842959617;
assign addr[28539] = 825338484;
assign addr[28540] = 807651907;
assign addr[28541] = 789901288;
assign addr[28542] = 772088034;
assign addr[28543] = 754213559;
assign addr[28544] = 736279279;
assign addr[28545] = 718286617;
assign addr[28546] = 700236999;
assign addr[28547] = 682131857;
assign addr[28548] = 663972625;
assign addr[28549] = 645760745;
assign addr[28550] = 627497660;
assign addr[28551] = 609184818;
assign addr[28552] = 590823671;
assign addr[28553] = 572415676;
assign addr[28554] = 553962291;
assign addr[28555] = 535464981;
assign addr[28556] = 516925212;
assign addr[28557] = 498344454;
assign addr[28558] = 479724180;
assign addr[28559] = 461065866;
assign addr[28560] = 442370993;
assign addr[28561] = 423641043;
assign addr[28562] = 404877501;
assign addr[28563] = 386081854;
assign addr[28564] = 367255594;
assign addr[28565] = 348400212;
assign addr[28566] = 329517204;
assign addr[28567] = 310608068;
assign addr[28568] = 291674302;
assign addr[28569] = 272717408;
assign addr[28570] = 253738890;
assign addr[28571] = 234740251;
assign addr[28572] = 215722999;
assign addr[28573] = 196688642;
assign addr[28574] = 177638688;
assign addr[28575] = 158574649;
assign addr[28576] = 139498035;
assign addr[28577] = 120410361;
assign addr[28578] = 101313138;
assign addr[28579] = 82207882;
assign addr[28580] = 63096108;
assign addr[28581] = 43979330;
assign addr[28582] = 24859065;
assign addr[28583] = 5736829;
assign addr[28584] = -13385863;
assign addr[28585] = -32507492;
assign addr[28586] = -51626544;
assign addr[28587] = -70741503;
assign addr[28588] = -89850852;
assign addr[28589] = -108953076;
assign addr[28590] = -128046661;
assign addr[28591] = -147130093;
assign addr[28592] = -166201858;
assign addr[28593] = -185260444;
assign addr[28594] = -204304341;
assign addr[28595] = -223332037;
assign addr[28596] = -242342025;
assign addr[28597] = -261332796;
assign addr[28598] = -280302845;
assign addr[28599] = -299250668;
assign addr[28600] = -318174762;
assign addr[28601] = -337073627;
assign addr[28602] = -355945764;
assign addr[28603] = -374789676;
assign addr[28604] = -393603870;
assign addr[28605] = -412386854;
assign addr[28606] = -431137138;
assign addr[28607] = -449853235;
assign addr[28608] = -468533662;
assign addr[28609] = -487176937;
assign addr[28610] = -505781581;
assign addr[28611] = -524346121;
assign addr[28612] = -542869083;
assign addr[28613] = -561348998;
assign addr[28614] = -579784402;
assign addr[28615] = -598173833;
assign addr[28616] = -616515832;
assign addr[28617] = -634808946;
assign addr[28618] = -653051723;
assign addr[28619] = -671242716;
assign addr[28620] = -689380485;
assign addr[28621] = -707463589;
assign addr[28622] = -725490597;
assign addr[28623] = -743460077;
assign addr[28624] = -761370605;
assign addr[28625] = -779220762;
assign addr[28626] = -797009130;
assign addr[28627] = -814734301;
assign addr[28628] = -832394869;
assign addr[28629] = -849989433;
assign addr[28630] = -867516597;
assign addr[28631] = -884974973;
assign addr[28632] = -902363176;
assign addr[28633] = -919679827;
assign addr[28634] = -936923553;
assign addr[28635] = -954092986;
assign addr[28636] = -971186766;
assign addr[28637] = -988203537;
assign addr[28638] = -1005141949;
assign addr[28639] = -1022000660;
assign addr[28640] = -1038778332;
assign addr[28641] = -1055473635;
assign addr[28642] = -1072085246;
assign addr[28643] = -1088611847;
assign addr[28644] = -1105052128;
assign addr[28645] = -1121404785;
assign addr[28646] = -1137668521;
assign addr[28647] = -1153842047;
assign addr[28648] = -1169924081;
assign addr[28649] = -1185913346;
assign addr[28650] = -1201808576;
assign addr[28651] = -1217608510;
assign addr[28652] = -1233311895;
assign addr[28653] = -1248917486;
assign addr[28654] = -1264424045;
assign addr[28655] = -1279830344;
assign addr[28656] = -1295135159;
assign addr[28657] = -1310337279;
assign addr[28658] = -1325435496;
assign addr[28659] = -1340428615;
assign addr[28660] = -1355315445;
assign addr[28661] = -1370094808;
assign addr[28662] = -1384765530;
assign addr[28663] = -1399326449;
assign addr[28664] = -1413776410;
assign addr[28665] = -1428114267;
assign addr[28666] = -1442338884;
assign addr[28667] = -1456449131;
assign addr[28668] = -1470443891;
assign addr[28669] = -1484322054;
assign addr[28670] = -1498082520;
assign addr[28671] = -1511724196;
assign addr[28672] = -1525246002;
assign addr[28673] = -1538646865;
assign addr[28674] = -1551925723;
assign addr[28675] = -1565081523;
assign addr[28676] = -1578113222;
assign addr[28677] = -1591019785;
assign addr[28678] = -1603800191;
assign addr[28679] = -1616453425;
assign addr[28680] = -1628978484;
assign addr[28681] = -1641374375;
assign addr[28682] = -1653640115;
assign addr[28683] = -1665774731;
assign addr[28684] = -1677777262;
assign addr[28685] = -1689646755;
assign addr[28686] = -1701382270;
assign addr[28687] = -1712982875;
assign addr[28688] = -1724447652;
assign addr[28689] = -1735775690;
assign addr[28690] = -1746966091;
assign addr[28691] = -1758017969;
assign addr[28692] = -1768930447;
assign addr[28693] = -1779702660;
assign addr[28694] = -1790333753;
assign addr[28695] = -1800822883;
assign addr[28696] = -1811169220;
assign addr[28697] = -1821371941;
assign addr[28698] = -1831430239;
assign addr[28699] = -1841343316;
assign addr[28700] = -1851110385;
assign addr[28701] = -1860730673;
assign addr[28702] = -1870203416;
assign addr[28703] = -1879527863;
assign addr[28704] = -1888703276;
assign addr[28705] = -1897728925;
assign addr[28706] = -1906604097;
assign addr[28707] = -1915328086;
assign addr[28708] = -1923900201;
assign addr[28709] = -1932319763;
assign addr[28710] = -1940586104;
assign addr[28711] = -1948698568;
assign addr[28712] = -1956656513;
assign addr[28713] = -1964459306;
assign addr[28714] = -1972106330;
assign addr[28715] = -1979596978;
assign addr[28716] = -1986930656;
assign addr[28717] = -1994106782;
assign addr[28718] = -2001124788;
assign addr[28719] = -2007984117;
assign addr[28720] = -2014684225;
assign addr[28721] = -2021224581;
assign addr[28722] = -2027604666;
assign addr[28723] = -2033823974;
assign addr[28724] = -2039882013;
assign addr[28725] = -2045778302;
assign addr[28726] = -2051512372;
assign addr[28727] = -2057083771;
assign addr[28728] = -2062492055;
assign addr[28729] = -2067736796;
assign addr[28730] = -2072817579;
assign addr[28731] = -2077733999;
assign addr[28732] = -2082485668;
assign addr[28733] = -2087072209;
assign addr[28734] = -2091493257;
assign addr[28735] = -2095748463;
assign addr[28736] = -2099837489;
assign addr[28737] = -2103760010;
assign addr[28738] = -2107515716;
assign addr[28739] = -2111104309;
assign addr[28740] = -2114525505;
assign addr[28741] = -2117779031;
assign addr[28742] = -2120864631;
assign addr[28743] = -2123782059;
assign addr[28744] = -2126531084;
assign addr[28745] = -2129111488;
assign addr[28746] = -2131523066;
assign addr[28747] = -2133765628;
assign addr[28748] = -2135838995;
assign addr[28749] = -2137743003;
assign addr[28750] = -2139477502;
assign addr[28751] = -2141042352;
assign addr[28752] = -2142437431;
assign addr[28753] = -2143662628;
assign addr[28754] = -2144717846;
assign addr[28755] = -2145603001;
assign addr[28756] = -2146318022;
assign addr[28757] = -2146862854;
assign addr[28758] = -2147237452;
assign addr[28759] = -2147441787;
assign addr[28760] = -2147475844;
assign addr[28761] = -2147339619;
assign addr[28762] = -2147033123;
assign addr[28763] = -2146556380;
assign addr[28764] = -2145909429;
assign addr[28765] = -2145092320;
assign addr[28766] = -2144105118;
assign addr[28767] = -2142947902;
assign addr[28768] = -2141620763;
assign addr[28769] = -2140123807;
assign addr[28770] = -2138457152;
assign addr[28771] = -2136620930;
assign addr[28772] = -2134615288;
assign addr[28773] = -2132440383;
assign addr[28774] = -2130096389;
assign addr[28775] = -2127583492;
assign addr[28776] = -2124901890;
assign addr[28777] = -2122051796;
assign addr[28778] = -2119033436;
assign addr[28779] = -2115847050;
assign addr[28780] = -2112492891;
assign addr[28781] = -2108971223;
assign addr[28782] = -2105282327;
assign addr[28783] = -2101426496;
assign addr[28784] = -2097404033;
assign addr[28785] = -2093215260;
assign addr[28786] = -2088860507;
assign addr[28787] = -2084340120;
assign addr[28788] = -2079654458;
assign addr[28789] = -2074803892;
assign addr[28790] = -2069788807;
assign addr[28791] = -2064609600;
assign addr[28792] = -2059266683;
assign addr[28793] = -2053760478;
assign addr[28794] = -2048091422;
assign addr[28795] = -2042259965;
assign addr[28796] = -2036266570;
assign addr[28797] = -2030111710;
assign addr[28798] = -2023795876;
assign addr[28799] = -2017319567;
assign addr[28800] = -2010683297;
assign addr[28801] = -2003887591;
assign addr[28802] = -1996932990;
assign addr[28803] = -1989820044;
assign addr[28804] = -1982549318;
assign addr[28805] = -1975121388;
assign addr[28806] = -1967536842;
assign addr[28807] = -1959796283;
assign addr[28808] = -1951900324;
assign addr[28809] = -1943849591;
assign addr[28810] = -1935644723;
assign addr[28811] = -1927286370;
assign addr[28812] = -1918775195;
assign addr[28813] = -1910111873;
assign addr[28814] = -1901297091;
assign addr[28815] = -1892331547;
assign addr[28816] = -1883215953;
assign addr[28817] = -1873951032;
assign addr[28818] = -1864537518;
assign addr[28819] = -1854976157;
assign addr[28820] = -1845267708;
assign addr[28821] = -1835412941;
assign addr[28822] = -1825412636;
assign addr[28823] = -1815267588;
assign addr[28824] = -1804978599;
assign addr[28825] = -1794546487;
assign addr[28826] = -1783972079;
assign addr[28827] = -1773256212;
assign addr[28828] = -1762399737;
assign addr[28829] = -1751403515;
assign addr[28830] = -1740268417;
assign addr[28831] = -1728995326;
assign addr[28832] = -1717585136;
assign addr[28833] = -1706038753;
assign addr[28834] = -1694357091;
assign addr[28835] = -1682541077;
assign addr[28836] = -1670591647;
assign addr[28837] = -1658509750;
assign addr[28838] = -1646296344;
assign addr[28839] = -1633952396;
assign addr[28840] = -1621478885;
assign addr[28841] = -1608876801;
assign addr[28842] = -1596147143;
assign addr[28843] = -1583290921;
assign addr[28844] = -1570309153;
assign addr[28845] = -1557202869;
assign addr[28846] = -1543973108;
assign addr[28847] = -1530620920;
assign addr[28848] = -1517147363;
assign addr[28849] = -1503553506;
assign addr[28850] = -1489840425;
assign addr[28851] = -1476009210;
assign addr[28852] = -1462060956;
assign addr[28853] = -1447996770;
assign addr[28854] = -1433817766;
assign addr[28855] = -1419525069;
assign addr[28856] = -1405119813;
assign addr[28857] = -1390603139;
assign addr[28858] = -1375976199;
assign addr[28859] = -1361240152;
assign addr[28860] = -1346396168;
assign addr[28861] = -1331445422;
assign addr[28862] = -1316389101;
assign addr[28863] = -1301228398;
assign addr[28864] = -1285964516;
assign addr[28865] = -1270598665;
assign addr[28866] = -1255132063;
assign addr[28867] = -1239565936;
assign addr[28868] = -1223901520;
assign addr[28869] = -1208140056;
assign addr[28870] = -1192282793;
assign addr[28871] = -1176330990;
assign addr[28872] = -1160285911;
assign addr[28873] = -1144148829;
assign addr[28874] = -1127921022;
assign addr[28875] = -1111603778;
assign addr[28876] = -1095198391;
assign addr[28877] = -1078706161;
assign addr[28878] = -1062128397;
assign addr[28879] = -1045466412;
assign addr[28880] = -1028721528;
assign addr[28881] = -1011895073;
assign addr[28882] = -994988380;
assign addr[28883] = -978002791;
assign addr[28884] = -960939653;
assign addr[28885] = -943800318;
assign addr[28886] = -926586145;
assign addr[28887] = -909298500;
assign addr[28888] = -891938752;
assign addr[28889] = -874508280;
assign addr[28890] = -857008464;
assign addr[28891] = -839440693;
assign addr[28892] = -821806359;
assign addr[28893] = -804106861;
assign addr[28894] = -786343603;
assign addr[28895] = -768517992;
assign addr[28896] = -750631442;
assign addr[28897] = -732685372;
assign addr[28898] = -714681204;
assign addr[28899] = -696620367;
assign addr[28900] = -678504291;
assign addr[28901] = -660334415;
assign addr[28902] = -642112178;
assign addr[28903] = -623839025;
assign addr[28904] = -605516406;
assign addr[28905] = -587145773;
assign addr[28906] = -568728583;
assign addr[28907] = -550266296;
assign addr[28908] = -531760377;
assign addr[28909] = -513212292;
assign addr[28910] = -494623513;
assign addr[28911] = -475995513;
assign addr[28912] = -457329769;
assign addr[28913] = -438627762;
assign addr[28914] = -419890975;
assign addr[28915] = -401120892;
assign addr[28916] = -382319004;
assign addr[28917] = -363486799;
assign addr[28918] = -344625773;
assign addr[28919] = -325737419;
assign addr[28920] = -306823237;
assign addr[28921] = -287884725;
assign addr[28922] = -268923386;
assign addr[28923] = -249940723;
assign addr[28924] = -230938242;
assign addr[28925] = -211917448;
assign addr[28926] = -192879850;
assign addr[28927] = -173826959;
assign addr[28928] = -154760284;
assign addr[28929] = -135681337;
assign addr[28930] = -116591632;
assign addr[28931] = -97492681;
assign addr[28932] = -78386000;
assign addr[28933] = -59273104;
assign addr[28934] = -40155507;
assign addr[28935] = -21034727;
assign addr[28936] = -1912278;
assign addr[28937] = 17210322;
assign addr[28938] = 36331557;
assign addr[28939] = 55449912;
assign addr[28940] = 74563870;
assign addr[28941] = 93671915;
assign addr[28942] = 112772533;
assign addr[28943] = 131864208;
assign addr[28944] = 150945428;
assign addr[28945] = 170014678;
assign addr[28946] = 189070447;
assign addr[28947] = 208111224;
assign addr[28948] = 227135500;
assign addr[28949] = 246141764;
assign addr[28950] = 265128512;
assign addr[28951] = 284094236;
assign addr[28952] = 303037433;
assign addr[28953] = 321956601;
assign addr[28954] = 340850240;
assign addr[28955] = 359716852;
assign addr[28956] = 378554940;
assign addr[28957] = 397363011;
assign addr[28958] = 416139574;
assign addr[28959] = 434883140;
assign addr[28960] = 453592221;
assign addr[28961] = 472265336;
assign addr[28962] = 490901003;
assign addr[28963] = 509497745;
assign addr[28964] = 528054086;
assign addr[28965] = 546568556;
assign addr[28966] = 565039687;
assign addr[28967] = 583466013;
assign addr[28968] = 601846074;
assign addr[28969] = 620178412;
assign addr[28970] = 638461574;
assign addr[28971] = 656694110;
assign addr[28972] = 674874574;
assign addr[28973] = 693001525;
assign addr[28974] = 711073524;
assign addr[28975] = 729089140;
assign addr[28976] = 747046944;
assign addr[28977] = 764945512;
assign addr[28978] = 782783424;
assign addr[28979] = 800559266;
assign addr[28980] = 818271628;
assign addr[28981] = 835919107;
assign addr[28982] = 853500302;
assign addr[28983] = 871013820;
assign addr[28984] = 888458272;
assign addr[28985] = 905832274;
assign addr[28986] = 923134450;
assign addr[28987] = 940363427;
assign addr[28988] = 957517838;
assign addr[28989] = 974596324;
assign addr[28990] = 991597531;
assign addr[28991] = 1008520110;
assign addr[28992] = 1025362720;
assign addr[28993] = 1042124025;
assign addr[28994] = 1058802695;
assign addr[28995] = 1075397409;
assign addr[28996] = 1091906851;
assign addr[28997] = 1108329711;
assign addr[28998] = 1124664687;
assign addr[28999] = 1140910484;
assign addr[29000] = 1157065814;
assign addr[29001] = 1173129396;
assign addr[29002] = 1189099956;
assign addr[29003] = 1204976227;
assign addr[29004] = 1220756951;
assign addr[29005] = 1236440877;
assign addr[29006] = 1252026760;
assign addr[29007] = 1267513365;
assign addr[29008] = 1282899464;
assign addr[29009] = 1298183838;
assign addr[29010] = 1313365273;
assign addr[29011] = 1328442566;
assign addr[29012] = 1343414522;
assign addr[29013] = 1358279953;
assign addr[29014] = 1373037681;
assign addr[29015] = 1387686535;
assign addr[29016] = 1402225355;
assign addr[29017] = 1416652986;
assign addr[29018] = 1430968286;
assign addr[29019] = 1445170118;
assign addr[29020] = 1459257358;
assign addr[29021] = 1473228887;
assign addr[29022] = 1487083598;
assign addr[29023] = 1500820393;
assign addr[29024] = 1514438181;
assign addr[29025] = 1527935884;
assign addr[29026] = 1541312431;
assign addr[29027] = 1554566762;
assign addr[29028] = 1567697824;
assign addr[29029] = 1580704578;
assign addr[29030] = 1593585992;
assign addr[29031] = 1606341043;
assign addr[29032] = 1618968722;
assign addr[29033] = 1631468027;
assign addr[29034] = 1643837966;
assign addr[29035] = 1656077559;
assign addr[29036] = 1668185835;
assign addr[29037] = 1680161834;
assign addr[29038] = 1692004606;
assign addr[29039] = 1703713213;
assign addr[29040] = 1715286726;
assign addr[29041] = 1726724227;
assign addr[29042] = 1738024810;
assign addr[29043] = 1749187577;
assign addr[29044] = 1760211645;
assign addr[29045] = 1771096139;
assign addr[29046] = 1781840195;
assign addr[29047] = 1792442963;
assign addr[29048] = 1802903601;
assign addr[29049] = 1813221279;
assign addr[29050] = 1823395180;
assign addr[29051] = 1833424497;
assign addr[29052] = 1843308435;
assign addr[29053] = 1853046210;
assign addr[29054] = 1862637049;
assign addr[29055] = 1872080193;
assign addr[29056] = 1881374892;
assign addr[29057] = 1890520410;
assign addr[29058] = 1899516021;
assign addr[29059] = 1908361011;
assign addr[29060] = 1917054681;
assign addr[29061] = 1925596340;
assign addr[29062] = 1933985310;
assign addr[29063] = 1942220928;
assign addr[29064] = 1950302539;
assign addr[29065] = 1958229503;
assign addr[29066] = 1966001192;
assign addr[29067] = 1973616989;
assign addr[29068] = 1981076290;
assign addr[29069] = 1988378503;
assign addr[29070] = 1995523051;
assign addr[29071] = 2002509365;
assign addr[29072] = 2009336893;
assign addr[29073] = 2016005093;
assign addr[29074] = 2022513436;
assign addr[29075] = 2028861406;
assign addr[29076] = 2035048499;
assign addr[29077] = 2041074226;
assign addr[29078] = 2046938108;
assign addr[29079] = 2052639680;
assign addr[29080] = 2058178491;
assign addr[29081] = 2063554100;
assign addr[29082] = 2068766083;
assign addr[29083] = 2073814024;
assign addr[29084] = 2078697525;
assign addr[29085] = 2083416198;
assign addr[29086] = 2087969669;
assign addr[29087] = 2092357577;
assign addr[29088] = 2096579573;
assign addr[29089] = 2100635323;
assign addr[29090] = 2104524506;
assign addr[29091] = 2108246813;
assign addr[29092] = 2111801949;
assign addr[29093] = 2115189632;
assign addr[29094] = 2118409593;
assign addr[29095] = 2121461578;
assign addr[29096] = 2124345343;
assign addr[29097] = 2127060661;
assign addr[29098] = 2129607316;
assign addr[29099] = 2131985106;
assign addr[29100] = 2134193842;
assign addr[29101] = 2136233350;
assign addr[29102] = 2138103468;
assign addr[29103] = 2139804048;
assign addr[29104] = 2141334954;
assign addr[29105] = 2142696065;
assign addr[29106] = 2143887273;
assign addr[29107] = 2144908484;
assign addr[29108] = 2145759618;
assign addr[29109] = 2146440605;
assign addr[29110] = 2146951393;
assign addr[29111] = 2147291941;
assign addr[29112] = 2147462221;
assign addr[29113] = 2147462221;
assign addr[29114] = 2147291941;
assign addr[29115] = 2146951393;
assign addr[29116] = 2146440605;
assign addr[29117] = 2145759618;
assign addr[29118] = 2144908484;
assign addr[29119] = 2143887273;
assign addr[29120] = 2142696065;
assign addr[29121] = 2141334954;
assign addr[29122] = 2139804048;
assign addr[29123] = 2138103468;
assign addr[29124] = 2136233350;
assign addr[29125] = 2134193842;
assign addr[29126] = 2131985106;
assign addr[29127] = 2129607316;
assign addr[29128] = 2127060661;
assign addr[29129] = 2124345343;
assign addr[29130] = 2121461578;
assign addr[29131] = 2118409593;
assign addr[29132] = 2115189632;
assign addr[29133] = 2111801949;
assign addr[29134] = 2108246813;
assign addr[29135] = 2104524506;
assign addr[29136] = 2100635323;
assign addr[29137] = 2096579573;
assign addr[29138] = 2092357577;
assign addr[29139] = 2087969669;
assign addr[29140] = 2083416198;
assign addr[29141] = 2078697525;
assign addr[29142] = 2073814024;
assign addr[29143] = 2068766083;
assign addr[29144] = 2063554100;
assign addr[29145] = 2058178491;
assign addr[29146] = 2052639680;
assign addr[29147] = 2046938108;
assign addr[29148] = 2041074226;
assign addr[29149] = 2035048499;
assign addr[29150] = 2028861406;
assign addr[29151] = 2022513436;
assign addr[29152] = 2016005093;
assign addr[29153] = 2009336893;
assign addr[29154] = 2002509365;
assign addr[29155] = 1995523051;
assign addr[29156] = 1988378503;
assign addr[29157] = 1981076290;
assign addr[29158] = 1973616989;
assign addr[29159] = 1966001192;
assign addr[29160] = 1958229503;
assign addr[29161] = 1950302539;
assign addr[29162] = 1942220928;
assign addr[29163] = 1933985310;
assign addr[29164] = 1925596340;
assign addr[29165] = 1917054681;
assign addr[29166] = 1908361011;
assign addr[29167] = 1899516021;
assign addr[29168] = 1890520410;
assign addr[29169] = 1881374892;
assign addr[29170] = 1872080193;
assign addr[29171] = 1862637049;
assign addr[29172] = 1853046210;
assign addr[29173] = 1843308435;
assign addr[29174] = 1833424497;
assign addr[29175] = 1823395180;
assign addr[29176] = 1813221279;
assign addr[29177] = 1802903601;
assign addr[29178] = 1792442963;
assign addr[29179] = 1781840195;
assign addr[29180] = 1771096139;
assign addr[29181] = 1760211645;
assign addr[29182] = 1749187577;
assign addr[29183] = 1738024810;
assign addr[29184] = 1726724227;
assign addr[29185] = 1715286726;
assign addr[29186] = 1703713213;
assign addr[29187] = 1692004606;
assign addr[29188] = 1680161834;
assign addr[29189] = 1668185835;
assign addr[29190] = 1656077559;
assign addr[29191] = 1643837966;
assign addr[29192] = 1631468027;
assign addr[29193] = 1618968722;
assign addr[29194] = 1606341043;
assign addr[29195] = 1593585992;
assign addr[29196] = 1580704578;
assign addr[29197] = 1567697824;
assign addr[29198] = 1554566762;
assign addr[29199] = 1541312431;
assign addr[29200] = 1527935884;
assign addr[29201] = 1514438181;
assign addr[29202] = 1500820393;
assign addr[29203] = 1487083598;
assign addr[29204] = 1473228887;
assign addr[29205] = 1459257358;
assign addr[29206] = 1445170118;
assign addr[29207] = 1430968286;
assign addr[29208] = 1416652986;
assign addr[29209] = 1402225355;
assign addr[29210] = 1387686535;
assign addr[29211] = 1373037681;
assign addr[29212] = 1358279953;
assign addr[29213] = 1343414522;
assign addr[29214] = 1328442566;
assign addr[29215] = 1313365273;
assign addr[29216] = 1298183838;
assign addr[29217] = 1282899464;
assign addr[29218] = 1267513365;
assign addr[29219] = 1252026760;
assign addr[29220] = 1236440877;
assign addr[29221] = 1220756951;
assign addr[29222] = 1204976227;
assign addr[29223] = 1189099956;
assign addr[29224] = 1173129396;
assign addr[29225] = 1157065814;
assign addr[29226] = 1140910484;
assign addr[29227] = 1124664687;
assign addr[29228] = 1108329711;
assign addr[29229] = 1091906851;
assign addr[29230] = 1075397409;
assign addr[29231] = 1058802695;
assign addr[29232] = 1042124025;
assign addr[29233] = 1025362720;
assign addr[29234] = 1008520110;
assign addr[29235] = 991597531;
assign addr[29236] = 974596324;
assign addr[29237] = 957517838;
assign addr[29238] = 940363427;
assign addr[29239] = 923134450;
assign addr[29240] = 905832274;
assign addr[29241] = 888458272;
assign addr[29242] = 871013820;
assign addr[29243] = 853500302;
assign addr[29244] = 835919107;
assign addr[29245] = 818271628;
assign addr[29246] = 800559266;
assign addr[29247] = 782783424;
assign addr[29248] = 764945512;
assign addr[29249] = 747046944;
assign addr[29250] = 729089140;
assign addr[29251] = 711073524;
assign addr[29252] = 693001525;
assign addr[29253] = 674874574;
assign addr[29254] = 656694110;
assign addr[29255] = 638461574;
assign addr[29256] = 620178412;
assign addr[29257] = 601846074;
assign addr[29258] = 583466013;
assign addr[29259] = 565039687;
assign addr[29260] = 546568556;
assign addr[29261] = 528054086;
assign addr[29262] = 509497745;
assign addr[29263] = 490901003;
assign addr[29264] = 472265336;
assign addr[29265] = 453592221;
assign addr[29266] = 434883140;
assign addr[29267] = 416139574;
assign addr[29268] = 397363011;
assign addr[29269] = 378554940;
assign addr[29270] = 359716852;
assign addr[29271] = 340850240;
assign addr[29272] = 321956601;
assign addr[29273] = 303037433;
assign addr[29274] = 284094236;
assign addr[29275] = 265128512;
assign addr[29276] = 246141764;
assign addr[29277] = 227135500;
assign addr[29278] = 208111224;
assign addr[29279] = 189070447;
assign addr[29280] = 170014678;
assign addr[29281] = 150945428;
assign addr[29282] = 131864208;
assign addr[29283] = 112772533;
assign addr[29284] = 93671915;
assign addr[29285] = 74563870;
assign addr[29286] = 55449912;
assign addr[29287] = 36331557;
assign addr[29288] = 17210322;
assign addr[29289] = -1912278;
assign addr[29290] = -21034727;
assign addr[29291] = -40155507;
assign addr[29292] = -59273104;
assign addr[29293] = -78386000;
assign addr[29294] = -97492681;
assign addr[29295] = -116591632;
assign addr[29296] = -135681337;
assign addr[29297] = -154760284;
assign addr[29298] = -173826959;
assign addr[29299] = -192879850;
assign addr[29300] = -211917448;
assign addr[29301] = -230938242;
assign addr[29302] = -249940723;
assign addr[29303] = -268923386;
assign addr[29304] = -287884725;
assign addr[29305] = -306823237;
assign addr[29306] = -325737419;
assign addr[29307] = -344625773;
assign addr[29308] = -363486799;
assign addr[29309] = -382319004;
assign addr[29310] = -401120892;
assign addr[29311] = -419890975;
assign addr[29312] = -438627762;
assign addr[29313] = -457329769;
assign addr[29314] = -475995513;
assign addr[29315] = -494623513;
assign addr[29316] = -513212292;
assign addr[29317] = -531760377;
assign addr[29318] = -550266296;
assign addr[29319] = -568728583;
assign addr[29320] = -587145773;
assign addr[29321] = -605516406;
assign addr[29322] = -623839025;
assign addr[29323] = -642112178;
assign addr[29324] = -660334415;
assign addr[29325] = -678504291;
assign addr[29326] = -696620367;
assign addr[29327] = -714681204;
assign addr[29328] = -732685372;
assign addr[29329] = -750631442;
assign addr[29330] = -768517992;
assign addr[29331] = -786343603;
assign addr[29332] = -804106861;
assign addr[29333] = -821806359;
assign addr[29334] = -839440693;
assign addr[29335] = -857008464;
assign addr[29336] = -874508280;
assign addr[29337] = -891938752;
assign addr[29338] = -909298500;
assign addr[29339] = -926586145;
assign addr[29340] = -943800318;
assign addr[29341] = -960939653;
assign addr[29342] = -978002791;
assign addr[29343] = -994988380;
assign addr[29344] = -1011895073;
assign addr[29345] = -1028721528;
assign addr[29346] = -1045466412;
assign addr[29347] = -1062128397;
assign addr[29348] = -1078706161;
assign addr[29349] = -1095198391;
assign addr[29350] = -1111603778;
assign addr[29351] = -1127921022;
assign addr[29352] = -1144148829;
assign addr[29353] = -1160285911;
assign addr[29354] = -1176330990;
assign addr[29355] = -1192282793;
assign addr[29356] = -1208140056;
assign addr[29357] = -1223901520;
assign addr[29358] = -1239565936;
assign addr[29359] = -1255132063;
assign addr[29360] = -1270598665;
assign addr[29361] = -1285964516;
assign addr[29362] = -1301228398;
assign addr[29363] = -1316389101;
assign addr[29364] = -1331445422;
assign addr[29365] = -1346396168;
assign addr[29366] = -1361240152;
assign addr[29367] = -1375976199;
assign addr[29368] = -1390603139;
assign addr[29369] = -1405119813;
assign addr[29370] = -1419525069;
assign addr[29371] = -1433817766;
assign addr[29372] = -1447996770;
assign addr[29373] = -1462060956;
assign addr[29374] = -1476009210;
assign addr[29375] = -1489840425;
assign addr[29376] = -1503553506;
assign addr[29377] = -1517147363;
assign addr[29378] = -1530620920;
assign addr[29379] = -1543973108;
assign addr[29380] = -1557202869;
assign addr[29381] = -1570309153;
assign addr[29382] = -1583290921;
assign addr[29383] = -1596147143;
assign addr[29384] = -1608876801;
assign addr[29385] = -1621478885;
assign addr[29386] = -1633952396;
assign addr[29387] = -1646296344;
assign addr[29388] = -1658509750;
assign addr[29389] = -1670591647;
assign addr[29390] = -1682541077;
assign addr[29391] = -1694357091;
assign addr[29392] = -1706038753;
assign addr[29393] = -1717585136;
assign addr[29394] = -1728995326;
assign addr[29395] = -1740268417;
assign addr[29396] = -1751403515;
assign addr[29397] = -1762399737;
assign addr[29398] = -1773256212;
assign addr[29399] = -1783972079;
assign addr[29400] = -1794546487;
assign addr[29401] = -1804978599;
assign addr[29402] = -1815267588;
assign addr[29403] = -1825412636;
assign addr[29404] = -1835412941;
assign addr[29405] = -1845267708;
assign addr[29406] = -1854976157;
assign addr[29407] = -1864537518;
assign addr[29408] = -1873951032;
assign addr[29409] = -1883215953;
assign addr[29410] = -1892331547;
assign addr[29411] = -1901297091;
assign addr[29412] = -1910111873;
assign addr[29413] = -1918775195;
assign addr[29414] = -1927286370;
assign addr[29415] = -1935644723;
assign addr[29416] = -1943849591;
assign addr[29417] = -1951900324;
assign addr[29418] = -1959796283;
assign addr[29419] = -1967536842;
assign addr[29420] = -1975121388;
assign addr[29421] = -1982549318;
assign addr[29422] = -1989820044;
assign addr[29423] = -1996932990;
assign addr[29424] = -2003887591;
assign addr[29425] = -2010683297;
assign addr[29426] = -2017319567;
assign addr[29427] = -2023795876;
assign addr[29428] = -2030111710;
assign addr[29429] = -2036266570;
assign addr[29430] = -2042259965;
assign addr[29431] = -2048091422;
assign addr[29432] = -2053760478;
assign addr[29433] = -2059266683;
assign addr[29434] = -2064609600;
assign addr[29435] = -2069788807;
assign addr[29436] = -2074803892;
assign addr[29437] = -2079654458;
assign addr[29438] = -2084340120;
assign addr[29439] = -2088860507;
assign addr[29440] = -2093215260;
assign addr[29441] = -2097404033;
assign addr[29442] = -2101426496;
assign addr[29443] = -2105282327;
assign addr[29444] = -2108971223;
assign addr[29445] = -2112492891;
assign addr[29446] = -2115847050;
assign addr[29447] = -2119033436;
assign addr[29448] = -2122051796;
assign addr[29449] = -2124901890;
assign addr[29450] = -2127583492;
assign addr[29451] = -2130096389;
assign addr[29452] = -2132440383;
assign addr[29453] = -2134615288;
assign addr[29454] = -2136620930;
assign addr[29455] = -2138457152;
assign addr[29456] = -2140123807;
assign addr[29457] = -2141620763;
assign addr[29458] = -2142947902;
assign addr[29459] = -2144105118;
assign addr[29460] = -2145092320;
assign addr[29461] = -2145909429;
assign addr[29462] = -2146556380;
assign addr[29463] = -2147033123;
assign addr[29464] = -2147339619;
assign addr[29465] = -2147475844;
assign addr[29466] = -2147441787;
assign addr[29467] = -2147237452;
assign addr[29468] = -2146862854;
assign addr[29469] = -2146318022;
assign addr[29470] = -2145603001;
assign addr[29471] = -2144717846;
assign addr[29472] = -2143662628;
assign addr[29473] = -2142437431;
assign addr[29474] = -2141042352;
assign addr[29475] = -2139477502;
assign addr[29476] = -2137743003;
assign addr[29477] = -2135838995;
assign addr[29478] = -2133765628;
assign addr[29479] = -2131523066;
assign addr[29480] = -2129111488;
assign addr[29481] = -2126531084;
assign addr[29482] = -2123782059;
assign addr[29483] = -2120864631;
assign addr[29484] = -2117779031;
assign addr[29485] = -2114525505;
assign addr[29486] = -2111104309;
assign addr[29487] = -2107515716;
assign addr[29488] = -2103760010;
assign addr[29489] = -2099837489;
assign addr[29490] = -2095748463;
assign addr[29491] = -2091493257;
assign addr[29492] = -2087072209;
assign addr[29493] = -2082485668;
assign addr[29494] = -2077733999;
assign addr[29495] = -2072817579;
assign addr[29496] = -2067736796;
assign addr[29497] = -2062492055;
assign addr[29498] = -2057083771;
assign addr[29499] = -2051512372;
assign addr[29500] = -2045778302;
assign addr[29501] = -2039882013;
assign addr[29502] = -2033823974;
assign addr[29503] = -2027604666;
assign addr[29504] = -2021224581;
assign addr[29505] = -2014684225;
assign addr[29506] = -2007984117;
assign addr[29507] = -2001124788;
assign addr[29508] = -1994106782;
assign addr[29509] = -1986930656;
assign addr[29510] = -1979596978;
assign addr[29511] = -1972106330;
assign addr[29512] = -1964459306;
assign addr[29513] = -1956656513;
assign addr[29514] = -1948698568;
assign addr[29515] = -1940586104;
assign addr[29516] = -1932319763;
assign addr[29517] = -1923900201;
assign addr[29518] = -1915328086;
assign addr[29519] = -1906604097;
assign addr[29520] = -1897728925;
assign addr[29521] = -1888703276;
assign addr[29522] = -1879527863;
assign addr[29523] = -1870203416;
assign addr[29524] = -1860730673;
assign addr[29525] = -1851110385;
assign addr[29526] = -1841343316;
assign addr[29527] = -1831430239;
assign addr[29528] = -1821371941;
assign addr[29529] = -1811169220;
assign addr[29530] = -1800822883;
assign addr[29531] = -1790333753;
assign addr[29532] = -1779702660;
assign addr[29533] = -1768930447;
assign addr[29534] = -1758017969;
assign addr[29535] = -1746966091;
assign addr[29536] = -1735775690;
assign addr[29537] = -1724447652;
assign addr[29538] = -1712982875;
assign addr[29539] = -1701382270;
assign addr[29540] = -1689646755;
assign addr[29541] = -1677777262;
assign addr[29542] = -1665774731;
assign addr[29543] = -1653640115;
assign addr[29544] = -1641374375;
assign addr[29545] = -1628978484;
assign addr[29546] = -1616453425;
assign addr[29547] = -1603800191;
assign addr[29548] = -1591019785;
assign addr[29549] = -1578113222;
assign addr[29550] = -1565081523;
assign addr[29551] = -1551925723;
assign addr[29552] = -1538646865;
assign addr[29553] = -1525246002;
assign addr[29554] = -1511724196;
assign addr[29555] = -1498082520;
assign addr[29556] = -1484322054;
assign addr[29557] = -1470443891;
assign addr[29558] = -1456449131;
assign addr[29559] = -1442338884;
assign addr[29560] = -1428114267;
assign addr[29561] = -1413776410;
assign addr[29562] = -1399326449;
assign addr[29563] = -1384765530;
assign addr[29564] = -1370094808;
assign addr[29565] = -1355315445;
assign addr[29566] = -1340428615;
assign addr[29567] = -1325435496;
assign addr[29568] = -1310337279;
assign addr[29569] = -1295135159;
assign addr[29570] = -1279830344;
assign addr[29571] = -1264424045;
assign addr[29572] = -1248917486;
assign addr[29573] = -1233311895;
assign addr[29574] = -1217608510;
assign addr[29575] = -1201808576;
assign addr[29576] = -1185913346;
assign addr[29577] = -1169924081;
assign addr[29578] = -1153842047;
assign addr[29579] = -1137668521;
assign addr[29580] = -1121404785;
assign addr[29581] = -1105052128;
assign addr[29582] = -1088611847;
assign addr[29583] = -1072085246;
assign addr[29584] = -1055473635;
assign addr[29585] = -1038778332;
assign addr[29586] = -1022000660;
assign addr[29587] = -1005141949;
assign addr[29588] = -988203537;
assign addr[29589] = -971186766;
assign addr[29590] = -954092986;
assign addr[29591] = -936923553;
assign addr[29592] = -919679827;
assign addr[29593] = -902363176;
assign addr[29594] = -884974973;
assign addr[29595] = -867516597;
assign addr[29596] = -849989433;
assign addr[29597] = -832394869;
assign addr[29598] = -814734301;
assign addr[29599] = -797009130;
assign addr[29600] = -779220762;
assign addr[29601] = -761370605;
assign addr[29602] = -743460077;
assign addr[29603] = -725490597;
assign addr[29604] = -707463589;
assign addr[29605] = -689380485;
assign addr[29606] = -671242716;
assign addr[29607] = -653051723;
assign addr[29608] = -634808946;
assign addr[29609] = -616515832;
assign addr[29610] = -598173833;
assign addr[29611] = -579784402;
assign addr[29612] = -561348998;
assign addr[29613] = -542869083;
assign addr[29614] = -524346121;
assign addr[29615] = -505781581;
assign addr[29616] = -487176937;
assign addr[29617] = -468533662;
assign addr[29618] = -449853235;
assign addr[29619] = -431137138;
assign addr[29620] = -412386854;
assign addr[29621] = -393603870;
assign addr[29622] = -374789676;
assign addr[29623] = -355945764;
assign addr[29624] = -337073627;
assign addr[29625] = -318174762;
assign addr[29626] = -299250668;
assign addr[29627] = -280302845;
assign addr[29628] = -261332796;
assign addr[29629] = -242342025;
assign addr[29630] = -223332037;
assign addr[29631] = -204304341;
assign addr[29632] = -185260444;
assign addr[29633] = -166201858;
assign addr[29634] = -147130093;
assign addr[29635] = -128046661;
assign addr[29636] = -108953076;
assign addr[29637] = -89850852;
assign addr[29638] = -70741503;
assign addr[29639] = -51626544;
assign addr[29640] = -32507492;
assign addr[29641] = -13385863;
assign addr[29642] = 5736829;
assign addr[29643] = 24859065;
assign addr[29644] = 43979330;
assign addr[29645] = 63096108;
assign addr[29646] = 82207882;
assign addr[29647] = 101313138;
assign addr[29648] = 120410361;
assign addr[29649] = 139498035;
assign addr[29650] = 158574649;
assign addr[29651] = 177638688;
assign addr[29652] = 196688642;
assign addr[29653] = 215722999;
assign addr[29654] = 234740251;
assign addr[29655] = 253738890;
assign addr[29656] = 272717408;
assign addr[29657] = 291674302;
assign addr[29658] = 310608068;
assign addr[29659] = 329517204;
assign addr[29660] = 348400212;
assign addr[29661] = 367255594;
assign addr[29662] = 386081854;
assign addr[29663] = 404877501;
assign addr[29664] = 423641043;
assign addr[29665] = 442370993;
assign addr[29666] = 461065866;
assign addr[29667] = 479724180;
assign addr[29668] = 498344454;
assign addr[29669] = 516925212;
assign addr[29670] = 535464981;
assign addr[29671] = 553962291;
assign addr[29672] = 572415676;
assign addr[29673] = 590823671;
assign addr[29674] = 609184818;
assign addr[29675] = 627497660;
assign addr[29676] = 645760745;
assign addr[29677] = 663972625;
assign addr[29678] = 682131857;
assign addr[29679] = 700236999;
assign addr[29680] = 718286617;
assign addr[29681] = 736279279;
assign addr[29682] = 754213559;
assign addr[29683] = 772088034;
assign addr[29684] = 789901288;
assign addr[29685] = 807651907;
assign addr[29686] = 825338484;
assign addr[29687] = 842959617;
assign addr[29688] = 860513908;
assign addr[29689] = 877999966;
assign addr[29690] = 895416404;
assign addr[29691] = 912761841;
assign addr[29692] = 930034901;
assign addr[29693] = 947234215;
assign addr[29694] = 964358420;
assign addr[29695] = 981406156;
assign addr[29696] = 998376073;
assign addr[29697] = 1015266825;
assign addr[29698] = 1032077073;
assign addr[29699] = 1048805483;
assign addr[29700] = 1065450729;
assign addr[29701] = 1082011492;
assign addr[29702] = 1098486458;
assign addr[29703] = 1114874320;
assign addr[29704] = 1131173780;
assign addr[29705] = 1147383544;
assign addr[29706] = 1163502328;
assign addr[29707] = 1179528853;
assign addr[29708] = 1195461849;
assign addr[29709] = 1211300053;
assign addr[29710] = 1227042207;
assign addr[29711] = 1242687064;
assign addr[29712] = 1258233384;
assign addr[29713] = 1273679934;
assign addr[29714] = 1289025489;
assign addr[29715] = 1304268832;
assign addr[29716] = 1319408754;
assign addr[29717] = 1334444055;
assign addr[29718] = 1349373543;
assign addr[29719] = 1364196034;
assign addr[29720] = 1378910353;
assign addr[29721] = 1393515332;
assign addr[29722] = 1408009814;
assign addr[29723] = 1422392650;
assign addr[29724] = 1436662698;
assign addr[29725] = 1450818828;
assign addr[29726] = 1464859917;
assign addr[29727] = 1478784851;
assign addr[29728] = 1492592527;
assign addr[29729] = 1506281850;
assign addr[29730] = 1519851733;
assign addr[29731] = 1533301101;
assign addr[29732] = 1546628888;
assign addr[29733] = 1559834037;
assign addr[29734] = 1572915501;
assign addr[29735] = 1585872242;
assign addr[29736] = 1598703233;
assign addr[29737] = 1611407456;
assign addr[29738] = 1623983905;
assign addr[29739] = 1636431582;
assign addr[29740] = 1648749499;
assign addr[29741] = 1660936681;
assign addr[29742] = 1672992161;
assign addr[29743] = 1684914983;
assign addr[29744] = 1696704201;
assign addr[29745] = 1708358881;
assign addr[29746] = 1719878099;
assign addr[29747] = 1731260941;
assign addr[29748] = 1742506504;
assign addr[29749] = 1753613897;
assign addr[29750] = 1764582240;
assign addr[29751] = 1775410662;
assign addr[29752] = 1786098304;
assign addr[29753] = 1796644320;
assign addr[29754] = 1807047873;
assign addr[29755] = 1817308138;
assign addr[29756] = 1827424302;
assign addr[29757] = 1837395562;
assign addr[29758] = 1847221128;
assign addr[29759] = 1856900221;
assign addr[29760] = 1866432072;
assign addr[29761] = 1875815927;
assign addr[29762] = 1885051042;
assign addr[29763] = 1894136683;
assign addr[29764] = 1903072131;
assign addr[29765] = 1911856677;
assign addr[29766] = 1920489624;
assign addr[29767] = 1928970288;
assign addr[29768] = 1937297997;
assign addr[29769] = 1945472089;
assign addr[29770] = 1953491918;
assign addr[29771] = 1961356847;
assign addr[29772] = 1969066252;
assign addr[29773] = 1976619522;
assign addr[29774] = 1984016058;
assign addr[29775] = 1991255274;
assign addr[29776] = 1998336596;
assign addr[29777] = 2005259462;
assign addr[29778] = 2012023322;
assign addr[29779] = 2018627642;
assign addr[29780] = 2025071897;
assign addr[29781] = 2031355576;
assign addr[29782] = 2037478181;
assign addr[29783] = 2043439226;
assign addr[29784] = 2049238240;
assign addr[29785] = 2054874761;
assign addr[29786] = 2060348343;
assign addr[29787] = 2065658552;
assign addr[29788] = 2070804967;
assign addr[29789] = 2075787180;
assign addr[29790] = 2080604795;
assign addr[29791] = 2085257431;
assign addr[29792] = 2089744719;
assign addr[29793] = 2094066304;
assign addr[29794] = 2098221841;
assign addr[29795] = 2102211002;
assign addr[29796] = 2106033471;
assign addr[29797] = 2109688944;
assign addr[29798] = 2113177132;
assign addr[29799] = 2116497758;
assign addr[29800] = 2119650558;
assign addr[29801] = 2122635283;
assign addr[29802] = 2125451696;
assign addr[29803] = 2128099574;
assign addr[29804] = 2130578706;
assign addr[29805] = 2132888897;
assign addr[29806] = 2135029962;
assign addr[29807] = 2137001733;
assign addr[29808] = 2138804053;
assign addr[29809] = 2140436778;
assign addr[29810] = 2141899780;
assign addr[29811] = 2143192942;
assign addr[29812] = 2144316162;
assign addr[29813] = 2145269351;
assign addr[29814] = 2146052433;
assign addr[29815] = 2146665347;
assign addr[29816] = 2147108043;
assign addr[29817] = 2147380486;
assign addr[29818] = 2147482655;
assign addr[29819] = 2147414542;
assign addr[29820] = 2147176152;
assign addr[29821] = 2146767505;
assign addr[29822] = 2146188631;
assign addr[29823] = 2145439578;
assign addr[29824] = 2144520405;
assign addr[29825] = 2143431184;
assign addr[29826] = 2142172003;
assign addr[29827] = 2140742960;
assign addr[29828] = 2139144169;
assign addr[29829] = 2137375758;
assign addr[29830] = 2135437865;
assign addr[29831] = 2133330646;
assign addr[29832] = 2131054266;
assign addr[29833] = 2128608907;
assign addr[29834] = 2125994762;
assign addr[29835] = 2123212038;
assign addr[29836] = 2120260957;
assign addr[29837] = 2117141752;
assign addr[29838] = 2113854671;
assign addr[29839] = 2110399974;
assign addr[29840] = 2106777935;
assign addr[29841] = 2102988841;
assign addr[29842] = 2099032994;
assign addr[29843] = 2094910706;
assign addr[29844] = 2090622304;
assign addr[29845] = 2086168128;
assign addr[29846] = 2081548533;
assign addr[29847] = 2076763883;
assign addr[29848] = 2071814558;
assign addr[29849] = 2066700952;
assign addr[29850] = 2061423468;
assign addr[29851] = 2055982526;
assign addr[29852] = 2050378558;
assign addr[29853] = 2044612007;
assign addr[29854] = 2038683330;
assign addr[29855] = 2032592999;
assign addr[29856] = 2026341495;
assign addr[29857] = 2019929315;
assign addr[29858] = 2013356967;
assign addr[29859] = 2006624971;
assign addr[29860] = 1999733863;
assign addr[29861] = 1992684188;
assign addr[29862] = 1985476506;
assign addr[29863] = 1978111387;
assign addr[29864] = 1970589416;
assign addr[29865] = 1962911189;
assign addr[29866] = 1955077316;
assign addr[29867] = 1947088417;
assign addr[29868] = 1938945125;
assign addr[29869] = 1930648088;
assign addr[29870] = 1922197961;
assign addr[29871] = 1913595416;
assign addr[29872] = 1904841135;
assign addr[29873] = 1895935811;
assign addr[29874] = 1886880151;
assign addr[29875] = 1877674873;
assign addr[29876] = 1868320707;
assign addr[29877] = 1858818395;
assign addr[29878] = 1849168689;
assign addr[29879] = 1839372356;
assign addr[29880] = 1829430172;
assign addr[29881] = 1819342925;
assign addr[29882] = 1809111415;
assign addr[29883] = 1798736454;
assign addr[29884] = 1788218865;
assign addr[29885] = 1777559480;
assign addr[29886] = 1766759146;
assign addr[29887] = 1755818718;
assign addr[29888] = 1744739065;
assign addr[29889] = 1733521064;
assign addr[29890] = 1722165606;
assign addr[29891] = 1710673591;
assign addr[29892] = 1699045930;
assign addr[29893] = 1687283545;
assign addr[29894] = 1675387369;
assign addr[29895] = 1663358344;
assign addr[29896] = 1651197426;
assign addr[29897] = 1638905577;
assign addr[29898] = 1626483774;
assign addr[29899] = 1613933000;
assign addr[29900] = 1601254251;
assign addr[29901] = 1588448533;
assign addr[29902] = 1575516860;
assign addr[29903] = 1562460258;
assign addr[29904] = 1549279763;
assign addr[29905] = 1535976419;
assign addr[29906] = 1522551282;
assign addr[29907] = 1509005416;
assign addr[29908] = 1495339895;
assign addr[29909] = 1481555802;
assign addr[29910] = 1467654232;
assign addr[29911] = 1453636285;
assign addr[29912] = 1439503074;
assign addr[29913] = 1425255719;
assign addr[29914] = 1410895350;
assign addr[29915] = 1396423105;
assign addr[29916] = 1381840133;
assign addr[29917] = 1367147589;
assign addr[29918] = 1352346639;
assign addr[29919] = 1337438456;
assign addr[29920] = 1322424222;
assign addr[29921] = 1307305128;
assign addr[29922] = 1292082373;
assign addr[29923] = 1276757164;
assign addr[29924] = 1261330715;
assign addr[29925] = 1245804251;
assign addr[29926] = 1230179002;
assign addr[29927] = 1214456207;
assign addr[29928] = 1198637114;
assign addr[29929] = 1182722976;
assign addr[29930] = 1166715055;
assign addr[29931] = 1150614620;
assign addr[29932] = 1134422949;
assign addr[29933] = 1118141326;
assign addr[29934] = 1101771040;
assign addr[29935] = 1085313391;
assign addr[29936] = 1068769683;
assign addr[29937] = 1052141228;
assign addr[29938] = 1035429345;
assign addr[29939] = 1018635358;
assign addr[29940] = 1001760600;
assign addr[29941] = 984806408;
assign addr[29942] = 967774128;
assign addr[29943] = 950665109;
assign addr[29944] = 933480707;
assign addr[29945] = 916222287;
assign addr[29946] = 898891215;
assign addr[29947] = 881488868;
assign addr[29948] = 864016623;
assign addr[29949] = 846475867;
assign addr[29950] = 828867991;
assign addr[29951] = 811194391;
assign addr[29952] = 793456467;
assign addr[29953] = 775655628;
assign addr[29954] = 757793284;
assign addr[29955] = 739870851;
assign addr[29956] = 721889752;
assign addr[29957] = 703851410;
assign addr[29958] = 685757258;
assign addr[29959] = 667608730;
assign addr[29960] = 649407264;
assign addr[29961] = 631154304;
assign addr[29962] = 612851297;
assign addr[29963] = 594499695;
assign addr[29964] = 576100953;
assign addr[29965] = 557656529;
assign addr[29966] = 539167887;
assign addr[29967] = 520636492;
assign addr[29968] = 502063814;
assign addr[29969] = 483451325;
assign addr[29970] = 464800501;
assign addr[29971] = 446112822;
assign addr[29972] = 427389768;
assign addr[29973] = 408632825;
assign addr[29974] = 389843480;
assign addr[29975] = 371023223;
assign addr[29976] = 352173546;
assign addr[29977] = 333295944;
assign addr[29978] = 314391913;
assign addr[29979] = 295462954;
assign addr[29980] = 276510565;
assign addr[29981] = 257536251;
assign addr[29982] = 238541516;
assign addr[29983] = 219527866;
assign addr[29984] = 200496809;
assign addr[29985] = 181449854;
assign addr[29986] = 162388511;
assign addr[29987] = 143314291;
assign addr[29988] = 124228708;
assign addr[29989] = 105133274;
assign addr[29990] = 86029503;
assign addr[29991] = 66918911;
assign addr[29992] = 47803013;
assign addr[29993] = 28683324;
assign addr[29994] = 9561361;
assign addr[29995] = -9561361;
assign addr[29996] = -28683324;
assign addr[29997] = -47803013;
assign addr[29998] = -66918911;
assign addr[29999] = -86029503;
assign addr[30000] = -105133274;
assign addr[30001] = -124228708;
assign addr[30002] = -143314291;
assign addr[30003] = -162388511;
assign addr[30004] = -181449854;
assign addr[30005] = -200496809;
assign addr[30006] = -219527866;
assign addr[30007] = -238541516;
assign addr[30008] = -257536251;
assign addr[30009] = -276510565;
assign addr[30010] = -295462954;
assign addr[30011] = -314391913;
assign addr[30012] = -333295944;
assign addr[30013] = -352173546;
assign addr[30014] = -371023223;
assign addr[30015] = -389843480;
assign addr[30016] = -408632825;
assign addr[30017] = -427389768;
assign addr[30018] = -446112822;
assign addr[30019] = -464800501;
assign addr[30020] = -483451325;
assign addr[30021] = -502063814;
assign addr[30022] = -520636492;
assign addr[30023] = -539167887;
assign addr[30024] = -557656529;
assign addr[30025] = -576100953;
assign addr[30026] = -594499695;
assign addr[30027] = -612851297;
assign addr[30028] = -631154304;
assign addr[30029] = -649407264;
assign addr[30030] = -667608730;
assign addr[30031] = -685757258;
assign addr[30032] = -703851410;
assign addr[30033] = -721889752;
assign addr[30034] = -739870851;
assign addr[30035] = -757793284;
assign addr[30036] = -775655628;
assign addr[30037] = -793456467;
assign addr[30038] = -811194391;
assign addr[30039] = -828867991;
assign addr[30040] = -846475867;
assign addr[30041] = -864016623;
assign addr[30042] = -881488868;
assign addr[30043] = -898891215;
assign addr[30044] = -916222287;
assign addr[30045] = -933480707;
assign addr[30046] = -950665109;
assign addr[30047] = -967774128;
assign addr[30048] = -984806408;
assign addr[30049] = -1001760600;
assign addr[30050] = -1018635358;
assign addr[30051] = -1035429345;
assign addr[30052] = -1052141228;
assign addr[30053] = -1068769683;
assign addr[30054] = -1085313391;
assign addr[30055] = -1101771040;
assign addr[30056] = -1118141326;
assign addr[30057] = -1134422949;
assign addr[30058] = -1150614620;
assign addr[30059] = -1166715055;
assign addr[30060] = -1182722976;
assign addr[30061] = -1198637114;
assign addr[30062] = -1214456207;
assign addr[30063] = -1230179002;
assign addr[30064] = -1245804251;
assign addr[30065] = -1261330715;
assign addr[30066] = -1276757164;
assign addr[30067] = -1292082373;
assign addr[30068] = -1307305128;
assign addr[30069] = -1322424222;
assign addr[30070] = -1337438456;
assign addr[30071] = -1352346639;
assign addr[30072] = -1367147589;
assign addr[30073] = -1381840133;
assign addr[30074] = -1396423105;
assign addr[30075] = -1410895350;
assign addr[30076] = -1425255719;
assign addr[30077] = -1439503074;
assign addr[30078] = -1453636285;
assign addr[30079] = -1467654232;
assign addr[30080] = -1481555802;
assign addr[30081] = -1495339895;
assign addr[30082] = -1509005416;
assign addr[30083] = -1522551282;
assign addr[30084] = -1535976419;
assign addr[30085] = -1549279763;
assign addr[30086] = -1562460258;
assign addr[30087] = -1575516860;
assign addr[30088] = -1588448533;
assign addr[30089] = -1601254251;
assign addr[30090] = -1613933000;
assign addr[30091] = -1626483774;
assign addr[30092] = -1638905577;
assign addr[30093] = -1651197426;
assign addr[30094] = -1663358344;
assign addr[30095] = -1675387369;
assign addr[30096] = -1687283545;
assign addr[30097] = -1699045930;
assign addr[30098] = -1710673591;
assign addr[30099] = -1722165606;
assign addr[30100] = -1733521064;
assign addr[30101] = -1744739065;
assign addr[30102] = -1755818718;
assign addr[30103] = -1766759146;
assign addr[30104] = -1777559480;
assign addr[30105] = -1788218865;
assign addr[30106] = -1798736454;
assign addr[30107] = -1809111415;
assign addr[30108] = -1819342925;
assign addr[30109] = -1829430172;
assign addr[30110] = -1839372356;
assign addr[30111] = -1849168689;
assign addr[30112] = -1858818395;
assign addr[30113] = -1868320707;
assign addr[30114] = -1877674873;
assign addr[30115] = -1886880151;
assign addr[30116] = -1895935811;
assign addr[30117] = -1904841135;
assign addr[30118] = -1913595416;
assign addr[30119] = -1922197961;
assign addr[30120] = -1930648088;
assign addr[30121] = -1938945125;
assign addr[30122] = -1947088417;
assign addr[30123] = -1955077316;
assign addr[30124] = -1962911189;
assign addr[30125] = -1970589416;
assign addr[30126] = -1978111387;
assign addr[30127] = -1985476506;
assign addr[30128] = -1992684188;
assign addr[30129] = -1999733863;
assign addr[30130] = -2006624971;
assign addr[30131] = -2013356967;
assign addr[30132] = -2019929315;
assign addr[30133] = -2026341495;
assign addr[30134] = -2032592999;
assign addr[30135] = -2038683330;
assign addr[30136] = -2044612007;
assign addr[30137] = -2050378558;
assign addr[30138] = -2055982526;
assign addr[30139] = -2061423468;
assign addr[30140] = -2066700952;
assign addr[30141] = -2071814558;
assign addr[30142] = -2076763883;
assign addr[30143] = -2081548533;
assign addr[30144] = -2086168128;
assign addr[30145] = -2090622304;
assign addr[30146] = -2094910706;
assign addr[30147] = -2099032994;
assign addr[30148] = -2102988841;
assign addr[30149] = -2106777935;
assign addr[30150] = -2110399974;
assign addr[30151] = -2113854671;
assign addr[30152] = -2117141752;
assign addr[30153] = -2120260957;
assign addr[30154] = -2123212038;
assign addr[30155] = -2125994762;
assign addr[30156] = -2128608907;
assign addr[30157] = -2131054266;
assign addr[30158] = -2133330646;
assign addr[30159] = -2135437865;
assign addr[30160] = -2137375758;
assign addr[30161] = -2139144169;
assign addr[30162] = -2140742960;
assign addr[30163] = -2142172003;
assign addr[30164] = -2143431184;
assign addr[30165] = -2144520405;
assign addr[30166] = -2145439578;
assign addr[30167] = -2146188631;
assign addr[30168] = -2146767505;
assign addr[30169] = -2147176152;
assign addr[30170] = -2147414542;
assign addr[30171] = -2147482655;
assign addr[30172] = -2147380486;
assign addr[30173] = -2147108043;
assign addr[30174] = -2146665347;
assign addr[30175] = -2146052433;
assign addr[30176] = -2145269351;
assign addr[30177] = -2144316162;
assign addr[30178] = -2143192942;
assign addr[30179] = -2141899780;
assign addr[30180] = -2140436778;
assign addr[30181] = -2138804053;
assign addr[30182] = -2137001733;
assign addr[30183] = -2135029962;
assign addr[30184] = -2132888897;
assign addr[30185] = -2130578706;
assign addr[30186] = -2128099574;
assign addr[30187] = -2125451696;
assign addr[30188] = -2122635283;
assign addr[30189] = -2119650558;
assign addr[30190] = -2116497758;
assign addr[30191] = -2113177132;
assign addr[30192] = -2109688944;
assign addr[30193] = -2106033471;
assign addr[30194] = -2102211002;
assign addr[30195] = -2098221841;
assign addr[30196] = -2094066304;
assign addr[30197] = -2089744719;
assign addr[30198] = -2085257431;
assign addr[30199] = -2080604795;
assign addr[30200] = -2075787180;
assign addr[30201] = -2070804967;
assign addr[30202] = -2065658552;
assign addr[30203] = -2060348343;
assign addr[30204] = -2054874761;
assign addr[30205] = -2049238240;
assign addr[30206] = -2043439226;
assign addr[30207] = -2037478181;
assign addr[30208] = -2031355576;
assign addr[30209] = -2025071897;
assign addr[30210] = -2018627642;
assign addr[30211] = -2012023322;
assign addr[30212] = -2005259462;
assign addr[30213] = -1998336596;
assign addr[30214] = -1991255274;
assign addr[30215] = -1984016058;
assign addr[30216] = -1976619522;
assign addr[30217] = -1969066252;
assign addr[30218] = -1961356847;
assign addr[30219] = -1953491918;
assign addr[30220] = -1945472089;
assign addr[30221] = -1937297997;
assign addr[30222] = -1928970288;
assign addr[30223] = -1920489624;
assign addr[30224] = -1911856677;
assign addr[30225] = -1903072131;
assign addr[30226] = -1894136683;
assign addr[30227] = -1885051042;
assign addr[30228] = -1875815927;
assign addr[30229] = -1866432072;
assign addr[30230] = -1856900221;
assign addr[30231] = -1847221128;
assign addr[30232] = -1837395562;
assign addr[30233] = -1827424302;
assign addr[30234] = -1817308138;
assign addr[30235] = -1807047873;
assign addr[30236] = -1796644320;
assign addr[30237] = -1786098304;
assign addr[30238] = -1775410662;
assign addr[30239] = -1764582240;
assign addr[30240] = -1753613897;
assign addr[30241] = -1742506504;
assign addr[30242] = -1731260941;
assign addr[30243] = -1719878099;
assign addr[30244] = -1708358881;
assign addr[30245] = -1696704201;
assign addr[30246] = -1684914983;
assign addr[30247] = -1672992161;
assign addr[30248] = -1660936681;
assign addr[30249] = -1648749499;
assign addr[30250] = -1636431582;
assign addr[30251] = -1623983905;
assign addr[30252] = -1611407456;
assign addr[30253] = -1598703233;
assign addr[30254] = -1585872242;
assign addr[30255] = -1572915501;
assign addr[30256] = -1559834037;
assign addr[30257] = -1546628888;
assign addr[30258] = -1533301101;
assign addr[30259] = -1519851733;
assign addr[30260] = -1506281850;
assign addr[30261] = -1492592527;
assign addr[30262] = -1478784851;
assign addr[30263] = -1464859917;
assign addr[30264] = -1450818828;
assign addr[30265] = -1436662698;
assign addr[30266] = -1422392650;
assign addr[30267] = -1408009814;
assign addr[30268] = -1393515332;
assign addr[30269] = -1378910353;
assign addr[30270] = -1364196034;
assign addr[30271] = -1349373543;
assign addr[30272] = -1334444055;
assign addr[30273] = -1319408754;
assign addr[30274] = -1304268832;
assign addr[30275] = -1289025489;
assign addr[30276] = -1273679934;
assign addr[30277] = -1258233384;
assign addr[30278] = -1242687064;
assign addr[30279] = -1227042207;
assign addr[30280] = -1211300053;
assign addr[30281] = -1195461849;
assign addr[30282] = -1179528853;
assign addr[30283] = -1163502328;
assign addr[30284] = -1147383544;
assign addr[30285] = -1131173780;
assign addr[30286] = -1114874320;
assign addr[30287] = -1098486458;
assign addr[30288] = -1082011492;
assign addr[30289] = -1065450729;
assign addr[30290] = -1048805483;
assign addr[30291] = -1032077073;
assign addr[30292] = -1015266825;
assign addr[30293] = -998376073;
assign addr[30294] = -981406156;
assign addr[30295] = -964358420;
assign addr[30296] = -947234215;
assign addr[30297] = -930034901;
assign addr[30298] = -912761841;
assign addr[30299] = -895416404;
assign addr[30300] = -877999966;
assign addr[30301] = -860513908;
assign addr[30302] = -842959617;
assign addr[30303] = -825338484;
assign addr[30304] = -807651907;
assign addr[30305] = -789901288;
assign addr[30306] = -772088034;
assign addr[30307] = -754213559;
assign addr[30308] = -736279279;
assign addr[30309] = -718286617;
assign addr[30310] = -700236999;
assign addr[30311] = -682131857;
assign addr[30312] = -663972625;
assign addr[30313] = -645760745;
assign addr[30314] = -627497660;
assign addr[30315] = -609184818;
assign addr[30316] = -590823671;
assign addr[30317] = -572415676;
assign addr[30318] = -553962291;
assign addr[30319] = -535464981;
assign addr[30320] = -516925212;
assign addr[30321] = -498344454;
assign addr[30322] = -479724180;
assign addr[30323] = -461065866;
assign addr[30324] = -442370993;
assign addr[30325] = -423641043;
assign addr[30326] = -404877501;
assign addr[30327] = -386081854;
assign addr[30328] = -367255594;
assign addr[30329] = -348400212;
assign addr[30330] = -329517204;
assign addr[30331] = -310608068;
assign addr[30332] = -291674302;
assign addr[30333] = -272717408;
assign addr[30334] = -253738890;
assign addr[30335] = -234740251;
assign addr[30336] = -215722999;
assign addr[30337] = -196688642;
assign addr[30338] = -177638688;
assign addr[30339] = -158574649;
assign addr[30340] = -139498035;
assign addr[30341] = -120410361;
assign addr[30342] = -101313138;
assign addr[30343] = -82207882;
assign addr[30344] = -63096108;
assign addr[30345] = -43979330;
assign addr[30346] = -24859065;
assign addr[30347] = -5736829;
assign addr[30348] = 13385863;
assign addr[30349] = 32507492;
assign addr[30350] = 51626544;
assign addr[30351] = 70741503;
assign addr[30352] = 89850852;
assign addr[30353] = 108953076;
assign addr[30354] = 128046661;
assign addr[30355] = 147130093;
assign addr[30356] = 166201858;
assign addr[30357] = 185260444;
assign addr[30358] = 204304341;
assign addr[30359] = 223332037;
assign addr[30360] = 242342025;
assign addr[30361] = 261332796;
assign addr[30362] = 280302845;
assign addr[30363] = 299250668;
assign addr[30364] = 318174762;
assign addr[30365] = 337073627;
assign addr[30366] = 355945764;
assign addr[30367] = 374789676;
assign addr[30368] = 393603870;
assign addr[30369] = 412386854;
assign addr[30370] = 431137138;
assign addr[30371] = 449853235;
assign addr[30372] = 468533662;
assign addr[30373] = 487176937;
assign addr[30374] = 505781581;
assign addr[30375] = 524346121;
assign addr[30376] = 542869083;
assign addr[30377] = 561348998;
assign addr[30378] = 579784402;
assign addr[30379] = 598173833;
assign addr[30380] = 616515832;
assign addr[30381] = 634808946;
assign addr[30382] = 653051723;
assign addr[30383] = 671242716;
assign addr[30384] = 689380485;
assign addr[30385] = 707463589;
assign addr[30386] = 725490597;
assign addr[30387] = 743460077;
assign addr[30388] = 761370605;
assign addr[30389] = 779220762;
assign addr[30390] = 797009130;
assign addr[30391] = 814734301;
assign addr[30392] = 832394869;
assign addr[30393] = 849989433;
assign addr[30394] = 867516597;
assign addr[30395] = 884974973;
assign addr[30396] = 902363176;
assign addr[30397] = 919679827;
assign addr[30398] = 936923553;
assign addr[30399] = 954092986;
assign addr[30400] = 971186766;
assign addr[30401] = 988203537;
assign addr[30402] = 1005141949;
assign addr[30403] = 1022000660;
assign addr[30404] = 1038778332;
assign addr[30405] = 1055473635;
assign addr[30406] = 1072085246;
assign addr[30407] = 1088611847;
assign addr[30408] = 1105052128;
assign addr[30409] = 1121404785;
assign addr[30410] = 1137668521;
assign addr[30411] = 1153842047;
assign addr[30412] = 1169924081;
assign addr[30413] = 1185913346;
assign addr[30414] = 1201808576;
assign addr[30415] = 1217608510;
assign addr[30416] = 1233311895;
assign addr[30417] = 1248917486;
assign addr[30418] = 1264424045;
assign addr[30419] = 1279830344;
assign addr[30420] = 1295135159;
assign addr[30421] = 1310337279;
assign addr[30422] = 1325435496;
assign addr[30423] = 1340428615;
assign addr[30424] = 1355315445;
assign addr[30425] = 1370094808;
assign addr[30426] = 1384765530;
assign addr[30427] = 1399326449;
assign addr[30428] = 1413776410;
assign addr[30429] = 1428114267;
assign addr[30430] = 1442338884;
assign addr[30431] = 1456449131;
assign addr[30432] = 1470443891;
assign addr[30433] = 1484322054;
assign addr[30434] = 1498082520;
assign addr[30435] = 1511724196;
assign addr[30436] = 1525246002;
assign addr[30437] = 1538646865;
assign addr[30438] = 1551925723;
assign addr[30439] = 1565081523;
assign addr[30440] = 1578113222;
assign addr[30441] = 1591019785;
assign addr[30442] = 1603800191;
assign addr[30443] = 1616453425;
assign addr[30444] = 1628978484;
assign addr[30445] = 1641374375;
assign addr[30446] = 1653640115;
assign addr[30447] = 1665774731;
assign addr[30448] = 1677777262;
assign addr[30449] = 1689646755;
assign addr[30450] = 1701382270;
assign addr[30451] = 1712982875;
assign addr[30452] = 1724447652;
assign addr[30453] = 1735775690;
assign addr[30454] = 1746966091;
assign addr[30455] = 1758017969;
assign addr[30456] = 1768930447;
assign addr[30457] = 1779702660;
assign addr[30458] = 1790333753;
assign addr[30459] = 1800822883;
assign addr[30460] = 1811169220;
assign addr[30461] = 1821371941;
assign addr[30462] = 1831430239;
assign addr[30463] = 1841343316;
assign addr[30464] = 1851110385;
assign addr[30465] = 1860730673;
assign addr[30466] = 1870203416;
assign addr[30467] = 1879527863;
assign addr[30468] = 1888703276;
assign addr[30469] = 1897728925;
assign addr[30470] = 1906604097;
assign addr[30471] = 1915328086;
assign addr[30472] = 1923900201;
assign addr[30473] = 1932319763;
assign addr[30474] = 1940586104;
assign addr[30475] = 1948698568;
assign addr[30476] = 1956656513;
assign addr[30477] = 1964459306;
assign addr[30478] = 1972106330;
assign addr[30479] = 1979596978;
assign addr[30480] = 1986930656;
assign addr[30481] = 1994106782;
assign addr[30482] = 2001124788;
assign addr[30483] = 2007984117;
assign addr[30484] = 2014684225;
assign addr[30485] = 2021224581;
assign addr[30486] = 2027604666;
assign addr[30487] = 2033823974;
assign addr[30488] = 2039882013;
assign addr[30489] = 2045778302;
assign addr[30490] = 2051512372;
assign addr[30491] = 2057083771;
assign addr[30492] = 2062492055;
assign addr[30493] = 2067736796;
assign addr[30494] = 2072817579;
assign addr[30495] = 2077733999;
assign addr[30496] = 2082485668;
assign addr[30497] = 2087072209;
assign addr[30498] = 2091493257;
assign addr[30499] = 2095748463;
assign addr[30500] = 2099837489;
assign addr[30501] = 2103760010;
assign addr[30502] = 2107515716;
assign addr[30503] = 2111104309;
assign addr[30504] = 2114525505;
assign addr[30505] = 2117779031;
assign addr[30506] = 2120864631;
assign addr[30507] = 2123782059;
assign addr[30508] = 2126531084;
assign addr[30509] = 2129111488;
assign addr[30510] = 2131523066;
assign addr[30511] = 2133765628;
assign addr[30512] = 2135838995;
assign addr[30513] = 2137743003;
assign addr[30514] = 2139477502;
assign addr[30515] = 2141042352;
assign addr[30516] = 2142437431;
assign addr[30517] = 2143662628;
assign addr[30518] = 2144717846;
assign addr[30519] = 2145603001;
assign addr[30520] = 2146318022;
assign addr[30521] = 2146862854;
assign addr[30522] = 2147237452;
assign addr[30523] = 2147441787;
assign addr[30524] = 2147475844;
assign addr[30525] = 2147339619;
assign addr[30526] = 2147033123;
assign addr[30527] = 2146556380;
assign addr[30528] = 2145909429;
assign addr[30529] = 2145092320;
assign addr[30530] = 2144105118;
assign addr[30531] = 2142947902;
assign addr[30532] = 2141620763;
assign addr[30533] = 2140123807;
assign addr[30534] = 2138457152;
assign addr[30535] = 2136620930;
assign addr[30536] = 2134615288;
assign addr[30537] = 2132440383;
assign addr[30538] = 2130096389;
assign addr[30539] = 2127583492;
assign addr[30540] = 2124901890;
assign addr[30541] = 2122051796;
assign addr[30542] = 2119033436;
assign addr[30543] = 2115847050;
assign addr[30544] = 2112492891;
assign addr[30545] = 2108971223;
assign addr[30546] = 2105282327;
assign addr[30547] = 2101426496;
assign addr[30548] = 2097404033;
assign addr[30549] = 2093215260;
assign addr[30550] = 2088860507;
assign addr[30551] = 2084340120;
assign addr[30552] = 2079654458;
assign addr[30553] = 2074803892;
assign addr[30554] = 2069788807;
assign addr[30555] = 2064609600;
assign addr[30556] = 2059266683;
assign addr[30557] = 2053760478;
assign addr[30558] = 2048091422;
assign addr[30559] = 2042259965;
assign addr[30560] = 2036266570;
assign addr[30561] = 2030111710;
assign addr[30562] = 2023795876;
assign addr[30563] = 2017319567;
assign addr[30564] = 2010683297;
assign addr[30565] = 2003887591;
assign addr[30566] = 1996932990;
assign addr[30567] = 1989820044;
assign addr[30568] = 1982549318;
assign addr[30569] = 1975121388;
assign addr[30570] = 1967536842;
assign addr[30571] = 1959796283;
assign addr[30572] = 1951900324;
assign addr[30573] = 1943849591;
assign addr[30574] = 1935644723;
assign addr[30575] = 1927286370;
assign addr[30576] = 1918775195;
assign addr[30577] = 1910111873;
assign addr[30578] = 1901297091;
assign addr[30579] = 1892331547;
assign addr[30580] = 1883215953;
assign addr[30581] = 1873951032;
assign addr[30582] = 1864537518;
assign addr[30583] = 1854976157;
assign addr[30584] = 1845267708;
assign addr[30585] = 1835412941;
assign addr[30586] = 1825412636;
assign addr[30587] = 1815267588;
assign addr[30588] = 1804978599;
assign addr[30589] = 1794546487;
assign addr[30590] = 1783972079;
assign addr[30591] = 1773256212;
assign addr[30592] = 1762399737;
assign addr[30593] = 1751403515;
assign addr[30594] = 1740268417;
assign addr[30595] = 1728995326;
assign addr[30596] = 1717585136;
assign addr[30597] = 1706038753;
assign addr[30598] = 1694357091;
assign addr[30599] = 1682541077;
assign addr[30600] = 1670591647;
assign addr[30601] = 1658509750;
assign addr[30602] = 1646296344;
assign addr[30603] = 1633952396;
assign addr[30604] = 1621478885;
assign addr[30605] = 1608876801;
assign addr[30606] = 1596147143;
assign addr[30607] = 1583290921;
assign addr[30608] = 1570309153;
assign addr[30609] = 1557202869;
assign addr[30610] = 1543973108;
assign addr[30611] = 1530620920;
assign addr[30612] = 1517147363;
assign addr[30613] = 1503553506;
assign addr[30614] = 1489840425;
assign addr[30615] = 1476009210;
assign addr[30616] = 1462060956;
assign addr[30617] = 1447996770;
assign addr[30618] = 1433817766;
assign addr[30619] = 1419525069;
assign addr[30620] = 1405119813;
assign addr[30621] = 1390603139;
assign addr[30622] = 1375976199;
assign addr[30623] = 1361240152;
assign addr[30624] = 1346396168;
assign addr[30625] = 1331445422;
assign addr[30626] = 1316389101;
assign addr[30627] = 1301228398;
assign addr[30628] = 1285964516;
assign addr[30629] = 1270598665;
assign addr[30630] = 1255132063;
assign addr[30631] = 1239565936;
assign addr[30632] = 1223901520;
assign addr[30633] = 1208140056;
assign addr[30634] = 1192282793;
assign addr[30635] = 1176330990;
assign addr[30636] = 1160285911;
assign addr[30637] = 1144148829;
assign addr[30638] = 1127921022;
assign addr[30639] = 1111603778;
assign addr[30640] = 1095198391;
assign addr[30641] = 1078706161;
assign addr[30642] = 1062128397;
assign addr[30643] = 1045466412;
assign addr[30644] = 1028721528;
assign addr[30645] = 1011895073;
assign addr[30646] = 994988380;
assign addr[30647] = 978002791;
assign addr[30648] = 960939653;
assign addr[30649] = 943800318;
assign addr[30650] = 926586145;
assign addr[30651] = 909298500;
assign addr[30652] = 891938752;
assign addr[30653] = 874508280;
assign addr[30654] = 857008464;
assign addr[30655] = 839440693;
assign addr[30656] = 821806359;
assign addr[30657] = 804106861;
assign addr[30658] = 786343603;
assign addr[30659] = 768517992;
assign addr[30660] = 750631442;
assign addr[30661] = 732685372;
assign addr[30662] = 714681204;
assign addr[30663] = 696620367;
assign addr[30664] = 678504291;
assign addr[30665] = 660334415;
assign addr[30666] = 642112178;
assign addr[30667] = 623839025;
assign addr[30668] = 605516406;
assign addr[30669] = 587145773;
assign addr[30670] = 568728583;
assign addr[30671] = 550266296;
assign addr[30672] = 531760377;
assign addr[30673] = 513212292;
assign addr[30674] = 494623513;
assign addr[30675] = 475995513;
assign addr[30676] = 457329769;
assign addr[30677] = 438627762;
assign addr[30678] = 419890975;
assign addr[30679] = 401120892;
assign addr[30680] = 382319004;
assign addr[30681] = 363486799;
assign addr[30682] = 344625773;
assign addr[30683] = 325737419;
assign addr[30684] = 306823237;
assign addr[30685] = 287884725;
assign addr[30686] = 268923386;
assign addr[30687] = 249940723;
assign addr[30688] = 230938242;
assign addr[30689] = 211917448;
assign addr[30690] = 192879850;
assign addr[30691] = 173826959;
assign addr[30692] = 154760284;
assign addr[30693] = 135681337;
assign addr[30694] = 116591632;
assign addr[30695] = 97492681;
assign addr[30696] = 78386000;
assign addr[30697] = 59273104;
assign addr[30698] = 40155507;
assign addr[30699] = 21034727;
assign addr[30700] = 1912278;
assign addr[30701] = -17210322;
assign addr[30702] = -36331557;
assign addr[30703] = -55449912;
assign addr[30704] = -74563870;
assign addr[30705] = -93671915;
assign addr[30706] = -112772533;
assign addr[30707] = -131864208;
assign addr[30708] = -150945428;
assign addr[30709] = -170014678;
assign addr[30710] = -189070447;
assign addr[30711] = -208111224;
assign addr[30712] = -227135500;
assign addr[30713] = -246141764;
assign addr[30714] = -265128512;
assign addr[30715] = -284094236;
assign addr[30716] = -303037433;
assign addr[30717] = -321956601;
assign addr[30718] = -340850240;
assign addr[30719] = -359716852;
assign addr[30720] = -378554940;
assign addr[30721] = -397363011;
assign addr[30722] = -416139574;
assign addr[30723] = -434883140;
assign addr[30724] = -453592221;
assign addr[30725] = -472265336;
assign addr[30726] = -490901003;
assign addr[30727] = -509497745;
assign addr[30728] = -528054086;
assign addr[30729] = -546568556;
assign addr[30730] = -565039687;
assign addr[30731] = -583466013;
assign addr[30732] = -601846074;
assign addr[30733] = -620178412;
assign addr[30734] = -638461574;
assign addr[30735] = -656694110;
assign addr[30736] = -674874574;
assign addr[30737] = -693001525;
assign addr[30738] = -711073524;
assign addr[30739] = -729089140;
assign addr[30740] = -747046944;
assign addr[30741] = -764945512;
assign addr[30742] = -782783424;
assign addr[30743] = -800559266;
assign addr[30744] = -818271628;
assign addr[30745] = -835919107;
assign addr[30746] = -853500302;
assign addr[30747] = -871013820;
assign addr[30748] = -888458272;
assign addr[30749] = -905832274;
assign addr[30750] = -923134450;
assign addr[30751] = -940363427;
assign addr[30752] = -957517838;
assign addr[30753] = -974596324;
assign addr[30754] = -991597531;
assign addr[30755] = -1008520110;
assign addr[30756] = -1025362720;
assign addr[30757] = -1042124025;
assign addr[30758] = -1058802695;
assign addr[30759] = -1075397409;
assign addr[30760] = -1091906851;
assign addr[30761] = -1108329711;
assign addr[30762] = -1124664687;
assign addr[30763] = -1140910484;
assign addr[30764] = -1157065814;
assign addr[30765] = -1173129396;
assign addr[30766] = -1189099956;
assign addr[30767] = -1204976227;
assign addr[30768] = -1220756951;
assign addr[30769] = -1236440877;
assign addr[30770] = -1252026760;
assign addr[30771] = -1267513365;
assign addr[30772] = -1282899464;
assign addr[30773] = -1298183838;
assign addr[30774] = -1313365273;
assign addr[30775] = -1328442566;
assign addr[30776] = -1343414522;
assign addr[30777] = -1358279953;
assign addr[30778] = -1373037681;
assign addr[30779] = -1387686535;
assign addr[30780] = -1402225355;
assign addr[30781] = -1416652986;
assign addr[30782] = -1430968286;
assign addr[30783] = -1445170118;
assign addr[30784] = -1459257358;
assign addr[30785] = -1473228887;
assign addr[30786] = -1487083598;
assign addr[30787] = -1500820393;
assign addr[30788] = -1514438181;
assign addr[30789] = -1527935884;
assign addr[30790] = -1541312431;
assign addr[30791] = -1554566762;
assign addr[30792] = -1567697824;
assign addr[30793] = -1580704578;
assign addr[30794] = -1593585992;
assign addr[30795] = -1606341043;
assign addr[30796] = -1618968722;
assign addr[30797] = -1631468027;
assign addr[30798] = -1643837966;
assign addr[30799] = -1656077559;
assign addr[30800] = -1668185835;
assign addr[30801] = -1680161834;
assign addr[30802] = -1692004606;
assign addr[30803] = -1703713213;
assign addr[30804] = -1715286726;
assign addr[30805] = -1726724227;
assign addr[30806] = -1738024810;
assign addr[30807] = -1749187577;
assign addr[30808] = -1760211645;
assign addr[30809] = -1771096139;
assign addr[30810] = -1781840195;
assign addr[30811] = -1792442963;
assign addr[30812] = -1802903601;
assign addr[30813] = -1813221279;
assign addr[30814] = -1823395180;
assign addr[30815] = -1833424497;
assign addr[30816] = -1843308435;
assign addr[30817] = -1853046210;
assign addr[30818] = -1862637049;
assign addr[30819] = -1872080193;
assign addr[30820] = -1881374892;
assign addr[30821] = -1890520410;
assign addr[30822] = -1899516021;
assign addr[30823] = -1908361011;
assign addr[30824] = -1917054681;
assign addr[30825] = -1925596340;
assign addr[30826] = -1933985310;
assign addr[30827] = -1942220928;
assign addr[30828] = -1950302539;
assign addr[30829] = -1958229503;
assign addr[30830] = -1966001192;
assign addr[30831] = -1973616989;
assign addr[30832] = -1981076290;
assign addr[30833] = -1988378503;
assign addr[30834] = -1995523051;
assign addr[30835] = -2002509365;
assign addr[30836] = -2009336893;
assign addr[30837] = -2016005093;
assign addr[30838] = -2022513436;
assign addr[30839] = -2028861406;
assign addr[30840] = -2035048499;
assign addr[30841] = -2041074226;
assign addr[30842] = -2046938108;
assign addr[30843] = -2052639680;
assign addr[30844] = -2058178491;
assign addr[30845] = -2063554100;
assign addr[30846] = -2068766083;
assign addr[30847] = -2073814024;
assign addr[30848] = -2078697525;
assign addr[30849] = -2083416198;
assign addr[30850] = -2087969669;
assign addr[30851] = -2092357577;
assign addr[30852] = -2096579573;
assign addr[30853] = -2100635323;
assign addr[30854] = -2104524506;
assign addr[30855] = -2108246813;
assign addr[30856] = -2111801949;
assign addr[30857] = -2115189632;
assign addr[30858] = -2118409593;
assign addr[30859] = -2121461578;
assign addr[30860] = -2124345343;
assign addr[30861] = -2127060661;
assign addr[30862] = -2129607316;
assign addr[30863] = -2131985106;
assign addr[30864] = -2134193842;
assign addr[30865] = -2136233350;
assign addr[30866] = -2138103468;
assign addr[30867] = -2139804048;
assign addr[30868] = -2141334954;
assign addr[30869] = -2142696065;
assign addr[30870] = -2143887273;
assign addr[30871] = -2144908484;
assign addr[30872] = -2145759618;
assign addr[30873] = -2146440605;
assign addr[30874] = -2146951393;
assign addr[30875] = -2147291941;
assign addr[30876] = -2147462221;
assign addr[30877] = -2147462221;
assign addr[30878] = -2147291941;
assign addr[30879] = -2146951393;
assign addr[30880] = -2146440605;
assign addr[30881] = -2145759618;
assign addr[30882] = -2144908484;
assign addr[30883] = -2143887273;
assign addr[30884] = -2142696065;
assign addr[30885] = -2141334954;
assign addr[30886] = -2139804048;
assign addr[30887] = -2138103468;
assign addr[30888] = -2136233350;
assign addr[30889] = -2134193842;
assign addr[30890] = -2131985106;
assign addr[30891] = -2129607316;
assign addr[30892] = -2127060661;
assign addr[30893] = -2124345343;
assign addr[30894] = -2121461578;
assign addr[30895] = -2118409593;
assign addr[30896] = -2115189632;
assign addr[30897] = -2111801949;
assign addr[30898] = -2108246813;
assign addr[30899] = -2104524506;
assign addr[30900] = -2100635323;
assign addr[30901] = -2096579573;
assign addr[30902] = -2092357577;
assign addr[30903] = -2087969669;
assign addr[30904] = -2083416198;
assign addr[30905] = -2078697525;
assign addr[30906] = -2073814024;
assign addr[30907] = -2068766083;
assign addr[30908] = -2063554100;
assign addr[30909] = -2058178491;
assign addr[30910] = -2052639680;
assign addr[30911] = -2046938108;
assign addr[30912] = -2041074226;
assign addr[30913] = -2035048499;
assign addr[30914] = -2028861406;
assign addr[30915] = -2022513436;
assign addr[30916] = -2016005093;
assign addr[30917] = -2009336893;
assign addr[30918] = -2002509365;
assign addr[30919] = -1995523051;
assign addr[30920] = -1988378503;
assign addr[30921] = -1981076290;
assign addr[30922] = -1973616989;
assign addr[30923] = -1966001192;
assign addr[30924] = -1958229503;
assign addr[30925] = -1950302539;
assign addr[30926] = -1942220928;
assign addr[30927] = -1933985310;
assign addr[30928] = -1925596340;
assign addr[30929] = -1917054681;
assign addr[30930] = -1908361011;
assign addr[30931] = -1899516021;
assign addr[30932] = -1890520410;
assign addr[30933] = -1881374892;
assign addr[30934] = -1872080193;
assign addr[30935] = -1862637049;
assign addr[30936] = -1853046210;
assign addr[30937] = -1843308435;
assign addr[30938] = -1833424497;
assign addr[30939] = -1823395180;
assign addr[30940] = -1813221279;
assign addr[30941] = -1802903601;
assign addr[30942] = -1792442963;
assign addr[30943] = -1781840195;
assign addr[30944] = -1771096139;
assign addr[30945] = -1760211645;
assign addr[30946] = -1749187577;
assign addr[30947] = -1738024810;
assign addr[30948] = -1726724227;
assign addr[30949] = -1715286726;
assign addr[30950] = -1703713213;
assign addr[30951] = -1692004606;
assign addr[30952] = -1680161834;
assign addr[30953] = -1668185835;
assign addr[30954] = -1656077559;
assign addr[30955] = -1643837966;
assign addr[30956] = -1631468027;
assign addr[30957] = -1618968722;
assign addr[30958] = -1606341043;
assign addr[30959] = -1593585992;
assign addr[30960] = -1580704578;
assign addr[30961] = -1567697824;
assign addr[30962] = -1554566762;
assign addr[30963] = -1541312431;
assign addr[30964] = -1527935884;
assign addr[30965] = -1514438181;
assign addr[30966] = -1500820393;
assign addr[30967] = -1487083598;
assign addr[30968] = -1473228887;
assign addr[30969] = -1459257358;
assign addr[30970] = -1445170118;
assign addr[30971] = -1430968286;
assign addr[30972] = -1416652986;
assign addr[30973] = -1402225355;
assign addr[30974] = -1387686535;
assign addr[30975] = -1373037681;
assign addr[30976] = -1358279953;
assign addr[30977] = -1343414522;
assign addr[30978] = -1328442566;
assign addr[30979] = -1313365273;
assign addr[30980] = -1298183838;
assign addr[30981] = -1282899464;
assign addr[30982] = -1267513365;
assign addr[30983] = -1252026760;
assign addr[30984] = -1236440877;
assign addr[30985] = -1220756951;
assign addr[30986] = -1204976227;
assign addr[30987] = -1189099956;
assign addr[30988] = -1173129396;
assign addr[30989] = -1157065814;
assign addr[30990] = -1140910484;
assign addr[30991] = -1124664687;
assign addr[30992] = -1108329711;
assign addr[30993] = -1091906851;
assign addr[30994] = -1075397409;
assign addr[30995] = -1058802695;
assign addr[30996] = -1042124025;
assign addr[30997] = -1025362720;
assign addr[30998] = -1008520110;
assign addr[30999] = -991597531;
assign addr[31000] = -974596324;
assign addr[31001] = -957517838;
assign addr[31002] = -940363427;
assign addr[31003] = -923134450;
assign addr[31004] = -905832274;
assign addr[31005] = -888458272;
assign addr[31006] = -871013820;
assign addr[31007] = -853500302;
assign addr[31008] = -835919107;
assign addr[31009] = -818271628;
assign addr[31010] = -800559266;
assign addr[31011] = -782783424;
assign addr[31012] = -764945512;
assign addr[31013] = -747046944;
assign addr[31014] = -729089140;
assign addr[31015] = -711073524;
assign addr[31016] = -693001525;
assign addr[31017] = -674874574;
assign addr[31018] = -656694110;
assign addr[31019] = -638461574;
assign addr[31020] = -620178412;
assign addr[31021] = -601846074;
assign addr[31022] = -583466013;
assign addr[31023] = -565039687;
assign addr[31024] = -546568556;
assign addr[31025] = -528054086;
assign addr[31026] = -509497745;
assign addr[31027] = -490901003;
assign addr[31028] = -472265336;
assign addr[31029] = -453592221;
assign addr[31030] = -434883140;
assign addr[31031] = -416139574;
assign addr[31032] = -397363011;
assign addr[31033] = -378554940;
assign addr[31034] = -359716852;
assign addr[31035] = -340850240;
assign addr[31036] = -321956601;
assign addr[31037] = -303037433;
assign addr[31038] = -284094236;
assign addr[31039] = -265128512;
assign addr[31040] = -246141764;
assign addr[31041] = -227135500;
assign addr[31042] = -208111224;
assign addr[31043] = -189070447;
assign addr[31044] = -170014678;
assign addr[31045] = -150945428;
assign addr[31046] = -131864208;
assign addr[31047] = -112772533;
assign addr[31048] = -93671915;
assign addr[31049] = -74563870;
assign addr[31050] = -55449912;
assign addr[31051] = -36331557;
assign addr[31052] = -17210322;
assign addr[31053] = 1912278;
assign addr[31054] = 21034727;
assign addr[31055] = 40155507;
assign addr[31056] = 59273104;
assign addr[31057] = 78386000;
assign addr[31058] = 97492681;
assign addr[31059] = 116591632;
assign addr[31060] = 135681337;
assign addr[31061] = 154760284;
assign addr[31062] = 173826959;
assign addr[31063] = 192879850;
assign addr[31064] = 211917448;
assign addr[31065] = 230938242;
assign addr[31066] = 249940723;
assign addr[31067] = 268923386;
assign addr[31068] = 287884725;
assign addr[31069] = 306823237;
assign addr[31070] = 325737419;
assign addr[31071] = 344625773;
assign addr[31072] = 363486799;
assign addr[31073] = 382319004;
assign addr[31074] = 401120892;
assign addr[31075] = 419890975;
assign addr[31076] = 438627762;
assign addr[31077] = 457329769;
assign addr[31078] = 475995513;
assign addr[31079] = 494623513;
assign addr[31080] = 513212292;
assign addr[31081] = 531760377;
assign addr[31082] = 550266296;
assign addr[31083] = 568728583;
assign addr[31084] = 587145773;
assign addr[31085] = 605516406;
assign addr[31086] = 623839025;
assign addr[31087] = 642112178;
assign addr[31088] = 660334415;
assign addr[31089] = 678504291;
assign addr[31090] = 696620367;
assign addr[31091] = 714681204;
assign addr[31092] = 732685372;
assign addr[31093] = 750631442;
assign addr[31094] = 768517992;
assign addr[31095] = 786343603;
assign addr[31096] = 804106861;
assign addr[31097] = 821806359;
assign addr[31098] = 839440693;
assign addr[31099] = 857008464;
assign addr[31100] = 874508280;
assign addr[31101] = 891938752;
assign addr[31102] = 909298500;
assign addr[31103] = 926586145;
assign addr[31104] = 943800318;
assign addr[31105] = 960939653;
assign addr[31106] = 978002791;
assign addr[31107] = 994988380;
assign addr[31108] = 1011895073;
assign addr[31109] = 1028721528;
assign addr[31110] = 1045466412;
assign addr[31111] = 1062128397;
assign addr[31112] = 1078706161;
assign addr[31113] = 1095198391;
assign addr[31114] = 1111603778;
assign addr[31115] = 1127921022;
assign addr[31116] = 1144148829;
assign addr[31117] = 1160285911;
assign addr[31118] = 1176330990;
assign addr[31119] = 1192282793;
assign addr[31120] = 1208140056;
assign addr[31121] = 1223901520;
assign addr[31122] = 1239565936;
assign addr[31123] = 1255132063;
assign addr[31124] = 1270598665;
assign addr[31125] = 1285964516;
assign addr[31126] = 1301228398;
assign addr[31127] = 1316389101;
assign addr[31128] = 1331445422;
assign addr[31129] = 1346396168;
assign addr[31130] = 1361240152;
assign addr[31131] = 1375976199;
assign addr[31132] = 1390603139;
assign addr[31133] = 1405119813;
assign addr[31134] = 1419525069;
assign addr[31135] = 1433817766;
assign addr[31136] = 1447996770;
assign addr[31137] = 1462060956;
assign addr[31138] = 1476009210;
assign addr[31139] = 1489840425;
assign addr[31140] = 1503553506;
assign addr[31141] = 1517147363;
assign addr[31142] = 1530620920;
assign addr[31143] = 1543973108;
assign addr[31144] = 1557202869;
assign addr[31145] = 1570309153;
assign addr[31146] = 1583290921;
assign addr[31147] = 1596147143;
assign addr[31148] = 1608876801;
assign addr[31149] = 1621478885;
assign addr[31150] = 1633952396;
assign addr[31151] = 1646296344;
assign addr[31152] = 1658509750;
assign addr[31153] = 1670591647;
assign addr[31154] = 1682541077;
assign addr[31155] = 1694357091;
assign addr[31156] = 1706038753;
assign addr[31157] = 1717585136;
assign addr[31158] = 1728995326;
assign addr[31159] = 1740268417;
assign addr[31160] = 1751403515;
assign addr[31161] = 1762399737;
assign addr[31162] = 1773256212;
assign addr[31163] = 1783972079;
assign addr[31164] = 1794546487;
assign addr[31165] = 1804978599;
assign addr[31166] = 1815267588;
assign addr[31167] = 1825412636;
assign addr[31168] = 1835412941;
assign addr[31169] = 1845267708;
assign addr[31170] = 1854976157;
assign addr[31171] = 1864537518;
assign addr[31172] = 1873951032;
assign addr[31173] = 1883215953;
assign addr[31174] = 1892331547;
assign addr[31175] = 1901297091;
assign addr[31176] = 1910111873;
assign addr[31177] = 1918775195;
assign addr[31178] = 1927286370;
assign addr[31179] = 1935644723;
assign addr[31180] = 1943849591;
assign addr[31181] = 1951900324;
assign addr[31182] = 1959796283;
assign addr[31183] = 1967536842;
assign addr[31184] = 1975121388;
assign addr[31185] = 1982549318;
assign addr[31186] = 1989820044;
assign addr[31187] = 1996932990;
assign addr[31188] = 2003887591;
assign addr[31189] = 2010683297;
assign addr[31190] = 2017319567;
assign addr[31191] = 2023795876;
assign addr[31192] = 2030111710;
assign addr[31193] = 2036266570;
assign addr[31194] = 2042259965;
assign addr[31195] = 2048091422;
assign addr[31196] = 2053760478;
assign addr[31197] = 2059266683;
assign addr[31198] = 2064609600;
assign addr[31199] = 2069788807;
assign addr[31200] = 2074803892;
assign addr[31201] = 2079654458;
assign addr[31202] = 2084340120;
assign addr[31203] = 2088860507;
assign addr[31204] = 2093215260;
assign addr[31205] = 2097404033;
assign addr[31206] = 2101426496;
assign addr[31207] = 2105282327;
assign addr[31208] = 2108971223;
assign addr[31209] = 2112492891;
assign addr[31210] = 2115847050;
assign addr[31211] = 2119033436;
assign addr[31212] = 2122051796;
assign addr[31213] = 2124901890;
assign addr[31214] = 2127583492;
assign addr[31215] = 2130096389;
assign addr[31216] = 2132440383;
assign addr[31217] = 2134615288;
assign addr[31218] = 2136620930;
assign addr[31219] = 2138457152;
assign addr[31220] = 2140123807;
assign addr[31221] = 2141620763;
assign addr[31222] = 2142947902;
assign addr[31223] = 2144105118;
assign addr[31224] = 2145092320;
assign addr[31225] = 2145909429;
assign addr[31226] = 2146556380;
assign addr[31227] = 2147033123;
assign addr[31228] = 2147339619;
assign addr[31229] = 2147475844;
assign addr[31230] = 2147441787;
assign addr[31231] = 2147237452;
assign addr[31232] = 2146862854;
assign addr[31233] = 2146318022;
assign addr[31234] = 2145603001;
assign addr[31235] = 2144717846;
assign addr[31236] = 2143662628;
assign addr[31237] = 2142437431;
assign addr[31238] = 2141042352;
assign addr[31239] = 2139477502;
assign addr[31240] = 2137743003;
assign addr[31241] = 2135838995;
assign addr[31242] = 2133765628;
assign addr[31243] = 2131523066;
assign addr[31244] = 2129111488;
assign addr[31245] = 2126531084;
assign addr[31246] = 2123782059;
assign addr[31247] = 2120864631;
assign addr[31248] = 2117779031;
assign addr[31249] = 2114525505;
assign addr[31250] = 2111104309;
assign addr[31251] = 2107515716;
assign addr[31252] = 2103760010;
assign addr[31253] = 2099837489;
assign addr[31254] = 2095748463;
assign addr[31255] = 2091493257;
assign addr[31256] = 2087072209;
assign addr[31257] = 2082485668;
assign addr[31258] = 2077733999;
assign addr[31259] = 2072817579;
assign addr[31260] = 2067736796;
assign addr[31261] = 2062492055;
assign addr[31262] = 2057083771;
assign addr[31263] = 2051512372;
assign addr[31264] = 2045778302;
assign addr[31265] = 2039882013;
assign addr[31266] = 2033823974;
assign addr[31267] = 2027604666;
assign addr[31268] = 2021224581;
assign addr[31269] = 2014684225;
assign addr[31270] = 2007984117;
assign addr[31271] = 2001124788;
assign addr[31272] = 1994106782;
assign addr[31273] = 1986930656;
assign addr[31274] = 1979596978;
assign addr[31275] = 1972106330;
assign addr[31276] = 1964459306;
assign addr[31277] = 1956656513;
assign addr[31278] = 1948698568;
assign addr[31279] = 1940586104;
assign addr[31280] = 1932319763;
assign addr[31281] = 1923900201;
assign addr[31282] = 1915328086;
assign addr[31283] = 1906604097;
assign addr[31284] = 1897728925;
assign addr[31285] = 1888703276;
assign addr[31286] = 1879527863;
assign addr[31287] = 1870203416;
assign addr[31288] = 1860730673;
assign addr[31289] = 1851110385;
assign addr[31290] = 1841343316;
assign addr[31291] = 1831430239;
assign addr[31292] = 1821371941;
assign addr[31293] = 1811169220;
assign addr[31294] = 1800822883;
assign addr[31295] = 1790333753;
assign addr[31296] = 1779702660;
assign addr[31297] = 1768930447;
assign addr[31298] = 1758017969;
assign addr[31299] = 1746966091;
assign addr[31300] = 1735775690;
assign addr[31301] = 1724447652;
assign addr[31302] = 1712982875;
assign addr[31303] = 1701382270;
assign addr[31304] = 1689646755;
assign addr[31305] = 1677777262;
assign addr[31306] = 1665774731;
assign addr[31307] = 1653640115;
assign addr[31308] = 1641374375;
assign addr[31309] = 1628978484;
assign addr[31310] = 1616453425;
assign addr[31311] = 1603800191;
assign addr[31312] = 1591019785;
assign addr[31313] = 1578113222;
assign addr[31314] = 1565081523;
assign addr[31315] = 1551925723;
assign addr[31316] = 1538646865;
assign addr[31317] = 1525246002;
assign addr[31318] = 1511724196;
assign addr[31319] = 1498082520;
assign addr[31320] = 1484322054;
assign addr[31321] = 1470443891;
assign addr[31322] = 1456449131;
assign addr[31323] = 1442338884;
assign addr[31324] = 1428114267;
assign addr[31325] = 1413776410;
assign addr[31326] = 1399326449;
assign addr[31327] = 1384765530;
assign addr[31328] = 1370094808;
assign addr[31329] = 1355315445;
assign addr[31330] = 1340428615;
assign addr[31331] = 1325435496;
assign addr[31332] = 1310337279;
assign addr[31333] = 1295135159;
assign addr[31334] = 1279830344;
assign addr[31335] = 1264424045;
assign addr[31336] = 1248917486;
assign addr[31337] = 1233311895;
assign addr[31338] = 1217608510;
assign addr[31339] = 1201808576;
assign addr[31340] = 1185913346;
assign addr[31341] = 1169924081;
assign addr[31342] = 1153842047;
assign addr[31343] = 1137668521;
assign addr[31344] = 1121404785;
assign addr[31345] = 1105052128;
assign addr[31346] = 1088611847;
assign addr[31347] = 1072085246;
assign addr[31348] = 1055473635;
assign addr[31349] = 1038778332;
assign addr[31350] = 1022000660;
assign addr[31351] = 1005141949;
assign addr[31352] = 988203537;
assign addr[31353] = 971186766;
assign addr[31354] = 954092986;
assign addr[31355] = 936923553;
assign addr[31356] = 919679827;
assign addr[31357] = 902363176;
assign addr[31358] = 884974973;
assign addr[31359] = 867516597;
assign addr[31360] = 849989433;
assign addr[31361] = 832394869;
assign addr[31362] = 814734301;
assign addr[31363] = 797009130;
assign addr[31364] = 779220762;
assign addr[31365] = 761370605;
assign addr[31366] = 743460077;
assign addr[31367] = 725490597;
assign addr[31368] = 707463589;
assign addr[31369] = 689380485;
assign addr[31370] = 671242716;
assign addr[31371] = 653051723;
assign addr[31372] = 634808946;
assign addr[31373] = 616515832;
assign addr[31374] = 598173833;
assign addr[31375] = 579784402;
assign addr[31376] = 561348998;
assign addr[31377] = 542869083;
assign addr[31378] = 524346121;
assign addr[31379] = 505781581;
assign addr[31380] = 487176937;
assign addr[31381] = 468533662;
assign addr[31382] = 449853235;
assign addr[31383] = 431137138;
assign addr[31384] = 412386854;
assign addr[31385] = 393603870;
assign addr[31386] = 374789676;
assign addr[31387] = 355945764;
assign addr[31388] = 337073627;
assign addr[31389] = 318174762;
assign addr[31390] = 299250668;
assign addr[31391] = 280302845;
assign addr[31392] = 261332796;
assign addr[31393] = 242342025;
assign addr[31394] = 223332037;
assign addr[31395] = 204304341;
assign addr[31396] = 185260444;
assign addr[31397] = 166201858;
assign addr[31398] = 147130093;
assign addr[31399] = 128046661;
assign addr[31400] = 108953076;
assign addr[31401] = 89850852;
assign addr[31402] = 70741503;
assign addr[31403] = 51626544;
assign addr[31404] = 32507492;
assign addr[31405] = 13385863;
assign addr[31406] = -5736829;
assign addr[31407] = -24859065;
assign addr[31408] = -43979330;
assign addr[31409] = -63096108;
assign addr[31410] = -82207882;
assign addr[31411] = -101313138;
assign addr[31412] = -120410361;
assign addr[31413] = -139498035;
assign addr[31414] = -158574649;
assign addr[31415] = -177638688;
assign addr[31416] = -196688642;
assign addr[31417] = -215722999;
assign addr[31418] = -234740251;
assign addr[31419] = -253738890;
assign addr[31420] = -272717408;
assign addr[31421] = -291674302;
assign addr[31422] = -310608068;
assign addr[31423] = -329517204;
assign addr[31424] = -348400212;
assign addr[31425] = -367255594;
assign addr[31426] = -386081854;
assign addr[31427] = -404877501;
assign addr[31428] = -423641043;
assign addr[31429] = -442370993;
assign addr[31430] = -461065866;
assign addr[31431] = -479724180;
assign addr[31432] = -498344454;
assign addr[31433] = -516925212;
assign addr[31434] = -535464981;
assign addr[31435] = -553962291;
assign addr[31436] = -572415676;
assign addr[31437] = -590823671;
assign addr[31438] = -609184818;
assign addr[31439] = -627497660;
assign addr[31440] = -645760745;
assign addr[31441] = -663972625;
assign addr[31442] = -682131857;
assign addr[31443] = -700236999;
assign addr[31444] = -718286617;
assign addr[31445] = -736279279;
assign addr[31446] = -754213559;
assign addr[31447] = -772088034;
assign addr[31448] = -789901288;
assign addr[31449] = -807651907;
assign addr[31450] = -825338484;
assign addr[31451] = -842959617;
assign addr[31452] = -860513908;
assign addr[31453] = -877999966;
assign addr[31454] = -895416404;
assign addr[31455] = -912761841;
assign addr[31456] = -930034901;
assign addr[31457] = -947234215;
assign addr[31458] = -964358420;
assign addr[31459] = -981406156;
assign addr[31460] = -998376073;
assign addr[31461] = -1015266825;
assign addr[31462] = -1032077073;
assign addr[31463] = -1048805483;
assign addr[31464] = -1065450729;
assign addr[31465] = -1082011492;
assign addr[31466] = -1098486458;
assign addr[31467] = -1114874320;
assign addr[31468] = -1131173780;
assign addr[31469] = -1147383544;
assign addr[31470] = -1163502328;
assign addr[31471] = -1179528853;
assign addr[31472] = -1195461849;
assign addr[31473] = -1211300053;
assign addr[31474] = -1227042207;
assign addr[31475] = -1242687064;
assign addr[31476] = -1258233384;
assign addr[31477] = -1273679934;
assign addr[31478] = -1289025489;
assign addr[31479] = -1304268832;
assign addr[31480] = -1319408754;
assign addr[31481] = -1334444055;
assign addr[31482] = -1349373543;
assign addr[31483] = -1364196034;
assign addr[31484] = -1378910353;
assign addr[31485] = -1393515332;
assign addr[31486] = -1408009814;
assign addr[31487] = -1422392650;
assign addr[31488] = -1436662698;
assign addr[31489] = -1450818828;
assign addr[31490] = -1464859917;
assign addr[31491] = -1478784851;
assign addr[31492] = -1492592527;
assign addr[31493] = -1506281850;
assign addr[31494] = -1519851733;
assign addr[31495] = -1533301101;
assign addr[31496] = -1546628888;
assign addr[31497] = -1559834037;
assign addr[31498] = -1572915501;
assign addr[31499] = -1585872242;
assign addr[31500] = -1598703233;
assign addr[31501] = -1611407456;
assign addr[31502] = -1623983905;
assign addr[31503] = -1636431582;
assign addr[31504] = -1648749499;
assign addr[31505] = -1660936681;
assign addr[31506] = -1672992161;
assign addr[31507] = -1684914983;
assign addr[31508] = -1696704201;
assign addr[31509] = -1708358881;
assign addr[31510] = -1719878099;
assign addr[31511] = -1731260941;
assign addr[31512] = -1742506504;
assign addr[31513] = -1753613897;
assign addr[31514] = -1764582240;
assign addr[31515] = -1775410662;
assign addr[31516] = -1786098304;
assign addr[31517] = -1796644320;
assign addr[31518] = -1807047873;
assign addr[31519] = -1817308138;
assign addr[31520] = -1827424302;
assign addr[31521] = -1837395562;
assign addr[31522] = -1847221128;
assign addr[31523] = -1856900221;
assign addr[31524] = -1866432072;
assign addr[31525] = -1875815927;
assign addr[31526] = -1885051042;
assign addr[31527] = -1894136683;
assign addr[31528] = -1903072131;
assign addr[31529] = -1911856677;
assign addr[31530] = -1920489624;
assign addr[31531] = -1928970288;
assign addr[31532] = -1937297997;
assign addr[31533] = -1945472089;
assign addr[31534] = -1953491918;
assign addr[31535] = -1961356847;
assign addr[31536] = -1969066252;
assign addr[31537] = -1976619522;
assign addr[31538] = -1984016058;
assign addr[31539] = -1991255274;
assign addr[31540] = -1998336596;
assign addr[31541] = -2005259462;
assign addr[31542] = -2012023322;
assign addr[31543] = -2018627642;
assign addr[31544] = -2025071897;
assign addr[31545] = -2031355576;
assign addr[31546] = -2037478181;
assign addr[31547] = -2043439226;
assign addr[31548] = -2049238240;
assign addr[31549] = -2054874761;
assign addr[31550] = -2060348343;
assign addr[31551] = -2065658552;
assign addr[31552] = -2070804967;
assign addr[31553] = -2075787180;
assign addr[31554] = -2080604795;
assign addr[31555] = -2085257431;
assign addr[31556] = -2089744719;
assign addr[31557] = -2094066304;
assign addr[31558] = -2098221841;
assign addr[31559] = -2102211002;
assign addr[31560] = -2106033471;
assign addr[31561] = -2109688944;
assign addr[31562] = -2113177132;
assign addr[31563] = -2116497758;
assign addr[31564] = -2119650558;
assign addr[31565] = -2122635283;
assign addr[31566] = -2125451696;
assign addr[31567] = -2128099574;
assign addr[31568] = -2130578706;
assign addr[31569] = -2132888897;
assign addr[31570] = -2135029962;
assign addr[31571] = -2137001733;
assign addr[31572] = -2138804053;
assign addr[31573] = -2140436778;
assign addr[31574] = -2141899780;
assign addr[31575] = -2143192942;
assign addr[31576] = -2144316162;
assign addr[31577] = -2145269351;
assign addr[31578] = -2146052433;
assign addr[31579] = -2146665347;
assign addr[31580] = -2147108043;
assign addr[31581] = -2147380486;
assign addr[31582] = -2147482655;
assign addr[31583] = -2147414542;
assign addr[31584] = -2147176152;
assign addr[31585] = -2146767505;
assign addr[31586] = -2146188631;
assign addr[31587] = -2145439578;
assign addr[31588] = -2144520405;
assign addr[31589] = -2143431184;
assign addr[31590] = -2142172003;
assign addr[31591] = -2140742960;
assign addr[31592] = -2139144169;
assign addr[31593] = -2137375758;
assign addr[31594] = -2135437865;
assign addr[31595] = -2133330646;
assign addr[31596] = -2131054266;
assign addr[31597] = -2128608907;
assign addr[31598] = -2125994762;
assign addr[31599] = -2123212038;
assign addr[31600] = -2120260957;
assign addr[31601] = -2117141752;
assign addr[31602] = -2113854671;
assign addr[31603] = -2110399974;
assign addr[31604] = -2106777935;
assign addr[31605] = -2102988841;
assign addr[31606] = -2099032994;
assign addr[31607] = -2094910706;
assign addr[31608] = -2090622304;
assign addr[31609] = -2086168128;
assign addr[31610] = -2081548533;
assign addr[31611] = -2076763883;
assign addr[31612] = -2071814558;
assign addr[31613] = -2066700952;
assign addr[31614] = -2061423468;
assign addr[31615] = -2055982526;
assign addr[31616] = -2050378558;
assign addr[31617] = -2044612007;
assign addr[31618] = -2038683330;
assign addr[31619] = -2032592999;
assign addr[31620] = -2026341495;
assign addr[31621] = -2019929315;
assign addr[31622] = -2013356967;
assign addr[31623] = -2006624971;
assign addr[31624] = -1999733863;
assign addr[31625] = -1992684188;
assign addr[31626] = -1985476506;
assign addr[31627] = -1978111387;
assign addr[31628] = -1970589416;
assign addr[31629] = -1962911189;
assign addr[31630] = -1955077316;
assign addr[31631] = -1947088417;
assign addr[31632] = -1938945125;
assign addr[31633] = -1930648088;
assign addr[31634] = -1922197961;
assign addr[31635] = -1913595416;
assign addr[31636] = -1904841135;
assign addr[31637] = -1895935811;
assign addr[31638] = -1886880151;
assign addr[31639] = -1877674873;
assign addr[31640] = -1868320707;
assign addr[31641] = -1858818395;
assign addr[31642] = -1849168689;
assign addr[31643] = -1839372356;
assign addr[31644] = -1829430172;
assign addr[31645] = -1819342925;
assign addr[31646] = -1809111415;
assign addr[31647] = -1798736454;
assign addr[31648] = -1788218865;
assign addr[31649] = -1777559480;
assign addr[31650] = -1766759146;
assign addr[31651] = -1755818718;
assign addr[31652] = -1744739065;
assign addr[31653] = -1733521064;
assign addr[31654] = -1722165606;
assign addr[31655] = -1710673591;
assign addr[31656] = -1699045930;
assign addr[31657] = -1687283545;
assign addr[31658] = -1675387369;
assign addr[31659] = -1663358344;
assign addr[31660] = -1651197426;
assign addr[31661] = -1638905577;
assign addr[31662] = -1626483774;
assign addr[31663] = -1613933000;
assign addr[31664] = -1601254251;
assign addr[31665] = -1588448533;
assign addr[31666] = -1575516860;
assign addr[31667] = -1562460258;
assign addr[31668] = -1549279763;
assign addr[31669] = -1535976419;
assign addr[31670] = -1522551282;
assign addr[31671] = -1509005416;
assign addr[31672] = -1495339895;
assign addr[31673] = -1481555802;
assign addr[31674] = -1467654232;
assign addr[31675] = -1453636285;
assign addr[31676] = -1439503074;
assign addr[31677] = -1425255719;
assign addr[31678] = -1410895350;
assign addr[31679] = -1396423105;
assign addr[31680] = -1381840133;
assign addr[31681] = -1367147589;
assign addr[31682] = -1352346639;
assign addr[31683] = -1337438456;
assign addr[31684] = -1322424222;
assign addr[31685] = -1307305128;
assign addr[31686] = -1292082373;
assign addr[31687] = -1276757164;
assign addr[31688] = -1261330715;
assign addr[31689] = -1245804251;
assign addr[31690] = -1230179002;
assign addr[31691] = -1214456207;
assign addr[31692] = -1198637114;
assign addr[31693] = -1182722976;
assign addr[31694] = -1166715055;
assign addr[31695] = -1150614620;
assign addr[31696] = -1134422949;
assign addr[31697] = -1118141326;
assign addr[31698] = -1101771040;
assign addr[31699] = -1085313391;
assign addr[31700] = -1068769683;
assign addr[31701] = -1052141228;
assign addr[31702] = -1035429345;
assign addr[31703] = -1018635358;
assign addr[31704] = -1001760600;
assign addr[31705] = -984806408;
assign addr[31706] = -967774128;
assign addr[31707] = -950665109;
assign addr[31708] = -933480707;
assign addr[31709] = -916222287;
assign addr[31710] = -898891215;
assign addr[31711] = -881488868;
assign addr[31712] = -864016623;
assign addr[31713] = -846475867;
assign addr[31714] = -828867991;
assign addr[31715] = -811194391;
assign addr[31716] = -793456467;
assign addr[31717] = -775655628;
assign addr[31718] = -757793284;
assign addr[31719] = -739870851;
assign addr[31720] = -721889752;
assign addr[31721] = -703851410;
assign addr[31722] = -685757258;
assign addr[31723] = -667608730;
assign addr[31724] = -649407264;
assign addr[31725] = -631154304;
assign addr[31726] = -612851297;
assign addr[31727] = -594499695;
assign addr[31728] = -576100953;
assign addr[31729] = -557656529;
assign addr[31730] = -539167887;
assign addr[31731] = -520636492;
assign addr[31732] = -502063814;
assign addr[31733] = -483451325;
assign addr[31734] = -464800501;
assign addr[31735] = -446112822;
assign addr[31736] = -427389768;
assign addr[31737] = -408632825;
assign addr[31738] = -389843480;
assign addr[31739] = -371023223;
assign addr[31740] = -352173546;
assign addr[31741] = -333295944;
assign addr[31742] = -314391913;
assign addr[31743] = -295462954;
assign addr[31744] = -276510565;
assign addr[31745] = -257536251;
assign addr[31746] = -238541516;
assign addr[31747] = -219527866;
assign addr[31748] = -200496809;
assign addr[31749] = -181449854;
assign addr[31750] = -162388511;
assign addr[31751] = -143314291;
assign addr[31752] = -124228708;
assign addr[31753] = -105133274;
assign addr[31754] = -86029503;
assign addr[31755] = -66918911;
assign addr[31756] = -47803013;
assign addr[31757] = -28683324;
assign addr[31758] = -9561361;
assign addr[31759] = 9561361;
assign addr[31760] = 28683324;
assign addr[31761] = 47803013;
assign addr[31762] = 66918911;
assign addr[31763] = 86029503;
assign addr[31764] = 105133274;
assign addr[31765] = 124228708;
assign addr[31766] = 143314291;
assign addr[31767] = 162388511;
assign addr[31768] = 181449854;
assign addr[31769] = 200496809;
assign addr[31770] = 219527866;
assign addr[31771] = 238541516;
assign addr[31772] = 257536251;
assign addr[31773] = 276510565;
assign addr[31774] = 295462954;
assign addr[31775] = 314391913;
assign addr[31776] = 333295944;
assign addr[31777] = 352173546;
assign addr[31778] = 371023223;
assign addr[31779] = 389843480;
assign addr[31780] = 408632825;
assign addr[31781] = 427389768;
assign addr[31782] = 446112822;
assign addr[31783] = 464800501;
assign addr[31784] = 483451325;
assign addr[31785] = 502063814;
assign addr[31786] = 520636492;
assign addr[31787] = 539167887;
assign addr[31788] = 557656529;
assign addr[31789] = 576100953;
assign addr[31790] = 594499695;
assign addr[31791] = 612851297;
assign addr[31792] = 631154304;
assign addr[31793] = 649407264;
assign addr[31794] = 667608730;
assign addr[31795] = 685757258;
assign addr[31796] = 703851410;
assign addr[31797] = 721889752;
assign addr[31798] = 739870851;
assign addr[31799] = 757793284;
assign addr[31800] = 775655628;
assign addr[31801] = 793456467;
assign addr[31802] = 811194391;
assign addr[31803] = 828867991;
assign addr[31804] = 846475867;
assign addr[31805] = 864016623;
assign addr[31806] = 881488868;
assign addr[31807] = 898891215;
assign addr[31808] = 916222287;
assign addr[31809] = 933480707;
assign addr[31810] = 950665109;
assign addr[31811] = 967774128;
assign addr[31812] = 984806408;
assign addr[31813] = 1001760600;
assign addr[31814] = 1018635358;
assign addr[31815] = 1035429345;
assign addr[31816] = 1052141228;
assign addr[31817] = 1068769683;
assign addr[31818] = 1085313391;
assign addr[31819] = 1101771040;
assign addr[31820] = 1118141326;
assign addr[31821] = 1134422949;
assign addr[31822] = 1150614620;
assign addr[31823] = 1166715055;
assign addr[31824] = 1182722976;
assign addr[31825] = 1198637114;
assign addr[31826] = 1214456207;
assign addr[31827] = 1230179002;
assign addr[31828] = 1245804251;
assign addr[31829] = 1261330715;
assign addr[31830] = 1276757164;
assign addr[31831] = 1292082373;
assign addr[31832] = 1307305128;
assign addr[31833] = 1322424222;
assign addr[31834] = 1337438456;
assign addr[31835] = 1352346639;
assign addr[31836] = 1367147589;
assign addr[31837] = 1381840133;
assign addr[31838] = 1396423105;
assign addr[31839] = 1410895350;
assign addr[31840] = 1425255719;
assign addr[31841] = 1439503074;
assign addr[31842] = 1453636285;
assign addr[31843] = 1467654232;
assign addr[31844] = 1481555802;
assign addr[31845] = 1495339895;
assign addr[31846] = 1509005416;
assign addr[31847] = 1522551282;
assign addr[31848] = 1535976419;
assign addr[31849] = 1549279763;
assign addr[31850] = 1562460258;
assign addr[31851] = 1575516860;
assign addr[31852] = 1588448533;
assign addr[31853] = 1601254251;
assign addr[31854] = 1613933000;
assign addr[31855] = 1626483774;
assign addr[31856] = 1638905577;
assign addr[31857] = 1651197426;
assign addr[31858] = 1663358344;
assign addr[31859] = 1675387369;
assign addr[31860] = 1687283545;
assign addr[31861] = 1699045930;
assign addr[31862] = 1710673591;
assign addr[31863] = 1722165606;
assign addr[31864] = 1733521064;
assign addr[31865] = 1744739065;
assign addr[31866] = 1755818718;
assign addr[31867] = 1766759146;
assign addr[31868] = 1777559480;
assign addr[31869] = 1788218865;
assign addr[31870] = 1798736454;
assign addr[31871] = 1809111415;
assign addr[31872] = 1819342925;
assign addr[31873] = 1829430172;
assign addr[31874] = 1839372356;
assign addr[31875] = 1849168689;
assign addr[31876] = 1858818395;
assign addr[31877] = 1868320707;
assign addr[31878] = 1877674873;
assign addr[31879] = 1886880151;
assign addr[31880] = 1895935811;
assign addr[31881] = 1904841135;
assign addr[31882] = 1913595416;
assign addr[31883] = 1922197961;
assign addr[31884] = 1930648088;
assign addr[31885] = 1938945125;
assign addr[31886] = 1947088417;
assign addr[31887] = 1955077316;
assign addr[31888] = 1962911189;
assign addr[31889] = 1970589416;
assign addr[31890] = 1978111387;
assign addr[31891] = 1985476506;
assign addr[31892] = 1992684188;
assign addr[31893] = 1999733863;
assign addr[31894] = 2006624971;
assign addr[31895] = 2013356967;
assign addr[31896] = 2019929315;
assign addr[31897] = 2026341495;
assign addr[31898] = 2032592999;
assign addr[31899] = 2038683330;
assign addr[31900] = 2044612007;
assign addr[31901] = 2050378558;
assign addr[31902] = 2055982526;
assign addr[31903] = 2061423468;
assign addr[31904] = 2066700952;
assign addr[31905] = 2071814558;
assign addr[31906] = 2076763883;
assign addr[31907] = 2081548533;
assign addr[31908] = 2086168128;
assign addr[31909] = 2090622304;
assign addr[31910] = 2094910706;
assign addr[31911] = 2099032994;
assign addr[31912] = 2102988841;
assign addr[31913] = 2106777935;
assign addr[31914] = 2110399974;
assign addr[31915] = 2113854671;
assign addr[31916] = 2117141752;
assign addr[31917] = 2120260957;
assign addr[31918] = 2123212038;
assign addr[31919] = 2125994762;
assign addr[31920] = 2128608907;
assign addr[31921] = 2131054266;
assign addr[31922] = 2133330646;
assign addr[31923] = 2135437865;
assign addr[31924] = 2137375758;
assign addr[31925] = 2139144169;
assign addr[31926] = 2140742960;
assign addr[31927] = 2142172003;
assign addr[31928] = 2143431184;
assign addr[31929] = 2144520405;
assign addr[31930] = 2145439578;
assign addr[31931] = 2146188631;
assign addr[31932] = 2146767505;
assign addr[31933] = 2147176152;
assign addr[31934] = 2147414542;
assign addr[31935] = 2147482655;
assign addr[31936] = 2147380486;
assign addr[31937] = 2147108043;
assign addr[31938] = 2146665347;
assign addr[31939] = 2146052433;
assign addr[31940] = 2145269351;
assign addr[31941] = 2144316162;
assign addr[31942] = 2143192942;
assign addr[31943] = 2141899780;
assign addr[31944] = 2140436778;
assign addr[31945] = 2138804053;
assign addr[31946] = 2137001733;
assign addr[31947] = 2135029962;
assign addr[31948] = 2132888897;
assign addr[31949] = 2130578706;
assign addr[31950] = 2128099574;
assign addr[31951] = 2125451696;
assign addr[31952] = 2122635283;
assign addr[31953] = 2119650558;
assign addr[31954] = 2116497758;
assign addr[31955] = 2113177132;
assign addr[31956] = 2109688944;
assign addr[31957] = 2106033471;
assign addr[31958] = 2102211002;
assign addr[31959] = 2098221841;
assign addr[31960] = 2094066304;
assign addr[31961] = 2089744719;
assign addr[31962] = 2085257431;
assign addr[31963] = 2080604795;
assign addr[31964] = 2075787180;
assign addr[31965] = 2070804967;
assign addr[31966] = 2065658552;
assign addr[31967] = 2060348343;
assign addr[31968] = 2054874761;
assign addr[31969] = 2049238240;
assign addr[31970] = 2043439226;
assign addr[31971] = 2037478181;
assign addr[31972] = 2031355576;
assign addr[31973] = 2025071897;
assign addr[31974] = 2018627642;
assign addr[31975] = 2012023322;
assign addr[31976] = 2005259462;
assign addr[31977] = 1998336596;
assign addr[31978] = 1991255274;
assign addr[31979] = 1984016058;
assign addr[31980] = 1976619522;
assign addr[31981] = 1969066252;
assign addr[31982] = 1961356847;
assign addr[31983] = 1953491918;
assign addr[31984] = 1945472089;
assign addr[31985] = 1937297997;
assign addr[31986] = 1928970288;
assign addr[31987] = 1920489624;
assign addr[31988] = 1911856677;
assign addr[31989] = 1903072131;
assign addr[31990] = 1894136683;
assign addr[31991] = 1885051042;
assign addr[31992] = 1875815927;
assign addr[31993] = 1866432072;
assign addr[31994] = 1856900221;
assign addr[31995] = 1847221128;
assign addr[31996] = 1837395562;
assign addr[31997] = 1827424302;
assign addr[31998] = 1817308138;
assign addr[31999] = 1807047873;
assign addr[32000] = 1796644320;
assign addr[32001] = 1786098304;
assign addr[32002] = 1775410662;
assign addr[32003] = 1764582240;
assign addr[32004] = 1753613897;
assign addr[32005] = 1742506504;
assign addr[32006] = 1731260941;
assign addr[32007] = 1719878099;
assign addr[32008] = 1708358881;
assign addr[32009] = 1696704201;
assign addr[32010] = 1684914983;
assign addr[32011] = 1672992161;
assign addr[32012] = 1660936681;
assign addr[32013] = 1648749499;
assign addr[32014] = 1636431582;
assign addr[32015] = 1623983905;
assign addr[32016] = 1611407456;
assign addr[32017] = 1598703233;
assign addr[32018] = 1585872242;
assign addr[32019] = 1572915501;
assign addr[32020] = 1559834037;
assign addr[32021] = 1546628888;
assign addr[32022] = 1533301101;
assign addr[32023] = 1519851733;
assign addr[32024] = 1506281850;
assign addr[32025] = 1492592527;
assign addr[32026] = 1478784851;
assign addr[32027] = 1464859917;
assign addr[32028] = 1450818828;
assign addr[32029] = 1436662698;
assign addr[32030] = 1422392650;
assign addr[32031] = 1408009814;
assign addr[32032] = 1393515332;
assign addr[32033] = 1378910353;
assign addr[32034] = 1364196034;
assign addr[32035] = 1349373543;
assign addr[32036] = 1334444055;
assign addr[32037] = 1319408754;
assign addr[32038] = 1304268832;
assign addr[32039] = 1289025489;
assign addr[32040] = 1273679934;
assign addr[32041] = 1258233384;
assign addr[32042] = 1242687064;
assign addr[32043] = 1227042207;
assign addr[32044] = 1211300053;
assign addr[32045] = 1195461849;
assign addr[32046] = 1179528853;
assign addr[32047] = 1163502328;
assign addr[32048] = 1147383544;
assign addr[32049] = 1131173780;
assign addr[32050] = 1114874320;
assign addr[32051] = 1098486458;
assign addr[32052] = 1082011492;
assign addr[32053] = 1065450729;
assign addr[32054] = 1048805483;
assign addr[32055] = 1032077073;
assign addr[32056] = 1015266825;
assign addr[32057] = 998376073;
assign addr[32058] = 981406156;
assign addr[32059] = 964358420;
assign addr[32060] = 947234215;
assign addr[32061] = 930034901;
assign addr[32062] = 912761841;
assign addr[32063] = 895416404;
assign addr[32064] = 877999966;
assign addr[32065] = 860513908;
assign addr[32066] = 842959617;
assign addr[32067] = 825338484;
assign addr[32068] = 807651907;
assign addr[32069] = 789901288;
assign addr[32070] = 772088034;
assign addr[32071] = 754213559;
assign addr[32072] = 736279279;
assign addr[32073] = 718286617;
assign addr[32074] = 700236999;
assign addr[32075] = 682131857;
assign addr[32076] = 663972625;
assign addr[32077] = 645760745;
assign addr[32078] = 627497660;
assign addr[32079] = 609184818;
assign addr[32080] = 590823671;
assign addr[32081] = 572415676;
assign addr[32082] = 553962291;
assign addr[32083] = 535464981;
assign addr[32084] = 516925212;
assign addr[32085] = 498344454;
assign addr[32086] = 479724180;
assign addr[32087] = 461065866;
assign addr[32088] = 442370993;
assign addr[32089] = 423641043;
assign addr[32090] = 404877501;
assign addr[32091] = 386081854;
assign addr[32092] = 367255594;
assign addr[32093] = 348400212;
assign addr[32094] = 329517204;
assign addr[32095] = 310608068;
assign addr[32096] = 291674302;
assign addr[32097] = 272717408;
assign addr[32098] = 253738890;
assign addr[32099] = 234740251;
assign addr[32100] = 215722999;
assign addr[32101] = 196688642;
assign addr[32102] = 177638688;
assign addr[32103] = 158574649;
assign addr[32104] = 139498035;
assign addr[32105] = 120410361;
assign addr[32106] = 101313138;
assign addr[32107] = 82207882;
assign addr[32108] = 63096108;
assign addr[32109] = 43979330;
assign addr[32110] = 24859065;
assign addr[32111] = 5736829;
assign addr[32112] = -13385863;
assign addr[32113] = -32507492;
assign addr[32114] = -51626544;
assign addr[32115] = -70741503;
assign addr[32116] = -89850852;
assign addr[32117] = -108953076;
assign addr[32118] = -128046661;
assign addr[32119] = -147130093;
assign addr[32120] = -166201858;
assign addr[32121] = -185260444;
assign addr[32122] = -204304341;
assign addr[32123] = -223332037;
assign addr[32124] = -242342025;
assign addr[32125] = -261332796;
assign addr[32126] = -280302845;
assign addr[32127] = -299250668;
assign addr[32128] = -318174762;
assign addr[32129] = -337073627;
assign addr[32130] = -355945764;
assign addr[32131] = -374789676;
assign addr[32132] = -393603870;
assign addr[32133] = -412386854;
assign addr[32134] = -431137138;
assign addr[32135] = -449853235;
assign addr[32136] = -468533662;
assign addr[32137] = -487176937;
assign addr[32138] = -505781581;
assign addr[32139] = -524346121;
assign addr[32140] = -542869083;
assign addr[32141] = -561348998;
assign addr[32142] = -579784402;
assign addr[32143] = -598173833;
assign addr[32144] = -616515832;
assign addr[32145] = -634808946;
assign addr[32146] = -653051723;
assign addr[32147] = -671242716;
assign addr[32148] = -689380485;
assign addr[32149] = -707463589;
assign addr[32150] = -725490597;
assign addr[32151] = -743460077;
assign addr[32152] = -761370605;
assign addr[32153] = -779220762;
assign addr[32154] = -797009130;
assign addr[32155] = -814734301;
assign addr[32156] = -832394869;
assign addr[32157] = -849989433;
assign addr[32158] = -867516597;
assign addr[32159] = -884974973;
assign addr[32160] = -902363176;
assign addr[32161] = -919679827;
assign addr[32162] = -936923553;
assign addr[32163] = -954092986;
assign addr[32164] = -971186766;
assign addr[32165] = -988203537;
assign addr[32166] = -1005141949;
assign addr[32167] = -1022000660;
assign addr[32168] = -1038778332;
assign addr[32169] = -1055473635;
assign addr[32170] = -1072085246;
assign addr[32171] = -1088611847;
assign addr[32172] = -1105052128;
assign addr[32173] = -1121404785;
assign addr[32174] = -1137668521;
assign addr[32175] = -1153842047;
assign addr[32176] = -1169924081;
assign addr[32177] = -1185913346;
assign addr[32178] = -1201808576;
assign addr[32179] = -1217608510;
assign addr[32180] = -1233311895;
assign addr[32181] = -1248917486;
assign addr[32182] = -1264424045;
assign addr[32183] = -1279830344;
assign addr[32184] = -1295135159;
assign addr[32185] = -1310337279;
assign addr[32186] = -1325435496;
assign addr[32187] = -1340428615;
assign addr[32188] = -1355315445;
assign addr[32189] = -1370094808;
assign addr[32190] = -1384765530;
assign addr[32191] = -1399326449;
assign addr[32192] = -1413776410;
assign addr[32193] = -1428114267;
assign addr[32194] = -1442338884;
assign addr[32195] = -1456449131;
assign addr[32196] = -1470443891;
assign addr[32197] = -1484322054;
assign addr[32198] = -1498082520;
assign addr[32199] = -1511724196;
assign addr[32200] = -1525246002;
assign addr[32201] = -1538646865;
assign addr[32202] = -1551925723;
assign addr[32203] = -1565081523;
assign addr[32204] = -1578113222;
assign addr[32205] = -1591019785;
assign addr[32206] = -1603800191;
assign addr[32207] = -1616453425;
assign addr[32208] = -1628978484;
assign addr[32209] = -1641374375;
assign addr[32210] = -1653640115;
assign addr[32211] = -1665774731;
assign addr[32212] = -1677777262;
assign addr[32213] = -1689646755;
assign addr[32214] = -1701382270;
assign addr[32215] = -1712982875;
assign addr[32216] = -1724447652;
assign addr[32217] = -1735775690;
assign addr[32218] = -1746966091;
assign addr[32219] = -1758017969;
assign addr[32220] = -1768930447;
assign addr[32221] = -1779702660;
assign addr[32222] = -1790333753;
assign addr[32223] = -1800822883;
assign addr[32224] = -1811169220;
assign addr[32225] = -1821371941;
assign addr[32226] = -1831430239;
assign addr[32227] = -1841343316;
assign addr[32228] = -1851110385;
assign addr[32229] = -1860730673;
assign addr[32230] = -1870203416;
assign addr[32231] = -1879527863;
assign addr[32232] = -1888703276;
assign addr[32233] = -1897728925;
assign addr[32234] = -1906604097;
assign addr[32235] = -1915328086;
assign addr[32236] = -1923900201;
assign addr[32237] = -1932319763;
assign addr[32238] = -1940586104;
assign addr[32239] = -1948698568;
assign addr[32240] = -1956656513;
assign addr[32241] = -1964459306;
assign addr[32242] = -1972106330;
assign addr[32243] = -1979596978;
assign addr[32244] = -1986930656;
assign addr[32245] = -1994106782;
assign addr[32246] = -2001124788;
assign addr[32247] = -2007984117;
assign addr[32248] = -2014684225;
assign addr[32249] = -2021224581;
assign addr[32250] = -2027604666;
assign addr[32251] = -2033823974;
assign addr[32252] = -2039882013;
assign addr[32253] = -2045778302;
assign addr[32254] = -2051512372;
assign addr[32255] = -2057083771;
assign addr[32256] = -2062492055;
assign addr[32257] = -2067736796;
assign addr[32258] = -2072817579;
assign addr[32259] = -2077733999;
assign addr[32260] = -2082485668;
assign addr[32261] = -2087072209;
assign addr[32262] = -2091493257;
assign addr[32263] = -2095748463;
assign addr[32264] = -2099837489;
assign addr[32265] = -2103760010;
assign addr[32266] = -2107515716;
assign addr[32267] = -2111104309;
assign addr[32268] = -2114525505;
assign addr[32269] = -2117779031;
assign addr[32270] = -2120864631;
assign addr[32271] = -2123782059;
assign addr[32272] = -2126531084;
assign addr[32273] = -2129111488;
assign addr[32274] = -2131523066;
assign addr[32275] = -2133765628;
assign addr[32276] = -2135838995;
assign addr[32277] = -2137743003;
assign addr[32278] = -2139477502;
assign addr[32279] = -2141042352;
assign addr[32280] = -2142437431;
assign addr[32281] = -2143662628;
assign addr[32282] = -2144717846;
assign addr[32283] = -2145603001;
assign addr[32284] = -2146318022;
assign addr[32285] = -2146862854;
assign addr[32286] = -2147237452;
assign addr[32287] = -2147441787;
assign addr[32288] = -2147475844;
assign addr[32289] = -2147339619;
assign addr[32290] = -2147033123;
assign addr[32291] = -2146556380;
assign addr[32292] = -2145909429;
assign addr[32293] = -2145092320;
assign addr[32294] = -2144105118;
assign addr[32295] = -2142947902;
assign addr[32296] = -2141620763;
assign addr[32297] = -2140123807;
assign addr[32298] = -2138457152;
assign addr[32299] = -2136620930;
assign addr[32300] = -2134615288;
assign addr[32301] = -2132440383;
assign addr[32302] = -2130096389;
assign addr[32303] = -2127583492;
assign addr[32304] = -2124901890;
assign addr[32305] = -2122051796;
assign addr[32306] = -2119033436;
assign addr[32307] = -2115847050;
assign addr[32308] = -2112492891;
assign addr[32309] = -2108971223;
assign addr[32310] = -2105282327;
assign addr[32311] = -2101426496;
assign addr[32312] = -2097404033;
assign addr[32313] = -2093215260;
assign addr[32314] = -2088860507;
assign addr[32315] = -2084340120;
assign addr[32316] = -2079654458;
assign addr[32317] = -2074803892;
assign addr[32318] = -2069788807;
assign addr[32319] = -2064609600;
assign addr[32320] = -2059266683;
assign addr[32321] = -2053760478;
assign addr[32322] = -2048091422;
assign addr[32323] = -2042259965;
assign addr[32324] = -2036266570;
assign addr[32325] = -2030111710;
assign addr[32326] = -2023795876;
assign addr[32327] = -2017319567;
assign addr[32328] = -2010683297;
assign addr[32329] = -2003887591;
assign addr[32330] = -1996932990;
assign addr[32331] = -1989820044;
assign addr[32332] = -1982549318;
assign addr[32333] = -1975121388;
assign addr[32334] = -1967536842;
assign addr[32335] = -1959796283;
assign addr[32336] = -1951900324;
assign addr[32337] = -1943849591;
assign addr[32338] = -1935644723;
assign addr[32339] = -1927286370;
assign addr[32340] = -1918775195;
assign addr[32341] = -1910111873;
assign addr[32342] = -1901297091;
assign addr[32343] = -1892331547;
assign addr[32344] = -1883215953;
assign addr[32345] = -1873951032;
assign addr[32346] = -1864537518;
assign addr[32347] = -1854976157;
assign addr[32348] = -1845267708;
assign addr[32349] = -1835412941;
assign addr[32350] = -1825412636;
assign addr[32351] = -1815267588;
assign addr[32352] = -1804978599;
assign addr[32353] = -1794546487;
assign addr[32354] = -1783972079;
assign addr[32355] = -1773256212;
assign addr[32356] = -1762399737;
assign addr[32357] = -1751403515;
assign addr[32358] = -1740268417;
assign addr[32359] = -1728995326;
assign addr[32360] = -1717585136;
assign addr[32361] = -1706038753;
assign addr[32362] = -1694357091;
assign addr[32363] = -1682541077;
assign addr[32364] = -1670591647;
assign addr[32365] = -1658509750;
assign addr[32366] = -1646296344;
assign addr[32367] = -1633952396;
assign addr[32368] = -1621478885;
assign addr[32369] = -1608876801;
assign addr[32370] = -1596147143;
assign addr[32371] = -1583290921;
assign addr[32372] = -1570309153;
assign addr[32373] = -1557202869;
assign addr[32374] = -1543973108;
assign addr[32375] = -1530620920;
assign addr[32376] = -1517147363;
assign addr[32377] = -1503553506;
assign addr[32378] = -1489840425;
assign addr[32379] = -1476009210;
assign addr[32380] = -1462060956;
assign addr[32381] = -1447996770;
assign addr[32382] = -1433817766;
assign addr[32383] = -1419525069;
assign addr[32384] = -1405119813;
assign addr[32385] = -1390603139;
assign addr[32386] = -1375976199;
assign addr[32387] = -1361240152;
assign addr[32388] = -1346396168;
assign addr[32389] = -1331445422;
assign addr[32390] = -1316389101;
assign addr[32391] = -1301228398;
assign addr[32392] = -1285964516;
assign addr[32393] = -1270598665;
assign addr[32394] = -1255132063;
assign addr[32395] = -1239565936;
assign addr[32396] = -1223901520;
assign addr[32397] = -1208140056;
assign addr[32398] = -1192282793;
assign addr[32399] = -1176330990;
assign addr[32400] = -1160285911;
assign addr[32401] = -1144148829;
assign addr[32402] = -1127921022;
assign addr[32403] = -1111603778;
assign addr[32404] = -1095198391;
assign addr[32405] = -1078706161;
assign addr[32406] = -1062128397;
assign addr[32407] = -1045466412;
assign addr[32408] = -1028721528;
assign addr[32409] = -1011895073;
assign addr[32410] = -994988380;
assign addr[32411] = -978002791;
assign addr[32412] = -960939653;
assign addr[32413] = -943800318;
assign addr[32414] = -926586145;
assign addr[32415] = -909298500;
assign addr[32416] = -891938752;
assign addr[32417] = -874508280;
assign addr[32418] = -857008464;
assign addr[32419] = -839440693;
assign addr[32420] = -821806359;
assign addr[32421] = -804106861;
assign addr[32422] = -786343603;
assign addr[32423] = -768517992;
assign addr[32424] = -750631442;
assign addr[32425] = -732685372;
assign addr[32426] = -714681204;
assign addr[32427] = -696620367;
assign addr[32428] = -678504291;
assign addr[32429] = -660334415;
assign addr[32430] = -642112178;
assign addr[32431] = -623839025;
assign addr[32432] = -605516406;
assign addr[32433] = -587145773;
assign addr[32434] = -568728583;
assign addr[32435] = -550266296;
assign addr[32436] = -531760377;
assign addr[32437] = -513212292;
assign addr[32438] = -494623513;
assign addr[32439] = -475995513;
assign addr[32440] = -457329769;
assign addr[32441] = -438627762;
assign addr[32442] = -419890975;
assign addr[32443] = -401120892;
assign addr[32444] = -382319004;
assign addr[32445] = -363486799;
assign addr[32446] = -344625773;
assign addr[32447] = -325737419;
assign addr[32448] = -306823237;
assign addr[32449] = -287884725;
assign addr[32450] = -268923386;
assign addr[32451] = -249940723;
assign addr[32452] = -230938242;
assign addr[32453] = -211917448;
assign addr[32454] = -192879850;
assign addr[32455] = -173826959;
assign addr[32456] = -154760284;
assign addr[32457] = -135681337;
assign addr[32458] = -116591632;
assign addr[32459] = -97492681;
assign addr[32460] = -78386000;
assign addr[32461] = -59273104;
assign addr[32462] = -40155507;
assign addr[32463] = -21034727;
assign addr[32464] = -1912278;
assign addr[32465] = 17210322;
assign addr[32466] = 36331557;
assign addr[32467] = 55449912;
assign addr[32468] = 74563870;
assign addr[32469] = 93671915;
assign addr[32470] = 112772533;
assign addr[32471] = 131864208;
assign addr[32472] = 150945428;
assign addr[32473] = 170014678;
assign addr[32474] = 189070447;
assign addr[32475] = 208111224;
assign addr[32476] = 227135500;
assign addr[32477] = 246141764;
assign addr[32478] = 265128512;
assign addr[32479] = 284094236;
assign addr[32480] = 303037433;
assign addr[32481] = 321956601;
assign addr[32482] = 340850240;
assign addr[32483] = 359716852;
assign addr[32484] = 378554940;
assign addr[32485] = 397363011;
assign addr[32486] = 416139574;
assign addr[32487] = 434883140;
assign addr[32488] = 453592221;
assign addr[32489] = 472265336;
assign addr[32490] = 490901003;
assign addr[32491] = 509497745;
assign addr[32492] = 528054086;
assign addr[32493] = 546568556;
assign addr[32494] = 565039687;
assign addr[32495] = 583466013;
assign addr[32496] = 601846074;
assign addr[32497] = 620178412;
assign addr[32498] = 638461574;
assign addr[32499] = 656694110;
assign addr[32500] = 674874574;
assign addr[32501] = 693001525;
assign addr[32502] = 711073524;
assign addr[32503] = 729089140;
assign addr[32504] = 747046944;
assign addr[32505] = 764945512;
assign addr[32506] = 782783424;
assign addr[32507] = 800559266;
assign addr[32508] = 818271628;
assign addr[32509] = 835919107;
assign addr[32510] = 853500302;
assign addr[32511] = 871013820;
assign addr[32512] = 888458272;
assign addr[32513] = 905832274;
assign addr[32514] = 923134450;
assign addr[32515] = 940363427;
assign addr[32516] = 957517838;
assign addr[32517] = 974596324;
assign addr[32518] = 991597531;
assign addr[32519] = 1008520110;
assign addr[32520] = 1025362720;
assign addr[32521] = 1042124025;
assign addr[32522] = 1058802695;
assign addr[32523] = 1075397409;
assign addr[32524] = 1091906851;
assign addr[32525] = 1108329711;
assign addr[32526] = 1124664687;
assign addr[32527] = 1140910484;
assign addr[32528] = 1157065814;
assign addr[32529] = 1173129396;
assign addr[32530] = 1189099956;
assign addr[32531] = 1204976227;
assign addr[32532] = 1220756951;
assign addr[32533] = 1236440877;
assign addr[32534] = 1252026760;
assign addr[32535] = 1267513365;
assign addr[32536] = 1282899464;
assign addr[32537] = 1298183838;
assign addr[32538] = 1313365273;
assign addr[32539] = 1328442566;
assign addr[32540] = 1343414522;
assign addr[32541] = 1358279953;
assign addr[32542] = 1373037681;
assign addr[32543] = 1387686535;
assign addr[32544] = 1402225355;
assign addr[32545] = 1416652986;
assign addr[32546] = 1430968286;
assign addr[32547] = 1445170118;
assign addr[32548] = 1459257358;
assign addr[32549] = 1473228887;
assign addr[32550] = 1487083598;
assign addr[32551] = 1500820393;
assign addr[32552] = 1514438181;
assign addr[32553] = 1527935884;
assign addr[32554] = 1541312431;
assign addr[32555] = 1554566762;
assign addr[32556] = 1567697824;
assign addr[32557] = 1580704578;
assign addr[32558] = 1593585992;
assign addr[32559] = 1606341043;
assign addr[32560] = 1618968722;
assign addr[32561] = 1631468027;
assign addr[32562] = 1643837966;
assign addr[32563] = 1656077559;
assign addr[32564] = 1668185835;
assign addr[32565] = 1680161834;
assign addr[32566] = 1692004606;
assign addr[32567] = 1703713213;
assign addr[32568] = 1715286726;
assign addr[32569] = 1726724227;
assign addr[32570] = 1738024810;
assign addr[32571] = 1749187577;
assign addr[32572] = 1760211645;
assign addr[32573] = 1771096139;
assign addr[32574] = 1781840195;
assign addr[32575] = 1792442963;
assign addr[32576] = 1802903601;
assign addr[32577] = 1813221279;
assign addr[32578] = 1823395180;
assign addr[32579] = 1833424497;
assign addr[32580] = 1843308435;
assign addr[32581] = 1853046210;
assign addr[32582] = 1862637049;
assign addr[32583] = 1872080193;
assign addr[32584] = 1881374892;
assign addr[32585] = 1890520410;
assign addr[32586] = 1899516021;
assign addr[32587] = 1908361011;
assign addr[32588] = 1917054681;
assign addr[32589] = 1925596340;
assign addr[32590] = 1933985310;
assign addr[32591] = 1942220928;
assign addr[32592] = 1950302539;
assign addr[32593] = 1958229503;
assign addr[32594] = 1966001192;
assign addr[32595] = 1973616989;
assign addr[32596] = 1981076290;
assign addr[32597] = 1988378503;
assign addr[32598] = 1995523051;
assign addr[32599] = 2002509365;
assign addr[32600] = 2009336893;
assign addr[32601] = 2016005093;
assign addr[32602] = 2022513436;
assign addr[32603] = 2028861406;
assign addr[32604] = 2035048499;
assign addr[32605] = 2041074226;
assign addr[32606] = 2046938108;
assign addr[32607] = 2052639680;
assign addr[32608] = 2058178491;
assign addr[32609] = 2063554100;
assign addr[32610] = 2068766083;
assign addr[32611] = 2073814024;
assign addr[32612] = 2078697525;
assign addr[32613] = 2083416198;
assign addr[32614] = 2087969669;
assign addr[32615] = 2092357577;
assign addr[32616] = 2096579573;
assign addr[32617] = 2100635323;
assign addr[32618] = 2104524506;
assign addr[32619] = 2108246813;
assign addr[32620] = 2111801949;
assign addr[32621] = 2115189632;
assign addr[32622] = 2118409593;
assign addr[32623] = 2121461578;
assign addr[32624] = 2124345343;
assign addr[32625] = 2127060661;
assign addr[32626] = 2129607316;
assign addr[32627] = 2131985106;
assign addr[32628] = 2134193842;
assign addr[32629] = 2136233350;
assign addr[32630] = 2138103468;
assign addr[32631] = 2139804048;
assign addr[32632] = 2141334954;
assign addr[32633] = 2142696065;
assign addr[32634] = 2143887273;
assign addr[32635] = 2144908484;
assign addr[32636] = 2145759618;
assign addr[32637] = 2146440605;
assign addr[32638] = 2146951393;
assign addr[32639] = 2147291941;
assign addr[32640] = 2147462221;
assign addr[32641] = 2147462221;
assign addr[32642] = 2147291941;
assign addr[32643] = 2146951393;
assign addr[32644] = 2146440605;
assign addr[32645] = 2145759618;
assign addr[32646] = 2144908484;
assign addr[32647] = 2143887273;
assign addr[32648] = 2142696065;
assign addr[32649] = 2141334954;
assign addr[32650] = 2139804048;
assign addr[32651] = 2138103468;
assign addr[32652] = 2136233350;
assign addr[32653] = 2134193842;
assign addr[32654] = 2131985106;
assign addr[32655] = 2129607316;
assign addr[32656] = 2127060661;
assign addr[32657] = 2124345343;
assign addr[32658] = 2121461578;
assign addr[32659] = 2118409593;
assign addr[32660] = 2115189632;
assign addr[32661] = 2111801949;
assign addr[32662] = 2108246813;
assign addr[32663] = 2104524506;
assign addr[32664] = 2100635323;
assign addr[32665] = 2096579573;
assign addr[32666] = 2092357577;
assign addr[32667] = 2087969669;
assign addr[32668] = 2083416198;
assign addr[32669] = 2078697525;
assign addr[32670] = 2073814024;
assign addr[32671] = 2068766083;
assign addr[32672] = 2063554100;
assign addr[32673] = 2058178491;
assign addr[32674] = 2052639680;
assign addr[32675] = 2046938108;
assign addr[32676] = 2041074226;
assign addr[32677] = 2035048499;
assign addr[32678] = 2028861406;
assign addr[32679] = 2022513436;
assign addr[32680] = 2016005093;
assign addr[32681] = 2009336893;
assign addr[32682] = 2002509365;
assign addr[32683] = 1995523051;
assign addr[32684] = 1988378503;
assign addr[32685] = 1981076290;
assign addr[32686] = 1973616989;
assign addr[32687] = 1966001192;
assign addr[32688] = 1958229503;
assign addr[32689] = 1950302539;
assign addr[32690] = 1942220928;
assign addr[32691] = 1933985310;
assign addr[32692] = 1925596340;
assign addr[32693] = 1917054681;
assign addr[32694] = 1908361011;
assign addr[32695] = 1899516021;
assign addr[32696] = 1890520410;
assign addr[32697] = 1881374892;
assign addr[32698] = 1872080193;
assign addr[32699] = 1862637049;
assign addr[32700] = 1853046210;
assign addr[32701] = 1843308435;
assign addr[32702] = 1833424497;
assign addr[32703] = 1823395180;
assign addr[32704] = 1813221279;
assign addr[32705] = 1802903601;
assign addr[32706] = 1792442963;
assign addr[32707] = 1781840195;
assign addr[32708] = 1771096139;
assign addr[32709] = 1760211645;
assign addr[32710] = 1749187577;
assign addr[32711] = 1738024810;
assign addr[32712] = 1726724227;
assign addr[32713] = 1715286726;
assign addr[32714] = 1703713213;
assign addr[32715] = 1692004606;
assign addr[32716] = 1680161834;
assign addr[32717] = 1668185835;
assign addr[32718] = 1656077559;
assign addr[32719] = 1643837966;
assign addr[32720] = 1631468027;
assign addr[32721] = 1618968722;
assign addr[32722] = 1606341043;
assign addr[32723] = 1593585992;
assign addr[32724] = 1580704578;
assign addr[32725] = 1567697824;
assign addr[32726] = 1554566762;
assign addr[32727] = 1541312431;
assign addr[32728] = 1527935884;
assign addr[32729] = 1514438181;
assign addr[32730] = 1500820393;
assign addr[32731] = 1487083598;
assign addr[32732] = 1473228887;
assign addr[32733] = 1459257358;
assign addr[32734] = 1445170118;
assign addr[32735] = 1430968286;
assign addr[32736] = 1416652986;
assign addr[32737] = 1402225355;
assign addr[32738] = 1387686535;
assign addr[32739] = 1373037681;
assign addr[32740] = 1358279953;
assign addr[32741] = 1343414522;
assign addr[32742] = 1328442566;
assign addr[32743] = 1313365273;
assign addr[32744] = 1298183838;
assign addr[32745] = 1282899464;
assign addr[32746] = 1267513365;
assign addr[32747] = 1252026760;
assign addr[32748] = 1236440877;
assign addr[32749] = 1220756951;
assign addr[32750] = 1204976227;
assign addr[32751] = 1189099956;
assign addr[32752] = 1173129396;
assign addr[32753] = 1157065814;
assign addr[32754] = 1140910484;
assign addr[32755] = 1124664687;
assign addr[32756] = 1108329711;
assign addr[32757] = 1091906851;
assign addr[32758] = 1075397409;
assign addr[32759] = 1058802695;
assign addr[32760] = 1042124025;
assign addr[32761] = 1025362720;
assign addr[32762] = 1008520110;
assign addr[32763] = 991597531;
assign addr[32764] = 974596324;
assign addr[32765] = 957517838;
assign addr[32766] = 940363427;
assign addr[32767] = 923134450;
assign addr[32768] = 905832274;
assign addr[32769] = 888458272;
assign addr[32770] = 871013820;
assign addr[32771] = 853500302;
assign addr[32772] = 835919107;
assign addr[32773] = 818271628;
assign addr[32774] = 800559266;
assign addr[32775] = 782783424;
assign addr[32776] = 764945512;
assign addr[32777] = 747046944;
assign addr[32778] = 729089140;
assign addr[32779] = 711073524;
assign addr[32780] = 693001525;
assign addr[32781] = 674874574;
assign addr[32782] = 656694110;
assign addr[32783] = 638461574;
assign addr[32784] = 620178412;
assign addr[32785] = 601846074;
assign addr[32786] = 583466013;
assign addr[32787] = 565039687;
assign addr[32788] = 546568556;
assign addr[32789] = 528054086;
assign addr[32790] = 509497745;
assign addr[32791] = 490901003;
assign addr[32792] = 472265336;
assign addr[32793] = 453592221;
assign addr[32794] = 434883140;
assign addr[32795] = 416139574;
assign addr[32796] = 397363011;
assign addr[32797] = 378554940;
assign addr[32798] = 359716852;
assign addr[32799] = 340850240;
assign addr[32800] = 321956601;
assign addr[32801] = 303037433;
assign addr[32802] = 284094236;
assign addr[32803] = 265128512;
assign addr[32804] = 246141764;
assign addr[32805] = 227135500;
assign addr[32806] = 208111224;
assign addr[32807] = 189070447;
assign addr[32808] = 170014678;
assign addr[32809] = 150945428;
assign addr[32810] = 131864208;
assign addr[32811] = 112772533;
assign addr[32812] = 93671915;
assign addr[32813] = 74563870;
assign addr[32814] = 55449912;
assign addr[32815] = 36331557;
assign addr[32816] = 17210322;
assign addr[32817] = -1912278;
assign addr[32818] = -21034727;
assign addr[32819] = -40155507;
assign addr[32820] = -59273104;
assign addr[32821] = -78386000;
assign addr[32822] = -97492681;
assign addr[32823] = -116591632;
assign addr[32824] = -135681337;
assign addr[32825] = -154760284;
assign addr[32826] = -173826959;
assign addr[32827] = -192879850;
assign addr[32828] = -211917448;
assign addr[32829] = -230938242;
assign addr[32830] = -249940723;
assign addr[32831] = -268923386;
assign addr[32832] = -287884725;
assign addr[32833] = -306823237;
assign addr[32834] = -325737419;
assign addr[32835] = -344625773;
assign addr[32836] = -363486799;
assign addr[32837] = -382319004;
assign addr[32838] = -401120892;
assign addr[32839] = -419890975;
assign addr[32840] = -438627762;
assign addr[32841] = -457329769;
assign addr[32842] = -475995513;
assign addr[32843] = -494623513;
assign addr[32844] = -513212292;
assign addr[32845] = -531760377;
assign addr[32846] = -550266296;
assign addr[32847] = -568728583;
assign addr[32848] = -587145773;
assign addr[32849] = -605516406;
assign addr[32850] = -623839025;
assign addr[32851] = -642112178;
assign addr[32852] = -660334415;
assign addr[32853] = -678504291;
assign addr[32854] = -696620367;
assign addr[32855] = -714681204;
assign addr[32856] = -732685372;
assign addr[32857] = -750631442;
assign addr[32858] = -768517992;
assign addr[32859] = -786343603;
assign addr[32860] = -804106861;
assign addr[32861] = -821806359;
assign addr[32862] = -839440693;
assign addr[32863] = -857008464;
assign addr[32864] = -874508280;
assign addr[32865] = -891938752;
assign addr[32866] = -909298500;
assign addr[32867] = -926586145;
assign addr[32868] = -943800318;
assign addr[32869] = -960939653;
assign addr[32870] = -978002791;
assign addr[32871] = -994988380;
assign addr[32872] = -1011895073;
assign addr[32873] = -1028721528;
assign addr[32874] = -1045466412;
assign addr[32875] = -1062128397;
assign addr[32876] = -1078706161;
assign addr[32877] = -1095198391;
assign addr[32878] = -1111603778;
assign addr[32879] = -1127921022;
assign addr[32880] = -1144148829;
assign addr[32881] = -1160285911;
assign addr[32882] = -1176330990;
assign addr[32883] = -1192282793;
assign addr[32884] = -1208140056;
assign addr[32885] = -1223901520;
assign addr[32886] = -1239565936;
assign addr[32887] = -1255132063;
assign addr[32888] = -1270598665;
assign addr[32889] = -1285964516;
assign addr[32890] = -1301228398;
assign addr[32891] = -1316389101;
assign addr[32892] = -1331445422;
assign addr[32893] = -1346396168;
assign addr[32894] = -1361240152;
assign addr[32895] = -1375976199;
assign addr[32896] = -1390603139;
assign addr[32897] = -1405119813;
assign addr[32898] = -1419525069;
assign addr[32899] = -1433817766;
assign addr[32900] = -1447996770;
assign addr[32901] = -1462060956;
assign addr[32902] = -1476009210;
assign addr[32903] = -1489840425;
assign addr[32904] = -1503553506;
assign addr[32905] = -1517147363;
assign addr[32906] = -1530620920;
assign addr[32907] = -1543973108;
assign addr[32908] = -1557202869;
assign addr[32909] = -1570309153;
assign addr[32910] = -1583290921;
assign addr[32911] = -1596147143;
assign addr[32912] = -1608876801;
assign addr[32913] = -1621478885;
assign addr[32914] = -1633952396;
assign addr[32915] = -1646296344;
assign addr[32916] = -1658509750;
assign addr[32917] = -1670591647;
assign addr[32918] = -1682541077;
assign addr[32919] = -1694357091;
assign addr[32920] = -1706038753;
assign addr[32921] = -1717585136;
assign addr[32922] = -1728995326;
assign addr[32923] = -1740268417;
assign addr[32924] = -1751403515;
assign addr[32925] = -1762399737;
assign addr[32926] = -1773256212;
assign addr[32927] = -1783972079;
assign addr[32928] = -1794546487;
assign addr[32929] = -1804978599;
assign addr[32930] = -1815267588;
assign addr[32931] = -1825412636;
assign addr[32932] = -1835412941;
assign addr[32933] = -1845267708;
assign addr[32934] = -1854976157;
assign addr[32935] = -1864537518;
assign addr[32936] = -1873951032;
assign addr[32937] = -1883215953;
assign addr[32938] = -1892331547;
assign addr[32939] = -1901297091;
assign addr[32940] = -1910111873;
assign addr[32941] = -1918775195;
assign addr[32942] = -1927286370;
assign addr[32943] = -1935644723;
assign addr[32944] = -1943849591;
assign addr[32945] = -1951900324;
assign addr[32946] = -1959796283;
assign addr[32947] = -1967536842;
assign addr[32948] = -1975121388;
assign addr[32949] = -1982549318;
assign addr[32950] = -1989820044;
assign addr[32951] = -1996932990;
assign addr[32952] = -2003887591;
assign addr[32953] = -2010683297;
assign addr[32954] = -2017319567;
assign addr[32955] = -2023795876;
assign addr[32956] = -2030111710;
assign addr[32957] = -2036266570;
assign addr[32958] = -2042259965;
assign addr[32959] = -2048091422;
assign addr[32960] = -2053760478;
assign addr[32961] = -2059266683;
assign addr[32962] = -2064609600;
assign addr[32963] = -2069788807;
assign addr[32964] = -2074803892;
assign addr[32965] = -2079654458;
assign addr[32966] = -2084340120;
assign addr[32967] = -2088860507;
assign addr[32968] = -2093215260;
assign addr[32969] = -2097404033;
assign addr[32970] = -2101426496;
assign addr[32971] = -2105282327;
assign addr[32972] = -2108971223;
assign addr[32973] = -2112492891;
assign addr[32974] = -2115847050;
assign addr[32975] = -2119033436;
assign addr[32976] = -2122051796;
assign addr[32977] = -2124901890;
assign addr[32978] = -2127583492;
assign addr[32979] = -2130096389;
assign addr[32980] = -2132440383;
assign addr[32981] = -2134615288;
assign addr[32982] = -2136620930;
assign addr[32983] = -2138457152;
assign addr[32984] = -2140123807;
assign addr[32985] = -2141620763;
assign addr[32986] = -2142947902;
assign addr[32987] = -2144105118;
assign addr[32988] = -2145092320;
assign addr[32989] = -2145909429;
assign addr[32990] = -2146556380;
assign addr[32991] = -2147033123;
assign addr[32992] = -2147339619;
assign addr[32993] = -2147475844;
assign addr[32994] = -2147441787;
assign addr[32995] = -2147237452;
assign addr[32996] = -2146862854;
assign addr[32997] = -2146318022;
assign addr[32998] = -2145603001;
assign addr[32999] = -2144717846;
assign addr[33000] = -2143662628;
assign addr[33001] = -2142437431;
assign addr[33002] = -2141042352;
assign addr[33003] = -2139477502;
assign addr[33004] = -2137743003;
assign addr[33005] = -2135838995;
assign addr[33006] = -2133765628;
assign addr[33007] = -2131523066;
assign addr[33008] = -2129111488;
assign addr[33009] = -2126531084;
assign addr[33010] = -2123782059;
assign addr[33011] = -2120864631;
assign addr[33012] = -2117779031;
assign addr[33013] = -2114525505;
assign addr[33014] = -2111104309;
assign addr[33015] = -2107515716;
assign addr[33016] = -2103760010;
assign addr[33017] = -2099837489;
assign addr[33018] = -2095748463;
assign addr[33019] = -2091493257;
assign addr[33020] = -2087072209;
assign addr[33021] = -2082485668;
assign addr[33022] = -2077733999;
assign addr[33023] = -2072817579;
assign addr[33024] = -2067736796;
assign addr[33025] = -2062492055;
assign addr[33026] = -2057083771;
assign addr[33027] = -2051512372;
assign addr[33028] = -2045778302;
assign addr[33029] = -2039882013;
assign addr[33030] = -2033823974;
assign addr[33031] = -2027604666;
assign addr[33032] = -2021224581;
assign addr[33033] = -2014684225;
assign addr[33034] = -2007984117;
assign addr[33035] = -2001124788;
assign addr[33036] = -1994106782;
assign addr[33037] = -1986930656;
assign addr[33038] = -1979596978;
assign addr[33039] = -1972106330;
assign addr[33040] = -1964459306;
assign addr[33041] = -1956656513;
assign addr[33042] = -1948698568;
assign addr[33043] = -1940586104;
assign addr[33044] = -1932319763;
assign addr[33045] = -1923900201;
assign addr[33046] = -1915328086;
assign addr[33047] = -1906604097;
assign addr[33048] = -1897728925;
assign addr[33049] = -1888703276;
assign addr[33050] = -1879527863;
assign addr[33051] = -1870203416;
assign addr[33052] = -1860730673;
assign addr[33053] = -1851110385;
assign addr[33054] = -1841343316;
assign addr[33055] = -1831430239;
assign addr[33056] = -1821371941;
assign addr[33057] = -1811169220;
assign addr[33058] = -1800822883;
assign addr[33059] = -1790333753;
assign addr[33060] = -1779702660;
assign addr[33061] = -1768930447;
assign addr[33062] = -1758017969;
assign addr[33063] = -1746966091;
assign addr[33064] = -1735775690;
assign addr[33065] = -1724447652;
assign addr[33066] = -1712982875;
assign addr[33067] = -1701382270;
assign addr[33068] = -1689646755;
assign addr[33069] = -1677777262;
assign addr[33070] = -1665774731;
assign addr[33071] = -1653640115;
assign addr[33072] = -1641374375;
assign addr[33073] = -1628978484;
assign addr[33074] = -1616453425;
assign addr[33075] = -1603800191;
assign addr[33076] = -1591019785;
assign addr[33077] = -1578113222;
assign addr[33078] = -1565081523;
assign addr[33079] = -1551925723;
assign addr[33080] = -1538646865;
assign addr[33081] = -1525246002;
assign addr[33082] = -1511724196;
assign addr[33083] = -1498082520;
assign addr[33084] = -1484322054;
assign addr[33085] = -1470443891;
assign addr[33086] = -1456449131;
assign addr[33087] = -1442338884;
assign addr[33088] = -1428114267;
assign addr[33089] = -1413776410;
assign addr[33090] = -1399326449;
assign addr[33091] = -1384765530;
assign addr[33092] = -1370094808;
assign addr[33093] = -1355315445;
assign addr[33094] = -1340428615;
assign addr[33095] = -1325435496;
assign addr[33096] = -1310337279;
assign addr[33097] = -1295135159;
assign addr[33098] = -1279830344;
assign addr[33099] = -1264424045;
assign addr[33100] = -1248917486;
assign addr[33101] = -1233311895;
assign addr[33102] = -1217608510;
assign addr[33103] = -1201808576;
assign addr[33104] = -1185913346;
assign addr[33105] = -1169924081;
assign addr[33106] = -1153842047;
assign addr[33107] = -1137668521;
assign addr[33108] = -1121404785;
assign addr[33109] = -1105052128;
assign addr[33110] = -1088611847;
assign addr[33111] = -1072085246;
assign addr[33112] = -1055473635;
assign addr[33113] = -1038778332;
assign addr[33114] = -1022000660;
assign addr[33115] = -1005141949;
assign addr[33116] = -988203537;
assign addr[33117] = -971186766;
assign addr[33118] = -954092986;
assign addr[33119] = -936923553;
assign addr[33120] = -919679827;
assign addr[33121] = -902363176;
assign addr[33122] = -884974973;
assign addr[33123] = -867516597;
assign addr[33124] = -849989433;
assign addr[33125] = -832394869;
assign addr[33126] = -814734301;
assign addr[33127] = -797009130;
assign addr[33128] = -779220762;
assign addr[33129] = -761370605;
assign addr[33130] = -743460077;
assign addr[33131] = -725490597;
assign addr[33132] = -707463589;
assign addr[33133] = -689380485;
assign addr[33134] = -671242716;
assign addr[33135] = -653051723;
assign addr[33136] = -634808946;
assign addr[33137] = -616515832;
assign addr[33138] = -598173833;
assign addr[33139] = -579784402;
assign addr[33140] = -561348998;
assign addr[33141] = -542869083;
assign addr[33142] = -524346121;
assign addr[33143] = -505781581;
assign addr[33144] = -487176937;
assign addr[33145] = -468533662;
assign addr[33146] = -449853235;
assign addr[33147] = -431137138;
assign addr[33148] = -412386854;
assign addr[33149] = -393603870;
assign addr[33150] = -374789676;
assign addr[33151] = -355945764;
assign addr[33152] = -337073627;
assign addr[33153] = -318174762;
assign addr[33154] = -299250668;
assign addr[33155] = -280302845;
assign addr[33156] = -261332796;
assign addr[33157] = -242342025;
assign addr[33158] = -223332037;
assign addr[33159] = -204304341;
assign addr[33160] = -185260444;
assign addr[33161] = -166201858;
assign addr[33162] = -147130093;
assign addr[33163] = -128046661;
assign addr[33164] = -108953076;
assign addr[33165] = -89850852;
assign addr[33166] = -70741503;
assign addr[33167] = -51626544;
assign addr[33168] = -32507492;
assign addr[33169] = -13385863;
assign addr[33170] = 5736829;
assign addr[33171] = 24859065;
assign addr[33172] = 43979330;
assign addr[33173] = 63096108;
assign addr[33174] = 82207882;
assign addr[33175] = 101313138;
assign addr[33176] = 120410361;
assign addr[33177] = 139498035;
assign addr[33178] = 158574649;
assign addr[33179] = 177638688;
assign addr[33180] = 196688642;
assign addr[33181] = 215722999;
assign addr[33182] = 234740251;
assign addr[33183] = 253738890;
assign addr[33184] = 272717408;
assign addr[33185] = 291674302;
assign addr[33186] = 310608068;
assign addr[33187] = 329517204;
assign addr[33188] = 348400212;
assign addr[33189] = 367255594;
assign addr[33190] = 386081854;
assign addr[33191] = 404877501;
assign addr[33192] = 423641043;
assign addr[33193] = 442370993;
assign addr[33194] = 461065866;
assign addr[33195] = 479724180;
assign addr[33196] = 498344454;
assign addr[33197] = 516925212;
assign addr[33198] = 535464981;
assign addr[33199] = 553962291;
assign addr[33200] = 572415676;
assign addr[33201] = 590823671;
assign addr[33202] = 609184818;
assign addr[33203] = 627497660;
assign addr[33204] = 645760745;
assign addr[33205] = 663972625;
assign addr[33206] = 682131857;
assign addr[33207] = 700236999;
assign addr[33208] = 718286617;
assign addr[33209] = 736279279;
assign addr[33210] = 754213559;
assign addr[33211] = 772088034;
assign addr[33212] = 789901288;
assign addr[33213] = 807651907;
assign addr[33214] = 825338484;
assign addr[33215] = 842959617;
assign addr[33216] = 860513908;
assign addr[33217] = 877999966;
assign addr[33218] = 895416404;
assign addr[33219] = 912761841;
assign addr[33220] = 930034901;
assign addr[33221] = 947234215;
assign addr[33222] = 964358420;
assign addr[33223] = 981406156;
assign addr[33224] = 998376073;
assign addr[33225] = 1015266825;
assign addr[33226] = 1032077073;
assign addr[33227] = 1048805483;
assign addr[33228] = 1065450729;
assign addr[33229] = 1082011492;
assign addr[33230] = 1098486458;
assign addr[33231] = 1114874320;
assign addr[33232] = 1131173780;
assign addr[33233] = 1147383544;
assign addr[33234] = 1163502328;
assign addr[33235] = 1179528853;
assign addr[33236] = 1195461849;
assign addr[33237] = 1211300053;
assign addr[33238] = 1227042207;
assign addr[33239] = 1242687064;
assign addr[33240] = 1258233384;
assign addr[33241] = 1273679934;
assign addr[33242] = 1289025489;
assign addr[33243] = 1304268832;
assign addr[33244] = 1319408754;
assign addr[33245] = 1334444055;
assign addr[33246] = 1349373543;
assign addr[33247] = 1364196034;
assign addr[33248] = 1378910353;
assign addr[33249] = 1393515332;
assign addr[33250] = 1408009814;
assign addr[33251] = 1422392650;
assign addr[33252] = 1436662698;
assign addr[33253] = 1450818828;
assign addr[33254] = 1464859917;
assign addr[33255] = 1478784851;
assign addr[33256] = 1492592527;
assign addr[33257] = 1506281850;
assign addr[33258] = 1519851733;
assign addr[33259] = 1533301101;
assign addr[33260] = 1546628888;
assign addr[33261] = 1559834037;
assign addr[33262] = 1572915501;
assign addr[33263] = 1585872242;
assign addr[33264] = 1598703233;
assign addr[33265] = 1611407456;
assign addr[33266] = 1623983905;
assign addr[33267] = 1636431582;
assign addr[33268] = 1648749499;
assign addr[33269] = 1660936681;
assign addr[33270] = 1672992161;
assign addr[33271] = 1684914983;
assign addr[33272] = 1696704201;
assign addr[33273] = 1708358881;
assign addr[33274] = 1719878099;
assign addr[33275] = 1731260941;
assign addr[33276] = 1742506504;
assign addr[33277] = 1753613897;
assign addr[33278] = 1764582240;
assign addr[33279] = 1775410662;
assign addr[33280] = 1786098304;
assign addr[33281] = 1796644320;
assign addr[33282] = 1807047873;
assign addr[33283] = 1817308138;
assign addr[33284] = 1827424302;
assign addr[33285] = 1837395562;
assign addr[33286] = 1847221128;
assign addr[33287] = 1856900221;
assign addr[33288] = 1866432072;
assign addr[33289] = 1875815927;
assign addr[33290] = 1885051042;
assign addr[33291] = 1894136683;
assign addr[33292] = 1903072131;
assign addr[33293] = 1911856677;
assign addr[33294] = 1920489624;
assign addr[33295] = 1928970288;
assign addr[33296] = 1937297997;
assign addr[33297] = 1945472089;
assign addr[33298] = 1953491918;
assign addr[33299] = 1961356847;
assign addr[33300] = 1969066252;
assign addr[33301] = 1976619522;
assign addr[33302] = 1984016058;
assign addr[33303] = 1991255274;
assign addr[33304] = 1998336596;
assign addr[33305] = 2005259462;
assign addr[33306] = 2012023322;
assign addr[33307] = 2018627642;
assign addr[33308] = 2025071897;
assign addr[33309] = 2031355576;
assign addr[33310] = 2037478181;
assign addr[33311] = 2043439226;
assign addr[33312] = 2049238240;
assign addr[33313] = 2054874761;
assign addr[33314] = 2060348343;
assign addr[33315] = 2065658552;
assign addr[33316] = 2070804967;
assign addr[33317] = 2075787180;
assign addr[33318] = 2080604795;
assign addr[33319] = 2085257431;
assign addr[33320] = 2089744719;
assign addr[33321] = 2094066304;
assign addr[33322] = 2098221841;
assign addr[33323] = 2102211002;
assign addr[33324] = 2106033471;
assign addr[33325] = 2109688944;
assign addr[33326] = 2113177132;
assign addr[33327] = 2116497758;
assign addr[33328] = 2119650558;
assign addr[33329] = 2122635283;
assign addr[33330] = 2125451696;
assign addr[33331] = 2128099574;
assign addr[33332] = 2130578706;
assign addr[33333] = 2132888897;
assign addr[33334] = 2135029962;
assign addr[33335] = 2137001733;
assign addr[33336] = 2138804053;
assign addr[33337] = 2140436778;
assign addr[33338] = 2141899780;
assign addr[33339] = 2143192942;
assign addr[33340] = 2144316162;
assign addr[33341] = 2145269351;
assign addr[33342] = 2146052433;
assign addr[33343] = 2146665347;
assign addr[33344] = 2147108043;
assign addr[33345] = 2147380486;
assign addr[33346] = 2147482655;
assign addr[33347] = 2147414542;
assign addr[33348] = 2147176152;
assign addr[33349] = 2146767505;
assign addr[33350] = 2146188631;
assign addr[33351] = 2145439578;
assign addr[33352] = 2144520405;
assign addr[33353] = 2143431184;
assign addr[33354] = 2142172003;
assign addr[33355] = 2140742960;
assign addr[33356] = 2139144169;
assign addr[33357] = 2137375758;
assign addr[33358] = 2135437865;
assign addr[33359] = 2133330646;
assign addr[33360] = 2131054266;
assign addr[33361] = 2128608907;
assign addr[33362] = 2125994762;
assign addr[33363] = 2123212038;
assign addr[33364] = 2120260957;
assign addr[33365] = 2117141752;
assign addr[33366] = 2113854671;
assign addr[33367] = 2110399974;
assign addr[33368] = 2106777935;
assign addr[33369] = 2102988841;
assign addr[33370] = 2099032994;
assign addr[33371] = 2094910706;
assign addr[33372] = 2090622304;
assign addr[33373] = 2086168128;
assign addr[33374] = 2081548533;
assign addr[33375] = 2076763883;
assign addr[33376] = 2071814558;
assign addr[33377] = 2066700952;
assign addr[33378] = 2061423468;
assign addr[33379] = 2055982526;
assign addr[33380] = 2050378558;
assign addr[33381] = 2044612007;
assign addr[33382] = 2038683330;
assign addr[33383] = 2032592999;
assign addr[33384] = 2026341495;
assign addr[33385] = 2019929315;
assign addr[33386] = 2013356967;
assign addr[33387] = 2006624971;
assign addr[33388] = 1999733863;
assign addr[33389] = 1992684188;
assign addr[33390] = 1985476506;
assign addr[33391] = 1978111387;
assign addr[33392] = 1970589416;
assign addr[33393] = 1962911189;
assign addr[33394] = 1955077316;
assign addr[33395] = 1947088417;
assign addr[33396] = 1938945125;
assign addr[33397] = 1930648088;
assign addr[33398] = 1922197961;
assign addr[33399] = 1913595416;
assign addr[33400] = 1904841135;
assign addr[33401] = 1895935811;
assign addr[33402] = 1886880151;
assign addr[33403] = 1877674873;
assign addr[33404] = 1868320707;
assign addr[33405] = 1858818395;
assign addr[33406] = 1849168689;
assign addr[33407] = 1839372356;
assign addr[33408] = 1829430172;
assign addr[33409] = 1819342925;
assign addr[33410] = 1809111415;
assign addr[33411] = 1798736454;
assign addr[33412] = 1788218865;
assign addr[33413] = 1777559480;
assign addr[33414] = 1766759146;
assign addr[33415] = 1755818718;
assign addr[33416] = 1744739065;
assign addr[33417] = 1733521064;
assign addr[33418] = 1722165606;
assign addr[33419] = 1710673591;
assign addr[33420] = 1699045930;
assign addr[33421] = 1687283545;
assign addr[33422] = 1675387369;
assign addr[33423] = 1663358344;
assign addr[33424] = 1651197426;
assign addr[33425] = 1638905577;
assign addr[33426] = 1626483774;
assign addr[33427] = 1613933000;
assign addr[33428] = 1601254251;
assign addr[33429] = 1588448533;
assign addr[33430] = 1575516860;
assign addr[33431] = 1562460258;
assign addr[33432] = 1549279763;
assign addr[33433] = 1535976419;
assign addr[33434] = 1522551282;
assign addr[33435] = 1509005416;
assign addr[33436] = 1495339895;
assign addr[33437] = 1481555802;
assign addr[33438] = 1467654232;
assign addr[33439] = 1453636285;
assign addr[33440] = 1439503074;
assign addr[33441] = 1425255719;
assign addr[33442] = 1410895350;
assign addr[33443] = 1396423105;
assign addr[33444] = 1381840133;
assign addr[33445] = 1367147589;
assign addr[33446] = 1352346639;
assign addr[33447] = 1337438456;
assign addr[33448] = 1322424222;
assign addr[33449] = 1307305128;
assign addr[33450] = 1292082373;
assign addr[33451] = 1276757164;
assign addr[33452] = 1261330715;
assign addr[33453] = 1245804251;
assign addr[33454] = 1230179002;
assign addr[33455] = 1214456207;
assign addr[33456] = 1198637114;
assign addr[33457] = 1182722976;
assign addr[33458] = 1166715055;
assign addr[33459] = 1150614620;
assign addr[33460] = 1134422949;
assign addr[33461] = 1118141326;
assign addr[33462] = 1101771040;
assign addr[33463] = 1085313391;
assign addr[33464] = 1068769683;
assign addr[33465] = 1052141228;
assign addr[33466] = 1035429345;
assign addr[33467] = 1018635358;
assign addr[33468] = 1001760600;
assign addr[33469] = 984806408;
assign addr[33470] = 967774128;
assign addr[33471] = 950665109;
assign addr[33472] = 933480707;
assign addr[33473] = 916222287;
assign addr[33474] = 898891215;
assign addr[33475] = 881488868;
assign addr[33476] = 864016623;
assign addr[33477] = 846475867;
assign addr[33478] = 828867991;
assign addr[33479] = 811194391;
assign addr[33480] = 793456467;
assign addr[33481] = 775655628;
assign addr[33482] = 757793284;
assign addr[33483] = 739870851;
assign addr[33484] = 721889752;
assign addr[33485] = 703851410;
assign addr[33486] = 685757258;
assign addr[33487] = 667608730;
assign addr[33488] = 649407264;
assign addr[33489] = 631154304;
assign addr[33490] = 612851297;
assign addr[33491] = 594499695;
assign addr[33492] = 576100953;
assign addr[33493] = 557656529;
assign addr[33494] = 539167887;
assign addr[33495] = 520636492;
assign addr[33496] = 502063814;
assign addr[33497] = 483451325;
assign addr[33498] = 464800501;
assign addr[33499] = 446112822;
assign addr[33500] = 427389768;
assign addr[33501] = 408632825;
assign addr[33502] = 389843480;
assign addr[33503] = 371023223;
assign addr[33504] = 352173546;
assign addr[33505] = 333295944;
assign addr[33506] = 314391913;
assign addr[33507] = 295462954;
assign addr[33508] = 276510565;
assign addr[33509] = 257536251;
assign addr[33510] = 238541516;
assign addr[33511] = 219527866;
assign addr[33512] = 200496809;
assign addr[33513] = 181449854;
assign addr[33514] = 162388511;
assign addr[33515] = 143314291;
assign addr[33516] = 124228708;
assign addr[33517] = 105133274;
assign addr[33518] = 86029503;
assign addr[33519] = 66918911;
assign addr[33520] = 47803013;
assign addr[33521] = 28683324;
assign addr[33522] = 9561361;
assign addr[33523] = -9561361;
assign addr[33524] = -28683324;
assign addr[33525] = -47803013;
assign addr[33526] = -66918911;
assign addr[33527] = -86029503;
assign addr[33528] = -105133274;
assign addr[33529] = -124228708;
assign addr[33530] = -143314291;
assign addr[33531] = -162388511;
assign addr[33532] = -181449854;
assign addr[33533] = -200496809;
assign addr[33534] = -219527866;
assign addr[33535] = -238541516;
assign addr[33536] = -257536251;
assign addr[33537] = -276510565;
assign addr[33538] = -295462953;
assign addr[33539] = -314391913;
assign addr[33540] = -333295944;
assign addr[33541] = -352173546;
assign addr[33542] = -371023223;
assign addr[33543] = -389843480;
assign addr[33544] = -408632825;
assign addr[33545] = -427389768;
assign addr[33546] = -446112822;
assign addr[33547] = -464800501;
assign addr[33548] = -483451325;
assign addr[33549] = -502063814;
assign addr[33550] = -520636492;
assign addr[33551] = -539167887;
assign addr[33552] = -557656529;
assign addr[33553] = -576100953;
assign addr[33554] = -594499695;
assign addr[33555] = -612851297;
assign addr[33556] = -631154304;
assign addr[33557] = -649407264;
assign addr[33558] = -667608730;
assign addr[33559] = -685757258;
assign addr[33560] = -703851410;
assign addr[33561] = -721889752;
assign addr[33562] = -739870851;
assign addr[33563] = -757793284;
assign addr[33564] = -775655628;
assign addr[33565] = -793456467;
assign addr[33566] = -811194391;
assign addr[33567] = -828867991;
assign addr[33568] = -846475867;
assign addr[33569] = -864016623;
assign addr[33570] = -881488868;
assign addr[33571] = -898891215;
assign addr[33572] = -916222287;
assign addr[33573] = -933480707;
assign addr[33574] = -950665109;
assign addr[33575] = -967774128;
assign addr[33576] = -984806408;
assign addr[33577] = -1001760600;
assign addr[33578] = -1018635358;
assign addr[33579] = -1035429345;
assign addr[33580] = -1052141228;
assign addr[33581] = -1068769683;
assign addr[33582] = -1085313391;
assign addr[33583] = -1101771040;
assign addr[33584] = -1118141326;
assign addr[33585] = -1134422949;
assign addr[33586] = -1150614620;
assign addr[33587] = -1166715055;
assign addr[33588] = -1182722976;
assign addr[33589] = -1198637114;
assign addr[33590] = -1214456207;
assign addr[33591] = -1230179002;
assign addr[33592] = -1245804251;
assign addr[33593] = -1261330715;
assign addr[33594] = -1276757164;
assign addr[33595] = -1292082373;
assign addr[33596] = -1307305128;
assign addr[33597] = -1322424222;
assign addr[33598] = -1337438456;
assign addr[33599] = -1352346639;
assign addr[33600] = -1367147589;
assign addr[33601] = -1381840133;
assign addr[33602] = -1396423105;
assign addr[33603] = -1410895350;
assign addr[33604] = -1425255719;
assign addr[33605] = -1439503074;
assign addr[33606] = -1453636285;
assign addr[33607] = -1467654232;
assign addr[33608] = -1481555802;
assign addr[33609] = -1495339895;
assign addr[33610] = -1509005416;
assign addr[33611] = -1522551282;
assign addr[33612] = -1535976419;
assign addr[33613] = -1549279763;
assign addr[33614] = -1562460258;
assign addr[33615] = -1575516860;
assign addr[33616] = -1588448533;
assign addr[33617] = -1601254251;
assign addr[33618] = -1613933000;
assign addr[33619] = -1626483774;
assign addr[33620] = -1638905577;
assign addr[33621] = -1651197426;
assign addr[33622] = -1663358344;
assign addr[33623] = -1675387369;
assign addr[33624] = -1687283545;
assign addr[33625] = -1699045930;
assign addr[33626] = -1710673591;
assign addr[33627] = -1722165606;
assign addr[33628] = -1733521064;
assign addr[33629] = -1744739065;
assign addr[33630] = -1755818718;
assign addr[33631] = -1766759146;
assign addr[33632] = -1777559480;
assign addr[33633] = -1788218865;
assign addr[33634] = -1798736454;
assign addr[33635] = -1809111415;
assign addr[33636] = -1819342925;
assign addr[33637] = -1829430172;
assign addr[33638] = -1839372356;
assign addr[33639] = -1849168689;
assign addr[33640] = -1858818395;
assign addr[33641] = -1868320707;
assign addr[33642] = -1877674873;
assign addr[33643] = -1886880151;
assign addr[33644] = -1895935811;
assign addr[33645] = -1904841135;
assign addr[33646] = -1913595416;
assign addr[33647] = -1922197961;
assign addr[33648] = -1930648088;
assign addr[33649] = -1938945125;
assign addr[33650] = -1947088417;
assign addr[33651] = -1955077316;
assign addr[33652] = -1962911189;
assign addr[33653] = -1970589416;
assign addr[33654] = -1978111387;
assign addr[33655] = -1985476506;
assign addr[33656] = -1992684188;
assign addr[33657] = -1999733863;
assign addr[33658] = -2006624971;
assign addr[33659] = -2013356967;
assign addr[33660] = -2019929315;
assign addr[33661] = -2026341495;
assign addr[33662] = -2032592999;
assign addr[33663] = -2038683330;
assign addr[33664] = -2044612007;
assign addr[33665] = -2050378558;
assign addr[33666] = -2055982526;
assign addr[33667] = -2061423468;
assign addr[33668] = -2066700952;
assign addr[33669] = -2071814558;
assign addr[33670] = -2076763883;
assign addr[33671] = -2081548533;
assign addr[33672] = -2086168128;
assign addr[33673] = -2090622304;
assign addr[33674] = -2094910706;
assign addr[33675] = -2099032994;
assign addr[33676] = -2102988841;
assign addr[33677] = -2106777935;
assign addr[33678] = -2110399974;
assign addr[33679] = -2113854671;
assign addr[33680] = -2117141752;
assign addr[33681] = -2120260957;
assign addr[33682] = -2123212038;
assign addr[33683] = -2125994762;
assign addr[33684] = -2128608907;
assign addr[33685] = -2131054266;
assign addr[33686] = -2133330646;
assign addr[33687] = -2135437865;
assign addr[33688] = -2137375758;
assign addr[33689] = -2139144169;
assign addr[33690] = -2140742960;
assign addr[33691] = -2142172003;
assign addr[33692] = -2143431184;
assign addr[33693] = -2144520405;
assign addr[33694] = -2145439578;
assign addr[33695] = -2146188631;
assign addr[33696] = -2146767505;
assign addr[33697] = -2147176152;
assign addr[33698] = -2147414542;
assign addr[33699] = -2147482655;
assign addr[33700] = -2147380486;
assign addr[33701] = -2147108043;
assign addr[33702] = -2146665347;
assign addr[33703] = -2146052433;
assign addr[33704] = -2145269351;
assign addr[33705] = -2144316162;
assign addr[33706] = -2143192942;
assign addr[33707] = -2141899780;
assign addr[33708] = -2140436778;
assign addr[33709] = -2138804053;
assign addr[33710] = -2137001733;
assign addr[33711] = -2135029962;
assign addr[33712] = -2132888897;
assign addr[33713] = -2130578706;
assign addr[33714] = -2128099574;
assign addr[33715] = -2125451696;
assign addr[33716] = -2122635283;
assign addr[33717] = -2119650558;
assign addr[33718] = -2116497758;
assign addr[33719] = -2113177132;
assign addr[33720] = -2109688944;
assign addr[33721] = -2106033471;
assign addr[33722] = -2102211002;
assign addr[33723] = -2098221841;
assign addr[33724] = -2094066304;
assign addr[33725] = -2089744719;
assign addr[33726] = -2085257431;
assign addr[33727] = -2080604795;
assign addr[33728] = -2075787180;
assign addr[33729] = -2070804967;
assign addr[33730] = -2065658552;
assign addr[33731] = -2060348343;
assign addr[33732] = -2054874761;
assign addr[33733] = -2049238240;
assign addr[33734] = -2043439226;
assign addr[33735] = -2037478181;
assign addr[33736] = -2031355576;
assign addr[33737] = -2025071897;
assign addr[33738] = -2018627642;
assign addr[33739] = -2012023322;
assign addr[33740] = -2005259462;
assign addr[33741] = -1998336596;
assign addr[33742] = -1991255274;
assign addr[33743] = -1984016058;
assign addr[33744] = -1976619522;
assign addr[33745] = -1969066252;
assign addr[33746] = -1961356847;
assign addr[33747] = -1953491918;
assign addr[33748] = -1945472089;
assign addr[33749] = -1937297997;
assign addr[33750] = -1928970288;
assign addr[33751] = -1920489624;
assign addr[33752] = -1911856677;
assign addr[33753] = -1903072131;
assign addr[33754] = -1894136683;
assign addr[33755] = -1885051042;
assign addr[33756] = -1875815927;
assign addr[33757] = -1866432072;
assign addr[33758] = -1856900221;
assign addr[33759] = -1847221128;
assign addr[33760] = -1837395562;
assign addr[33761] = -1827424302;
assign addr[33762] = -1817308138;
assign addr[33763] = -1807047873;
assign addr[33764] = -1796644320;
assign addr[33765] = -1786098304;
assign addr[33766] = -1775410662;
assign addr[33767] = -1764582240;
assign addr[33768] = -1753613897;
assign addr[33769] = -1742506504;
assign addr[33770] = -1731260941;
assign addr[33771] = -1719878099;
assign addr[33772] = -1708358881;
assign addr[33773] = -1696704201;
assign addr[33774] = -1684914983;
assign addr[33775] = -1672992161;
assign addr[33776] = -1660936681;
assign addr[33777] = -1648749499;
assign addr[33778] = -1636431582;
assign addr[33779] = -1623983905;
assign addr[33780] = -1611407456;
assign addr[33781] = -1598703233;
assign addr[33782] = -1585872242;
assign addr[33783] = -1572915501;
assign addr[33784] = -1559834037;
assign addr[33785] = -1546628888;
assign addr[33786] = -1533301101;
assign addr[33787] = -1519851733;
assign addr[33788] = -1506281850;
assign addr[33789] = -1492592527;
assign addr[33790] = -1478784851;
assign addr[33791] = -1464859917;
assign addr[33792] = -1450818828;
assign addr[33793] = -1436662698;
assign addr[33794] = -1422392650;
assign addr[33795] = -1408009814;
assign addr[33796] = -1393515332;
assign addr[33797] = -1378910353;
assign addr[33798] = -1364196034;
assign addr[33799] = -1349373543;
assign addr[33800] = -1334444055;
assign addr[33801] = -1319408754;
assign addr[33802] = -1304268832;
assign addr[33803] = -1289025489;
assign addr[33804] = -1273679934;
assign addr[33805] = -1258233384;
assign addr[33806] = -1242687064;
assign addr[33807] = -1227042207;
assign addr[33808] = -1211300053;
assign addr[33809] = -1195461849;
assign addr[33810] = -1179528853;
assign addr[33811] = -1163502328;
assign addr[33812] = -1147383544;
assign addr[33813] = -1131173780;
assign addr[33814] = -1114874320;
assign addr[33815] = -1098486458;
assign addr[33816] = -1082011492;
assign addr[33817] = -1065450729;
assign addr[33818] = -1048805483;
assign addr[33819] = -1032077073;
assign addr[33820] = -1015266825;
assign addr[33821] = -998376073;
assign addr[33822] = -981406156;
assign addr[33823] = -964358420;
assign addr[33824] = -947234215;
assign addr[33825] = -930034901;
assign addr[33826] = -912761841;
assign addr[33827] = -895416404;
assign addr[33828] = -877999966;
assign addr[33829] = -860513908;
assign addr[33830] = -842959617;
assign addr[33831] = -825338484;
assign addr[33832] = -807651907;
assign addr[33833] = -789901288;
assign addr[33834] = -772088034;
assign addr[33835] = -754213559;
assign addr[33836] = -736279279;
assign addr[33837] = -718286617;
assign addr[33838] = -700236999;
assign addr[33839] = -682131857;
assign addr[33840] = -663972625;
assign addr[33841] = -645760745;
assign addr[33842] = -627497660;
assign addr[33843] = -609184818;
assign addr[33844] = -590823671;
assign addr[33845] = -572415676;
assign addr[33846] = -553962291;
assign addr[33847] = -535464981;
assign addr[33848] = -516925212;
assign addr[33849] = -498344454;
assign addr[33850] = -479724180;
assign addr[33851] = -461065866;
assign addr[33852] = -442370993;
assign addr[33853] = -423641043;
assign addr[33854] = -404877501;
assign addr[33855] = -386081854;
assign addr[33856] = -367255594;
assign addr[33857] = -348400212;
assign addr[33858] = -329517204;
assign addr[33859] = -310608068;
assign addr[33860] = -291674302;
assign addr[33861] = -272717408;
assign addr[33862] = -253738890;
assign addr[33863] = -234740251;
assign addr[33864] = -215722999;
assign addr[33865] = -196688642;
assign addr[33866] = -177638688;
assign addr[33867] = -158574649;
assign addr[33868] = -139498035;
assign addr[33869] = -120410361;
assign addr[33870] = -101313138;
assign addr[33871] = -82207882;
assign addr[33872] = -63096108;
assign addr[33873] = -43979330;
assign addr[33874] = -24859065;
assign addr[33875] = -5736829;
assign addr[33876] = 13385863;
assign addr[33877] = 32507492;
assign addr[33878] = 51626544;
assign addr[33879] = 70741503;
assign addr[33880] = 89850852;
assign addr[33881] = 108953076;
assign addr[33882] = 128046661;
assign addr[33883] = 147130093;
assign addr[33884] = 166201858;
assign addr[33885] = 185260444;
assign addr[33886] = 204304341;
assign addr[33887] = 223332037;
assign addr[33888] = 242342025;
assign addr[33889] = 261332796;
assign addr[33890] = 280302845;
assign addr[33891] = 299250668;
assign addr[33892] = 318174762;
assign addr[33893] = 337073627;
assign addr[33894] = 355945764;
assign addr[33895] = 374789676;
assign addr[33896] = 393603870;
assign addr[33897] = 412386854;
assign addr[33898] = 431137138;
assign addr[33899] = 449853235;
assign addr[33900] = 468533662;
assign addr[33901] = 487176937;
assign addr[33902] = 505781581;
assign addr[33903] = 524346121;
assign addr[33904] = 542869083;
assign addr[33905] = 561348998;
assign addr[33906] = 579784402;
assign addr[33907] = 598173833;
assign addr[33908] = 616515832;
assign addr[33909] = 634808946;
assign addr[33910] = 653051723;
assign addr[33911] = 671242716;
assign addr[33912] = 689380485;
assign addr[33913] = 707463589;
assign addr[33914] = 725490597;
assign addr[33915] = 743460077;
assign addr[33916] = 761370605;
assign addr[33917] = 779220762;
assign addr[33918] = 797009130;
assign addr[33919] = 814734301;
assign addr[33920] = 832394869;
assign addr[33921] = 849989433;
assign addr[33922] = 867516597;
assign addr[33923] = 884974973;
assign addr[33924] = 902363176;
assign addr[33925] = 919679827;
assign addr[33926] = 936923553;
assign addr[33927] = 954092986;
assign addr[33928] = 971186766;
assign addr[33929] = 988203537;
assign addr[33930] = 1005141949;
assign addr[33931] = 1022000660;
assign addr[33932] = 1038778332;
assign addr[33933] = 1055473635;
assign addr[33934] = 1072085246;
assign addr[33935] = 1088611847;
assign addr[33936] = 1105052128;
assign addr[33937] = 1121404785;
assign addr[33938] = 1137668521;
assign addr[33939] = 1153842047;
assign addr[33940] = 1169924081;
assign addr[33941] = 1185913346;
assign addr[33942] = 1201808576;
assign addr[33943] = 1217608510;
assign addr[33944] = 1233311895;
assign addr[33945] = 1248917486;
assign addr[33946] = 1264424045;
assign addr[33947] = 1279830344;
assign addr[33948] = 1295135159;
assign addr[33949] = 1310337279;
assign addr[33950] = 1325435496;
assign addr[33951] = 1340428615;
assign addr[33952] = 1355315445;
assign addr[33953] = 1370094808;
assign addr[33954] = 1384765530;
assign addr[33955] = 1399326449;
assign addr[33956] = 1413776410;
assign addr[33957] = 1428114267;
assign addr[33958] = 1442338884;
assign addr[33959] = 1456449131;
assign addr[33960] = 1470443891;
assign addr[33961] = 1484322054;
assign addr[33962] = 1498082520;
assign addr[33963] = 1511724196;
assign addr[33964] = 1525246002;
assign addr[33965] = 1538646865;
assign addr[33966] = 1551925723;
assign addr[33967] = 1565081523;
assign addr[33968] = 1578113222;
assign addr[33969] = 1591019785;
assign addr[33970] = 1603800191;
assign addr[33971] = 1616453425;
assign addr[33972] = 1628978484;
assign addr[33973] = 1641374375;
assign addr[33974] = 1653640115;
assign addr[33975] = 1665774731;
assign addr[33976] = 1677777262;
assign addr[33977] = 1689646755;
assign addr[33978] = 1701382270;
assign addr[33979] = 1712982875;
assign addr[33980] = 1724447652;
assign addr[33981] = 1735775690;
assign addr[33982] = 1746966091;
assign addr[33983] = 1758017969;
assign addr[33984] = 1768930447;
assign addr[33985] = 1779702660;
assign addr[33986] = 1790333753;
assign addr[33987] = 1800822883;
assign addr[33988] = 1811169220;
assign addr[33989] = 1821371941;
assign addr[33990] = 1831430239;
assign addr[33991] = 1841343316;
assign addr[33992] = 1851110385;
assign addr[33993] = 1860730673;
assign addr[33994] = 1870203416;
assign addr[33995] = 1879527863;
assign addr[33996] = 1888703276;
assign addr[33997] = 1897728925;
assign addr[33998] = 1906604097;
assign addr[33999] = 1915328086;
assign addr[34000] = 1923900201;
assign addr[34001] = 1932319763;
assign addr[34002] = 1940586104;
assign addr[34003] = 1948698568;
assign addr[34004] = 1956656513;
assign addr[34005] = 1964459306;
assign addr[34006] = 1972106330;
assign addr[34007] = 1979596978;
assign addr[34008] = 1986930656;
assign addr[34009] = 1994106782;
assign addr[34010] = 2001124788;
assign addr[34011] = 2007984117;
assign addr[34012] = 2014684225;
assign addr[34013] = 2021224581;
assign addr[34014] = 2027604666;
assign addr[34015] = 2033823974;
assign addr[34016] = 2039882013;
assign addr[34017] = 2045778302;
assign addr[34018] = 2051512372;
assign addr[34019] = 2057083771;
assign addr[34020] = 2062492055;
assign addr[34021] = 2067736796;
assign addr[34022] = 2072817579;
assign addr[34023] = 2077733999;
assign addr[34024] = 2082485668;
assign addr[34025] = 2087072209;
assign addr[34026] = 2091493257;
assign addr[34027] = 2095748463;
assign addr[34028] = 2099837489;
assign addr[34029] = 2103760010;
assign addr[34030] = 2107515716;
assign addr[34031] = 2111104309;
assign addr[34032] = 2114525505;
assign addr[34033] = 2117779031;
assign addr[34034] = 2120864631;
assign addr[34035] = 2123782059;
assign addr[34036] = 2126531084;
assign addr[34037] = 2129111488;
assign addr[34038] = 2131523066;
assign addr[34039] = 2133765628;
assign addr[34040] = 2135838995;
assign addr[34041] = 2137743003;
assign addr[34042] = 2139477502;
assign addr[34043] = 2141042352;
assign addr[34044] = 2142437431;
assign addr[34045] = 2143662628;
assign addr[34046] = 2144717846;
assign addr[34047] = 2145603001;
assign addr[34048] = 2146318022;
assign addr[34049] = 2146862854;
assign addr[34050] = 2147237452;
assign addr[34051] = 2147441787;
assign addr[34052] = 2147475844;
assign addr[34053] = 2147339619;
assign addr[34054] = 2147033123;
assign addr[34055] = 2146556380;
assign addr[34056] = 2145909429;
assign addr[34057] = 2145092320;
assign addr[34058] = 2144105118;
assign addr[34059] = 2142947902;
assign addr[34060] = 2141620763;
assign addr[34061] = 2140123807;
assign addr[34062] = 2138457152;
assign addr[34063] = 2136620930;
assign addr[34064] = 2134615288;
assign addr[34065] = 2132440383;
assign addr[34066] = 2130096389;
assign addr[34067] = 2127583492;
assign addr[34068] = 2124901890;
assign addr[34069] = 2122051796;
assign addr[34070] = 2119033436;
assign addr[34071] = 2115847050;
assign addr[34072] = 2112492891;
assign addr[34073] = 2108971223;
assign addr[34074] = 2105282327;
assign addr[34075] = 2101426496;
assign addr[34076] = 2097404033;
assign addr[34077] = 2093215260;
assign addr[34078] = 2088860507;
assign addr[34079] = 2084340120;
assign addr[34080] = 2079654458;
assign addr[34081] = 2074803892;
assign addr[34082] = 2069788807;
assign addr[34083] = 2064609600;
assign addr[34084] = 2059266683;
assign addr[34085] = 2053760478;
assign addr[34086] = 2048091422;
assign addr[34087] = 2042259965;
assign addr[34088] = 2036266570;
assign addr[34089] = 2030111710;
assign addr[34090] = 2023795876;
assign addr[34091] = 2017319567;
assign addr[34092] = 2010683297;
assign addr[34093] = 2003887591;
assign addr[34094] = 1996932990;
assign addr[34095] = 1989820044;
assign addr[34096] = 1982549318;
assign addr[34097] = 1975121388;
assign addr[34098] = 1967536842;
assign addr[34099] = 1959796283;
assign addr[34100] = 1951900324;
assign addr[34101] = 1943849591;
assign addr[34102] = 1935644723;
assign addr[34103] = 1927286370;
assign addr[34104] = 1918775195;
assign addr[34105] = 1910111873;
assign addr[34106] = 1901297091;
assign addr[34107] = 1892331547;
assign addr[34108] = 1883215953;
assign addr[34109] = 1873951032;
assign addr[34110] = 1864537518;
assign addr[34111] = 1854976157;
assign addr[34112] = 1845267708;
assign addr[34113] = 1835412941;
assign addr[34114] = 1825412636;
assign addr[34115] = 1815267588;
assign addr[34116] = 1804978599;
assign addr[34117] = 1794546487;
assign addr[34118] = 1783972079;
assign addr[34119] = 1773256212;
assign addr[34120] = 1762399737;
assign addr[34121] = 1751403515;
assign addr[34122] = 1740268417;
assign addr[34123] = 1728995326;
assign addr[34124] = 1717585136;
assign addr[34125] = 1706038753;
assign addr[34126] = 1694357091;
assign addr[34127] = 1682541077;
assign addr[34128] = 1670591647;
assign addr[34129] = 1658509750;
assign addr[34130] = 1646296344;
assign addr[34131] = 1633952396;
assign addr[34132] = 1621478885;
assign addr[34133] = 1608876801;
assign addr[34134] = 1596147143;
assign addr[34135] = 1583290921;
assign addr[34136] = 1570309153;
assign addr[34137] = 1557202869;
assign addr[34138] = 1543973108;
assign addr[34139] = 1530620920;
assign addr[34140] = 1517147363;
assign addr[34141] = 1503553506;
assign addr[34142] = 1489840425;
assign addr[34143] = 1476009210;
assign addr[34144] = 1462060956;
assign addr[34145] = 1447996770;
assign addr[34146] = 1433817766;
assign addr[34147] = 1419525069;
assign addr[34148] = 1405119813;
assign addr[34149] = 1390603139;
assign addr[34150] = 1375976199;
assign addr[34151] = 1361240152;
assign addr[34152] = 1346396168;
assign addr[34153] = 1331445422;
assign addr[34154] = 1316389101;
assign addr[34155] = 1301228398;
assign addr[34156] = 1285964516;
assign addr[34157] = 1270598665;
assign addr[34158] = 1255132063;
assign addr[34159] = 1239565936;
assign addr[34160] = 1223901520;
assign addr[34161] = 1208140056;
assign addr[34162] = 1192282793;
assign addr[34163] = 1176330990;
assign addr[34164] = 1160285911;
assign addr[34165] = 1144148829;
assign addr[34166] = 1127921022;
assign addr[34167] = 1111603778;
assign addr[34168] = 1095198391;
assign addr[34169] = 1078706161;
assign addr[34170] = 1062128397;
assign addr[34171] = 1045466412;
assign addr[34172] = 1028721528;
assign addr[34173] = 1011895073;
assign addr[34174] = 994988380;
assign addr[34175] = 978002791;
assign addr[34176] = 960939653;
assign addr[34177] = 943800318;
assign addr[34178] = 926586145;
assign addr[34179] = 909298500;
assign addr[34180] = 891938752;
assign addr[34181] = 874508280;
assign addr[34182] = 857008464;
assign addr[34183] = 839440693;
assign addr[34184] = 821806359;
assign addr[34185] = 804106861;
assign addr[34186] = 786343603;
assign addr[34187] = 768517992;
assign addr[34188] = 750631442;
assign addr[34189] = 732685372;
assign addr[34190] = 714681204;
assign addr[34191] = 696620367;
assign addr[34192] = 678504291;
assign addr[34193] = 660334415;
assign addr[34194] = 642112178;
assign addr[34195] = 623839025;
assign addr[34196] = 605516406;
assign addr[34197] = 587145773;
assign addr[34198] = 568728583;
assign addr[34199] = 550266296;
assign addr[34200] = 531760377;
assign addr[34201] = 513212292;
assign addr[34202] = 494623513;
assign addr[34203] = 475995513;
assign addr[34204] = 457329769;
assign addr[34205] = 438627762;
assign addr[34206] = 419890975;
assign addr[34207] = 401120892;
assign addr[34208] = 382319004;
assign addr[34209] = 363486799;
assign addr[34210] = 344625773;
assign addr[34211] = 325737419;
assign addr[34212] = 306823237;
assign addr[34213] = 287884725;
assign addr[34214] = 268923386;
assign addr[34215] = 249940723;
assign addr[34216] = 230938242;
assign addr[34217] = 211917448;
assign addr[34218] = 192879850;
assign addr[34219] = 173826959;
assign addr[34220] = 154760284;
assign addr[34221] = 135681337;
assign addr[34222] = 116591632;
assign addr[34223] = 97492681;
assign addr[34224] = 78386000;
assign addr[34225] = 59273104;
assign addr[34226] = 40155507;
assign addr[34227] = 21034727;
assign addr[34228] = 1912278;
assign addr[34229] = -17210322;
assign addr[34230] = -36331557;
assign addr[34231] = -55449912;
assign addr[34232] = -74563870;
assign addr[34233] = -93671915;
assign addr[34234] = -112772533;
assign addr[34235] = -131864208;
assign addr[34236] = -150945428;
assign addr[34237] = -170014678;
assign addr[34238] = -189070447;
assign addr[34239] = -208111224;
assign addr[34240] = -227135500;
assign addr[34241] = -246141764;
assign addr[34242] = -265128512;
assign addr[34243] = -284094236;
assign addr[34244] = -303037433;
assign addr[34245] = -321956601;
assign addr[34246] = -340850240;
assign addr[34247] = -359716852;
assign addr[34248] = -378554940;
assign addr[34249] = -397363011;
assign addr[34250] = -416139574;
assign addr[34251] = -434883140;
assign addr[34252] = -453592221;
assign addr[34253] = -472265336;
assign addr[34254] = -490901003;
assign addr[34255] = -509497745;
assign addr[34256] = -528054086;
assign addr[34257] = -546568556;
assign addr[34258] = -565039687;
assign addr[34259] = -583466013;
assign addr[34260] = -601846074;
assign addr[34261] = -620178412;
assign addr[34262] = -638461574;
assign addr[34263] = -656694110;
assign addr[34264] = -674874574;
assign addr[34265] = -693001525;
assign addr[34266] = -711073524;
assign addr[34267] = -729089140;
assign addr[34268] = -747046944;
assign addr[34269] = -764945512;
assign addr[34270] = -782783424;
assign addr[34271] = -800559266;
assign addr[34272] = -818271628;
assign addr[34273] = -835919107;
assign addr[34274] = -853500302;
assign addr[34275] = -871013820;
assign addr[34276] = -888458272;
assign addr[34277] = -905832274;
assign addr[34278] = -923134450;
assign addr[34279] = -940363427;
assign addr[34280] = -957517838;
assign addr[34281] = -974596324;
assign addr[34282] = -991597531;
assign addr[34283] = -1008520110;
assign addr[34284] = -1025362720;
assign addr[34285] = -1042124025;
assign addr[34286] = -1058802695;
assign addr[34287] = -1075397409;
assign addr[34288] = -1091906851;
assign addr[34289] = -1108329711;
assign addr[34290] = -1124664687;
assign addr[34291] = -1140910484;
assign addr[34292] = -1157065814;
assign addr[34293] = -1173129396;
assign addr[34294] = -1189099956;
assign addr[34295] = -1204976227;
assign addr[34296] = -1220756951;
assign addr[34297] = -1236440877;
assign addr[34298] = -1252026760;
assign addr[34299] = -1267513365;
assign addr[34300] = -1282899464;
assign addr[34301] = -1298183838;
assign addr[34302] = -1313365273;
assign addr[34303] = -1328442566;
assign addr[34304] = -1343414522;
assign addr[34305] = -1358279953;
assign addr[34306] = -1373037681;
assign addr[34307] = -1387686535;
assign addr[34308] = -1402225355;
assign addr[34309] = -1416652986;
assign addr[34310] = -1430968286;
assign addr[34311] = -1445170118;
assign addr[34312] = -1459257358;
assign addr[34313] = -1473228887;
assign addr[34314] = -1487083598;
assign addr[34315] = -1500820393;
assign addr[34316] = -1514438181;
assign addr[34317] = -1527935884;
assign addr[34318] = -1541312431;
assign addr[34319] = -1554566762;
assign addr[34320] = -1567697824;
assign addr[34321] = -1580704578;
assign addr[34322] = -1593585992;
assign addr[34323] = -1606341043;
assign addr[34324] = -1618968722;
assign addr[34325] = -1631468027;
assign addr[34326] = -1643837966;
assign addr[34327] = -1656077559;
assign addr[34328] = -1668185835;
assign addr[34329] = -1680161834;
assign addr[34330] = -1692004606;
assign addr[34331] = -1703713213;
assign addr[34332] = -1715286726;
assign addr[34333] = -1726724227;
assign addr[34334] = -1738024810;
assign addr[34335] = -1749187577;
assign addr[34336] = -1760211645;
assign addr[34337] = -1771096139;
assign addr[34338] = -1781840195;
assign addr[34339] = -1792442963;
assign addr[34340] = -1802903601;
assign addr[34341] = -1813221279;
assign addr[34342] = -1823395180;
assign addr[34343] = -1833424497;
assign addr[34344] = -1843308435;
assign addr[34345] = -1853046210;
assign addr[34346] = -1862637049;
assign addr[34347] = -1872080193;
assign addr[34348] = -1881374892;
assign addr[34349] = -1890520410;
assign addr[34350] = -1899516021;
assign addr[34351] = -1908361011;
assign addr[34352] = -1917054681;
assign addr[34353] = -1925596340;
assign addr[34354] = -1933985310;
assign addr[34355] = -1942220928;
assign addr[34356] = -1950302539;
assign addr[34357] = -1958229503;
assign addr[34358] = -1966001192;
assign addr[34359] = -1973616989;
assign addr[34360] = -1981076290;
assign addr[34361] = -1988378503;
assign addr[34362] = -1995523051;
assign addr[34363] = -2002509365;
assign addr[34364] = -2009336893;
assign addr[34365] = -2016005093;
assign addr[34366] = -2022513436;
assign addr[34367] = -2028861406;
assign addr[34368] = -2035048499;
assign addr[34369] = -2041074226;
assign addr[34370] = -2046938108;
assign addr[34371] = -2052639680;
assign addr[34372] = -2058178491;
assign addr[34373] = -2063554100;
assign addr[34374] = -2068766083;
assign addr[34375] = -2073814024;
assign addr[34376] = -2078697525;
assign addr[34377] = -2083416198;
assign addr[34378] = -2087969669;
assign addr[34379] = -2092357577;
assign addr[34380] = -2096579573;
assign addr[34381] = -2100635323;
assign addr[34382] = -2104524506;
assign addr[34383] = -2108246813;
assign addr[34384] = -2111801949;
assign addr[34385] = -2115189632;
assign addr[34386] = -2118409593;
assign addr[34387] = -2121461578;
assign addr[34388] = -2124345343;
assign addr[34389] = -2127060661;
assign addr[34390] = -2129607316;
assign addr[34391] = -2131985106;
assign addr[34392] = -2134193842;
assign addr[34393] = -2136233350;
assign addr[34394] = -2138103468;
assign addr[34395] = -2139804048;
assign addr[34396] = -2141334954;
assign addr[34397] = -2142696065;
assign addr[34398] = -2143887273;
assign addr[34399] = -2144908484;
assign addr[34400] = -2145759618;
assign addr[34401] = -2146440605;
assign addr[34402] = -2146951393;
assign addr[34403] = -2147291941;
assign addr[34404] = -2147462221;
assign addr[34405] = -2147462221;
assign addr[34406] = -2147291941;
assign addr[34407] = -2146951393;
assign addr[34408] = -2146440605;
assign addr[34409] = -2145759618;
assign addr[34410] = -2144908484;
assign addr[34411] = -2143887273;
assign addr[34412] = -2142696065;
assign addr[34413] = -2141334954;
assign addr[34414] = -2139804048;
assign addr[34415] = -2138103468;
assign addr[34416] = -2136233350;
assign addr[34417] = -2134193842;
assign addr[34418] = -2131985106;
assign addr[34419] = -2129607316;
assign addr[34420] = -2127060661;
assign addr[34421] = -2124345343;
assign addr[34422] = -2121461578;
assign addr[34423] = -2118409593;
assign addr[34424] = -2115189632;
assign addr[34425] = -2111801949;
assign addr[34426] = -2108246813;
assign addr[34427] = -2104524506;
assign addr[34428] = -2100635323;
assign addr[34429] = -2096579573;
assign addr[34430] = -2092357577;
assign addr[34431] = -2087969669;
assign addr[34432] = -2083416198;
assign addr[34433] = -2078697525;
assign addr[34434] = -2073814024;
assign addr[34435] = -2068766083;
assign addr[34436] = -2063554100;
assign addr[34437] = -2058178491;
assign addr[34438] = -2052639680;
assign addr[34439] = -2046938108;
assign addr[34440] = -2041074226;
assign addr[34441] = -2035048499;
assign addr[34442] = -2028861406;
assign addr[34443] = -2022513436;
assign addr[34444] = -2016005093;
assign addr[34445] = -2009336893;
assign addr[34446] = -2002509365;
assign addr[34447] = -1995523051;
assign addr[34448] = -1988378503;
assign addr[34449] = -1981076290;
assign addr[34450] = -1973616989;
assign addr[34451] = -1966001192;
assign addr[34452] = -1958229503;
assign addr[34453] = -1950302539;
assign addr[34454] = -1942220928;
assign addr[34455] = -1933985310;
assign addr[34456] = -1925596340;
assign addr[34457] = -1917054681;
assign addr[34458] = -1908361011;
assign addr[34459] = -1899516021;
assign addr[34460] = -1890520410;
assign addr[34461] = -1881374892;
assign addr[34462] = -1872080193;
assign addr[34463] = -1862637049;
assign addr[34464] = -1853046210;
assign addr[34465] = -1843308435;
assign addr[34466] = -1833424497;
assign addr[34467] = -1823395180;
assign addr[34468] = -1813221279;
assign addr[34469] = -1802903601;
assign addr[34470] = -1792442963;
assign addr[34471] = -1781840195;
assign addr[34472] = -1771096139;
assign addr[34473] = -1760211645;
assign addr[34474] = -1749187577;
assign addr[34475] = -1738024810;
assign addr[34476] = -1726724227;
assign addr[34477] = -1715286726;
assign addr[34478] = -1703713213;
assign addr[34479] = -1692004606;
assign addr[34480] = -1680161834;
assign addr[34481] = -1668185835;
assign addr[34482] = -1656077559;
assign addr[34483] = -1643837966;
assign addr[34484] = -1631468027;
assign addr[34485] = -1618968722;
assign addr[34486] = -1606341043;
assign addr[34487] = -1593585992;
assign addr[34488] = -1580704578;
assign addr[34489] = -1567697824;
assign addr[34490] = -1554566762;
assign addr[34491] = -1541312431;
assign addr[34492] = -1527935884;
assign addr[34493] = -1514438181;
assign addr[34494] = -1500820393;
assign addr[34495] = -1487083598;
assign addr[34496] = -1473228887;
assign addr[34497] = -1459257358;
assign addr[34498] = -1445170118;
assign addr[34499] = -1430968286;
assign addr[34500] = -1416652986;
assign addr[34501] = -1402225355;
assign addr[34502] = -1387686535;
assign addr[34503] = -1373037681;
assign addr[34504] = -1358279953;
assign addr[34505] = -1343414522;
assign addr[34506] = -1328442566;
assign addr[34507] = -1313365273;
assign addr[34508] = -1298183838;
assign addr[34509] = -1282899464;
assign addr[34510] = -1267513365;
assign addr[34511] = -1252026760;
assign addr[34512] = -1236440877;
assign addr[34513] = -1220756951;
assign addr[34514] = -1204976227;
assign addr[34515] = -1189099956;
assign addr[34516] = -1173129396;
assign addr[34517] = -1157065814;
assign addr[34518] = -1140910484;
assign addr[34519] = -1124664687;
assign addr[34520] = -1108329711;
assign addr[34521] = -1091906851;
assign addr[34522] = -1075397409;
assign addr[34523] = -1058802695;
assign addr[34524] = -1042124025;
assign addr[34525] = -1025362720;
assign addr[34526] = -1008520110;
assign addr[34527] = -991597531;
assign addr[34528] = -974596324;
assign addr[34529] = -957517838;
assign addr[34530] = -940363427;
assign addr[34531] = -923134450;
assign addr[34532] = -905832274;
assign addr[34533] = -888458272;
assign addr[34534] = -871013820;
assign addr[34535] = -853500302;
assign addr[34536] = -835919107;
assign addr[34537] = -818271628;
assign addr[34538] = -800559266;
assign addr[34539] = -782783424;
assign addr[34540] = -764945512;
assign addr[34541] = -747046944;
assign addr[34542] = -729089140;
assign addr[34543] = -711073524;
assign addr[34544] = -693001525;
assign addr[34545] = -674874574;
assign addr[34546] = -656694110;
assign addr[34547] = -638461574;
assign addr[34548] = -620178412;
assign addr[34549] = -601846074;
assign addr[34550] = -583466013;
assign addr[34551] = -565039687;
assign addr[34552] = -546568556;
assign addr[34553] = -528054086;
assign addr[34554] = -509497745;
assign addr[34555] = -490901003;
assign addr[34556] = -472265336;
assign addr[34557] = -453592221;
assign addr[34558] = -434883140;
assign addr[34559] = -416139574;
assign addr[34560] = -397363011;
assign addr[34561] = -378554940;
assign addr[34562] = -359716852;
assign addr[34563] = -340850240;
assign addr[34564] = -321956601;
assign addr[34565] = -303037433;
assign addr[34566] = -284094236;
assign addr[34567] = -265128512;
assign addr[34568] = -246141764;
assign addr[34569] = -227135500;
assign addr[34570] = -208111224;
assign addr[34571] = -189070447;
assign addr[34572] = -170014678;
assign addr[34573] = -150945428;
assign addr[34574] = -131864208;
assign addr[34575] = -112772533;
assign addr[34576] = -93671915;
assign addr[34577] = -74563870;
assign addr[34578] = -55449912;
assign addr[34579] = -36331557;
assign addr[34580] = -17210322;
assign addr[34581] = 1912278;
assign addr[34582] = 21034727;
assign addr[34583] = 40155507;
assign addr[34584] = 59273104;
assign addr[34585] = 78386000;
assign addr[34586] = 97492681;
assign addr[34587] = 116591632;
assign addr[34588] = 135681337;
assign addr[34589] = 154760284;
assign addr[34590] = 173826959;
assign addr[34591] = 192879850;
assign addr[34592] = 211917448;
assign addr[34593] = 230938242;
assign addr[34594] = 249940723;
assign addr[34595] = 268923386;
assign addr[34596] = 287884725;
assign addr[34597] = 306823237;
assign addr[34598] = 325737419;
assign addr[34599] = 344625773;
assign addr[34600] = 363486799;
assign addr[34601] = 382319004;
assign addr[34602] = 401120892;
assign addr[34603] = 419890975;
assign addr[34604] = 438627762;
assign addr[34605] = 457329769;
assign addr[34606] = 475995513;
assign addr[34607] = 494623513;
assign addr[34608] = 513212292;
assign addr[34609] = 531760377;
assign addr[34610] = 550266296;
assign addr[34611] = 568728583;
assign addr[34612] = 587145773;
assign addr[34613] = 605516406;
assign addr[34614] = 623839025;
assign addr[34615] = 642112178;
assign addr[34616] = 660334415;
assign addr[34617] = 678504291;
assign addr[34618] = 696620367;
assign addr[34619] = 714681204;
assign addr[34620] = 732685372;
assign addr[34621] = 750631442;
assign addr[34622] = 768517992;
assign addr[34623] = 786343603;
assign addr[34624] = 804106861;
assign addr[34625] = 821806359;
assign addr[34626] = 839440693;
assign addr[34627] = 857008464;
assign addr[34628] = 874508280;
assign addr[34629] = 891938752;
assign addr[34630] = 909298500;
assign addr[34631] = 926586145;
assign addr[34632] = 943800318;
assign addr[34633] = 960939653;
assign addr[34634] = 978002791;
assign addr[34635] = 994988380;
assign addr[34636] = 1011895073;
assign addr[34637] = 1028721528;
assign addr[34638] = 1045466412;
assign addr[34639] = 1062128397;
assign addr[34640] = 1078706161;
assign addr[34641] = 1095198391;
assign addr[34642] = 1111603778;
assign addr[34643] = 1127921022;
assign addr[34644] = 1144148829;
assign addr[34645] = 1160285911;
assign addr[34646] = 1176330990;
assign addr[34647] = 1192282793;
assign addr[34648] = 1208140056;
assign addr[34649] = 1223901520;
assign addr[34650] = 1239565936;
assign addr[34651] = 1255132063;
assign addr[34652] = 1270598665;
assign addr[34653] = 1285964516;
assign addr[34654] = 1301228398;
assign addr[34655] = 1316389101;
assign addr[34656] = 1331445422;
assign addr[34657] = 1346396168;
assign addr[34658] = 1361240152;
assign addr[34659] = 1375976199;
assign addr[34660] = 1390603139;
assign addr[34661] = 1405119813;
assign addr[34662] = 1419525069;
assign addr[34663] = 1433817766;
assign addr[34664] = 1447996770;
assign addr[34665] = 1462060956;
assign addr[34666] = 1476009210;
assign addr[34667] = 1489840425;
assign addr[34668] = 1503553506;
assign addr[34669] = 1517147363;
assign addr[34670] = 1530620920;
assign addr[34671] = 1543973108;
assign addr[34672] = 1557202869;
assign addr[34673] = 1570309153;
assign addr[34674] = 1583290921;
assign addr[34675] = 1596147143;
assign addr[34676] = 1608876801;
assign addr[34677] = 1621478885;
assign addr[34678] = 1633952396;
assign addr[34679] = 1646296344;
assign addr[34680] = 1658509750;
assign addr[34681] = 1670591647;
assign addr[34682] = 1682541077;
assign addr[34683] = 1694357091;
assign addr[34684] = 1706038753;
assign addr[34685] = 1717585136;
assign addr[34686] = 1728995326;
assign addr[34687] = 1740268417;
assign addr[34688] = 1751403515;
assign addr[34689] = 1762399737;
assign addr[34690] = 1773256212;
assign addr[34691] = 1783972079;
assign addr[34692] = 1794546487;
assign addr[34693] = 1804978599;
assign addr[34694] = 1815267588;
assign addr[34695] = 1825412636;
assign addr[34696] = 1835412941;
assign addr[34697] = 1845267708;
assign addr[34698] = 1854976157;
assign addr[34699] = 1864537518;
assign addr[34700] = 1873951032;
assign addr[34701] = 1883215953;
assign addr[34702] = 1892331547;
assign addr[34703] = 1901297091;
assign addr[34704] = 1910111873;
assign addr[34705] = 1918775195;
assign addr[34706] = 1927286370;
assign addr[34707] = 1935644723;
assign addr[34708] = 1943849591;
assign addr[34709] = 1951900324;
assign addr[34710] = 1959796283;
assign addr[34711] = 1967536842;
assign addr[34712] = 1975121388;
assign addr[34713] = 1982549318;
assign addr[34714] = 1989820044;
assign addr[34715] = 1996932990;
assign addr[34716] = 2003887591;
assign addr[34717] = 2010683297;
assign addr[34718] = 2017319567;
assign addr[34719] = 2023795876;
assign addr[34720] = 2030111710;
assign addr[34721] = 2036266570;
assign addr[34722] = 2042259965;
assign addr[34723] = 2048091422;
assign addr[34724] = 2053760478;
assign addr[34725] = 2059266683;
assign addr[34726] = 2064609600;
assign addr[34727] = 2069788807;
assign addr[34728] = 2074803892;
assign addr[34729] = 2079654458;
assign addr[34730] = 2084340120;
assign addr[34731] = 2088860507;
assign addr[34732] = 2093215260;
assign addr[34733] = 2097404033;
assign addr[34734] = 2101426496;
assign addr[34735] = 2105282327;
assign addr[34736] = 2108971223;
assign addr[34737] = 2112492891;
assign addr[34738] = 2115847050;
assign addr[34739] = 2119033436;
assign addr[34740] = 2122051796;
assign addr[34741] = 2124901890;
assign addr[34742] = 2127583492;
assign addr[34743] = 2130096389;
assign addr[34744] = 2132440383;
assign addr[34745] = 2134615288;
assign addr[34746] = 2136620930;
assign addr[34747] = 2138457152;
assign addr[34748] = 2140123807;
assign addr[34749] = 2141620763;
assign addr[34750] = 2142947902;
assign addr[34751] = 2144105118;
assign addr[34752] = 2145092320;
assign addr[34753] = 2145909429;
assign addr[34754] = 2146556380;
assign addr[34755] = 2147033123;
assign addr[34756] = 2147339619;
assign addr[34757] = 2147475844;
assign addr[34758] = 2147441787;
assign addr[34759] = 2147237452;
assign addr[34760] = 2146862854;
assign addr[34761] = 2146318022;
assign addr[34762] = 2145603001;
assign addr[34763] = 2144717846;
assign addr[34764] = 2143662628;
assign addr[34765] = 2142437431;
assign addr[34766] = 2141042352;
assign addr[34767] = 2139477502;
assign addr[34768] = 2137743003;
assign addr[34769] = 2135838995;
assign addr[34770] = 2133765628;
assign addr[34771] = 2131523066;
assign addr[34772] = 2129111488;
assign addr[34773] = 2126531084;
assign addr[34774] = 2123782059;
assign addr[34775] = 2120864631;
assign addr[34776] = 2117779031;
assign addr[34777] = 2114525505;
assign addr[34778] = 2111104309;
assign addr[34779] = 2107515716;
assign addr[34780] = 2103760010;
assign addr[34781] = 2099837489;
assign addr[34782] = 2095748463;
assign addr[34783] = 2091493257;
assign addr[34784] = 2087072209;
assign addr[34785] = 2082485668;
assign addr[34786] = 2077733999;
assign addr[34787] = 2072817579;
assign addr[34788] = 2067736796;
assign addr[34789] = 2062492055;
assign addr[34790] = 2057083771;
assign addr[34791] = 2051512372;
assign addr[34792] = 2045778302;
assign addr[34793] = 2039882013;
assign addr[34794] = 2033823974;
assign addr[34795] = 2027604666;
assign addr[34796] = 2021224581;
assign addr[34797] = 2014684225;
assign addr[34798] = 2007984117;
assign addr[34799] = 2001124788;
assign addr[34800] = 1994106782;
assign addr[34801] = 1986930656;
assign addr[34802] = 1979596978;
assign addr[34803] = 1972106330;
assign addr[34804] = 1964459306;
assign addr[34805] = 1956656513;
assign addr[34806] = 1948698568;
assign addr[34807] = 1940586104;
assign addr[34808] = 1932319763;
assign addr[34809] = 1923900201;
assign addr[34810] = 1915328086;
assign addr[34811] = 1906604097;
assign addr[34812] = 1897728925;
assign addr[34813] = 1888703276;
assign addr[34814] = 1879527863;
assign addr[34815] = 1870203416;
assign addr[34816] = 1860730673;
assign addr[34817] = 1851110385;
assign addr[34818] = 1841343316;
assign addr[34819] = 1831430239;
assign addr[34820] = 1821371941;
assign addr[34821] = 1811169220;
assign addr[34822] = 1800822883;
assign addr[34823] = 1790333753;
assign addr[34824] = 1779702660;
assign addr[34825] = 1768930447;
assign addr[34826] = 1758017969;
assign addr[34827] = 1746966091;
assign addr[34828] = 1735775690;
assign addr[34829] = 1724447652;
assign addr[34830] = 1712982875;
assign addr[34831] = 1701382270;
assign addr[34832] = 1689646755;
assign addr[34833] = 1677777262;
assign addr[34834] = 1665774731;
assign addr[34835] = 1653640115;
assign addr[34836] = 1641374375;
assign addr[34837] = 1628978484;
assign addr[34838] = 1616453425;
assign addr[34839] = 1603800191;
assign addr[34840] = 1591019785;
assign addr[34841] = 1578113222;
assign addr[34842] = 1565081523;
assign addr[34843] = 1551925723;
assign addr[34844] = 1538646865;
assign addr[34845] = 1525246002;
assign addr[34846] = 1511724196;
assign addr[34847] = 1498082520;
assign addr[34848] = 1484322054;
assign addr[34849] = 1470443891;
assign addr[34850] = 1456449131;
assign addr[34851] = 1442338884;
assign addr[34852] = 1428114267;
assign addr[34853] = 1413776410;
assign addr[34854] = 1399326449;
assign addr[34855] = 1384765530;
assign addr[34856] = 1370094808;
assign addr[34857] = 1355315445;
assign addr[34858] = 1340428615;
assign addr[34859] = 1325435496;
assign addr[34860] = 1310337279;
assign addr[34861] = 1295135159;
assign addr[34862] = 1279830344;
assign addr[34863] = 1264424045;
assign addr[34864] = 1248917486;
assign addr[34865] = 1233311895;
assign addr[34866] = 1217608510;
assign addr[34867] = 1201808576;
assign addr[34868] = 1185913346;
assign addr[34869] = 1169924081;
assign addr[34870] = 1153842047;
assign addr[34871] = 1137668521;
assign addr[34872] = 1121404785;
assign addr[34873] = 1105052128;
assign addr[34874] = 1088611847;
assign addr[34875] = 1072085246;
assign addr[34876] = 1055473635;
assign addr[34877] = 1038778332;
assign addr[34878] = 1022000660;
assign addr[34879] = 1005141949;
assign addr[34880] = 988203537;
assign addr[34881] = 971186766;
assign addr[34882] = 954092986;
assign addr[34883] = 936923553;
assign addr[34884] = 919679827;
assign addr[34885] = 902363176;
assign addr[34886] = 884974973;
assign addr[34887] = 867516597;
assign addr[34888] = 849989433;
assign addr[34889] = 832394869;
assign addr[34890] = 814734301;
assign addr[34891] = 797009130;
assign addr[34892] = 779220762;
assign addr[34893] = 761370605;
assign addr[34894] = 743460077;
assign addr[34895] = 725490597;
assign addr[34896] = 707463589;
assign addr[34897] = 689380485;
assign addr[34898] = 671242716;
assign addr[34899] = 653051723;
assign addr[34900] = 634808946;
assign addr[34901] = 616515832;
assign addr[34902] = 598173833;
assign addr[34903] = 579784402;
assign addr[34904] = 561348998;
assign addr[34905] = 542869083;
assign addr[34906] = 524346121;
assign addr[34907] = 505781581;
assign addr[34908] = 487176937;
assign addr[34909] = 468533662;
assign addr[34910] = 449853235;
assign addr[34911] = 431137138;
assign addr[34912] = 412386854;
assign addr[34913] = 393603870;
assign addr[34914] = 374789676;
assign addr[34915] = 355945764;
assign addr[34916] = 337073627;
assign addr[34917] = 318174762;
assign addr[34918] = 299250668;
assign addr[34919] = 280302845;
assign addr[34920] = 261332796;
assign addr[34921] = 242342025;
assign addr[34922] = 223332037;
assign addr[34923] = 204304341;
assign addr[34924] = 185260444;
assign addr[34925] = 166201858;
assign addr[34926] = 147130093;
assign addr[34927] = 128046661;
assign addr[34928] = 108953076;
assign addr[34929] = 89850852;
assign addr[34930] = 70741503;
assign addr[34931] = 51626544;
assign addr[34932] = 32507492;
assign addr[34933] = 13385863;
assign addr[34934] = -5736829;
assign addr[34935] = -24859065;
assign addr[34936] = -43979330;
assign addr[34937] = -63096108;
assign addr[34938] = -82207882;
assign addr[34939] = -101313138;
assign addr[34940] = -120410361;
assign addr[34941] = -139498035;
assign addr[34942] = -158574649;
assign addr[34943] = -177638688;
assign addr[34944] = -196688642;
assign addr[34945] = -215722999;
assign addr[34946] = -234740251;
assign addr[34947] = -253738890;
assign addr[34948] = -272717408;
assign addr[34949] = -291674302;
assign addr[34950] = -310608068;
assign addr[34951] = -329517204;
assign addr[34952] = -348400212;
assign addr[34953] = -367255594;
assign addr[34954] = -386081854;
assign addr[34955] = -404877501;
assign addr[34956] = -423641043;
assign addr[34957] = -442370993;
assign addr[34958] = -461065866;
assign addr[34959] = -479724180;
assign addr[34960] = -498344454;
assign addr[34961] = -516925212;
assign addr[34962] = -535464981;
assign addr[34963] = -553962291;
assign addr[34964] = -572415676;
assign addr[34965] = -590823671;
assign addr[34966] = -609184818;
assign addr[34967] = -627497660;
assign addr[34968] = -645760745;
assign addr[34969] = -663972625;
assign addr[34970] = -682131857;
assign addr[34971] = -700236999;
assign addr[34972] = -718286617;
assign addr[34973] = -736279279;
assign addr[34974] = -754213559;
assign addr[34975] = -772088034;
assign addr[34976] = -789901288;
assign addr[34977] = -807651907;
assign addr[34978] = -825338484;
assign addr[34979] = -842959617;
assign addr[34980] = -860513908;
assign addr[34981] = -877999966;
assign addr[34982] = -895416404;
assign addr[34983] = -912761841;
assign addr[34984] = -930034901;
assign addr[34985] = -947234215;
assign addr[34986] = -964358420;
assign addr[34987] = -981406156;
assign addr[34988] = -998376073;
assign addr[34989] = -1015266825;
assign addr[34990] = -1032077073;
assign addr[34991] = -1048805483;
assign addr[34992] = -1065450729;
assign addr[34993] = -1082011492;
assign addr[34994] = -1098486458;
assign addr[34995] = -1114874320;
assign addr[34996] = -1131173780;
assign addr[34997] = -1147383544;
assign addr[34998] = -1163502328;
assign addr[34999] = -1179528853;
assign addr[35000] = -1195461849;
assign addr[35001] = -1211300053;
assign addr[35002] = -1227042207;
assign addr[35003] = -1242687064;
assign addr[35004] = -1258233384;
assign addr[35005] = -1273679934;
assign addr[35006] = -1289025489;
assign addr[35007] = -1304268832;
assign addr[35008] = -1319408754;
assign addr[35009] = -1334444055;
assign addr[35010] = -1349373543;
assign addr[35011] = -1364196034;
assign addr[35012] = -1378910353;
assign addr[35013] = -1393515332;
assign addr[35014] = -1408009814;
assign addr[35015] = -1422392650;
assign addr[35016] = -1436662698;
assign addr[35017] = -1450818828;
assign addr[35018] = -1464859917;
assign addr[35019] = -1478784851;
assign addr[35020] = -1492592527;
assign addr[35021] = -1506281850;
assign addr[35022] = -1519851733;
assign addr[35023] = -1533301101;
assign addr[35024] = -1546628888;
assign addr[35025] = -1559834037;
assign addr[35026] = -1572915501;
assign addr[35027] = -1585872242;
assign addr[35028] = -1598703233;
assign addr[35029] = -1611407456;
assign addr[35030] = -1623983905;
assign addr[35031] = -1636431582;
assign addr[35032] = -1648749499;
assign addr[35033] = -1660936681;
assign addr[35034] = -1672992161;
assign addr[35035] = -1684914983;
assign addr[35036] = -1696704201;
assign addr[35037] = -1708358881;
assign addr[35038] = -1719878099;
assign addr[35039] = -1731260941;
assign addr[35040] = -1742506504;
assign addr[35041] = -1753613897;
assign addr[35042] = -1764582240;
assign addr[35043] = -1775410662;
assign addr[35044] = -1786098304;
assign addr[35045] = -1796644320;
assign addr[35046] = -1807047873;
assign addr[35047] = -1817308138;
assign addr[35048] = -1827424302;
assign addr[35049] = -1837395562;
assign addr[35050] = -1847221128;
assign addr[35051] = -1856900221;
assign addr[35052] = -1866432072;
assign addr[35053] = -1875815927;
assign addr[35054] = -1885051042;
assign addr[35055] = -1894136683;
assign addr[35056] = -1903072131;
assign addr[35057] = -1911856677;
assign addr[35058] = -1920489624;
assign addr[35059] = -1928970288;
assign addr[35060] = -1937297997;
assign addr[35061] = -1945472089;
assign addr[35062] = -1953491918;
assign addr[35063] = -1961356847;
assign addr[35064] = -1969066252;
assign addr[35065] = -1976619522;
assign addr[35066] = -1984016058;
assign addr[35067] = -1991255274;
assign addr[35068] = -1998336596;
assign addr[35069] = -2005259462;
assign addr[35070] = -2012023322;
assign addr[35071] = -2018627642;
assign addr[35072] = -2025071897;
assign addr[35073] = -2031355576;
assign addr[35074] = -2037478181;
assign addr[35075] = -2043439226;
assign addr[35076] = -2049238240;
assign addr[35077] = -2054874761;
assign addr[35078] = -2060348343;
assign addr[35079] = -2065658552;
assign addr[35080] = -2070804967;
assign addr[35081] = -2075787180;
assign addr[35082] = -2080604795;
assign addr[35083] = -2085257431;
assign addr[35084] = -2089744719;
assign addr[35085] = -2094066304;
assign addr[35086] = -2098221841;
assign addr[35087] = -2102211002;
assign addr[35088] = -2106033471;
assign addr[35089] = -2109688944;
assign addr[35090] = -2113177132;
assign addr[35091] = -2116497758;
assign addr[35092] = -2119650558;
assign addr[35093] = -2122635283;
assign addr[35094] = -2125451696;
assign addr[35095] = -2128099574;
assign addr[35096] = -2130578706;
assign addr[35097] = -2132888897;
assign addr[35098] = -2135029962;
assign addr[35099] = -2137001733;
assign addr[35100] = -2138804053;
assign addr[35101] = -2140436778;
assign addr[35102] = -2141899780;
assign addr[35103] = -2143192942;
assign addr[35104] = -2144316162;
assign addr[35105] = -2145269351;
assign addr[35106] = -2146052433;
assign addr[35107] = -2146665347;
assign addr[35108] = -2147108043;
assign addr[35109] = -2147380486;
assign addr[35110] = -2147482655;
assign addr[35111] = -2147414542;
assign addr[35112] = -2147176152;
assign addr[35113] = -2146767505;
assign addr[35114] = -2146188631;
assign addr[35115] = -2145439578;
assign addr[35116] = -2144520405;
assign addr[35117] = -2143431184;
assign addr[35118] = -2142172003;
assign addr[35119] = -2140742960;
assign addr[35120] = -2139144169;
assign addr[35121] = -2137375758;
assign addr[35122] = -2135437865;
assign addr[35123] = -2133330646;
assign addr[35124] = -2131054266;
assign addr[35125] = -2128608907;
assign addr[35126] = -2125994762;
assign addr[35127] = -2123212038;
assign addr[35128] = -2120260957;
assign addr[35129] = -2117141752;
assign addr[35130] = -2113854671;
assign addr[35131] = -2110399974;
assign addr[35132] = -2106777935;
assign addr[35133] = -2102988841;
assign addr[35134] = -2099032994;
assign addr[35135] = -2094910706;
assign addr[35136] = -2090622304;
assign addr[35137] = -2086168128;
assign addr[35138] = -2081548533;
assign addr[35139] = -2076763883;
assign addr[35140] = -2071814558;
assign addr[35141] = -2066700952;
assign addr[35142] = -2061423468;
assign addr[35143] = -2055982526;
assign addr[35144] = -2050378558;
assign addr[35145] = -2044612007;
assign addr[35146] = -2038683330;
assign addr[35147] = -2032592999;
assign addr[35148] = -2026341495;
assign addr[35149] = -2019929315;
assign addr[35150] = -2013356967;
assign addr[35151] = -2006624971;
assign addr[35152] = -1999733863;
assign addr[35153] = -1992684188;
assign addr[35154] = -1985476506;
assign addr[35155] = -1978111387;
assign addr[35156] = -1970589416;
assign addr[35157] = -1962911189;
assign addr[35158] = -1955077316;
assign addr[35159] = -1947088417;
assign addr[35160] = -1938945125;
assign addr[35161] = -1930648088;
assign addr[35162] = -1922197961;
assign addr[35163] = -1913595416;
assign addr[35164] = -1904841135;
assign addr[35165] = -1895935811;
assign addr[35166] = -1886880151;
assign addr[35167] = -1877674873;
assign addr[35168] = -1868320707;
assign addr[35169] = -1858818395;
assign addr[35170] = -1849168689;
assign addr[35171] = -1839372356;
assign addr[35172] = -1829430172;
assign addr[35173] = -1819342925;
assign addr[35174] = -1809111415;
assign addr[35175] = -1798736454;
assign addr[35176] = -1788218865;
assign addr[35177] = -1777559480;
assign addr[35178] = -1766759146;
assign addr[35179] = -1755818718;
assign addr[35180] = -1744739065;
assign addr[35181] = -1733521064;
assign addr[35182] = -1722165606;
assign addr[35183] = -1710673591;
assign addr[35184] = -1699045930;
assign addr[35185] = -1687283545;
assign addr[35186] = -1675387369;
assign addr[35187] = -1663358344;
assign addr[35188] = -1651197426;
assign addr[35189] = -1638905577;
assign addr[35190] = -1626483774;
assign addr[35191] = -1613933000;
assign addr[35192] = -1601254251;
assign addr[35193] = -1588448533;
assign addr[35194] = -1575516860;
assign addr[35195] = -1562460258;
assign addr[35196] = -1549279763;
assign addr[35197] = -1535976419;
assign addr[35198] = -1522551282;
assign addr[35199] = -1509005416;
assign addr[35200] = -1495339895;
assign addr[35201] = -1481555802;
assign addr[35202] = -1467654232;
assign addr[35203] = -1453636285;
assign addr[35204] = -1439503074;
assign addr[35205] = -1425255719;
assign addr[35206] = -1410895350;
assign addr[35207] = -1396423105;
assign addr[35208] = -1381840133;
assign addr[35209] = -1367147589;
assign addr[35210] = -1352346639;
assign addr[35211] = -1337438456;
assign addr[35212] = -1322424222;
assign addr[35213] = -1307305128;
assign addr[35214] = -1292082373;
assign addr[35215] = -1276757164;
assign addr[35216] = -1261330715;
assign addr[35217] = -1245804251;
assign addr[35218] = -1230179002;
assign addr[35219] = -1214456207;
assign addr[35220] = -1198637114;
assign addr[35221] = -1182722976;
assign addr[35222] = -1166715055;
assign addr[35223] = -1150614620;
assign addr[35224] = -1134422949;
assign addr[35225] = -1118141326;
assign addr[35226] = -1101771040;
assign addr[35227] = -1085313391;
assign addr[35228] = -1068769683;
assign addr[35229] = -1052141228;
assign addr[35230] = -1035429345;
assign addr[35231] = -1018635358;
assign addr[35232] = -1001760600;
assign addr[35233] = -984806408;
assign addr[35234] = -967774128;
assign addr[35235] = -950665109;
assign addr[35236] = -933480707;
assign addr[35237] = -916222287;
assign addr[35238] = -898891215;
assign addr[35239] = -881488868;
assign addr[35240] = -864016623;
assign addr[35241] = -846475867;
assign addr[35242] = -828867991;
assign addr[35243] = -811194391;
assign addr[35244] = -793456467;
assign addr[35245] = -775655628;
assign addr[35246] = -757793284;
assign addr[35247] = -739870851;
assign addr[35248] = -721889752;
assign addr[35249] = -703851410;
assign addr[35250] = -685757258;
assign addr[35251] = -667608730;
assign addr[35252] = -649407264;
assign addr[35253] = -631154304;
assign addr[35254] = -612851297;
assign addr[35255] = -594499695;
assign addr[35256] = -576100953;
assign addr[35257] = -557656529;
assign addr[35258] = -539167887;
assign addr[35259] = -520636492;
assign addr[35260] = -502063814;
assign addr[35261] = -483451325;
assign addr[35262] = -464800501;
assign addr[35263] = -446112822;
assign addr[35264] = -427389768;
assign addr[35265] = -408632825;
assign addr[35266] = -389843480;
assign addr[35267] = -371023223;
assign addr[35268] = -352173546;
assign addr[35269] = -333295944;
assign addr[35270] = -314391913;
assign addr[35271] = -295462954;
assign addr[35272] = -276510565;
assign addr[35273] = -257536251;
assign addr[35274] = -238541516;
assign addr[35275] = -219527866;
assign addr[35276] = -200496809;
assign addr[35277] = -181449854;
assign addr[35278] = -162388511;
assign addr[35279] = -143314291;
assign addr[35280] = -124228708;
assign addr[35281] = -105133274;
assign addr[35282] = -86029503;
assign addr[35283] = -66918911;
assign addr[35284] = -47803013;
assign addr[35285] = -28683324;
assign addr[35286] = -9561361;
assign addr[35287] = 9561361;
assign addr[35288] = 28683324;
assign addr[35289] = 47803013;
assign addr[35290] = 66918911;
assign addr[35291] = 86029503;
assign addr[35292] = 105133274;
assign addr[35293] = 124228708;
assign addr[35294] = 143314291;
assign addr[35295] = 162388511;
assign addr[35296] = 181449854;
assign addr[35297] = 200496809;
assign addr[35298] = 219527866;
assign addr[35299] = 238541516;
assign addr[35300] = 257536251;
assign addr[35301] = 276510565;
assign addr[35302] = 295462953;
assign addr[35303] = 314391913;
assign addr[35304] = 333295944;
assign addr[35305] = 352173546;
assign addr[35306] = 371023223;
assign addr[35307] = 389843480;
assign addr[35308] = 408632825;
assign addr[35309] = 427389768;
assign addr[35310] = 446112822;
assign addr[35311] = 464800501;
assign addr[35312] = 483451325;
assign addr[35313] = 502063814;
assign addr[35314] = 520636492;
assign addr[35315] = 539167887;
assign addr[35316] = 557656529;
assign addr[35317] = 576100953;
assign addr[35318] = 594499695;
assign addr[35319] = 612851297;
assign addr[35320] = 631154304;
assign addr[35321] = 649407264;
assign addr[35322] = 667608730;
assign addr[35323] = 685757258;
assign addr[35324] = 703851410;
assign addr[35325] = 721889752;
assign addr[35326] = 739870851;
assign addr[35327] = 757793284;
assign addr[35328] = 775655628;
assign addr[35329] = 793456467;
assign addr[35330] = 811194391;
assign addr[35331] = 828867991;
assign addr[35332] = 846475867;
assign addr[35333] = 864016623;
assign addr[35334] = 881488868;
assign addr[35335] = 898891215;
assign addr[35336] = 916222287;
assign addr[35337] = 933480707;
assign addr[35338] = 950665109;
assign addr[35339] = 967774128;
assign addr[35340] = 984806408;
assign addr[35341] = 1001760600;
assign addr[35342] = 1018635358;
assign addr[35343] = 1035429345;
assign addr[35344] = 1052141228;
assign addr[35345] = 1068769683;
assign addr[35346] = 1085313391;
assign addr[35347] = 1101771040;
assign addr[35348] = 1118141326;
assign addr[35349] = 1134422949;
assign addr[35350] = 1150614620;
assign addr[35351] = 1166715055;
assign addr[35352] = 1182722976;
assign addr[35353] = 1198637114;
assign addr[35354] = 1214456207;
assign addr[35355] = 1230179002;
assign addr[35356] = 1245804251;
assign addr[35357] = 1261330715;
assign addr[35358] = 1276757164;
assign addr[35359] = 1292082373;
assign addr[35360] = 1307305128;
assign addr[35361] = 1322424222;
assign addr[35362] = 1337438456;
assign addr[35363] = 1352346639;
assign addr[35364] = 1367147589;
assign addr[35365] = 1381840133;
assign addr[35366] = 1396423105;
assign addr[35367] = 1410895350;
assign addr[35368] = 1425255719;
assign addr[35369] = 1439503074;
assign addr[35370] = 1453636285;
assign addr[35371] = 1467654232;
assign addr[35372] = 1481555802;
assign addr[35373] = 1495339895;
assign addr[35374] = 1509005416;
assign addr[35375] = 1522551282;
assign addr[35376] = 1535976419;
assign addr[35377] = 1549279763;
assign addr[35378] = 1562460258;
assign addr[35379] = 1575516860;
assign addr[35380] = 1588448533;
assign addr[35381] = 1601254251;
assign addr[35382] = 1613933000;
assign addr[35383] = 1626483774;
assign addr[35384] = 1638905577;
assign addr[35385] = 1651197426;
assign addr[35386] = 1663358344;
assign addr[35387] = 1675387369;
assign addr[35388] = 1687283545;
assign addr[35389] = 1699045930;
assign addr[35390] = 1710673591;
assign addr[35391] = 1722165606;
assign addr[35392] = 1733521064;
assign addr[35393] = 1744739065;
assign addr[35394] = 1755818718;
assign addr[35395] = 1766759146;
assign addr[35396] = 1777559480;
assign addr[35397] = 1788218865;
assign addr[35398] = 1798736454;
assign addr[35399] = 1809111415;
assign addr[35400] = 1819342925;
assign addr[35401] = 1829430172;
assign addr[35402] = 1839372356;
assign addr[35403] = 1849168689;
assign addr[35404] = 1858818395;
assign addr[35405] = 1868320707;
assign addr[35406] = 1877674873;
assign addr[35407] = 1886880151;
assign addr[35408] = 1895935811;
assign addr[35409] = 1904841135;
assign addr[35410] = 1913595416;
assign addr[35411] = 1922197961;
assign addr[35412] = 1930648088;
assign addr[35413] = 1938945125;
assign addr[35414] = 1947088417;
assign addr[35415] = 1955077316;
assign addr[35416] = 1962911189;
assign addr[35417] = 1970589416;
assign addr[35418] = 1978111387;
assign addr[35419] = 1985476506;
assign addr[35420] = 1992684188;
assign addr[35421] = 1999733863;
assign addr[35422] = 2006624971;
assign addr[35423] = 2013356967;
assign addr[35424] = 2019929315;
assign addr[35425] = 2026341495;
assign addr[35426] = 2032592999;
assign addr[35427] = 2038683330;
assign addr[35428] = 2044612007;
assign addr[35429] = 2050378558;
assign addr[35430] = 2055982526;
assign addr[35431] = 2061423468;
assign addr[35432] = 2066700952;
assign addr[35433] = 2071814558;
assign addr[35434] = 2076763883;
assign addr[35435] = 2081548533;
assign addr[35436] = 2086168128;
assign addr[35437] = 2090622304;
assign addr[35438] = 2094910706;
assign addr[35439] = 2099032994;
assign addr[35440] = 2102988841;
assign addr[35441] = 2106777935;
assign addr[35442] = 2110399974;
assign addr[35443] = 2113854671;
assign addr[35444] = 2117141752;
assign addr[35445] = 2120260957;
assign addr[35446] = 2123212038;
assign addr[35447] = 2125994762;
assign addr[35448] = 2128608907;
assign addr[35449] = 2131054266;
assign addr[35450] = 2133330646;
assign addr[35451] = 2135437865;
assign addr[35452] = 2137375758;
assign addr[35453] = 2139144169;
assign addr[35454] = 2140742960;
assign addr[35455] = 2142172003;
assign addr[35456] = 2143431184;
assign addr[35457] = 2144520405;
assign addr[35458] = 2145439578;
assign addr[35459] = 2146188631;
assign addr[35460] = 2146767505;
assign addr[35461] = 2147176152;
assign addr[35462] = 2147414542;
assign addr[35463] = 2147482655;
assign addr[35464] = 2147380486;
assign addr[35465] = 2147108043;
assign addr[35466] = 2146665347;
assign addr[35467] = 2146052433;
assign addr[35468] = 2145269351;
assign addr[35469] = 2144316162;
assign addr[35470] = 2143192942;
assign addr[35471] = 2141899780;
assign addr[35472] = 2140436778;
assign addr[35473] = 2138804053;
assign addr[35474] = 2137001733;
assign addr[35475] = 2135029962;
assign addr[35476] = 2132888897;
assign addr[35477] = 2130578706;
assign addr[35478] = 2128099574;
assign addr[35479] = 2125451696;
assign addr[35480] = 2122635283;
assign addr[35481] = 2119650558;
assign addr[35482] = 2116497758;
assign addr[35483] = 2113177132;
assign addr[35484] = 2109688944;
assign addr[35485] = 2106033471;
assign addr[35486] = 2102211002;
assign addr[35487] = 2098221841;
assign addr[35488] = 2094066304;
assign addr[35489] = 2089744719;
assign addr[35490] = 2085257431;
assign addr[35491] = 2080604795;
assign addr[35492] = 2075787180;
assign addr[35493] = 2070804967;
assign addr[35494] = 2065658552;
assign addr[35495] = 2060348343;
assign addr[35496] = 2054874761;
assign addr[35497] = 2049238240;
assign addr[35498] = 2043439226;
assign addr[35499] = 2037478181;
assign addr[35500] = 2031355576;
assign addr[35501] = 2025071897;
assign addr[35502] = 2018627642;
assign addr[35503] = 2012023322;
assign addr[35504] = 2005259462;
assign addr[35505] = 1998336596;
assign addr[35506] = 1991255274;
assign addr[35507] = 1984016058;
assign addr[35508] = 1976619522;
assign addr[35509] = 1969066252;
assign addr[35510] = 1961356847;
assign addr[35511] = 1953491918;
assign addr[35512] = 1945472089;
assign addr[35513] = 1937297997;
assign addr[35514] = 1928970288;
assign addr[35515] = 1920489624;
assign addr[35516] = 1911856677;
assign addr[35517] = 1903072131;
assign addr[35518] = 1894136683;
assign addr[35519] = 1885051042;
assign addr[35520] = 1875815927;
assign addr[35521] = 1866432072;
assign addr[35522] = 1856900221;
assign addr[35523] = 1847221128;
assign addr[35524] = 1837395562;
assign addr[35525] = 1827424302;
assign addr[35526] = 1817308138;
assign addr[35527] = 1807047873;
assign addr[35528] = 1796644320;
assign addr[35529] = 1786098304;
assign addr[35530] = 1775410662;
assign addr[35531] = 1764582240;
assign addr[35532] = 1753613897;
assign addr[35533] = 1742506504;
assign addr[35534] = 1731260941;
assign addr[35535] = 1719878099;
assign addr[35536] = 1708358881;
assign addr[35537] = 1696704201;
assign addr[35538] = 1684914983;
assign addr[35539] = 1672992161;
assign addr[35540] = 1660936681;
assign addr[35541] = 1648749499;
assign addr[35542] = 1636431582;
assign addr[35543] = 1623983905;
assign addr[35544] = 1611407456;
assign addr[35545] = 1598703233;
assign addr[35546] = 1585872242;
assign addr[35547] = 1572915501;
assign addr[35548] = 1559834037;
assign addr[35549] = 1546628888;
assign addr[35550] = 1533301101;
assign addr[35551] = 1519851733;
assign addr[35552] = 1506281850;
assign addr[35553] = 1492592527;
assign addr[35554] = 1478784851;
assign addr[35555] = 1464859917;
assign addr[35556] = 1450818828;
assign addr[35557] = 1436662698;
assign addr[35558] = 1422392650;
assign addr[35559] = 1408009814;
assign addr[35560] = 1393515332;
assign addr[35561] = 1378910353;
assign addr[35562] = 1364196034;
assign addr[35563] = 1349373543;
assign addr[35564] = 1334444055;
assign addr[35565] = 1319408754;
assign addr[35566] = 1304268832;
assign addr[35567] = 1289025489;
assign addr[35568] = 1273679934;
assign addr[35569] = 1258233384;
assign addr[35570] = 1242687064;
assign addr[35571] = 1227042207;
assign addr[35572] = 1211300053;
assign addr[35573] = 1195461849;
assign addr[35574] = 1179528853;
assign addr[35575] = 1163502328;
assign addr[35576] = 1147383544;
assign addr[35577] = 1131173780;
assign addr[35578] = 1114874320;
assign addr[35579] = 1098486458;
assign addr[35580] = 1082011492;
assign addr[35581] = 1065450729;
assign addr[35582] = 1048805483;
assign addr[35583] = 1032077073;
assign addr[35584] = 1015266825;
assign addr[35585] = 998376073;
assign addr[35586] = 981406156;
assign addr[35587] = 964358420;
assign addr[35588] = 947234215;
assign addr[35589] = 930034901;
assign addr[35590] = 912761841;
assign addr[35591] = 895416404;
assign addr[35592] = 877999966;
assign addr[35593] = 860513908;
assign addr[35594] = 842959617;
assign addr[35595] = 825338484;
assign addr[35596] = 807651907;
assign addr[35597] = 789901288;
assign addr[35598] = 772088034;
assign addr[35599] = 754213559;
assign addr[35600] = 736279279;
assign addr[35601] = 718286617;
assign addr[35602] = 700236999;
assign addr[35603] = 682131857;
assign addr[35604] = 663972625;
assign addr[35605] = 645760745;
assign addr[35606] = 627497660;
assign addr[35607] = 609184818;
assign addr[35608] = 590823671;
assign addr[35609] = 572415676;
assign addr[35610] = 553962291;
assign addr[35611] = 535464981;
assign addr[35612] = 516925212;
assign addr[35613] = 498344454;
assign addr[35614] = 479724180;
assign addr[35615] = 461065866;
assign addr[35616] = 442370993;
assign addr[35617] = 423641043;
assign addr[35618] = 404877501;
assign addr[35619] = 386081854;
assign addr[35620] = 367255594;
assign addr[35621] = 348400212;
assign addr[35622] = 329517204;
assign addr[35623] = 310608068;
assign addr[35624] = 291674302;
assign addr[35625] = 272717408;
assign addr[35626] = 253738890;
assign addr[35627] = 234740251;
assign addr[35628] = 215722999;
assign addr[35629] = 196688642;
assign addr[35630] = 177638688;
assign addr[35631] = 158574649;
assign addr[35632] = 139498035;
assign addr[35633] = 120410361;
assign addr[35634] = 101313138;
assign addr[35635] = 82207882;
assign addr[35636] = 63096108;
assign addr[35637] = 43979330;
assign addr[35638] = 24859065;
assign addr[35639] = 5736829;
assign addr[35640] = -13385863;
assign addr[35641] = -32507492;
assign addr[35642] = -51626544;
assign addr[35643] = -70741503;
assign addr[35644] = -89850852;
assign addr[35645] = -108953076;
assign addr[35646] = -128046661;
assign addr[35647] = -147130093;
assign addr[35648] = -166201858;
assign addr[35649] = -185260444;
assign addr[35650] = -204304341;
assign addr[35651] = -223332037;
assign addr[35652] = -242342025;
assign addr[35653] = -261332796;
assign addr[35654] = -280302845;
assign addr[35655] = -299250668;
assign addr[35656] = -318174762;
assign addr[35657] = -337073627;
assign addr[35658] = -355945764;
assign addr[35659] = -374789676;
assign addr[35660] = -393603870;
assign addr[35661] = -412386854;
assign addr[35662] = -431137138;
assign addr[35663] = -449853235;
assign addr[35664] = -468533662;
assign addr[35665] = -487176937;
assign addr[35666] = -505781581;
assign addr[35667] = -524346121;
assign addr[35668] = -542869083;
assign addr[35669] = -561348998;
assign addr[35670] = -579784402;
assign addr[35671] = -598173833;
assign addr[35672] = -616515832;
assign addr[35673] = -634808946;
assign addr[35674] = -653051723;
assign addr[35675] = -671242716;
assign addr[35676] = -689380485;
assign addr[35677] = -707463589;
assign addr[35678] = -725490597;
assign addr[35679] = -743460077;
assign addr[35680] = -761370605;
assign addr[35681] = -779220762;
assign addr[35682] = -797009130;
assign addr[35683] = -814734301;
assign addr[35684] = -832394869;
assign addr[35685] = -849989433;
assign addr[35686] = -867516597;
assign addr[35687] = -884974973;
assign addr[35688] = -902363176;
assign addr[35689] = -919679827;
assign addr[35690] = -936923553;
assign addr[35691] = -954092986;
assign addr[35692] = -971186766;
assign addr[35693] = -988203537;
assign addr[35694] = -1005141949;
assign addr[35695] = -1022000660;
assign addr[35696] = -1038778332;
assign addr[35697] = -1055473635;
assign addr[35698] = -1072085246;
assign addr[35699] = -1088611847;
assign addr[35700] = -1105052128;
assign addr[35701] = -1121404785;
assign addr[35702] = -1137668521;
assign addr[35703] = -1153842047;
assign addr[35704] = -1169924081;
assign addr[35705] = -1185913346;
assign addr[35706] = -1201808576;
assign addr[35707] = -1217608510;
assign addr[35708] = -1233311895;
assign addr[35709] = -1248917486;
assign addr[35710] = -1264424045;
assign addr[35711] = -1279830344;
assign addr[35712] = -1295135159;
assign addr[35713] = -1310337279;
assign addr[35714] = -1325435496;
assign addr[35715] = -1340428615;
assign addr[35716] = -1355315445;
assign addr[35717] = -1370094808;
assign addr[35718] = -1384765530;
assign addr[35719] = -1399326449;
assign addr[35720] = -1413776410;
assign addr[35721] = -1428114267;
assign addr[35722] = -1442338884;
assign addr[35723] = -1456449131;
assign addr[35724] = -1470443891;
assign addr[35725] = -1484322054;
assign addr[35726] = -1498082520;
assign addr[35727] = -1511724196;
assign addr[35728] = -1525246002;
assign addr[35729] = -1538646865;
assign addr[35730] = -1551925723;
assign addr[35731] = -1565081523;
assign addr[35732] = -1578113222;
assign addr[35733] = -1591019785;
assign addr[35734] = -1603800191;
assign addr[35735] = -1616453425;
assign addr[35736] = -1628978484;
assign addr[35737] = -1641374375;
assign addr[35738] = -1653640115;
assign addr[35739] = -1665774731;
assign addr[35740] = -1677777262;
assign addr[35741] = -1689646755;
assign addr[35742] = -1701382270;
assign addr[35743] = -1712982875;
assign addr[35744] = -1724447652;
assign addr[35745] = -1735775690;
assign addr[35746] = -1746966091;
assign addr[35747] = -1758017969;
assign addr[35748] = -1768930447;
assign addr[35749] = -1779702660;
assign addr[35750] = -1790333753;
assign addr[35751] = -1800822883;
assign addr[35752] = -1811169220;
assign addr[35753] = -1821371941;
assign addr[35754] = -1831430239;
assign addr[35755] = -1841343316;
assign addr[35756] = -1851110385;
assign addr[35757] = -1860730673;
assign addr[35758] = -1870203416;
assign addr[35759] = -1879527863;
assign addr[35760] = -1888703276;
assign addr[35761] = -1897728925;
assign addr[35762] = -1906604097;
assign addr[35763] = -1915328086;
assign addr[35764] = -1923900201;
assign addr[35765] = -1932319763;
assign addr[35766] = -1940586104;
assign addr[35767] = -1948698568;
assign addr[35768] = -1956656513;
assign addr[35769] = -1964459306;
assign addr[35770] = -1972106330;
assign addr[35771] = -1979596978;
assign addr[35772] = -1986930656;
assign addr[35773] = -1994106782;
assign addr[35774] = -2001124788;
assign addr[35775] = -2007984117;
assign addr[35776] = -2014684225;
assign addr[35777] = -2021224581;
assign addr[35778] = -2027604666;
assign addr[35779] = -2033823974;
assign addr[35780] = -2039882013;
assign addr[35781] = -2045778302;
assign addr[35782] = -2051512372;
assign addr[35783] = -2057083771;
assign addr[35784] = -2062492055;
assign addr[35785] = -2067736796;
assign addr[35786] = -2072817579;
assign addr[35787] = -2077733999;
assign addr[35788] = -2082485668;
assign addr[35789] = -2087072209;
assign addr[35790] = -2091493257;
assign addr[35791] = -2095748463;
assign addr[35792] = -2099837489;
assign addr[35793] = -2103760010;
assign addr[35794] = -2107515716;
assign addr[35795] = -2111104309;
assign addr[35796] = -2114525505;
assign addr[35797] = -2117779031;
assign addr[35798] = -2120864631;
assign addr[35799] = -2123782059;
assign addr[35800] = -2126531084;
assign addr[35801] = -2129111488;
assign addr[35802] = -2131523066;
assign addr[35803] = -2133765628;
assign addr[35804] = -2135838995;
assign addr[35805] = -2137743003;
assign addr[35806] = -2139477502;
assign addr[35807] = -2141042352;
assign addr[35808] = -2142437431;
assign addr[35809] = -2143662628;
assign addr[35810] = -2144717846;
assign addr[35811] = -2145603001;
assign addr[35812] = -2146318022;
assign addr[35813] = -2146862854;
assign addr[35814] = -2147237452;
assign addr[35815] = -2147441787;
assign addr[35816] = -2147475844;
assign addr[35817] = -2147339619;
assign addr[35818] = -2147033123;
assign addr[35819] = -2146556380;
assign addr[35820] = -2145909429;
assign addr[35821] = -2145092320;
assign addr[35822] = -2144105118;
assign addr[35823] = -2142947902;
assign addr[35824] = -2141620763;
assign addr[35825] = -2140123807;
assign addr[35826] = -2138457152;
assign addr[35827] = -2136620930;
assign addr[35828] = -2134615288;
assign addr[35829] = -2132440383;
assign addr[35830] = -2130096389;
assign addr[35831] = -2127583492;
assign addr[35832] = -2124901890;
assign addr[35833] = -2122051796;
assign addr[35834] = -2119033436;
assign addr[35835] = -2115847050;
assign addr[35836] = -2112492891;
assign addr[35837] = -2108971223;
assign addr[35838] = -2105282327;
assign addr[35839] = -2101426496;
assign addr[35840] = -2097404033;
assign addr[35841] = -2093215260;
assign addr[35842] = -2088860507;
assign addr[35843] = -2084340120;
assign addr[35844] = -2079654458;
assign addr[35845] = -2074803892;
assign addr[35846] = -2069788807;
assign addr[35847] = -2064609600;
assign addr[35848] = -2059266683;
assign addr[35849] = -2053760478;
assign addr[35850] = -2048091422;
assign addr[35851] = -2042259965;
assign addr[35852] = -2036266570;
assign addr[35853] = -2030111710;
assign addr[35854] = -2023795876;
assign addr[35855] = -2017319567;
assign addr[35856] = -2010683297;
assign addr[35857] = -2003887591;
assign addr[35858] = -1996932990;
assign addr[35859] = -1989820044;
assign addr[35860] = -1982549318;
assign addr[35861] = -1975121388;
assign addr[35862] = -1967536842;
assign addr[35863] = -1959796283;
assign addr[35864] = -1951900324;
assign addr[35865] = -1943849591;
assign addr[35866] = -1935644723;
assign addr[35867] = -1927286370;
assign addr[35868] = -1918775195;
assign addr[35869] = -1910111873;
assign addr[35870] = -1901297091;
assign addr[35871] = -1892331547;
assign addr[35872] = -1883215953;
assign addr[35873] = -1873951032;
assign addr[35874] = -1864537518;
assign addr[35875] = -1854976157;
assign addr[35876] = -1845267708;
assign addr[35877] = -1835412941;
assign addr[35878] = -1825412636;
assign addr[35879] = -1815267588;
assign addr[35880] = -1804978599;
assign addr[35881] = -1794546487;
assign addr[35882] = -1783972079;
assign addr[35883] = -1773256212;
assign addr[35884] = -1762399737;
assign addr[35885] = -1751403515;
assign addr[35886] = -1740268417;
assign addr[35887] = -1728995326;
assign addr[35888] = -1717585136;
assign addr[35889] = -1706038753;
assign addr[35890] = -1694357091;
assign addr[35891] = -1682541077;
assign addr[35892] = -1670591647;
assign addr[35893] = -1658509750;
assign addr[35894] = -1646296344;
assign addr[35895] = -1633952396;
assign addr[35896] = -1621478885;
assign addr[35897] = -1608876801;
assign addr[35898] = -1596147143;
assign addr[35899] = -1583290921;
assign addr[35900] = -1570309153;
assign addr[35901] = -1557202869;
assign addr[35902] = -1543973108;
assign addr[35903] = -1530620920;
assign addr[35904] = -1517147363;
assign addr[35905] = -1503553506;
assign addr[35906] = -1489840425;
assign addr[35907] = -1476009210;
assign addr[35908] = -1462060956;
assign addr[35909] = -1447996770;
assign addr[35910] = -1433817766;
assign addr[35911] = -1419525069;
assign addr[35912] = -1405119813;
assign addr[35913] = -1390603139;
assign addr[35914] = -1375976199;
assign addr[35915] = -1361240152;
assign addr[35916] = -1346396168;
assign addr[35917] = -1331445422;
assign addr[35918] = -1316389101;
assign addr[35919] = -1301228398;
assign addr[35920] = -1285964516;
assign addr[35921] = -1270598665;
assign addr[35922] = -1255132063;
assign addr[35923] = -1239565936;
assign addr[35924] = -1223901520;
assign addr[35925] = -1208140056;
assign addr[35926] = -1192282793;
assign addr[35927] = -1176330990;
assign addr[35928] = -1160285911;
assign addr[35929] = -1144148829;
assign addr[35930] = -1127921022;
assign addr[35931] = -1111603778;
assign addr[35932] = -1095198391;
assign addr[35933] = -1078706161;
assign addr[35934] = -1062128397;
assign addr[35935] = -1045466412;
assign addr[35936] = -1028721528;
assign addr[35937] = -1011895073;
assign addr[35938] = -994988380;
assign addr[35939] = -978002791;
assign addr[35940] = -960939653;
assign addr[35941] = -943800318;
assign addr[35942] = -926586145;
assign addr[35943] = -909298500;
assign addr[35944] = -891938752;
assign addr[35945] = -874508280;
assign addr[35946] = -857008464;
assign addr[35947] = -839440693;
assign addr[35948] = -821806359;
assign addr[35949] = -804106861;
assign addr[35950] = -786343603;
assign addr[35951] = -768517992;
assign addr[35952] = -750631442;
assign addr[35953] = -732685372;
assign addr[35954] = -714681204;
assign addr[35955] = -696620367;
assign addr[35956] = -678504291;
assign addr[35957] = -660334415;
assign addr[35958] = -642112178;
assign addr[35959] = -623839025;
assign addr[35960] = -605516406;
assign addr[35961] = -587145773;
assign addr[35962] = -568728583;
assign addr[35963] = -550266296;
assign addr[35964] = -531760377;
assign addr[35965] = -513212292;
assign addr[35966] = -494623513;
assign addr[35967] = -475995513;
assign addr[35968] = -457329769;
assign addr[35969] = -438627762;
assign addr[35970] = -419890975;
assign addr[35971] = -401120892;
assign addr[35972] = -382319004;
assign addr[35973] = -363486799;
assign addr[35974] = -344625773;
assign addr[35975] = -325737419;
assign addr[35976] = -306823237;
assign addr[35977] = -287884725;
assign addr[35978] = -268923386;
assign addr[35979] = -249940723;
assign addr[35980] = -230938242;
assign addr[35981] = -211917448;
assign addr[35982] = -192879850;
assign addr[35983] = -173826959;
assign addr[35984] = -154760284;
assign addr[35985] = -135681337;
assign addr[35986] = -116591632;
assign addr[35987] = -97492681;
assign addr[35988] = -78386000;
assign addr[35989] = -59273104;
assign addr[35990] = -40155507;
assign addr[35991] = -21034727;
assign addr[35992] = -1912278;
assign addr[35993] = 17210322;
assign addr[35994] = 36331557;
assign addr[35995] = 55449912;
assign addr[35996] = 74563870;
assign addr[35997] = 93671915;
assign addr[35998] = 112772533;
assign addr[35999] = 131864208;
assign addr[36000] = 150945428;
assign addr[36001] = 170014678;
assign addr[36002] = 189070447;
assign addr[36003] = 208111224;
assign addr[36004] = 227135500;
assign addr[36005] = 246141764;
assign addr[36006] = 265128512;
assign addr[36007] = 284094236;
assign addr[36008] = 303037433;
assign addr[36009] = 321956601;
assign addr[36010] = 340850240;
assign addr[36011] = 359716852;
assign addr[36012] = 378554940;
assign addr[36013] = 397363011;
assign addr[36014] = 416139574;
assign addr[36015] = 434883140;
assign addr[36016] = 453592221;
assign addr[36017] = 472265336;
assign addr[36018] = 490901003;
assign addr[36019] = 509497745;
assign addr[36020] = 528054086;
assign addr[36021] = 546568556;
assign addr[36022] = 565039687;
assign addr[36023] = 583466013;
assign addr[36024] = 601846074;
assign addr[36025] = 620178412;
assign addr[36026] = 638461574;
assign addr[36027] = 656694110;
assign addr[36028] = 674874574;
assign addr[36029] = 693001525;
assign addr[36030] = 711073524;
assign addr[36031] = 729089140;
assign addr[36032] = 747046944;
assign addr[36033] = 764945512;
assign addr[36034] = 782783424;
assign addr[36035] = 800559266;
assign addr[36036] = 818271628;
assign addr[36037] = 835919107;
assign addr[36038] = 853500302;
assign addr[36039] = 871013820;
assign addr[36040] = 888458272;
assign addr[36041] = 905832274;
assign addr[36042] = 923134450;
assign addr[36043] = 940363427;
assign addr[36044] = 957517838;
assign addr[36045] = 974596324;
assign addr[36046] = 991597531;
assign addr[36047] = 1008520110;
assign addr[36048] = 1025362720;
assign addr[36049] = 1042124025;
assign addr[36050] = 1058802695;
assign addr[36051] = 1075397409;
assign addr[36052] = 1091906851;
assign addr[36053] = 1108329711;
assign addr[36054] = 1124664687;
assign addr[36055] = 1140910484;
assign addr[36056] = 1157065814;
assign addr[36057] = 1173129396;
assign addr[36058] = 1189099956;
assign addr[36059] = 1204976227;
assign addr[36060] = 1220756951;
assign addr[36061] = 1236440877;
assign addr[36062] = 1252026760;
assign addr[36063] = 1267513365;
assign addr[36064] = 1282899464;
assign addr[36065] = 1298183838;
assign addr[36066] = 1313365273;
assign addr[36067] = 1328442566;
assign addr[36068] = 1343414522;
assign addr[36069] = 1358279953;
assign addr[36070] = 1373037681;
assign addr[36071] = 1387686535;
assign addr[36072] = 1402225355;
assign addr[36073] = 1416652986;
assign addr[36074] = 1430968286;
assign addr[36075] = 1445170118;
assign addr[36076] = 1459257358;
assign addr[36077] = 1473228887;
assign addr[36078] = 1487083598;
assign addr[36079] = 1500820393;
assign addr[36080] = 1514438181;
assign addr[36081] = 1527935884;
assign addr[36082] = 1541312431;
assign addr[36083] = 1554566762;
assign addr[36084] = 1567697824;
assign addr[36085] = 1580704578;
assign addr[36086] = 1593585992;
assign addr[36087] = 1606341043;
assign addr[36088] = 1618968722;
assign addr[36089] = 1631468027;
assign addr[36090] = 1643837966;
assign addr[36091] = 1656077559;
assign addr[36092] = 1668185835;
assign addr[36093] = 1680161834;
assign addr[36094] = 1692004606;
assign addr[36095] = 1703713213;
assign addr[36096] = 1715286726;
assign addr[36097] = 1726724227;
assign addr[36098] = 1738024810;
assign addr[36099] = 1749187577;
assign addr[36100] = 1760211645;
assign addr[36101] = 1771096139;
assign addr[36102] = 1781840195;
assign addr[36103] = 1792442963;
assign addr[36104] = 1802903601;
assign addr[36105] = 1813221279;
assign addr[36106] = 1823395180;
assign addr[36107] = 1833424497;
assign addr[36108] = 1843308435;
assign addr[36109] = 1853046210;
assign addr[36110] = 1862637049;
assign addr[36111] = 1872080193;
assign addr[36112] = 1881374892;
assign addr[36113] = 1890520410;
assign addr[36114] = 1899516021;
assign addr[36115] = 1908361011;
assign addr[36116] = 1917054681;
assign addr[36117] = 1925596340;
assign addr[36118] = 1933985310;
assign addr[36119] = 1942220928;
assign addr[36120] = 1950302539;
assign addr[36121] = 1958229503;
assign addr[36122] = 1966001192;
assign addr[36123] = 1973616989;
assign addr[36124] = 1981076290;
assign addr[36125] = 1988378503;
assign addr[36126] = 1995523051;
assign addr[36127] = 2002509365;
assign addr[36128] = 2009336893;
assign addr[36129] = 2016005093;
assign addr[36130] = 2022513436;
assign addr[36131] = 2028861406;
assign addr[36132] = 2035048499;
assign addr[36133] = 2041074226;
assign addr[36134] = 2046938108;
assign addr[36135] = 2052639680;
assign addr[36136] = 2058178491;
assign addr[36137] = 2063554100;
assign addr[36138] = 2068766083;
assign addr[36139] = 2073814024;
assign addr[36140] = 2078697525;
assign addr[36141] = 2083416198;
assign addr[36142] = 2087969669;
assign addr[36143] = 2092357577;
assign addr[36144] = 2096579573;
assign addr[36145] = 2100635323;
assign addr[36146] = 2104524506;
assign addr[36147] = 2108246813;
assign addr[36148] = 2111801949;
assign addr[36149] = 2115189632;
assign addr[36150] = 2118409593;
assign addr[36151] = 2121461578;
assign addr[36152] = 2124345343;
assign addr[36153] = 2127060661;
assign addr[36154] = 2129607316;
assign addr[36155] = 2131985106;
assign addr[36156] = 2134193842;
assign addr[36157] = 2136233350;
assign addr[36158] = 2138103468;
assign addr[36159] = 2139804048;
assign addr[36160] = 2141334954;
assign addr[36161] = 2142696065;
assign addr[36162] = 2143887273;
assign addr[36163] = 2144908484;
assign addr[36164] = 2145759618;
assign addr[36165] = 2146440605;
assign addr[36166] = 2146951393;
assign addr[36167] = 2147291941;
assign addr[36168] = 2147462221;
assign addr[36169] = 2147462221;
assign addr[36170] = 2147291941;
assign addr[36171] = 2146951393;
assign addr[36172] = 2146440605;
assign addr[36173] = 2145759618;
assign addr[36174] = 2144908484;
assign addr[36175] = 2143887273;
assign addr[36176] = 2142696065;
assign addr[36177] = 2141334954;
assign addr[36178] = 2139804048;
assign addr[36179] = 2138103468;
assign addr[36180] = 2136233350;
assign addr[36181] = 2134193842;
assign addr[36182] = 2131985106;
assign addr[36183] = 2129607316;
assign addr[36184] = 2127060661;
assign addr[36185] = 2124345343;
assign addr[36186] = 2121461578;
assign addr[36187] = 2118409593;
assign addr[36188] = 2115189632;
assign addr[36189] = 2111801949;
assign addr[36190] = 2108246813;
assign addr[36191] = 2104524506;
assign addr[36192] = 2100635323;
assign addr[36193] = 2096579573;
assign addr[36194] = 2092357577;
assign addr[36195] = 2087969669;
assign addr[36196] = 2083416198;
assign addr[36197] = 2078697525;
assign addr[36198] = 2073814024;
assign addr[36199] = 2068766083;
assign addr[36200] = 2063554100;
assign addr[36201] = 2058178491;
assign addr[36202] = 2052639680;
assign addr[36203] = 2046938108;
assign addr[36204] = 2041074226;
assign addr[36205] = 2035048499;
assign addr[36206] = 2028861406;
assign addr[36207] = 2022513436;
assign addr[36208] = 2016005093;
assign addr[36209] = 2009336893;
assign addr[36210] = 2002509365;
assign addr[36211] = 1995523051;
assign addr[36212] = 1988378503;
assign addr[36213] = 1981076290;
assign addr[36214] = 1973616989;
assign addr[36215] = 1966001192;
assign addr[36216] = 1958229503;
assign addr[36217] = 1950302539;
assign addr[36218] = 1942220928;
assign addr[36219] = 1933985310;
assign addr[36220] = 1925596340;
assign addr[36221] = 1917054681;
assign addr[36222] = 1908361011;
assign addr[36223] = 1899516021;
assign addr[36224] = 1890520410;
assign addr[36225] = 1881374892;
assign addr[36226] = 1872080193;
assign addr[36227] = 1862637049;
assign addr[36228] = 1853046210;
assign addr[36229] = 1843308435;
assign addr[36230] = 1833424497;
assign addr[36231] = 1823395180;
assign addr[36232] = 1813221279;
assign addr[36233] = 1802903601;
assign addr[36234] = 1792442963;
assign addr[36235] = 1781840195;
assign addr[36236] = 1771096139;
assign addr[36237] = 1760211645;
assign addr[36238] = 1749187577;
assign addr[36239] = 1738024810;
assign addr[36240] = 1726724227;
assign addr[36241] = 1715286726;
assign addr[36242] = 1703713213;
assign addr[36243] = 1692004606;
assign addr[36244] = 1680161834;
assign addr[36245] = 1668185835;
assign addr[36246] = 1656077559;
assign addr[36247] = 1643837966;
assign addr[36248] = 1631468027;
assign addr[36249] = 1618968722;
assign addr[36250] = 1606341043;
assign addr[36251] = 1593585992;
assign addr[36252] = 1580704578;
assign addr[36253] = 1567697824;
assign addr[36254] = 1554566762;
assign addr[36255] = 1541312431;
assign addr[36256] = 1527935884;
assign addr[36257] = 1514438181;
assign addr[36258] = 1500820393;
assign addr[36259] = 1487083598;
assign addr[36260] = 1473228887;
assign addr[36261] = 1459257358;
assign addr[36262] = 1445170118;
assign addr[36263] = 1430968286;
assign addr[36264] = 1416652986;
assign addr[36265] = 1402225355;
assign addr[36266] = 1387686535;
assign addr[36267] = 1373037681;
assign addr[36268] = 1358279953;
assign addr[36269] = 1343414522;
assign addr[36270] = 1328442566;
assign addr[36271] = 1313365273;
assign addr[36272] = 1298183838;
assign addr[36273] = 1282899464;
assign addr[36274] = 1267513365;
assign addr[36275] = 1252026760;
assign addr[36276] = 1236440877;
assign addr[36277] = 1220756951;
assign addr[36278] = 1204976227;
assign addr[36279] = 1189099956;
assign addr[36280] = 1173129396;
assign addr[36281] = 1157065814;
assign addr[36282] = 1140910484;
assign addr[36283] = 1124664687;
assign addr[36284] = 1108329711;
assign addr[36285] = 1091906851;
assign addr[36286] = 1075397409;
assign addr[36287] = 1058802695;
assign addr[36288] = 1042124025;
assign addr[36289] = 1025362720;
assign addr[36290] = 1008520110;
assign addr[36291] = 991597531;
assign addr[36292] = 974596324;
assign addr[36293] = 957517838;
assign addr[36294] = 940363427;
assign addr[36295] = 923134450;
assign addr[36296] = 905832274;
assign addr[36297] = 888458272;
assign addr[36298] = 871013820;
assign addr[36299] = 853500302;
assign addr[36300] = 835919107;
assign addr[36301] = 818271628;
assign addr[36302] = 800559266;
assign addr[36303] = 782783424;
assign addr[36304] = 764945512;
assign addr[36305] = 747046944;
assign addr[36306] = 729089140;
assign addr[36307] = 711073524;
assign addr[36308] = 693001525;
assign addr[36309] = 674874574;
assign addr[36310] = 656694110;
assign addr[36311] = 638461574;
assign addr[36312] = 620178412;
assign addr[36313] = 601846074;
assign addr[36314] = 583466013;
assign addr[36315] = 565039687;
assign addr[36316] = 546568556;
assign addr[36317] = 528054086;
assign addr[36318] = 509497745;
assign addr[36319] = 490901003;
assign addr[36320] = 472265336;
assign addr[36321] = 453592221;
assign addr[36322] = 434883140;
assign addr[36323] = 416139574;
assign addr[36324] = 397363011;
assign addr[36325] = 378554940;
assign addr[36326] = 359716852;
assign addr[36327] = 340850240;
assign addr[36328] = 321956601;
assign addr[36329] = 303037433;
assign addr[36330] = 284094236;
assign addr[36331] = 265128512;
assign addr[36332] = 246141764;
assign addr[36333] = 227135500;
assign addr[36334] = 208111224;
assign addr[36335] = 189070447;
assign addr[36336] = 170014678;
assign addr[36337] = 150945428;
assign addr[36338] = 131864208;
assign addr[36339] = 112772533;
assign addr[36340] = 93671915;
assign addr[36341] = 74563870;
assign addr[36342] = 55449912;
assign addr[36343] = 36331557;
assign addr[36344] = 17210322;
assign addr[36345] = -1912278;
assign addr[36346] = -21034727;
assign addr[36347] = -40155507;
assign addr[36348] = -59273104;
assign addr[36349] = -78386000;
assign addr[36350] = -97492681;
assign addr[36351] = -116591632;
assign addr[36352] = -135681337;
assign addr[36353] = -154760284;
assign addr[36354] = -173826959;
assign addr[36355] = -192879850;
assign addr[36356] = -211917448;
assign addr[36357] = -230938242;
assign addr[36358] = -249940723;
assign addr[36359] = -268923386;
assign addr[36360] = -287884725;
assign addr[36361] = -306823237;
assign addr[36362] = -325737419;
assign addr[36363] = -344625773;
assign addr[36364] = -363486799;
assign addr[36365] = -382319004;
assign addr[36366] = -401120892;
assign addr[36367] = -419890975;
assign addr[36368] = -438627762;
assign addr[36369] = -457329769;
assign addr[36370] = -475995513;
assign addr[36371] = -494623513;
assign addr[36372] = -513212292;
assign addr[36373] = -531760377;
assign addr[36374] = -550266296;
assign addr[36375] = -568728583;
assign addr[36376] = -587145773;
assign addr[36377] = -605516406;
assign addr[36378] = -623839025;
assign addr[36379] = -642112178;
assign addr[36380] = -660334415;
assign addr[36381] = -678504291;
assign addr[36382] = -696620367;
assign addr[36383] = -714681204;
assign addr[36384] = -732685372;
assign addr[36385] = -750631442;
assign addr[36386] = -768517992;
assign addr[36387] = -786343603;
assign addr[36388] = -804106861;
assign addr[36389] = -821806359;
assign addr[36390] = -839440693;
assign addr[36391] = -857008464;
assign addr[36392] = -874508280;
assign addr[36393] = -891938752;
assign addr[36394] = -909298500;
assign addr[36395] = -926586145;
assign addr[36396] = -943800318;
assign addr[36397] = -960939653;
assign addr[36398] = -978002791;
assign addr[36399] = -994988380;
assign addr[36400] = -1011895073;
assign addr[36401] = -1028721528;
assign addr[36402] = -1045466412;
assign addr[36403] = -1062128397;
assign addr[36404] = -1078706161;
assign addr[36405] = -1095198391;
assign addr[36406] = -1111603778;
assign addr[36407] = -1127921022;
assign addr[36408] = -1144148829;
assign addr[36409] = -1160285911;
assign addr[36410] = -1176330990;
assign addr[36411] = -1192282793;
assign addr[36412] = -1208140056;
assign addr[36413] = -1223901520;
assign addr[36414] = -1239565936;
assign addr[36415] = -1255132063;
assign addr[36416] = -1270598665;
assign addr[36417] = -1285964516;
assign addr[36418] = -1301228398;
assign addr[36419] = -1316389101;
assign addr[36420] = -1331445422;
assign addr[36421] = -1346396168;
assign addr[36422] = -1361240152;
assign addr[36423] = -1375976199;
assign addr[36424] = -1390603139;
assign addr[36425] = -1405119813;
assign addr[36426] = -1419525069;
assign addr[36427] = -1433817766;
assign addr[36428] = -1447996770;
assign addr[36429] = -1462060956;
assign addr[36430] = -1476009210;
assign addr[36431] = -1489840425;
assign addr[36432] = -1503553506;
assign addr[36433] = -1517147363;
assign addr[36434] = -1530620920;
assign addr[36435] = -1543973108;
assign addr[36436] = -1557202869;
assign addr[36437] = -1570309153;
assign addr[36438] = -1583290921;
assign addr[36439] = -1596147143;
assign addr[36440] = -1608876801;
assign addr[36441] = -1621478885;
assign addr[36442] = -1633952396;
assign addr[36443] = -1646296344;
assign addr[36444] = -1658509750;
assign addr[36445] = -1670591647;
assign addr[36446] = -1682541077;
assign addr[36447] = -1694357091;
assign addr[36448] = -1706038753;
assign addr[36449] = -1717585136;
assign addr[36450] = -1728995326;
assign addr[36451] = -1740268417;
assign addr[36452] = -1751403515;
assign addr[36453] = -1762399737;
assign addr[36454] = -1773256212;
assign addr[36455] = -1783972079;
assign addr[36456] = -1794546487;
assign addr[36457] = -1804978599;
assign addr[36458] = -1815267588;
assign addr[36459] = -1825412636;
assign addr[36460] = -1835412941;
assign addr[36461] = -1845267708;
assign addr[36462] = -1854976157;
assign addr[36463] = -1864537518;
assign addr[36464] = -1873951032;
assign addr[36465] = -1883215953;
assign addr[36466] = -1892331547;
assign addr[36467] = -1901297091;
assign addr[36468] = -1910111873;
assign addr[36469] = -1918775195;
assign addr[36470] = -1927286370;
assign addr[36471] = -1935644723;
assign addr[36472] = -1943849591;
assign addr[36473] = -1951900324;
assign addr[36474] = -1959796283;
assign addr[36475] = -1967536842;
assign addr[36476] = -1975121388;
assign addr[36477] = -1982549318;
assign addr[36478] = -1989820044;
assign addr[36479] = -1996932990;
assign addr[36480] = -2003887591;
assign addr[36481] = -2010683297;
assign addr[36482] = -2017319567;
assign addr[36483] = -2023795876;
assign addr[36484] = -2030111710;
assign addr[36485] = -2036266570;
assign addr[36486] = -2042259965;
assign addr[36487] = -2048091422;
assign addr[36488] = -2053760478;
assign addr[36489] = -2059266683;
assign addr[36490] = -2064609600;
assign addr[36491] = -2069788807;
assign addr[36492] = -2074803892;
assign addr[36493] = -2079654458;
assign addr[36494] = -2084340120;
assign addr[36495] = -2088860507;
assign addr[36496] = -2093215260;
assign addr[36497] = -2097404033;
assign addr[36498] = -2101426496;
assign addr[36499] = -2105282327;
assign addr[36500] = -2108971223;
assign addr[36501] = -2112492891;
assign addr[36502] = -2115847050;
assign addr[36503] = -2119033436;
assign addr[36504] = -2122051796;
assign addr[36505] = -2124901890;
assign addr[36506] = -2127583492;
assign addr[36507] = -2130096389;
assign addr[36508] = -2132440383;
assign addr[36509] = -2134615288;
assign addr[36510] = -2136620930;
assign addr[36511] = -2138457152;
assign addr[36512] = -2140123807;
assign addr[36513] = -2141620763;
assign addr[36514] = -2142947902;
assign addr[36515] = -2144105118;
assign addr[36516] = -2145092320;
assign addr[36517] = -2145909429;
assign addr[36518] = -2146556380;
assign addr[36519] = -2147033123;
assign addr[36520] = -2147339619;
assign addr[36521] = -2147475844;
assign addr[36522] = -2147441787;
assign addr[36523] = -2147237452;
assign addr[36524] = -2146862854;
assign addr[36525] = -2146318022;
assign addr[36526] = -2145603001;
assign addr[36527] = -2144717846;
assign addr[36528] = -2143662628;
assign addr[36529] = -2142437431;
assign addr[36530] = -2141042352;
assign addr[36531] = -2139477502;
assign addr[36532] = -2137743003;
assign addr[36533] = -2135838995;
assign addr[36534] = -2133765628;
assign addr[36535] = -2131523066;
assign addr[36536] = -2129111488;
assign addr[36537] = -2126531084;
assign addr[36538] = -2123782059;
assign addr[36539] = -2120864631;
assign addr[36540] = -2117779031;
assign addr[36541] = -2114525505;
assign addr[36542] = -2111104309;
assign addr[36543] = -2107515716;
assign addr[36544] = -2103760010;
assign addr[36545] = -2099837489;
assign addr[36546] = -2095748463;
assign addr[36547] = -2091493257;
assign addr[36548] = -2087072209;
assign addr[36549] = -2082485668;
assign addr[36550] = -2077733999;
assign addr[36551] = -2072817579;
assign addr[36552] = -2067736796;
assign addr[36553] = -2062492055;
assign addr[36554] = -2057083771;
assign addr[36555] = -2051512372;
assign addr[36556] = -2045778302;
assign addr[36557] = -2039882013;
assign addr[36558] = -2033823974;
assign addr[36559] = -2027604666;
assign addr[36560] = -2021224581;
assign addr[36561] = -2014684225;
assign addr[36562] = -2007984117;
assign addr[36563] = -2001124788;
assign addr[36564] = -1994106782;
assign addr[36565] = -1986930656;
assign addr[36566] = -1979596978;
assign addr[36567] = -1972106330;
assign addr[36568] = -1964459306;
assign addr[36569] = -1956656513;
assign addr[36570] = -1948698568;
assign addr[36571] = -1940586104;
assign addr[36572] = -1932319763;
assign addr[36573] = -1923900201;
assign addr[36574] = -1915328086;
assign addr[36575] = -1906604097;
assign addr[36576] = -1897728925;
assign addr[36577] = -1888703276;
assign addr[36578] = -1879527863;
assign addr[36579] = -1870203416;
assign addr[36580] = -1860730673;
assign addr[36581] = -1851110385;
assign addr[36582] = -1841343316;
assign addr[36583] = -1831430239;
assign addr[36584] = -1821371941;
assign addr[36585] = -1811169220;
assign addr[36586] = -1800822883;
assign addr[36587] = -1790333753;
assign addr[36588] = -1779702660;
assign addr[36589] = -1768930447;
assign addr[36590] = -1758017969;
assign addr[36591] = -1746966091;
assign addr[36592] = -1735775690;
assign addr[36593] = -1724447652;
assign addr[36594] = -1712982875;
assign addr[36595] = -1701382270;
assign addr[36596] = -1689646755;
assign addr[36597] = -1677777262;
assign addr[36598] = -1665774731;
assign addr[36599] = -1653640115;
assign addr[36600] = -1641374375;
assign addr[36601] = -1628978484;
assign addr[36602] = -1616453425;
assign addr[36603] = -1603800191;
assign addr[36604] = -1591019785;
assign addr[36605] = -1578113222;
assign addr[36606] = -1565081523;
assign addr[36607] = -1551925723;
assign addr[36608] = -1538646865;
assign addr[36609] = -1525246002;
assign addr[36610] = -1511724196;
assign addr[36611] = -1498082520;
assign addr[36612] = -1484322054;
assign addr[36613] = -1470443891;
assign addr[36614] = -1456449131;
assign addr[36615] = -1442338884;
assign addr[36616] = -1428114267;
assign addr[36617] = -1413776410;
assign addr[36618] = -1399326449;
assign addr[36619] = -1384765530;
assign addr[36620] = -1370094808;
assign addr[36621] = -1355315445;
assign addr[36622] = -1340428615;
assign addr[36623] = -1325435496;
assign addr[36624] = -1310337279;
assign addr[36625] = -1295135159;
assign addr[36626] = -1279830344;
assign addr[36627] = -1264424045;
assign addr[36628] = -1248917486;
assign addr[36629] = -1233311895;
assign addr[36630] = -1217608510;
assign addr[36631] = -1201808576;
assign addr[36632] = -1185913346;
assign addr[36633] = -1169924081;
assign addr[36634] = -1153842047;
assign addr[36635] = -1137668521;
assign addr[36636] = -1121404785;
assign addr[36637] = -1105052128;
assign addr[36638] = -1088611847;
assign addr[36639] = -1072085246;
assign addr[36640] = -1055473635;
assign addr[36641] = -1038778332;
assign addr[36642] = -1022000660;
assign addr[36643] = -1005141949;
assign addr[36644] = -988203537;
assign addr[36645] = -971186766;
assign addr[36646] = -954092986;
assign addr[36647] = -936923553;
assign addr[36648] = -919679827;
assign addr[36649] = -902363176;
assign addr[36650] = -884974973;
assign addr[36651] = -867516597;
assign addr[36652] = -849989433;
assign addr[36653] = -832394869;
assign addr[36654] = -814734301;
assign addr[36655] = -797009130;
assign addr[36656] = -779220762;
assign addr[36657] = -761370605;
assign addr[36658] = -743460077;
assign addr[36659] = -725490597;
assign addr[36660] = -707463589;
assign addr[36661] = -689380485;
assign addr[36662] = -671242716;
assign addr[36663] = -653051723;
assign addr[36664] = -634808946;
assign addr[36665] = -616515832;
assign addr[36666] = -598173833;
assign addr[36667] = -579784402;
assign addr[36668] = -561348998;
assign addr[36669] = -542869083;
assign addr[36670] = -524346121;
assign addr[36671] = -505781581;
assign addr[36672] = -487176937;
assign addr[36673] = -468533662;
assign addr[36674] = -449853235;
assign addr[36675] = -431137138;
assign addr[36676] = -412386854;
assign addr[36677] = -393603870;
assign addr[36678] = -374789676;
assign addr[36679] = -355945764;
assign addr[36680] = -337073627;
assign addr[36681] = -318174762;
assign addr[36682] = -299250668;
assign addr[36683] = -280302845;
assign addr[36684] = -261332796;
assign addr[36685] = -242342025;
assign addr[36686] = -223332037;
assign addr[36687] = -204304341;
assign addr[36688] = -185260444;
assign addr[36689] = -166201858;
assign addr[36690] = -147130093;
assign addr[36691] = -128046661;
assign addr[36692] = -108953076;
assign addr[36693] = -89850852;
assign addr[36694] = -70741503;
assign addr[36695] = -51626544;
assign addr[36696] = -32507492;
assign addr[36697] = -13385863;
assign addr[36698] = 5736829;
assign addr[36699] = 24859065;
assign addr[36700] = 43979330;
assign addr[36701] = 63096108;
assign addr[36702] = 82207882;
assign addr[36703] = 101313138;
assign addr[36704] = 120410361;
assign addr[36705] = 139498035;
assign addr[36706] = 158574649;
assign addr[36707] = 177638688;
assign addr[36708] = 196688642;
assign addr[36709] = 215722999;
assign addr[36710] = 234740251;
assign addr[36711] = 253738890;
assign addr[36712] = 272717408;
assign addr[36713] = 291674302;
assign addr[36714] = 310608068;
assign addr[36715] = 329517204;
assign addr[36716] = 348400212;
assign addr[36717] = 367255594;
assign addr[36718] = 386081854;
assign addr[36719] = 404877501;
assign addr[36720] = 423641043;
assign addr[36721] = 442370993;
assign addr[36722] = 461065866;
assign addr[36723] = 479724180;
assign addr[36724] = 498344454;
assign addr[36725] = 516925212;
assign addr[36726] = 535464981;
assign addr[36727] = 553962291;
assign addr[36728] = 572415676;
assign addr[36729] = 590823671;
assign addr[36730] = 609184818;
assign addr[36731] = 627497660;
assign addr[36732] = 645760745;
assign addr[36733] = 663972625;
assign addr[36734] = 682131857;
assign addr[36735] = 700236999;
assign addr[36736] = 718286617;
assign addr[36737] = 736279279;
assign addr[36738] = 754213559;
assign addr[36739] = 772088034;
assign addr[36740] = 789901288;
assign addr[36741] = 807651907;
assign addr[36742] = 825338484;
assign addr[36743] = 842959617;
assign addr[36744] = 860513908;
assign addr[36745] = 877999966;
assign addr[36746] = 895416404;
assign addr[36747] = 912761841;
assign addr[36748] = 930034901;
assign addr[36749] = 947234215;
assign addr[36750] = 964358420;
assign addr[36751] = 981406156;
assign addr[36752] = 998376073;
assign addr[36753] = 1015266825;
assign addr[36754] = 1032077073;
assign addr[36755] = 1048805483;
assign addr[36756] = 1065450729;
assign addr[36757] = 1082011492;
assign addr[36758] = 1098486458;
assign addr[36759] = 1114874320;
assign addr[36760] = 1131173780;
assign addr[36761] = 1147383544;
assign addr[36762] = 1163502328;
assign addr[36763] = 1179528853;
assign addr[36764] = 1195461849;
assign addr[36765] = 1211300053;
assign addr[36766] = 1227042207;
assign addr[36767] = 1242687064;
assign addr[36768] = 1258233384;
assign addr[36769] = 1273679934;
assign addr[36770] = 1289025489;
assign addr[36771] = 1304268832;
assign addr[36772] = 1319408754;
assign addr[36773] = 1334444055;
assign addr[36774] = 1349373543;
assign addr[36775] = 1364196034;
assign addr[36776] = 1378910353;
assign addr[36777] = 1393515332;
assign addr[36778] = 1408009814;
assign addr[36779] = 1422392650;
assign addr[36780] = 1436662698;
assign addr[36781] = 1450818828;
assign addr[36782] = 1464859917;
assign addr[36783] = 1478784851;
assign addr[36784] = 1492592527;
assign addr[36785] = 1506281850;
assign addr[36786] = 1519851733;
assign addr[36787] = 1533301101;
assign addr[36788] = 1546628888;
assign addr[36789] = 1559834037;
assign addr[36790] = 1572915501;
assign addr[36791] = 1585872242;
assign addr[36792] = 1598703233;
assign addr[36793] = 1611407456;
assign addr[36794] = 1623983905;
assign addr[36795] = 1636431582;
assign addr[36796] = 1648749499;
assign addr[36797] = 1660936681;
assign addr[36798] = 1672992161;
assign addr[36799] = 1684914983;
assign addr[36800] = 1696704201;
assign addr[36801] = 1708358881;
assign addr[36802] = 1719878099;
assign addr[36803] = 1731260941;
assign addr[36804] = 1742506504;
assign addr[36805] = 1753613897;
assign addr[36806] = 1764582240;
assign addr[36807] = 1775410662;
assign addr[36808] = 1786098304;
assign addr[36809] = 1796644320;
assign addr[36810] = 1807047873;
assign addr[36811] = 1817308138;
assign addr[36812] = 1827424302;
assign addr[36813] = 1837395562;
assign addr[36814] = 1847221128;
assign addr[36815] = 1856900221;
assign addr[36816] = 1866432072;
assign addr[36817] = 1875815927;
assign addr[36818] = 1885051042;
assign addr[36819] = 1894136683;
assign addr[36820] = 1903072131;
assign addr[36821] = 1911856677;
assign addr[36822] = 1920489624;
assign addr[36823] = 1928970288;
assign addr[36824] = 1937297997;
assign addr[36825] = 1945472089;
assign addr[36826] = 1953491918;
assign addr[36827] = 1961356847;
assign addr[36828] = 1969066252;
assign addr[36829] = 1976619522;
assign addr[36830] = 1984016058;
assign addr[36831] = 1991255274;
assign addr[36832] = 1998336596;
assign addr[36833] = 2005259462;
assign addr[36834] = 2012023322;
assign addr[36835] = 2018627642;
assign addr[36836] = 2025071897;
assign addr[36837] = 2031355576;
assign addr[36838] = 2037478181;
assign addr[36839] = 2043439226;
assign addr[36840] = 2049238240;
assign addr[36841] = 2054874761;
assign addr[36842] = 2060348343;
assign addr[36843] = 2065658552;
assign addr[36844] = 2070804967;
assign addr[36845] = 2075787180;
assign addr[36846] = 2080604795;
assign addr[36847] = 2085257431;
assign addr[36848] = 2089744719;
assign addr[36849] = 2094066304;
assign addr[36850] = 2098221841;
assign addr[36851] = 2102211002;
assign addr[36852] = 2106033471;
assign addr[36853] = 2109688944;
assign addr[36854] = 2113177132;
assign addr[36855] = 2116497758;
assign addr[36856] = 2119650558;
assign addr[36857] = 2122635283;
assign addr[36858] = 2125451696;
assign addr[36859] = 2128099574;
assign addr[36860] = 2130578706;
assign addr[36861] = 2132888897;
assign addr[36862] = 2135029962;
assign addr[36863] = 2137001733;
assign addr[36864] = 2138804053;
assign addr[36865] = 2140436778;
assign addr[36866] = 2141899780;
assign addr[36867] = 2143192942;
assign addr[36868] = 2144316162;
assign addr[36869] = 2145269351;
assign addr[36870] = 2146052433;
assign addr[36871] = 2146665347;
assign addr[36872] = 2147108043;
assign addr[36873] = 2147380486;
assign addr[36874] = 2147482655;
assign addr[36875] = 2147414542;
assign addr[36876] = 2147176152;
assign addr[36877] = 2146767505;
assign addr[36878] = 2146188631;
assign addr[36879] = 2145439578;
assign addr[36880] = 2144520405;
assign addr[36881] = 2143431184;
assign addr[36882] = 2142172003;
assign addr[36883] = 2140742960;
assign addr[36884] = 2139144169;
assign addr[36885] = 2137375758;
assign addr[36886] = 2135437865;
assign addr[36887] = 2133330646;
assign addr[36888] = 2131054266;
assign addr[36889] = 2128608907;
assign addr[36890] = 2125994762;
assign addr[36891] = 2123212038;
assign addr[36892] = 2120260957;
assign addr[36893] = 2117141752;
assign addr[36894] = 2113854671;
assign addr[36895] = 2110399974;
assign addr[36896] = 2106777935;
assign addr[36897] = 2102988841;
assign addr[36898] = 2099032994;
assign addr[36899] = 2094910706;
assign addr[36900] = 2090622304;
assign addr[36901] = 2086168128;
assign addr[36902] = 2081548533;
assign addr[36903] = 2076763883;
assign addr[36904] = 2071814558;
assign addr[36905] = 2066700952;
assign addr[36906] = 2061423468;
assign addr[36907] = 2055982526;
assign addr[36908] = 2050378558;
assign addr[36909] = 2044612007;
assign addr[36910] = 2038683330;
assign addr[36911] = 2032592999;
assign addr[36912] = 2026341495;
assign addr[36913] = 2019929315;
assign addr[36914] = 2013356967;
assign addr[36915] = 2006624971;
assign addr[36916] = 1999733863;
assign addr[36917] = 1992684188;
assign addr[36918] = 1985476506;
assign addr[36919] = 1978111387;
assign addr[36920] = 1970589416;
assign addr[36921] = 1962911189;
assign addr[36922] = 1955077316;
assign addr[36923] = 1947088417;
assign addr[36924] = 1938945125;
assign addr[36925] = 1930648088;
assign addr[36926] = 1922197961;
assign addr[36927] = 1913595416;
assign addr[36928] = 1904841135;
assign addr[36929] = 1895935811;
assign addr[36930] = 1886880151;
assign addr[36931] = 1877674873;
assign addr[36932] = 1868320707;
assign addr[36933] = 1858818395;
assign addr[36934] = 1849168689;
assign addr[36935] = 1839372356;
assign addr[36936] = 1829430172;
assign addr[36937] = 1819342925;
assign addr[36938] = 1809111415;
assign addr[36939] = 1798736454;
assign addr[36940] = 1788218865;
assign addr[36941] = 1777559480;
assign addr[36942] = 1766759146;
assign addr[36943] = 1755818718;
assign addr[36944] = 1744739065;
assign addr[36945] = 1733521064;
assign addr[36946] = 1722165606;
assign addr[36947] = 1710673591;
assign addr[36948] = 1699045930;
assign addr[36949] = 1687283545;
assign addr[36950] = 1675387369;
assign addr[36951] = 1663358344;
assign addr[36952] = 1651197426;
assign addr[36953] = 1638905577;
assign addr[36954] = 1626483774;
assign addr[36955] = 1613933000;
assign addr[36956] = 1601254251;
assign addr[36957] = 1588448533;
assign addr[36958] = 1575516860;
assign addr[36959] = 1562460258;
assign addr[36960] = 1549279763;
assign addr[36961] = 1535976419;
assign addr[36962] = 1522551282;
assign addr[36963] = 1509005416;
assign addr[36964] = 1495339895;
assign addr[36965] = 1481555802;
assign addr[36966] = 1467654232;
assign addr[36967] = 1453636285;
assign addr[36968] = 1439503074;
assign addr[36969] = 1425255719;
assign addr[36970] = 1410895350;
assign addr[36971] = 1396423105;
assign addr[36972] = 1381840133;
assign addr[36973] = 1367147589;
assign addr[36974] = 1352346639;
assign addr[36975] = 1337438456;
assign addr[36976] = 1322424222;
assign addr[36977] = 1307305128;
assign addr[36978] = 1292082373;
assign addr[36979] = 1276757164;
assign addr[36980] = 1261330715;
assign addr[36981] = 1245804251;
assign addr[36982] = 1230179002;
assign addr[36983] = 1214456207;
assign addr[36984] = 1198637114;
assign addr[36985] = 1182722976;
assign addr[36986] = 1166715055;
assign addr[36987] = 1150614620;
assign addr[36988] = 1134422949;
assign addr[36989] = 1118141326;
assign addr[36990] = 1101771040;
assign addr[36991] = 1085313391;
assign addr[36992] = 1068769683;
assign addr[36993] = 1052141228;
assign addr[36994] = 1035429345;
assign addr[36995] = 1018635358;
assign addr[36996] = 1001760600;
assign addr[36997] = 984806408;
assign addr[36998] = 967774128;
assign addr[36999] = 950665109;
assign addr[37000] = 933480707;
assign addr[37001] = 916222287;
assign addr[37002] = 898891215;
assign addr[37003] = 881488868;
assign addr[37004] = 864016623;
assign addr[37005] = 846475867;
assign addr[37006] = 828867991;
assign addr[37007] = 811194391;
assign addr[37008] = 793456467;
assign addr[37009] = 775655628;
assign addr[37010] = 757793284;
assign addr[37011] = 739870851;
assign addr[37012] = 721889752;
assign addr[37013] = 703851410;
assign addr[37014] = 685757258;
assign addr[37015] = 667608730;
assign addr[37016] = 649407264;
assign addr[37017] = 631154304;
assign addr[37018] = 612851297;
assign addr[37019] = 594499695;
assign addr[37020] = 576100953;
assign addr[37021] = 557656529;
assign addr[37022] = 539167887;
assign addr[37023] = 520636492;
assign addr[37024] = 502063814;
assign addr[37025] = 483451325;
assign addr[37026] = 464800501;
assign addr[37027] = 446112822;
assign addr[37028] = 427389768;
assign addr[37029] = 408632825;
assign addr[37030] = 389843480;
assign addr[37031] = 371023223;
assign addr[37032] = 352173546;
assign addr[37033] = 333295944;
assign addr[37034] = 314391913;
assign addr[37035] = 295462954;
assign addr[37036] = 276510565;
assign addr[37037] = 257536251;
assign addr[37038] = 238541516;
assign addr[37039] = 219527866;
assign addr[37040] = 200496809;
assign addr[37041] = 181449854;
assign addr[37042] = 162388511;
assign addr[37043] = 143314291;
assign addr[37044] = 124228708;
assign addr[37045] = 105133274;
assign addr[37046] = 86029503;
assign addr[37047] = 66918911;
assign addr[37048] = 47803013;
assign addr[37049] = 28683324;
assign addr[37050] = 9561361;
assign addr[37051] = -9561361;
assign addr[37052] = -28683324;
assign addr[37053] = -47803013;
assign addr[37054] = -66918911;
assign addr[37055] = -86029503;
assign addr[37056] = -105133274;
assign addr[37057] = -124228708;
assign addr[37058] = -143314291;
assign addr[37059] = -162388511;
assign addr[37060] = -181449854;
assign addr[37061] = -200496809;
assign addr[37062] = -219527866;
assign addr[37063] = -238541516;
assign addr[37064] = -257536251;
assign addr[37065] = -276510565;
assign addr[37066] = -295462954;
assign addr[37067] = -314391913;
assign addr[37068] = -333295944;
assign addr[37069] = -352173546;
assign addr[37070] = -371023223;
assign addr[37071] = -389843480;
assign addr[37072] = -408632825;
assign addr[37073] = -427389768;
assign addr[37074] = -446112822;
assign addr[37075] = -464800501;
assign addr[37076] = -483451325;
assign addr[37077] = -502063814;
assign addr[37078] = -520636492;
assign addr[37079] = -539167887;
assign addr[37080] = -557656529;
assign addr[37081] = -576100953;
assign addr[37082] = -594499695;
assign addr[37083] = -612851297;
assign addr[37084] = -631154304;
assign addr[37085] = -649407264;
assign addr[37086] = -667608730;
assign addr[37087] = -685757258;
assign addr[37088] = -703851410;
assign addr[37089] = -721889752;
assign addr[37090] = -739870851;
assign addr[37091] = -757793284;
assign addr[37092] = -775655628;
assign addr[37093] = -793456467;
assign addr[37094] = -811194391;
assign addr[37095] = -828867991;
assign addr[37096] = -846475867;
assign addr[37097] = -864016623;
assign addr[37098] = -881488868;
assign addr[37099] = -898891215;
assign addr[37100] = -916222287;
assign addr[37101] = -933480707;
assign addr[37102] = -950665109;
assign addr[37103] = -967774128;
assign addr[37104] = -984806408;
assign addr[37105] = -1001760600;
assign addr[37106] = -1018635358;
assign addr[37107] = -1035429345;
assign addr[37108] = -1052141228;
assign addr[37109] = -1068769683;
assign addr[37110] = -1085313391;
assign addr[37111] = -1101771040;
assign addr[37112] = -1118141326;
assign addr[37113] = -1134422949;
assign addr[37114] = -1150614620;
assign addr[37115] = -1166715055;
assign addr[37116] = -1182722976;
assign addr[37117] = -1198637114;
assign addr[37118] = -1214456207;
assign addr[37119] = -1230179002;
assign addr[37120] = -1245804251;
assign addr[37121] = -1261330715;
assign addr[37122] = -1276757164;
assign addr[37123] = -1292082373;
assign addr[37124] = -1307305128;
assign addr[37125] = -1322424222;
assign addr[37126] = -1337438456;
assign addr[37127] = -1352346639;
assign addr[37128] = -1367147589;
assign addr[37129] = -1381840133;
assign addr[37130] = -1396423105;
assign addr[37131] = -1410895350;
assign addr[37132] = -1425255719;
assign addr[37133] = -1439503074;
assign addr[37134] = -1453636285;
assign addr[37135] = -1467654232;
assign addr[37136] = -1481555802;
assign addr[37137] = -1495339895;
assign addr[37138] = -1509005416;
assign addr[37139] = -1522551282;
assign addr[37140] = -1535976419;
assign addr[37141] = -1549279763;
assign addr[37142] = -1562460258;
assign addr[37143] = -1575516860;
assign addr[37144] = -1588448533;
assign addr[37145] = -1601254251;
assign addr[37146] = -1613933000;
assign addr[37147] = -1626483774;
assign addr[37148] = -1638905577;
assign addr[37149] = -1651197426;
assign addr[37150] = -1663358344;
assign addr[37151] = -1675387369;
assign addr[37152] = -1687283545;
assign addr[37153] = -1699045930;
assign addr[37154] = -1710673591;
assign addr[37155] = -1722165606;
assign addr[37156] = -1733521064;
assign addr[37157] = -1744739065;
assign addr[37158] = -1755818718;
assign addr[37159] = -1766759146;
assign addr[37160] = -1777559480;
assign addr[37161] = -1788218865;
assign addr[37162] = -1798736454;
assign addr[37163] = -1809111415;
assign addr[37164] = -1819342925;
assign addr[37165] = -1829430172;
assign addr[37166] = -1839372356;
assign addr[37167] = -1849168689;
assign addr[37168] = -1858818395;
assign addr[37169] = -1868320707;
assign addr[37170] = -1877674873;
assign addr[37171] = -1886880151;
assign addr[37172] = -1895935811;
assign addr[37173] = -1904841135;
assign addr[37174] = -1913595416;
assign addr[37175] = -1922197961;
assign addr[37176] = -1930648088;
assign addr[37177] = -1938945125;
assign addr[37178] = -1947088417;
assign addr[37179] = -1955077316;
assign addr[37180] = -1962911189;
assign addr[37181] = -1970589416;
assign addr[37182] = -1978111387;
assign addr[37183] = -1985476506;
assign addr[37184] = -1992684188;
assign addr[37185] = -1999733863;
assign addr[37186] = -2006624971;
assign addr[37187] = -2013356967;
assign addr[37188] = -2019929315;
assign addr[37189] = -2026341495;
assign addr[37190] = -2032592999;
assign addr[37191] = -2038683330;
assign addr[37192] = -2044612007;
assign addr[37193] = -2050378558;
assign addr[37194] = -2055982526;
assign addr[37195] = -2061423468;
assign addr[37196] = -2066700952;
assign addr[37197] = -2071814558;
assign addr[37198] = -2076763883;
assign addr[37199] = -2081548533;
assign addr[37200] = -2086168128;
assign addr[37201] = -2090622304;
assign addr[37202] = -2094910706;
assign addr[37203] = -2099032994;
assign addr[37204] = -2102988841;
assign addr[37205] = -2106777935;
assign addr[37206] = -2110399974;
assign addr[37207] = -2113854671;
assign addr[37208] = -2117141752;
assign addr[37209] = -2120260957;
assign addr[37210] = -2123212038;
assign addr[37211] = -2125994762;
assign addr[37212] = -2128608907;
assign addr[37213] = -2131054266;
assign addr[37214] = -2133330646;
assign addr[37215] = -2135437865;
assign addr[37216] = -2137375758;
assign addr[37217] = -2139144169;
assign addr[37218] = -2140742960;
assign addr[37219] = -2142172003;
assign addr[37220] = -2143431184;
assign addr[37221] = -2144520405;
assign addr[37222] = -2145439578;
assign addr[37223] = -2146188631;
assign addr[37224] = -2146767505;
assign addr[37225] = -2147176152;
assign addr[37226] = -2147414542;
assign addr[37227] = -2147482655;
assign addr[37228] = -2147380486;
assign addr[37229] = -2147108043;
assign addr[37230] = -2146665347;
assign addr[37231] = -2146052433;
assign addr[37232] = -2145269351;
assign addr[37233] = -2144316162;
assign addr[37234] = -2143192942;
assign addr[37235] = -2141899780;
assign addr[37236] = -2140436778;
assign addr[37237] = -2138804053;
assign addr[37238] = -2137001733;
assign addr[37239] = -2135029962;
assign addr[37240] = -2132888897;
assign addr[37241] = -2130578706;
assign addr[37242] = -2128099574;
assign addr[37243] = -2125451696;
assign addr[37244] = -2122635283;
assign addr[37245] = -2119650558;
assign addr[37246] = -2116497758;
assign addr[37247] = -2113177132;
assign addr[37248] = -2109688944;
assign addr[37249] = -2106033471;
assign addr[37250] = -2102211002;
assign addr[37251] = -2098221841;
assign addr[37252] = -2094066304;
assign addr[37253] = -2089744719;
assign addr[37254] = -2085257431;
assign addr[37255] = -2080604795;
assign addr[37256] = -2075787180;
assign addr[37257] = -2070804967;
assign addr[37258] = -2065658552;
assign addr[37259] = -2060348343;
assign addr[37260] = -2054874761;
assign addr[37261] = -2049238240;
assign addr[37262] = -2043439226;
assign addr[37263] = -2037478181;
assign addr[37264] = -2031355576;
assign addr[37265] = -2025071897;
assign addr[37266] = -2018627642;
assign addr[37267] = -2012023322;
assign addr[37268] = -2005259462;
assign addr[37269] = -1998336596;
assign addr[37270] = -1991255274;
assign addr[37271] = -1984016058;
assign addr[37272] = -1976619522;
assign addr[37273] = -1969066252;
assign addr[37274] = -1961356847;
assign addr[37275] = -1953491918;
assign addr[37276] = -1945472089;
assign addr[37277] = -1937297997;
assign addr[37278] = -1928970288;
assign addr[37279] = -1920489624;
assign addr[37280] = -1911856677;
assign addr[37281] = -1903072131;
assign addr[37282] = -1894136683;
assign addr[37283] = -1885051042;
assign addr[37284] = -1875815927;
assign addr[37285] = -1866432072;
assign addr[37286] = -1856900221;
assign addr[37287] = -1847221128;
assign addr[37288] = -1837395562;
assign addr[37289] = -1827424302;
assign addr[37290] = -1817308138;
assign addr[37291] = -1807047873;
assign addr[37292] = -1796644320;
assign addr[37293] = -1786098304;
assign addr[37294] = -1775410662;
assign addr[37295] = -1764582240;
assign addr[37296] = -1753613897;
assign addr[37297] = -1742506504;
assign addr[37298] = -1731260941;
assign addr[37299] = -1719878099;
assign addr[37300] = -1708358881;
assign addr[37301] = -1696704201;
assign addr[37302] = -1684914983;
assign addr[37303] = -1672992161;
assign addr[37304] = -1660936681;
assign addr[37305] = -1648749499;
assign addr[37306] = -1636431582;
assign addr[37307] = -1623983905;
assign addr[37308] = -1611407456;
assign addr[37309] = -1598703233;
assign addr[37310] = -1585872242;
assign addr[37311] = -1572915501;
assign addr[37312] = -1559834037;
assign addr[37313] = -1546628888;
assign addr[37314] = -1533301101;
assign addr[37315] = -1519851733;
assign addr[37316] = -1506281850;
assign addr[37317] = -1492592527;
assign addr[37318] = -1478784851;
assign addr[37319] = -1464859917;
assign addr[37320] = -1450818828;
assign addr[37321] = -1436662698;
assign addr[37322] = -1422392650;
assign addr[37323] = -1408009814;
assign addr[37324] = -1393515332;
assign addr[37325] = -1378910353;
assign addr[37326] = -1364196034;
assign addr[37327] = -1349373543;
assign addr[37328] = -1334444055;
assign addr[37329] = -1319408754;
assign addr[37330] = -1304268832;
assign addr[37331] = -1289025489;
assign addr[37332] = -1273679934;
assign addr[37333] = -1258233384;
assign addr[37334] = -1242687064;
assign addr[37335] = -1227042207;
assign addr[37336] = -1211300053;
assign addr[37337] = -1195461849;
assign addr[37338] = -1179528853;
assign addr[37339] = -1163502328;
assign addr[37340] = -1147383544;
assign addr[37341] = -1131173780;
assign addr[37342] = -1114874320;
assign addr[37343] = -1098486458;
assign addr[37344] = -1082011492;
assign addr[37345] = -1065450729;
assign addr[37346] = -1048805483;
assign addr[37347] = -1032077073;
assign addr[37348] = -1015266825;
assign addr[37349] = -998376073;
assign addr[37350] = -981406156;
assign addr[37351] = -964358420;
assign addr[37352] = -947234215;
assign addr[37353] = -930034901;
assign addr[37354] = -912761841;
assign addr[37355] = -895416404;
assign addr[37356] = -877999966;
assign addr[37357] = -860513908;
assign addr[37358] = -842959617;
assign addr[37359] = -825338484;
assign addr[37360] = -807651907;
assign addr[37361] = -789901288;
assign addr[37362] = -772088034;
assign addr[37363] = -754213559;
assign addr[37364] = -736279279;
assign addr[37365] = -718286617;
assign addr[37366] = -700236999;
assign addr[37367] = -682131857;
assign addr[37368] = -663972625;
assign addr[37369] = -645760745;
assign addr[37370] = -627497660;
assign addr[37371] = -609184818;
assign addr[37372] = -590823671;
assign addr[37373] = -572415676;
assign addr[37374] = -553962291;
assign addr[37375] = -535464981;
assign addr[37376] = -516925212;
assign addr[37377] = -498344454;
assign addr[37378] = -479724180;
assign addr[37379] = -461065866;
assign addr[37380] = -442370993;
assign addr[37381] = -423641043;
assign addr[37382] = -404877501;
assign addr[37383] = -386081854;
assign addr[37384] = -367255594;
assign addr[37385] = -348400212;
assign addr[37386] = -329517204;
assign addr[37387] = -310608068;
assign addr[37388] = -291674302;
assign addr[37389] = -272717408;
assign addr[37390] = -253738890;
assign addr[37391] = -234740251;
assign addr[37392] = -215722999;
assign addr[37393] = -196688642;
assign addr[37394] = -177638688;
assign addr[37395] = -158574649;
assign addr[37396] = -139498035;
assign addr[37397] = -120410361;
assign addr[37398] = -101313138;
assign addr[37399] = -82207882;
assign addr[37400] = -63096108;
assign addr[37401] = -43979330;
assign addr[37402] = -24859065;
assign addr[37403] = -5736829;
assign addr[37404] = 13385863;
assign addr[37405] = 32507492;
assign addr[37406] = 51626544;
assign addr[37407] = 70741503;
assign addr[37408] = 89850852;
assign addr[37409] = 108953076;
assign addr[37410] = 128046661;
assign addr[37411] = 147130093;
assign addr[37412] = 166201858;
assign addr[37413] = 185260444;
assign addr[37414] = 204304341;
assign addr[37415] = 223332037;
assign addr[37416] = 242342025;
assign addr[37417] = 261332796;
assign addr[37418] = 280302845;
assign addr[37419] = 299250668;
assign addr[37420] = 318174762;
assign addr[37421] = 337073627;
assign addr[37422] = 355945764;
assign addr[37423] = 374789676;
assign addr[37424] = 393603870;
assign addr[37425] = 412386854;
assign addr[37426] = 431137138;
assign addr[37427] = 449853235;
assign addr[37428] = 468533662;
assign addr[37429] = 487176937;
assign addr[37430] = 505781581;
assign addr[37431] = 524346121;
assign addr[37432] = 542869083;
assign addr[37433] = 561348998;
assign addr[37434] = 579784402;
assign addr[37435] = 598173833;
assign addr[37436] = 616515832;
assign addr[37437] = 634808946;
assign addr[37438] = 653051723;
assign addr[37439] = 671242716;
assign addr[37440] = 689380485;
assign addr[37441] = 707463589;
assign addr[37442] = 725490597;
assign addr[37443] = 743460077;
assign addr[37444] = 761370605;
assign addr[37445] = 779220762;
assign addr[37446] = 797009130;
assign addr[37447] = 814734301;
assign addr[37448] = 832394869;
assign addr[37449] = 849989433;
assign addr[37450] = 867516597;
assign addr[37451] = 884974973;
assign addr[37452] = 902363176;
assign addr[37453] = 919679827;
assign addr[37454] = 936923553;
assign addr[37455] = 954092986;
assign addr[37456] = 971186766;
assign addr[37457] = 988203537;
assign addr[37458] = 1005141949;
assign addr[37459] = 1022000660;
assign addr[37460] = 1038778332;
assign addr[37461] = 1055473635;
assign addr[37462] = 1072085246;
assign addr[37463] = 1088611847;
assign addr[37464] = 1105052128;
assign addr[37465] = 1121404785;
assign addr[37466] = 1137668521;
assign addr[37467] = 1153842047;
assign addr[37468] = 1169924081;
assign addr[37469] = 1185913346;
assign addr[37470] = 1201808576;
assign addr[37471] = 1217608510;
assign addr[37472] = 1233311895;
assign addr[37473] = 1248917486;
assign addr[37474] = 1264424045;
assign addr[37475] = 1279830344;
assign addr[37476] = 1295135159;
assign addr[37477] = 1310337279;
assign addr[37478] = 1325435496;
assign addr[37479] = 1340428615;
assign addr[37480] = 1355315445;
assign addr[37481] = 1370094808;
assign addr[37482] = 1384765530;
assign addr[37483] = 1399326449;
assign addr[37484] = 1413776410;
assign addr[37485] = 1428114267;
assign addr[37486] = 1442338884;
assign addr[37487] = 1456449131;
assign addr[37488] = 1470443891;
assign addr[37489] = 1484322054;
assign addr[37490] = 1498082520;
assign addr[37491] = 1511724196;
assign addr[37492] = 1525246002;
assign addr[37493] = 1538646865;
assign addr[37494] = 1551925723;
assign addr[37495] = 1565081523;
assign addr[37496] = 1578113222;
assign addr[37497] = 1591019785;
assign addr[37498] = 1603800191;
assign addr[37499] = 1616453425;
assign addr[37500] = 1628978484;
assign addr[37501] = 1641374375;
assign addr[37502] = 1653640115;
assign addr[37503] = 1665774731;
assign addr[37504] = 1677777262;
assign addr[37505] = 1689646755;
assign addr[37506] = 1701382270;
assign addr[37507] = 1712982875;
assign addr[37508] = 1724447652;
assign addr[37509] = 1735775690;
assign addr[37510] = 1746966091;
assign addr[37511] = 1758017969;
assign addr[37512] = 1768930447;
assign addr[37513] = 1779702660;
assign addr[37514] = 1790333753;
assign addr[37515] = 1800822883;
assign addr[37516] = 1811169220;
assign addr[37517] = 1821371941;
assign addr[37518] = 1831430239;
assign addr[37519] = 1841343316;
assign addr[37520] = 1851110385;
assign addr[37521] = 1860730673;
assign addr[37522] = 1870203416;
assign addr[37523] = 1879527863;
assign addr[37524] = 1888703276;
assign addr[37525] = 1897728925;
assign addr[37526] = 1906604097;
assign addr[37527] = 1915328086;
assign addr[37528] = 1923900201;
assign addr[37529] = 1932319763;
assign addr[37530] = 1940586104;
assign addr[37531] = 1948698568;
assign addr[37532] = 1956656513;
assign addr[37533] = 1964459306;
assign addr[37534] = 1972106330;
assign addr[37535] = 1979596978;
assign addr[37536] = 1986930656;
assign addr[37537] = 1994106782;
assign addr[37538] = 2001124788;
assign addr[37539] = 2007984117;
assign addr[37540] = 2014684225;
assign addr[37541] = 2021224581;
assign addr[37542] = 2027604666;
assign addr[37543] = 2033823974;
assign addr[37544] = 2039882013;
assign addr[37545] = 2045778302;
assign addr[37546] = 2051512372;
assign addr[37547] = 2057083771;
assign addr[37548] = 2062492055;
assign addr[37549] = 2067736796;
assign addr[37550] = 2072817579;
assign addr[37551] = 2077733999;
assign addr[37552] = 2082485668;
assign addr[37553] = 2087072209;
assign addr[37554] = 2091493257;
assign addr[37555] = 2095748463;
assign addr[37556] = 2099837489;
assign addr[37557] = 2103760010;
assign addr[37558] = 2107515716;
assign addr[37559] = 2111104309;
assign addr[37560] = 2114525505;
assign addr[37561] = 2117779031;
assign addr[37562] = 2120864631;
assign addr[37563] = 2123782059;
assign addr[37564] = 2126531084;
assign addr[37565] = 2129111488;
assign addr[37566] = 2131523066;
assign addr[37567] = 2133765628;
assign addr[37568] = 2135838995;
assign addr[37569] = 2137743003;
assign addr[37570] = 2139477502;
assign addr[37571] = 2141042352;
assign addr[37572] = 2142437431;
assign addr[37573] = 2143662628;
assign addr[37574] = 2144717846;
assign addr[37575] = 2145603001;
assign addr[37576] = 2146318022;
assign addr[37577] = 2146862854;
assign addr[37578] = 2147237452;
assign addr[37579] = 2147441787;
assign addr[37580] = 2147475844;
assign addr[37581] = 2147339619;
assign addr[37582] = 2147033123;
assign addr[37583] = 2146556380;
assign addr[37584] = 2145909429;
assign addr[37585] = 2145092320;
assign addr[37586] = 2144105118;
assign addr[37587] = 2142947902;
assign addr[37588] = 2141620763;
assign addr[37589] = 2140123807;
assign addr[37590] = 2138457152;
assign addr[37591] = 2136620930;
assign addr[37592] = 2134615288;
assign addr[37593] = 2132440383;
assign addr[37594] = 2130096389;
assign addr[37595] = 2127583492;
assign addr[37596] = 2124901890;
assign addr[37597] = 2122051796;
assign addr[37598] = 2119033436;
assign addr[37599] = 2115847050;
assign addr[37600] = 2112492891;
assign addr[37601] = 2108971223;
assign addr[37602] = 2105282327;
assign addr[37603] = 2101426496;
assign addr[37604] = 2097404033;
assign addr[37605] = 2093215260;
assign addr[37606] = 2088860507;
assign addr[37607] = 2084340120;
assign addr[37608] = 2079654458;
assign addr[37609] = 2074803892;
assign addr[37610] = 2069788807;
assign addr[37611] = 2064609600;
assign addr[37612] = 2059266683;
assign addr[37613] = 2053760478;
assign addr[37614] = 2048091422;
assign addr[37615] = 2042259965;
assign addr[37616] = 2036266570;
assign addr[37617] = 2030111710;
assign addr[37618] = 2023795876;
assign addr[37619] = 2017319567;
assign addr[37620] = 2010683297;
assign addr[37621] = 2003887591;
assign addr[37622] = 1996932990;
assign addr[37623] = 1989820044;
assign addr[37624] = 1982549318;
assign addr[37625] = 1975121388;
assign addr[37626] = 1967536842;
assign addr[37627] = 1959796283;
assign addr[37628] = 1951900324;
assign addr[37629] = 1943849591;
assign addr[37630] = 1935644723;
assign addr[37631] = 1927286370;
assign addr[37632] = 1918775195;
assign addr[37633] = 1910111873;
assign addr[37634] = 1901297091;
assign addr[37635] = 1892331547;
assign addr[37636] = 1883215953;
assign addr[37637] = 1873951032;
assign addr[37638] = 1864537518;
assign addr[37639] = 1854976157;
assign addr[37640] = 1845267708;
assign addr[37641] = 1835412941;
assign addr[37642] = 1825412636;
assign addr[37643] = 1815267588;
assign addr[37644] = 1804978599;
assign addr[37645] = 1794546487;
assign addr[37646] = 1783972079;
assign addr[37647] = 1773256212;
assign addr[37648] = 1762399737;
assign addr[37649] = 1751403515;
assign addr[37650] = 1740268417;
assign addr[37651] = 1728995326;
assign addr[37652] = 1717585136;
assign addr[37653] = 1706038753;
assign addr[37654] = 1694357091;
assign addr[37655] = 1682541077;
assign addr[37656] = 1670591647;
assign addr[37657] = 1658509750;
assign addr[37658] = 1646296344;
assign addr[37659] = 1633952396;
assign addr[37660] = 1621478885;
assign addr[37661] = 1608876801;
assign addr[37662] = 1596147143;
assign addr[37663] = 1583290921;
assign addr[37664] = 1570309153;
assign addr[37665] = 1557202869;
assign addr[37666] = 1543973108;
assign addr[37667] = 1530620920;
assign addr[37668] = 1517147363;
assign addr[37669] = 1503553506;
assign addr[37670] = 1489840425;
assign addr[37671] = 1476009210;
assign addr[37672] = 1462060956;
assign addr[37673] = 1447996770;
assign addr[37674] = 1433817766;
assign addr[37675] = 1419525069;
assign addr[37676] = 1405119813;
assign addr[37677] = 1390603139;
assign addr[37678] = 1375976199;
assign addr[37679] = 1361240152;
assign addr[37680] = 1346396168;
assign addr[37681] = 1331445422;
assign addr[37682] = 1316389101;
assign addr[37683] = 1301228398;
assign addr[37684] = 1285964516;
assign addr[37685] = 1270598665;
assign addr[37686] = 1255132063;
assign addr[37687] = 1239565936;
assign addr[37688] = 1223901520;
assign addr[37689] = 1208140056;
assign addr[37690] = 1192282793;
assign addr[37691] = 1176330990;
assign addr[37692] = 1160285911;
assign addr[37693] = 1144148829;
assign addr[37694] = 1127921022;
assign addr[37695] = 1111603778;
assign addr[37696] = 1095198391;
assign addr[37697] = 1078706161;
assign addr[37698] = 1062128397;
assign addr[37699] = 1045466412;
assign addr[37700] = 1028721528;
assign addr[37701] = 1011895073;
assign addr[37702] = 994988380;
assign addr[37703] = 978002791;
assign addr[37704] = 960939653;
assign addr[37705] = 943800318;
assign addr[37706] = 926586145;
assign addr[37707] = 909298500;
assign addr[37708] = 891938752;
assign addr[37709] = 874508280;
assign addr[37710] = 857008464;
assign addr[37711] = 839440693;
assign addr[37712] = 821806359;
assign addr[37713] = 804106861;
assign addr[37714] = 786343603;
assign addr[37715] = 768517992;
assign addr[37716] = 750631442;
assign addr[37717] = 732685372;
assign addr[37718] = 714681204;
assign addr[37719] = 696620367;
assign addr[37720] = 678504291;
assign addr[37721] = 660334415;
assign addr[37722] = 642112178;
assign addr[37723] = 623839025;
assign addr[37724] = 605516406;
assign addr[37725] = 587145773;
assign addr[37726] = 568728583;
assign addr[37727] = 550266296;
assign addr[37728] = 531760377;
assign addr[37729] = 513212292;
assign addr[37730] = 494623513;
assign addr[37731] = 475995513;
assign addr[37732] = 457329769;
assign addr[37733] = 438627762;
assign addr[37734] = 419890975;
assign addr[37735] = 401120892;
assign addr[37736] = 382319004;
assign addr[37737] = 363486799;
assign addr[37738] = 344625773;
assign addr[37739] = 325737419;
assign addr[37740] = 306823237;
assign addr[37741] = 287884725;
assign addr[37742] = 268923386;
assign addr[37743] = 249940723;
assign addr[37744] = 230938242;
assign addr[37745] = 211917448;
assign addr[37746] = 192879850;
assign addr[37747] = 173826959;
assign addr[37748] = 154760284;
assign addr[37749] = 135681337;
assign addr[37750] = 116591632;
assign addr[37751] = 97492681;
assign addr[37752] = 78386000;
assign addr[37753] = 59273104;
assign addr[37754] = 40155507;
assign addr[37755] = 21034727;
assign addr[37756] = 1912278;
assign addr[37757] = -17210322;
assign addr[37758] = -36331557;
assign addr[37759] = -55449912;
assign addr[37760] = -74563870;
assign addr[37761] = -93671915;
assign addr[37762] = -112772533;
assign addr[37763] = -131864208;
assign addr[37764] = -150945428;
assign addr[37765] = -170014678;
assign addr[37766] = -189070447;
assign addr[37767] = -208111224;
assign addr[37768] = -227135500;
assign addr[37769] = -246141764;
assign addr[37770] = -265128512;
assign addr[37771] = -284094236;
assign addr[37772] = -303037433;
assign addr[37773] = -321956601;
assign addr[37774] = -340850240;
assign addr[37775] = -359716852;
assign addr[37776] = -378554940;
assign addr[37777] = -397363011;
assign addr[37778] = -416139574;
assign addr[37779] = -434883140;
assign addr[37780] = -453592221;
assign addr[37781] = -472265336;
assign addr[37782] = -490901003;
assign addr[37783] = -509497745;
assign addr[37784] = -528054086;
assign addr[37785] = -546568556;
assign addr[37786] = -565039687;
assign addr[37787] = -583466013;
assign addr[37788] = -601846074;
assign addr[37789] = -620178412;
assign addr[37790] = -638461574;
assign addr[37791] = -656694110;
assign addr[37792] = -674874574;
assign addr[37793] = -693001525;
assign addr[37794] = -711073524;
assign addr[37795] = -729089140;
assign addr[37796] = -747046944;
assign addr[37797] = -764945512;
assign addr[37798] = -782783424;
assign addr[37799] = -800559266;
assign addr[37800] = -818271628;
assign addr[37801] = -835919107;
assign addr[37802] = -853500302;
assign addr[37803] = -871013820;
assign addr[37804] = -888458272;
assign addr[37805] = -905832274;
assign addr[37806] = -923134450;
assign addr[37807] = -940363427;
assign addr[37808] = -957517838;
assign addr[37809] = -974596324;
assign addr[37810] = -991597531;
assign addr[37811] = -1008520110;
assign addr[37812] = -1025362720;
assign addr[37813] = -1042124025;
assign addr[37814] = -1058802695;
assign addr[37815] = -1075397409;
assign addr[37816] = -1091906851;
assign addr[37817] = -1108329711;
assign addr[37818] = -1124664687;
assign addr[37819] = -1140910484;
assign addr[37820] = -1157065814;
assign addr[37821] = -1173129396;
assign addr[37822] = -1189099956;
assign addr[37823] = -1204976227;
assign addr[37824] = -1220756951;
assign addr[37825] = -1236440877;
assign addr[37826] = -1252026760;
assign addr[37827] = -1267513365;
assign addr[37828] = -1282899464;
assign addr[37829] = -1298183838;
assign addr[37830] = -1313365273;
assign addr[37831] = -1328442566;
assign addr[37832] = -1343414522;
assign addr[37833] = -1358279953;
assign addr[37834] = -1373037681;
assign addr[37835] = -1387686535;
assign addr[37836] = -1402225355;
assign addr[37837] = -1416652986;
assign addr[37838] = -1430968286;
assign addr[37839] = -1445170118;
assign addr[37840] = -1459257358;
assign addr[37841] = -1473228887;
assign addr[37842] = -1487083598;
assign addr[37843] = -1500820393;
assign addr[37844] = -1514438181;
assign addr[37845] = -1527935884;
assign addr[37846] = -1541312431;
assign addr[37847] = -1554566762;
assign addr[37848] = -1567697824;
assign addr[37849] = -1580704578;
assign addr[37850] = -1593585992;
assign addr[37851] = -1606341043;
assign addr[37852] = -1618968722;
assign addr[37853] = -1631468027;
assign addr[37854] = -1643837966;
assign addr[37855] = -1656077559;
assign addr[37856] = -1668185835;
assign addr[37857] = -1680161834;
assign addr[37858] = -1692004606;
assign addr[37859] = -1703713213;
assign addr[37860] = -1715286726;
assign addr[37861] = -1726724227;
assign addr[37862] = -1738024810;
assign addr[37863] = -1749187577;
assign addr[37864] = -1760211645;
assign addr[37865] = -1771096139;
assign addr[37866] = -1781840195;
assign addr[37867] = -1792442963;
assign addr[37868] = -1802903601;
assign addr[37869] = -1813221279;
assign addr[37870] = -1823395180;
assign addr[37871] = -1833424497;
assign addr[37872] = -1843308435;
assign addr[37873] = -1853046210;
assign addr[37874] = -1862637049;
assign addr[37875] = -1872080193;
assign addr[37876] = -1881374892;
assign addr[37877] = -1890520410;
assign addr[37878] = -1899516021;
assign addr[37879] = -1908361011;
assign addr[37880] = -1917054681;
assign addr[37881] = -1925596340;
assign addr[37882] = -1933985310;
assign addr[37883] = -1942220928;
assign addr[37884] = -1950302539;
assign addr[37885] = -1958229503;
assign addr[37886] = -1966001192;
assign addr[37887] = -1973616989;
assign addr[37888] = -1981076290;
assign addr[37889] = -1988378503;
assign addr[37890] = -1995523051;
assign addr[37891] = -2002509365;
assign addr[37892] = -2009336893;
assign addr[37893] = -2016005093;
assign addr[37894] = -2022513436;
assign addr[37895] = -2028861406;
assign addr[37896] = -2035048499;
assign addr[37897] = -2041074226;
assign addr[37898] = -2046938108;
assign addr[37899] = -2052639680;
assign addr[37900] = -2058178491;
assign addr[37901] = -2063554100;
assign addr[37902] = -2068766083;
assign addr[37903] = -2073814024;
assign addr[37904] = -2078697525;
assign addr[37905] = -2083416198;
assign addr[37906] = -2087969669;
assign addr[37907] = -2092357577;
assign addr[37908] = -2096579573;
assign addr[37909] = -2100635323;
assign addr[37910] = -2104524506;
assign addr[37911] = -2108246813;
assign addr[37912] = -2111801949;
assign addr[37913] = -2115189632;
assign addr[37914] = -2118409593;
assign addr[37915] = -2121461578;
assign addr[37916] = -2124345343;
assign addr[37917] = -2127060661;
assign addr[37918] = -2129607316;
assign addr[37919] = -2131985106;
assign addr[37920] = -2134193842;
assign addr[37921] = -2136233350;
assign addr[37922] = -2138103468;
assign addr[37923] = -2139804048;
assign addr[37924] = -2141334954;
assign addr[37925] = -2142696065;
assign addr[37926] = -2143887273;
assign addr[37927] = -2144908484;
assign addr[37928] = -2145759618;
assign addr[37929] = -2146440605;
assign addr[37930] = -2146951393;
assign addr[37931] = -2147291941;
assign addr[37932] = -2147462221;
assign addr[37933] = -2147462221;
assign addr[37934] = -2147291941;
assign addr[37935] = -2146951393;
assign addr[37936] = -2146440605;
assign addr[37937] = -2145759618;
assign addr[37938] = -2144908484;
assign addr[37939] = -2143887273;
assign addr[37940] = -2142696065;
assign addr[37941] = -2141334954;
assign addr[37942] = -2139804048;
assign addr[37943] = -2138103468;
assign addr[37944] = -2136233350;
assign addr[37945] = -2134193842;
assign addr[37946] = -2131985106;
assign addr[37947] = -2129607316;
assign addr[37948] = -2127060661;
assign addr[37949] = -2124345343;
assign addr[37950] = -2121461578;
assign addr[37951] = -2118409593;
assign addr[37952] = -2115189632;
assign addr[37953] = -2111801949;
assign addr[37954] = -2108246813;
assign addr[37955] = -2104524506;
assign addr[37956] = -2100635323;
assign addr[37957] = -2096579573;
assign addr[37958] = -2092357577;
assign addr[37959] = -2087969669;
assign addr[37960] = -2083416198;
assign addr[37961] = -2078697525;
assign addr[37962] = -2073814024;
assign addr[37963] = -2068766083;
assign addr[37964] = -2063554100;
assign addr[37965] = -2058178491;
assign addr[37966] = -2052639680;
assign addr[37967] = -2046938108;
assign addr[37968] = -2041074226;
assign addr[37969] = -2035048499;
assign addr[37970] = -2028861406;
assign addr[37971] = -2022513436;
assign addr[37972] = -2016005093;
assign addr[37973] = -2009336893;
assign addr[37974] = -2002509365;
assign addr[37975] = -1995523051;
assign addr[37976] = -1988378503;
assign addr[37977] = -1981076290;
assign addr[37978] = -1973616989;
assign addr[37979] = -1966001192;
assign addr[37980] = -1958229503;
assign addr[37981] = -1950302539;
assign addr[37982] = -1942220928;
assign addr[37983] = -1933985310;
assign addr[37984] = -1925596340;
assign addr[37985] = -1917054681;
assign addr[37986] = -1908361011;
assign addr[37987] = -1899516021;
assign addr[37988] = -1890520410;
assign addr[37989] = -1881374892;
assign addr[37990] = -1872080193;
assign addr[37991] = -1862637049;
assign addr[37992] = -1853046210;
assign addr[37993] = -1843308435;
assign addr[37994] = -1833424497;
assign addr[37995] = -1823395180;
assign addr[37996] = -1813221279;
assign addr[37997] = -1802903601;
assign addr[37998] = -1792442963;
assign addr[37999] = -1781840195;
assign addr[38000] = -1771096139;
assign addr[38001] = -1760211645;
assign addr[38002] = -1749187577;
assign addr[38003] = -1738024810;
assign addr[38004] = -1726724227;
assign addr[38005] = -1715286726;
assign addr[38006] = -1703713213;
assign addr[38007] = -1692004606;
assign addr[38008] = -1680161834;
assign addr[38009] = -1668185835;
assign addr[38010] = -1656077559;
assign addr[38011] = -1643837966;
assign addr[38012] = -1631468027;
assign addr[38013] = -1618968722;
assign addr[38014] = -1606341043;
assign addr[38015] = -1593585992;
assign addr[38016] = -1580704578;
assign addr[38017] = -1567697824;
assign addr[38018] = -1554566762;
assign addr[38019] = -1541312431;
assign addr[38020] = -1527935884;
assign addr[38021] = -1514438181;
assign addr[38022] = -1500820393;
assign addr[38023] = -1487083598;
assign addr[38024] = -1473228887;
assign addr[38025] = -1459257358;
assign addr[38026] = -1445170118;
assign addr[38027] = -1430968286;
assign addr[38028] = -1416652986;
assign addr[38029] = -1402225355;
assign addr[38030] = -1387686535;
assign addr[38031] = -1373037681;
assign addr[38032] = -1358279953;
assign addr[38033] = -1343414522;
assign addr[38034] = -1328442566;
assign addr[38035] = -1313365273;
assign addr[38036] = -1298183838;
assign addr[38037] = -1282899464;
assign addr[38038] = -1267513365;
assign addr[38039] = -1252026760;
assign addr[38040] = -1236440877;
assign addr[38041] = -1220756951;
assign addr[38042] = -1204976227;
assign addr[38043] = -1189099956;
assign addr[38044] = -1173129396;
assign addr[38045] = -1157065814;
assign addr[38046] = -1140910484;
assign addr[38047] = -1124664687;
assign addr[38048] = -1108329711;
assign addr[38049] = -1091906851;
assign addr[38050] = -1075397409;
assign addr[38051] = -1058802695;
assign addr[38052] = -1042124025;
assign addr[38053] = -1025362720;
assign addr[38054] = -1008520110;
assign addr[38055] = -991597531;
assign addr[38056] = -974596324;
assign addr[38057] = -957517838;
assign addr[38058] = -940363427;
assign addr[38059] = -923134450;
assign addr[38060] = -905832274;
assign addr[38061] = -888458272;
assign addr[38062] = -871013820;
assign addr[38063] = -853500302;
assign addr[38064] = -835919107;
assign addr[38065] = -818271628;
assign addr[38066] = -800559266;
assign addr[38067] = -782783424;
assign addr[38068] = -764945512;
assign addr[38069] = -747046944;
assign addr[38070] = -729089140;
assign addr[38071] = -711073525;
assign addr[38072] = -693001525;
assign addr[38073] = -674874574;
assign addr[38074] = -656694110;
assign addr[38075] = -638461574;
assign addr[38076] = -620178412;
assign addr[38077] = -601846074;
assign addr[38078] = -583466013;
assign addr[38079] = -565039687;
assign addr[38080] = -546568556;
assign addr[38081] = -528054086;
assign addr[38082] = -509497745;
assign addr[38083] = -490901003;
assign addr[38084] = -472265336;
assign addr[38085] = -453592221;
assign addr[38086] = -434883140;
assign addr[38087] = -416139574;
assign addr[38088] = -397363011;
assign addr[38089] = -378554940;
assign addr[38090] = -359716852;
assign addr[38091] = -340850240;
assign addr[38092] = -321956601;
assign addr[38093] = -303037433;
assign addr[38094] = -284094236;
assign addr[38095] = -265128512;
assign addr[38096] = -246141764;
assign addr[38097] = -227135500;
assign addr[38098] = -208111224;
assign addr[38099] = -189070447;
assign addr[38100] = -170014678;
assign addr[38101] = -150945428;
assign addr[38102] = -131864208;
assign addr[38103] = -112772533;
assign addr[38104] = -93671915;
assign addr[38105] = -74563870;
assign addr[38106] = -55449912;
assign addr[38107] = -36331557;
assign addr[38108] = -17210322;
assign addr[38109] = 1912278;
assign addr[38110] = 21034727;
assign addr[38111] = 40155507;
assign addr[38112] = 59273104;
assign addr[38113] = 78386000;
assign addr[38114] = 97492681;
assign addr[38115] = 116591632;
assign addr[38116] = 135681337;
assign addr[38117] = 154760284;
assign addr[38118] = 173826959;
assign addr[38119] = 192879850;
assign addr[38120] = 211917448;
assign addr[38121] = 230938242;
assign addr[38122] = 249940723;
assign addr[38123] = 268923386;
assign addr[38124] = 287884725;
assign addr[38125] = 306823237;
assign addr[38126] = 325737419;
assign addr[38127] = 344625773;
assign addr[38128] = 363486799;
assign addr[38129] = 382319004;
assign addr[38130] = 401120892;
assign addr[38131] = 419890975;
assign addr[38132] = 438627762;
assign addr[38133] = 457329769;
assign addr[38134] = 475995513;
assign addr[38135] = 494623513;
assign addr[38136] = 513212292;
assign addr[38137] = 531760377;
assign addr[38138] = 550266296;
assign addr[38139] = 568728583;
assign addr[38140] = 587145773;
assign addr[38141] = 605516406;
assign addr[38142] = 623839025;
assign addr[38143] = 642112178;
assign addr[38144] = 660334415;
assign addr[38145] = 678504291;
assign addr[38146] = 696620367;
assign addr[38147] = 714681204;
assign addr[38148] = 732685372;
assign addr[38149] = 750631442;
assign addr[38150] = 768517992;
assign addr[38151] = 786343603;
assign addr[38152] = 804106861;
assign addr[38153] = 821806359;
assign addr[38154] = 839440693;
assign addr[38155] = 857008464;
assign addr[38156] = 874508280;
assign addr[38157] = 891938752;
assign addr[38158] = 909298500;
assign addr[38159] = 926586145;
assign addr[38160] = 943800318;
assign addr[38161] = 960939653;
assign addr[38162] = 978002791;
assign addr[38163] = 994988380;
assign addr[38164] = 1011895073;
assign addr[38165] = 1028721528;
assign addr[38166] = 1045466412;
assign addr[38167] = 1062128397;
assign addr[38168] = 1078706161;
assign addr[38169] = 1095198391;
assign addr[38170] = 1111603778;
assign addr[38171] = 1127921022;
assign addr[38172] = 1144148829;
assign addr[38173] = 1160285911;
assign addr[38174] = 1176330990;
assign addr[38175] = 1192282793;
assign addr[38176] = 1208140056;
assign addr[38177] = 1223901520;
assign addr[38178] = 1239565936;
assign addr[38179] = 1255132063;
assign addr[38180] = 1270598665;
assign addr[38181] = 1285964516;
assign addr[38182] = 1301228398;
assign addr[38183] = 1316389101;
assign addr[38184] = 1331445422;
assign addr[38185] = 1346396168;
assign addr[38186] = 1361240152;
assign addr[38187] = 1375976199;
assign addr[38188] = 1390603139;
assign addr[38189] = 1405119813;
assign addr[38190] = 1419525069;
assign addr[38191] = 1433817766;
assign addr[38192] = 1447996770;
assign addr[38193] = 1462060956;
assign addr[38194] = 1476009210;
assign addr[38195] = 1489840425;
assign addr[38196] = 1503553506;
assign addr[38197] = 1517147363;
assign addr[38198] = 1530620920;
assign addr[38199] = 1543973108;
assign addr[38200] = 1557202869;
assign addr[38201] = 1570309153;
assign addr[38202] = 1583290921;
assign addr[38203] = 1596147143;
assign addr[38204] = 1608876801;
assign addr[38205] = 1621478885;
assign addr[38206] = 1633952396;
assign addr[38207] = 1646296344;
assign addr[38208] = 1658509750;
assign addr[38209] = 1670591647;
assign addr[38210] = 1682541077;
assign addr[38211] = 1694357091;
assign addr[38212] = 1706038753;
assign addr[38213] = 1717585136;
assign addr[38214] = 1728995326;
assign addr[38215] = 1740268417;
assign addr[38216] = 1751403515;
assign addr[38217] = 1762399737;
assign addr[38218] = 1773256212;
assign addr[38219] = 1783972079;
assign addr[38220] = 1794546487;
assign addr[38221] = 1804978599;
assign addr[38222] = 1815267588;
assign addr[38223] = 1825412636;
assign addr[38224] = 1835412941;
assign addr[38225] = 1845267708;
assign addr[38226] = 1854976157;
assign addr[38227] = 1864537518;
assign addr[38228] = 1873951032;
assign addr[38229] = 1883215953;
assign addr[38230] = 1892331547;
assign addr[38231] = 1901297091;
assign addr[38232] = 1910111873;
assign addr[38233] = 1918775195;
assign addr[38234] = 1927286370;
assign addr[38235] = 1935644723;
assign addr[38236] = 1943849591;
assign addr[38237] = 1951900324;
assign addr[38238] = 1959796283;
assign addr[38239] = 1967536842;
assign addr[38240] = 1975121388;
assign addr[38241] = 1982549318;
assign addr[38242] = 1989820044;
assign addr[38243] = 1996932990;
assign addr[38244] = 2003887591;
assign addr[38245] = 2010683297;
assign addr[38246] = 2017319567;
assign addr[38247] = 2023795876;
assign addr[38248] = 2030111710;
assign addr[38249] = 2036266570;
assign addr[38250] = 2042259965;
assign addr[38251] = 2048091422;
assign addr[38252] = 2053760478;
assign addr[38253] = 2059266683;
assign addr[38254] = 2064609600;
assign addr[38255] = 2069788807;
assign addr[38256] = 2074803892;
assign addr[38257] = 2079654458;
assign addr[38258] = 2084340120;
assign addr[38259] = 2088860507;
assign addr[38260] = 2093215260;
assign addr[38261] = 2097404033;
assign addr[38262] = 2101426496;
assign addr[38263] = 2105282327;
assign addr[38264] = 2108971223;
assign addr[38265] = 2112492891;
assign addr[38266] = 2115847050;
assign addr[38267] = 2119033436;
assign addr[38268] = 2122051796;
assign addr[38269] = 2124901890;
assign addr[38270] = 2127583492;
assign addr[38271] = 2130096389;
assign addr[38272] = 2132440383;
assign addr[38273] = 2134615288;
assign addr[38274] = 2136620930;
assign addr[38275] = 2138457152;
assign addr[38276] = 2140123807;
assign addr[38277] = 2141620763;
assign addr[38278] = 2142947902;
assign addr[38279] = 2144105118;
assign addr[38280] = 2145092320;
assign addr[38281] = 2145909429;
assign addr[38282] = 2146556380;
assign addr[38283] = 2147033123;
assign addr[38284] = 2147339619;
assign addr[38285] = 2147475844;
assign addr[38286] = 2147441787;
assign addr[38287] = 2147237452;
assign addr[38288] = 2146862854;
assign addr[38289] = 2146318022;
assign addr[38290] = 2145603001;
assign addr[38291] = 2144717846;
assign addr[38292] = 2143662628;
assign addr[38293] = 2142437431;
assign addr[38294] = 2141042352;
assign addr[38295] = 2139477502;
assign addr[38296] = 2137743003;
assign addr[38297] = 2135838995;
assign addr[38298] = 2133765628;
assign addr[38299] = 2131523066;
assign addr[38300] = 2129111488;
assign addr[38301] = 2126531084;
assign addr[38302] = 2123782059;
assign addr[38303] = 2120864631;
assign addr[38304] = 2117779031;
assign addr[38305] = 2114525505;
assign addr[38306] = 2111104309;
assign addr[38307] = 2107515716;
assign addr[38308] = 2103760010;
assign addr[38309] = 2099837489;
assign addr[38310] = 2095748463;
assign addr[38311] = 2091493257;
assign addr[38312] = 2087072209;
assign addr[38313] = 2082485668;
assign addr[38314] = 2077733999;
assign addr[38315] = 2072817579;
assign addr[38316] = 2067736796;
assign addr[38317] = 2062492055;
assign addr[38318] = 2057083771;
assign addr[38319] = 2051512372;
assign addr[38320] = 2045778302;
assign addr[38321] = 2039882013;
assign addr[38322] = 2033823974;
assign addr[38323] = 2027604666;
assign addr[38324] = 2021224581;
assign addr[38325] = 2014684225;
assign addr[38326] = 2007984117;
assign addr[38327] = 2001124788;
assign addr[38328] = 1994106782;
assign addr[38329] = 1986930656;
assign addr[38330] = 1979596978;
assign addr[38331] = 1972106330;
assign addr[38332] = 1964459306;
assign addr[38333] = 1956656513;
assign addr[38334] = 1948698568;
assign addr[38335] = 1940586104;
assign addr[38336] = 1932319763;
assign addr[38337] = 1923900201;
assign addr[38338] = 1915328086;
assign addr[38339] = 1906604097;
assign addr[38340] = 1897728925;
assign addr[38341] = 1888703276;
assign addr[38342] = 1879527863;
assign addr[38343] = 1870203416;
assign addr[38344] = 1860730673;
assign addr[38345] = 1851110385;
assign addr[38346] = 1841343316;
assign addr[38347] = 1831430239;
assign addr[38348] = 1821371941;
assign addr[38349] = 1811169220;
assign addr[38350] = 1800822883;
assign addr[38351] = 1790333753;
assign addr[38352] = 1779702660;
assign addr[38353] = 1768930447;
assign addr[38354] = 1758017969;
assign addr[38355] = 1746966091;
assign addr[38356] = 1735775690;
assign addr[38357] = 1724447652;
assign addr[38358] = 1712982875;
assign addr[38359] = 1701382270;
assign addr[38360] = 1689646755;
assign addr[38361] = 1677777262;
assign addr[38362] = 1665774731;
assign addr[38363] = 1653640115;
assign addr[38364] = 1641374375;
assign addr[38365] = 1628978484;
assign addr[38366] = 1616453425;
assign addr[38367] = 1603800191;
assign addr[38368] = 1591019785;
assign addr[38369] = 1578113222;
assign addr[38370] = 1565081523;
assign addr[38371] = 1551925723;
assign addr[38372] = 1538646865;
assign addr[38373] = 1525246002;
assign addr[38374] = 1511724196;
assign addr[38375] = 1498082520;
assign addr[38376] = 1484322054;
assign addr[38377] = 1470443891;
assign addr[38378] = 1456449131;
assign addr[38379] = 1442338884;
assign addr[38380] = 1428114267;
assign addr[38381] = 1413776410;
assign addr[38382] = 1399326449;
assign addr[38383] = 1384765530;
assign addr[38384] = 1370094808;
assign addr[38385] = 1355315445;
assign addr[38386] = 1340428615;
assign addr[38387] = 1325435496;
assign addr[38388] = 1310337279;
assign addr[38389] = 1295135159;
assign addr[38390] = 1279830344;
assign addr[38391] = 1264424045;
assign addr[38392] = 1248917486;
assign addr[38393] = 1233311895;
assign addr[38394] = 1217608510;
assign addr[38395] = 1201808576;
assign addr[38396] = 1185913346;
assign addr[38397] = 1169924081;
assign addr[38398] = 1153842047;
assign addr[38399] = 1137668521;
assign addr[38400] = 1121404785;
assign addr[38401] = 1105052128;
assign addr[38402] = 1088611847;
assign addr[38403] = 1072085246;
assign addr[38404] = 1055473635;
assign addr[38405] = 1038778332;
assign addr[38406] = 1022000660;
assign addr[38407] = 1005141949;
assign addr[38408] = 988203537;
assign addr[38409] = 971186766;
assign addr[38410] = 954092986;
assign addr[38411] = 936923553;
assign addr[38412] = 919679827;
assign addr[38413] = 902363176;
assign addr[38414] = 884974973;
assign addr[38415] = 867516597;
assign addr[38416] = 849989433;
assign addr[38417] = 832394869;
assign addr[38418] = 814734301;
assign addr[38419] = 797009130;
assign addr[38420] = 779220762;
assign addr[38421] = 761370605;
assign addr[38422] = 743460077;
assign addr[38423] = 725490597;
assign addr[38424] = 707463589;
assign addr[38425] = 689380485;
assign addr[38426] = 671242716;
assign addr[38427] = 653051723;
assign addr[38428] = 634808946;
assign addr[38429] = 616515832;
assign addr[38430] = 598173833;
assign addr[38431] = 579784402;
assign addr[38432] = 561348998;
assign addr[38433] = 542869083;
assign addr[38434] = 524346121;
assign addr[38435] = 505781581;
assign addr[38436] = 487176937;
assign addr[38437] = 468533662;
assign addr[38438] = 449853235;
assign addr[38439] = 431137138;
assign addr[38440] = 412386854;
assign addr[38441] = 393603870;
assign addr[38442] = 374789676;
assign addr[38443] = 355945764;
assign addr[38444] = 337073627;
assign addr[38445] = 318174762;
assign addr[38446] = 299250668;
assign addr[38447] = 280302845;
assign addr[38448] = 261332796;
assign addr[38449] = 242342025;
assign addr[38450] = 223332037;
assign addr[38451] = 204304341;
assign addr[38452] = 185260444;
assign addr[38453] = 166201858;
assign addr[38454] = 147130093;
assign addr[38455] = 128046661;
assign addr[38456] = 108953076;
assign addr[38457] = 89850852;
assign addr[38458] = 70741503;
assign addr[38459] = 51626544;
assign addr[38460] = 32507492;
assign addr[38461] = 13385863;
assign addr[38462] = -5736829;
assign addr[38463] = -24859065;
assign addr[38464] = -43979330;
assign addr[38465] = -63096108;
assign addr[38466] = -82207882;
assign addr[38467] = -101313138;
assign addr[38468] = -120410361;
assign addr[38469] = -139498035;
assign addr[38470] = -158574649;
assign addr[38471] = -177638688;
assign addr[38472] = -196688642;
assign addr[38473] = -215722999;
assign addr[38474] = -234740251;
assign addr[38475] = -253738890;
assign addr[38476] = -272717408;
assign addr[38477] = -291674302;
assign addr[38478] = -310608068;
assign addr[38479] = -329517204;
assign addr[38480] = -348400212;
assign addr[38481] = -367255594;
assign addr[38482] = -386081854;
assign addr[38483] = -404877501;
assign addr[38484] = -423641043;
assign addr[38485] = -442370993;
assign addr[38486] = -461065866;
assign addr[38487] = -479724180;
assign addr[38488] = -498344454;
assign addr[38489] = -516925212;
assign addr[38490] = -535464981;
assign addr[38491] = -553962291;
assign addr[38492] = -572415676;
assign addr[38493] = -590823671;
assign addr[38494] = -609184818;
assign addr[38495] = -627497660;
assign addr[38496] = -645760745;
assign addr[38497] = -663972625;
assign addr[38498] = -682131857;
assign addr[38499] = -700236999;
assign addr[38500] = -718286617;
assign addr[38501] = -736279279;
assign addr[38502] = -754213559;
assign addr[38503] = -772088034;
assign addr[38504] = -789901288;
assign addr[38505] = -807651907;
assign addr[38506] = -825338484;
assign addr[38507] = -842959617;
assign addr[38508] = -860513908;
assign addr[38509] = -877999966;
assign addr[38510] = -895416404;
assign addr[38511] = -912761841;
assign addr[38512] = -930034901;
assign addr[38513] = -947234215;
assign addr[38514] = -964358420;
assign addr[38515] = -981406156;
assign addr[38516] = -998376073;
assign addr[38517] = -1015266825;
assign addr[38518] = -1032077073;
assign addr[38519] = -1048805483;
assign addr[38520] = -1065450729;
assign addr[38521] = -1082011492;
assign addr[38522] = -1098486458;
assign addr[38523] = -1114874320;
assign addr[38524] = -1131173780;
assign addr[38525] = -1147383544;
assign addr[38526] = -1163502328;
assign addr[38527] = -1179528853;
assign addr[38528] = -1195461849;
assign addr[38529] = -1211300053;
assign addr[38530] = -1227042207;
assign addr[38531] = -1242687064;
assign addr[38532] = -1258233384;
assign addr[38533] = -1273679934;
assign addr[38534] = -1289025489;
assign addr[38535] = -1304268832;
assign addr[38536] = -1319408754;
assign addr[38537] = -1334444055;
assign addr[38538] = -1349373543;
assign addr[38539] = -1364196034;
assign addr[38540] = -1378910353;
assign addr[38541] = -1393515332;
assign addr[38542] = -1408009814;
assign addr[38543] = -1422392650;
assign addr[38544] = -1436662698;
assign addr[38545] = -1450818828;
assign addr[38546] = -1464859917;
assign addr[38547] = -1478784851;
assign addr[38548] = -1492592527;
assign addr[38549] = -1506281850;
assign addr[38550] = -1519851733;
assign addr[38551] = -1533301101;
assign addr[38552] = -1546628888;
assign addr[38553] = -1559834037;
assign addr[38554] = -1572915501;
assign addr[38555] = -1585872242;
assign addr[38556] = -1598703233;
assign addr[38557] = -1611407456;
assign addr[38558] = -1623983905;
assign addr[38559] = -1636431582;
assign addr[38560] = -1648749499;
assign addr[38561] = -1660936681;
assign addr[38562] = -1672992161;
assign addr[38563] = -1684914983;
assign addr[38564] = -1696704201;
assign addr[38565] = -1708358881;
assign addr[38566] = -1719878099;
assign addr[38567] = -1731260941;
assign addr[38568] = -1742506504;
assign addr[38569] = -1753613897;
assign addr[38570] = -1764582240;
assign addr[38571] = -1775410662;
assign addr[38572] = -1786098304;
assign addr[38573] = -1796644320;
assign addr[38574] = -1807047873;
assign addr[38575] = -1817308138;
assign addr[38576] = -1827424302;
assign addr[38577] = -1837395562;
assign addr[38578] = -1847221128;
assign addr[38579] = -1856900221;
assign addr[38580] = -1866432072;
assign addr[38581] = -1875815927;
assign addr[38582] = -1885051042;
assign addr[38583] = -1894136683;
assign addr[38584] = -1903072131;
assign addr[38585] = -1911856677;
assign addr[38586] = -1920489624;
assign addr[38587] = -1928970288;
assign addr[38588] = -1937297997;
assign addr[38589] = -1945472089;
assign addr[38590] = -1953491918;
assign addr[38591] = -1961356847;
assign addr[38592] = -1969066252;
assign addr[38593] = -1976619522;
assign addr[38594] = -1984016058;
assign addr[38595] = -1991255274;
assign addr[38596] = -1998336596;
assign addr[38597] = -2005259462;
assign addr[38598] = -2012023322;
assign addr[38599] = -2018627642;
assign addr[38600] = -2025071897;
assign addr[38601] = -2031355576;
assign addr[38602] = -2037478181;
assign addr[38603] = -2043439226;
assign addr[38604] = -2049238240;
assign addr[38605] = -2054874761;
assign addr[38606] = -2060348343;
assign addr[38607] = -2065658552;
assign addr[38608] = -2070804967;
assign addr[38609] = -2075787180;
assign addr[38610] = -2080604795;
assign addr[38611] = -2085257431;
assign addr[38612] = -2089744719;
assign addr[38613] = -2094066304;
assign addr[38614] = -2098221841;
assign addr[38615] = -2102211002;
assign addr[38616] = -2106033471;
assign addr[38617] = -2109688944;
assign addr[38618] = -2113177132;
assign addr[38619] = -2116497758;
assign addr[38620] = -2119650558;
assign addr[38621] = -2122635283;
assign addr[38622] = -2125451696;
assign addr[38623] = -2128099574;
assign addr[38624] = -2130578706;
assign addr[38625] = -2132888897;
assign addr[38626] = -2135029962;
assign addr[38627] = -2137001733;
assign addr[38628] = -2138804053;
assign addr[38629] = -2140436778;
assign addr[38630] = -2141899780;
assign addr[38631] = -2143192942;
assign addr[38632] = -2144316162;
assign addr[38633] = -2145269351;
assign addr[38634] = -2146052433;
assign addr[38635] = -2146665347;
assign addr[38636] = -2147108043;
assign addr[38637] = -2147380486;
assign addr[38638] = -2147482655;
assign addr[38639] = -2147414542;
assign addr[38640] = -2147176152;
assign addr[38641] = -2146767505;
assign addr[38642] = -2146188631;
assign addr[38643] = -2145439578;
assign addr[38644] = -2144520405;
assign addr[38645] = -2143431184;
assign addr[38646] = -2142172003;
assign addr[38647] = -2140742960;
assign addr[38648] = -2139144169;
assign addr[38649] = -2137375758;
assign addr[38650] = -2135437865;
assign addr[38651] = -2133330646;
assign addr[38652] = -2131054266;
assign addr[38653] = -2128608907;
assign addr[38654] = -2125994762;
assign addr[38655] = -2123212038;
assign addr[38656] = -2120260957;
assign addr[38657] = -2117141752;
assign addr[38658] = -2113854671;
assign addr[38659] = -2110399974;
assign addr[38660] = -2106777935;
assign addr[38661] = -2102988841;
assign addr[38662] = -2099032994;
assign addr[38663] = -2094910706;
assign addr[38664] = -2090622304;
assign addr[38665] = -2086168128;
assign addr[38666] = -2081548533;
assign addr[38667] = -2076763883;
assign addr[38668] = -2071814558;
assign addr[38669] = -2066700952;
assign addr[38670] = -2061423468;
assign addr[38671] = -2055982526;
assign addr[38672] = -2050378558;
assign addr[38673] = -2044612007;
assign addr[38674] = -2038683330;
assign addr[38675] = -2032592999;
assign addr[38676] = -2026341495;
assign addr[38677] = -2019929315;
assign addr[38678] = -2013356967;
assign addr[38679] = -2006624971;
assign addr[38680] = -1999733863;
assign addr[38681] = -1992684188;
assign addr[38682] = -1985476506;
assign addr[38683] = -1978111387;
assign addr[38684] = -1970589416;
assign addr[38685] = -1962911189;
assign addr[38686] = -1955077316;
assign addr[38687] = -1947088417;
assign addr[38688] = -1938945125;
assign addr[38689] = -1930648088;
assign addr[38690] = -1922197961;
assign addr[38691] = -1913595416;
assign addr[38692] = -1904841135;
assign addr[38693] = -1895935811;
assign addr[38694] = -1886880151;
assign addr[38695] = -1877674873;
assign addr[38696] = -1868320707;
assign addr[38697] = -1858818395;
assign addr[38698] = -1849168689;
assign addr[38699] = -1839372356;
assign addr[38700] = -1829430172;
assign addr[38701] = -1819342925;
assign addr[38702] = -1809111415;
assign addr[38703] = -1798736454;
assign addr[38704] = -1788218865;
assign addr[38705] = -1777559480;
assign addr[38706] = -1766759146;
assign addr[38707] = -1755818718;
assign addr[38708] = -1744739065;
assign addr[38709] = -1733521064;
assign addr[38710] = -1722165606;
assign addr[38711] = -1710673591;
assign addr[38712] = -1699045930;
assign addr[38713] = -1687283545;
assign addr[38714] = -1675387369;
assign addr[38715] = -1663358344;
assign addr[38716] = -1651197426;
assign addr[38717] = -1638905577;
assign addr[38718] = -1626483774;
assign addr[38719] = -1613933000;
assign addr[38720] = -1601254251;
assign addr[38721] = -1588448533;
assign addr[38722] = -1575516860;
assign addr[38723] = -1562460258;
assign addr[38724] = -1549279763;
assign addr[38725] = -1535976419;
assign addr[38726] = -1522551282;
assign addr[38727] = -1509005416;
assign addr[38728] = -1495339895;
assign addr[38729] = -1481555802;
assign addr[38730] = -1467654232;
assign addr[38731] = -1453636285;
assign addr[38732] = -1439503074;
assign addr[38733] = -1425255719;
assign addr[38734] = -1410895350;
assign addr[38735] = -1396423105;
assign addr[38736] = -1381840133;
assign addr[38737] = -1367147589;
assign addr[38738] = -1352346639;
assign addr[38739] = -1337438456;
assign addr[38740] = -1322424222;
assign addr[38741] = -1307305128;
assign addr[38742] = -1292082373;
assign addr[38743] = -1276757164;
assign addr[38744] = -1261330715;
assign addr[38745] = -1245804251;
assign addr[38746] = -1230179002;
assign addr[38747] = -1214456207;
assign addr[38748] = -1198637114;
assign addr[38749] = -1182722976;
assign addr[38750] = -1166715055;
assign addr[38751] = -1150614620;
assign addr[38752] = -1134422949;
assign addr[38753] = -1118141326;
assign addr[38754] = -1101771040;
assign addr[38755] = -1085313391;
assign addr[38756] = -1068769683;
assign addr[38757] = -1052141228;
assign addr[38758] = -1035429345;
assign addr[38759] = -1018635358;
assign addr[38760] = -1001760600;
assign addr[38761] = -984806408;
assign addr[38762] = -967774128;
assign addr[38763] = -950665109;
assign addr[38764] = -933480707;
assign addr[38765] = -916222287;
assign addr[38766] = -898891215;
assign addr[38767] = -881488868;
assign addr[38768] = -864016623;
assign addr[38769] = -846475867;
assign addr[38770] = -828867991;
assign addr[38771] = -811194391;
assign addr[38772] = -793456467;
assign addr[38773] = -775655628;
assign addr[38774] = -757793284;
assign addr[38775] = -739870851;
assign addr[38776] = -721889752;
assign addr[38777] = -703851410;
assign addr[38778] = -685757258;
assign addr[38779] = -667608730;
assign addr[38780] = -649407264;
assign addr[38781] = -631154304;
assign addr[38782] = -612851297;
assign addr[38783] = -594499695;
assign addr[38784] = -576100953;
assign addr[38785] = -557656529;
assign addr[38786] = -539167887;
assign addr[38787] = -520636492;
assign addr[38788] = -502063814;
assign addr[38789] = -483451325;
assign addr[38790] = -464800501;
assign addr[38791] = -446112822;
assign addr[38792] = -427389768;
assign addr[38793] = -408632825;
assign addr[38794] = -389843480;
assign addr[38795] = -371023223;
assign addr[38796] = -352173546;
assign addr[38797] = -333295944;
assign addr[38798] = -314391913;
assign addr[38799] = -295462954;
assign addr[38800] = -276510565;
assign addr[38801] = -257536251;
assign addr[38802] = -238541516;
assign addr[38803] = -219527866;
assign addr[38804] = -200496809;
assign addr[38805] = -181449854;
assign addr[38806] = -162388511;
assign addr[38807] = -143314291;
assign addr[38808] = -124228708;
assign addr[38809] = -105133274;
assign addr[38810] = -86029503;
assign addr[38811] = -66918911;
assign addr[38812] = -47803013;
assign addr[38813] = -28683324;
assign addr[38814] = -9561361;
assign addr[38815] = 9561361;
assign addr[38816] = 28683324;
assign addr[38817] = 47803013;
assign addr[38818] = 66918911;
assign addr[38819] = 86029503;
assign addr[38820] = 105133274;
assign addr[38821] = 124228708;
assign addr[38822] = 143314291;
assign addr[38823] = 162388511;
assign addr[38824] = 181449854;
assign addr[38825] = 200496809;
assign addr[38826] = 219527866;
assign addr[38827] = 238541516;
assign addr[38828] = 257536251;
assign addr[38829] = 276510565;
assign addr[38830] = 295462953;
assign addr[38831] = 314391913;
assign addr[38832] = 333295944;
assign addr[38833] = 352173546;
assign addr[38834] = 371023223;
assign addr[38835] = 389843480;
assign addr[38836] = 408632825;
assign addr[38837] = 427389768;
assign addr[38838] = 446112822;
assign addr[38839] = 464800501;
assign addr[38840] = 483451325;
assign addr[38841] = 502063814;
assign addr[38842] = 520636492;
assign addr[38843] = 539167887;
assign addr[38844] = 557656529;
assign addr[38845] = 576100953;
assign addr[38846] = 594499695;
assign addr[38847] = 612851297;
assign addr[38848] = 631154304;
assign addr[38849] = 649407264;
assign addr[38850] = 667608730;
assign addr[38851] = 685757258;
assign addr[38852] = 703851410;
assign addr[38853] = 721889752;
assign addr[38854] = 739870851;
assign addr[38855] = 757793284;
assign addr[38856] = 775655628;
assign addr[38857] = 793456467;
assign addr[38858] = 811194391;
assign addr[38859] = 828867991;
assign addr[38860] = 846475867;
assign addr[38861] = 864016623;
assign addr[38862] = 881488868;
assign addr[38863] = 898891215;
assign addr[38864] = 916222287;
assign addr[38865] = 933480707;
assign addr[38866] = 950665109;
assign addr[38867] = 967774128;
assign addr[38868] = 984806408;
assign addr[38869] = 1001760600;
assign addr[38870] = 1018635358;
assign addr[38871] = 1035429345;
assign addr[38872] = 1052141228;
assign addr[38873] = 1068769683;
assign addr[38874] = 1085313391;
assign addr[38875] = 1101771040;
assign addr[38876] = 1118141326;
assign addr[38877] = 1134422949;
assign addr[38878] = 1150614620;
assign addr[38879] = 1166715055;
assign addr[38880] = 1182722976;
assign addr[38881] = 1198637114;
assign addr[38882] = 1214456207;
assign addr[38883] = 1230179002;
assign addr[38884] = 1245804251;
assign addr[38885] = 1261330715;
assign addr[38886] = 1276757164;
assign addr[38887] = 1292082373;
assign addr[38888] = 1307305128;
assign addr[38889] = 1322424222;
assign addr[38890] = 1337438456;
assign addr[38891] = 1352346639;
assign addr[38892] = 1367147589;
assign addr[38893] = 1381840133;
assign addr[38894] = 1396423105;
assign addr[38895] = 1410895350;
assign addr[38896] = 1425255719;
assign addr[38897] = 1439503074;
assign addr[38898] = 1453636285;
assign addr[38899] = 1467654232;
assign addr[38900] = 1481555802;
assign addr[38901] = 1495339895;
assign addr[38902] = 1509005416;
assign addr[38903] = 1522551282;
assign addr[38904] = 1535976419;
assign addr[38905] = 1549279763;
assign addr[38906] = 1562460258;
assign addr[38907] = 1575516860;
assign addr[38908] = 1588448533;
assign addr[38909] = 1601254251;
assign addr[38910] = 1613933000;
assign addr[38911] = 1626483774;
assign addr[38912] = 1638905577;
assign addr[38913] = 1651197426;
assign addr[38914] = 1663358344;
assign addr[38915] = 1675387369;
assign addr[38916] = 1687283545;
assign addr[38917] = 1699045930;
assign addr[38918] = 1710673591;
assign addr[38919] = 1722165606;
assign addr[38920] = 1733521064;
assign addr[38921] = 1744739065;
assign addr[38922] = 1755818718;
assign addr[38923] = 1766759146;
assign addr[38924] = 1777559480;
assign addr[38925] = 1788218865;
assign addr[38926] = 1798736454;
assign addr[38927] = 1809111415;
assign addr[38928] = 1819342925;
assign addr[38929] = 1829430172;
assign addr[38930] = 1839372356;
assign addr[38931] = 1849168689;
assign addr[38932] = 1858818395;
assign addr[38933] = 1868320707;
assign addr[38934] = 1877674873;
assign addr[38935] = 1886880151;
assign addr[38936] = 1895935811;
assign addr[38937] = 1904841135;
assign addr[38938] = 1913595416;
assign addr[38939] = 1922197961;
assign addr[38940] = 1930648088;
assign addr[38941] = 1938945125;
assign addr[38942] = 1947088417;
assign addr[38943] = 1955077316;
assign addr[38944] = 1962911189;
assign addr[38945] = 1970589416;
assign addr[38946] = 1978111387;
assign addr[38947] = 1985476506;
assign addr[38948] = 1992684188;
assign addr[38949] = 1999733863;
assign addr[38950] = 2006624971;
assign addr[38951] = 2013356967;
assign addr[38952] = 2019929315;
assign addr[38953] = 2026341495;
assign addr[38954] = 2032592999;
assign addr[38955] = 2038683330;
assign addr[38956] = 2044612007;
assign addr[38957] = 2050378558;
assign addr[38958] = 2055982526;
assign addr[38959] = 2061423468;
assign addr[38960] = 2066700952;
assign addr[38961] = 2071814558;
assign addr[38962] = 2076763883;
assign addr[38963] = 2081548533;
assign addr[38964] = 2086168128;
assign addr[38965] = 2090622304;
assign addr[38966] = 2094910706;
assign addr[38967] = 2099032994;
assign addr[38968] = 2102988841;
assign addr[38969] = 2106777935;
assign addr[38970] = 2110399974;
assign addr[38971] = 2113854671;
assign addr[38972] = 2117141752;
assign addr[38973] = 2120260957;
assign addr[38974] = 2123212038;
assign addr[38975] = 2125994762;
assign addr[38976] = 2128608907;
assign addr[38977] = 2131054266;
assign addr[38978] = 2133330646;
assign addr[38979] = 2135437865;
assign addr[38980] = 2137375758;
assign addr[38981] = 2139144169;
assign addr[38982] = 2140742960;
assign addr[38983] = 2142172003;
assign addr[38984] = 2143431184;
assign addr[38985] = 2144520405;
assign addr[38986] = 2145439578;
assign addr[38987] = 2146188631;
assign addr[38988] = 2146767505;
assign addr[38989] = 2147176152;
assign addr[38990] = 2147414542;
assign addr[38991] = 2147482655;
assign addr[38992] = 2147380486;
assign addr[38993] = 2147108043;
assign addr[38994] = 2146665347;
assign addr[38995] = 2146052433;
assign addr[38996] = 2145269351;
assign addr[38997] = 2144316162;
assign addr[38998] = 2143192942;
assign addr[38999] = 2141899780;
assign addr[39000] = 2140436778;
assign addr[39001] = 2138804053;
assign addr[39002] = 2137001733;
assign addr[39003] = 2135029962;
assign addr[39004] = 2132888897;
assign addr[39005] = 2130578706;
assign addr[39006] = 2128099574;
assign addr[39007] = 2125451696;
assign addr[39008] = 2122635283;
assign addr[39009] = 2119650558;
assign addr[39010] = 2116497758;
assign addr[39011] = 2113177132;
assign addr[39012] = 2109688944;
assign addr[39013] = 2106033471;
assign addr[39014] = 2102211002;
assign addr[39015] = 2098221841;
assign addr[39016] = 2094066304;
assign addr[39017] = 2089744719;
assign addr[39018] = 2085257431;
assign addr[39019] = 2080604795;
assign addr[39020] = 2075787180;
assign addr[39021] = 2070804967;
assign addr[39022] = 2065658552;
assign addr[39023] = 2060348343;
assign addr[39024] = 2054874761;
assign addr[39025] = 2049238240;
assign addr[39026] = 2043439226;
assign addr[39027] = 2037478181;
assign addr[39028] = 2031355576;
assign addr[39029] = 2025071897;
assign addr[39030] = 2018627642;
assign addr[39031] = 2012023322;
assign addr[39032] = 2005259462;
assign addr[39033] = 1998336596;
assign addr[39034] = 1991255274;
assign addr[39035] = 1984016058;
assign addr[39036] = 1976619522;
assign addr[39037] = 1969066252;
assign addr[39038] = 1961356847;
assign addr[39039] = 1953491918;
assign addr[39040] = 1945472089;
assign addr[39041] = 1937297997;
assign addr[39042] = 1928970288;
assign addr[39043] = 1920489624;
assign addr[39044] = 1911856677;
assign addr[39045] = 1903072131;
assign addr[39046] = 1894136683;
assign addr[39047] = 1885051042;
assign addr[39048] = 1875815927;
assign addr[39049] = 1866432072;
assign addr[39050] = 1856900221;
assign addr[39051] = 1847221128;
assign addr[39052] = 1837395562;
assign addr[39053] = 1827424302;
assign addr[39054] = 1817308138;
assign addr[39055] = 1807047873;
assign addr[39056] = 1796644320;
assign addr[39057] = 1786098304;
assign addr[39058] = 1775410662;
assign addr[39059] = 1764582240;
assign addr[39060] = 1753613897;
assign addr[39061] = 1742506504;
assign addr[39062] = 1731260941;
assign addr[39063] = 1719878099;
assign addr[39064] = 1708358881;
assign addr[39065] = 1696704201;
assign addr[39066] = 1684914983;
assign addr[39067] = 1672992161;
assign addr[39068] = 1660936681;
assign addr[39069] = 1648749499;
assign addr[39070] = 1636431582;
assign addr[39071] = 1623983905;
assign addr[39072] = 1611407456;
assign addr[39073] = 1598703233;
assign addr[39074] = 1585872242;
assign addr[39075] = 1572915501;
assign addr[39076] = 1559834037;
assign addr[39077] = 1546628888;
assign addr[39078] = 1533301101;
assign addr[39079] = 1519851733;
assign addr[39080] = 1506281850;
assign addr[39081] = 1492592527;
assign addr[39082] = 1478784851;
assign addr[39083] = 1464859917;
assign addr[39084] = 1450818828;
assign addr[39085] = 1436662698;
assign addr[39086] = 1422392650;
assign addr[39087] = 1408009814;
assign addr[39088] = 1393515332;
assign addr[39089] = 1378910353;
assign addr[39090] = 1364196034;
assign addr[39091] = 1349373543;
assign addr[39092] = 1334444055;
assign addr[39093] = 1319408754;
assign addr[39094] = 1304268832;
assign addr[39095] = 1289025489;
assign addr[39096] = 1273679934;
assign addr[39097] = 1258233384;
assign addr[39098] = 1242687064;
assign addr[39099] = 1227042207;
assign addr[39100] = 1211300053;
assign addr[39101] = 1195461849;
assign addr[39102] = 1179528853;
assign addr[39103] = 1163502328;
assign addr[39104] = 1147383544;
assign addr[39105] = 1131173780;
assign addr[39106] = 1114874320;
assign addr[39107] = 1098486458;
assign addr[39108] = 1082011492;
assign addr[39109] = 1065450729;
assign addr[39110] = 1048805483;
assign addr[39111] = 1032077073;
assign addr[39112] = 1015266825;
assign addr[39113] = 998376073;
assign addr[39114] = 981406156;
assign addr[39115] = 964358420;
assign addr[39116] = 947234215;
assign addr[39117] = 930034901;
assign addr[39118] = 912761841;
assign addr[39119] = 895416404;
assign addr[39120] = 877999966;
assign addr[39121] = 860513908;
assign addr[39122] = 842959617;
assign addr[39123] = 825338484;
assign addr[39124] = 807651907;
assign addr[39125] = 789901288;
assign addr[39126] = 772088034;
assign addr[39127] = 754213559;
assign addr[39128] = 736279279;
assign addr[39129] = 718286617;
assign addr[39130] = 700236999;
assign addr[39131] = 682131857;
assign addr[39132] = 663972625;
assign addr[39133] = 645760745;
assign addr[39134] = 627497660;
assign addr[39135] = 609184818;
assign addr[39136] = 590823671;
assign addr[39137] = 572415676;
assign addr[39138] = 553962291;
assign addr[39139] = 535464981;
assign addr[39140] = 516925212;
assign addr[39141] = 498344454;
assign addr[39142] = 479724180;
assign addr[39143] = 461065866;
assign addr[39144] = 442370993;
assign addr[39145] = 423641043;
assign addr[39146] = 404877501;
assign addr[39147] = 386081854;
assign addr[39148] = 367255594;
assign addr[39149] = 348400212;
assign addr[39150] = 329517204;
assign addr[39151] = 310608068;
assign addr[39152] = 291674302;
assign addr[39153] = 272717408;
assign addr[39154] = 253738890;
assign addr[39155] = 234740251;
assign addr[39156] = 215722999;
assign addr[39157] = 196688642;
assign addr[39158] = 177638688;
assign addr[39159] = 158574649;
assign addr[39160] = 139498035;
assign addr[39161] = 120410361;
assign addr[39162] = 101313138;
assign addr[39163] = 82207882;
assign addr[39164] = 63096108;
assign addr[39165] = 43979330;
assign addr[39166] = 24859065;
assign addr[39167] = 5736829;
assign addr[39168] = -13385863;
assign addr[39169] = -32507492;
assign addr[39170] = -51626544;
assign addr[39171] = -70741503;
assign addr[39172] = -89850852;
assign addr[39173] = -108953076;
assign addr[39174] = -128046661;
assign addr[39175] = -147130093;
assign addr[39176] = -166201858;
assign addr[39177] = -185260444;
assign addr[39178] = -204304341;
assign addr[39179] = -223332037;
assign addr[39180] = -242342025;
assign addr[39181] = -261332796;
assign addr[39182] = -280302845;
assign addr[39183] = -299250668;
assign addr[39184] = -318174762;
assign addr[39185] = -337073627;
assign addr[39186] = -355945764;
assign addr[39187] = -374789676;
assign addr[39188] = -393603870;
assign addr[39189] = -412386854;
assign addr[39190] = -431137138;
assign addr[39191] = -449853235;
assign addr[39192] = -468533662;
assign addr[39193] = -487176937;
assign addr[39194] = -505781581;
assign addr[39195] = -524346121;
assign addr[39196] = -542869083;
assign addr[39197] = -561348998;
assign addr[39198] = -579784402;
assign addr[39199] = -598173833;
assign addr[39200] = -616515832;
assign addr[39201] = -634808946;
assign addr[39202] = -653051723;
assign addr[39203] = -671242716;
assign addr[39204] = -689380485;
assign addr[39205] = -707463589;
assign addr[39206] = -725490597;
assign addr[39207] = -743460077;
assign addr[39208] = -761370605;
assign addr[39209] = -779220762;
assign addr[39210] = -797009130;
assign addr[39211] = -814734301;
assign addr[39212] = -832394869;
assign addr[39213] = -849989433;
assign addr[39214] = -867516597;
assign addr[39215] = -884974973;
assign addr[39216] = -902363176;
assign addr[39217] = -919679827;
assign addr[39218] = -936923553;
assign addr[39219] = -954092986;
assign addr[39220] = -971186766;
assign addr[39221] = -988203537;
assign addr[39222] = -1005141949;
assign addr[39223] = -1022000660;
assign addr[39224] = -1038778332;
assign addr[39225] = -1055473635;
assign addr[39226] = -1072085246;
assign addr[39227] = -1088611847;
assign addr[39228] = -1105052128;
assign addr[39229] = -1121404785;
assign addr[39230] = -1137668521;
assign addr[39231] = -1153842047;
assign addr[39232] = -1169924081;
assign addr[39233] = -1185913346;
assign addr[39234] = -1201808576;
assign addr[39235] = -1217608510;
assign addr[39236] = -1233311895;
assign addr[39237] = -1248917486;
assign addr[39238] = -1264424045;
assign addr[39239] = -1279830344;
assign addr[39240] = -1295135159;
assign addr[39241] = -1310337279;
assign addr[39242] = -1325435496;
assign addr[39243] = -1340428615;
assign addr[39244] = -1355315445;
assign addr[39245] = -1370094808;
assign addr[39246] = -1384765530;
assign addr[39247] = -1399326449;
assign addr[39248] = -1413776410;
assign addr[39249] = -1428114267;
assign addr[39250] = -1442338884;
assign addr[39251] = -1456449131;
assign addr[39252] = -1470443891;
assign addr[39253] = -1484322054;
assign addr[39254] = -1498082520;
assign addr[39255] = -1511724196;
assign addr[39256] = -1525246002;
assign addr[39257] = -1538646865;
assign addr[39258] = -1551925723;
assign addr[39259] = -1565081523;
assign addr[39260] = -1578113222;
assign addr[39261] = -1591019785;
assign addr[39262] = -1603800191;
assign addr[39263] = -1616453425;
assign addr[39264] = -1628978484;
assign addr[39265] = -1641374375;
assign addr[39266] = -1653640115;
assign addr[39267] = -1665774731;
assign addr[39268] = -1677777262;
assign addr[39269] = -1689646755;
assign addr[39270] = -1701382270;
assign addr[39271] = -1712982875;
assign addr[39272] = -1724447652;
assign addr[39273] = -1735775690;
assign addr[39274] = -1746966091;
assign addr[39275] = -1758017969;
assign addr[39276] = -1768930447;
assign addr[39277] = -1779702660;
assign addr[39278] = -1790333753;
assign addr[39279] = -1800822883;
assign addr[39280] = -1811169220;
assign addr[39281] = -1821371941;
assign addr[39282] = -1831430239;
assign addr[39283] = -1841343316;
assign addr[39284] = -1851110385;
assign addr[39285] = -1860730673;
assign addr[39286] = -1870203416;
assign addr[39287] = -1879527863;
assign addr[39288] = -1888703276;
assign addr[39289] = -1897728925;
assign addr[39290] = -1906604097;
assign addr[39291] = -1915328086;
assign addr[39292] = -1923900201;
assign addr[39293] = -1932319763;
assign addr[39294] = -1940586104;
assign addr[39295] = -1948698568;
assign addr[39296] = -1956656513;
assign addr[39297] = -1964459306;
assign addr[39298] = -1972106330;
assign addr[39299] = -1979596978;
assign addr[39300] = -1986930656;
assign addr[39301] = -1994106782;
assign addr[39302] = -2001124788;
assign addr[39303] = -2007984117;
assign addr[39304] = -2014684225;
assign addr[39305] = -2021224581;
assign addr[39306] = -2027604666;
assign addr[39307] = -2033823974;
assign addr[39308] = -2039882013;
assign addr[39309] = -2045778302;
assign addr[39310] = -2051512372;
assign addr[39311] = -2057083771;
assign addr[39312] = -2062492055;
assign addr[39313] = -2067736796;
assign addr[39314] = -2072817579;
assign addr[39315] = -2077733999;
assign addr[39316] = -2082485668;
assign addr[39317] = -2087072209;
assign addr[39318] = -2091493257;
assign addr[39319] = -2095748463;
assign addr[39320] = -2099837489;
assign addr[39321] = -2103760010;
assign addr[39322] = -2107515716;
assign addr[39323] = -2111104309;
assign addr[39324] = -2114525505;
assign addr[39325] = -2117779031;
assign addr[39326] = -2120864631;
assign addr[39327] = -2123782059;
assign addr[39328] = -2126531084;
assign addr[39329] = -2129111488;
assign addr[39330] = -2131523066;
assign addr[39331] = -2133765628;
assign addr[39332] = -2135838995;
assign addr[39333] = -2137743003;
assign addr[39334] = -2139477502;
assign addr[39335] = -2141042352;
assign addr[39336] = -2142437431;
assign addr[39337] = -2143662628;
assign addr[39338] = -2144717846;
assign addr[39339] = -2145603001;
assign addr[39340] = -2146318022;
assign addr[39341] = -2146862854;
assign addr[39342] = -2147237452;
assign addr[39343] = -2147441787;
assign addr[39344] = -2147475844;
assign addr[39345] = -2147339619;
assign addr[39346] = -2147033123;
assign addr[39347] = -2146556380;
assign addr[39348] = -2145909429;
assign addr[39349] = -2145092320;
assign addr[39350] = -2144105118;
assign addr[39351] = -2142947902;
assign addr[39352] = -2141620763;
assign addr[39353] = -2140123807;
assign addr[39354] = -2138457152;
assign addr[39355] = -2136620930;
assign addr[39356] = -2134615288;
assign addr[39357] = -2132440383;
assign addr[39358] = -2130096389;
assign addr[39359] = -2127583492;
assign addr[39360] = -2124901890;
assign addr[39361] = -2122051796;
assign addr[39362] = -2119033436;
assign addr[39363] = -2115847050;
assign addr[39364] = -2112492891;
assign addr[39365] = -2108971223;
assign addr[39366] = -2105282327;
assign addr[39367] = -2101426496;
assign addr[39368] = -2097404033;
assign addr[39369] = -2093215260;
assign addr[39370] = -2088860507;
assign addr[39371] = -2084340120;
assign addr[39372] = -2079654458;
assign addr[39373] = -2074803892;
assign addr[39374] = -2069788807;
assign addr[39375] = -2064609600;
assign addr[39376] = -2059266683;
assign addr[39377] = -2053760478;
assign addr[39378] = -2048091422;
assign addr[39379] = -2042259965;
assign addr[39380] = -2036266570;
assign addr[39381] = -2030111710;
assign addr[39382] = -2023795876;
assign addr[39383] = -2017319567;
assign addr[39384] = -2010683297;
assign addr[39385] = -2003887591;
assign addr[39386] = -1996932990;
assign addr[39387] = -1989820044;
assign addr[39388] = -1982549318;
assign addr[39389] = -1975121388;
assign addr[39390] = -1967536842;
assign addr[39391] = -1959796283;
assign addr[39392] = -1951900324;
assign addr[39393] = -1943849591;
assign addr[39394] = -1935644723;
assign addr[39395] = -1927286370;
assign addr[39396] = -1918775195;
assign addr[39397] = -1910111873;
assign addr[39398] = -1901297091;
assign addr[39399] = -1892331547;
assign addr[39400] = -1883215953;
assign addr[39401] = -1873951032;
assign addr[39402] = -1864537518;
assign addr[39403] = -1854976157;
assign addr[39404] = -1845267708;
assign addr[39405] = -1835412941;
assign addr[39406] = -1825412636;
assign addr[39407] = -1815267588;
assign addr[39408] = -1804978599;
assign addr[39409] = -1794546487;
assign addr[39410] = -1783972079;
assign addr[39411] = -1773256212;
assign addr[39412] = -1762399737;
assign addr[39413] = -1751403515;
assign addr[39414] = -1740268417;
assign addr[39415] = -1728995326;
assign addr[39416] = -1717585136;
assign addr[39417] = -1706038753;
assign addr[39418] = -1694357091;
assign addr[39419] = -1682541077;
assign addr[39420] = -1670591647;
assign addr[39421] = -1658509750;
assign addr[39422] = -1646296344;
assign addr[39423] = -1633952396;
assign addr[39424] = -1621478885;
assign addr[39425] = -1608876801;
assign addr[39426] = -1596147143;
assign addr[39427] = -1583290921;
assign addr[39428] = -1570309153;
assign addr[39429] = -1557202869;
assign addr[39430] = -1543973108;
assign addr[39431] = -1530620920;
assign addr[39432] = -1517147363;
assign addr[39433] = -1503553506;
assign addr[39434] = -1489840425;
assign addr[39435] = -1476009210;
assign addr[39436] = -1462060956;
assign addr[39437] = -1447996770;
assign addr[39438] = -1433817766;
assign addr[39439] = -1419525069;
assign addr[39440] = -1405119813;
assign addr[39441] = -1390603139;
assign addr[39442] = -1375976199;
assign addr[39443] = -1361240152;
assign addr[39444] = -1346396168;
assign addr[39445] = -1331445422;
assign addr[39446] = -1316389101;
assign addr[39447] = -1301228398;
assign addr[39448] = -1285964516;
assign addr[39449] = -1270598665;
assign addr[39450] = -1255132063;
assign addr[39451] = -1239565936;
assign addr[39452] = -1223901520;
assign addr[39453] = -1208140056;
assign addr[39454] = -1192282793;
assign addr[39455] = -1176330990;
assign addr[39456] = -1160285911;
assign addr[39457] = -1144148829;
assign addr[39458] = -1127921022;
assign addr[39459] = -1111603778;
assign addr[39460] = -1095198391;
assign addr[39461] = -1078706161;
assign addr[39462] = -1062128397;
assign addr[39463] = -1045466412;
assign addr[39464] = -1028721528;
assign addr[39465] = -1011895073;
assign addr[39466] = -994988380;
assign addr[39467] = -978002791;
assign addr[39468] = -960939653;
assign addr[39469] = -943800318;
assign addr[39470] = -926586145;
assign addr[39471] = -909298500;
assign addr[39472] = -891938752;
assign addr[39473] = -874508280;
assign addr[39474] = -857008464;
assign addr[39475] = -839440693;
assign addr[39476] = -821806359;
assign addr[39477] = -804106861;
assign addr[39478] = -786343603;
assign addr[39479] = -768517992;
assign addr[39480] = -750631442;
assign addr[39481] = -732685372;
assign addr[39482] = -714681204;
assign addr[39483] = -696620367;
assign addr[39484] = -678504291;
assign addr[39485] = -660334415;
assign addr[39486] = -642112178;
assign addr[39487] = -623839025;
assign addr[39488] = -605516406;
assign addr[39489] = -587145773;
assign addr[39490] = -568728583;
assign addr[39491] = -550266296;
assign addr[39492] = -531760377;
assign addr[39493] = -513212292;
assign addr[39494] = -494623513;
assign addr[39495] = -475995513;
assign addr[39496] = -457329769;
assign addr[39497] = -438627762;
assign addr[39498] = -419890975;
assign addr[39499] = -401120892;
assign addr[39500] = -382319004;
assign addr[39501] = -363486799;
assign addr[39502] = -344625773;
assign addr[39503] = -325737419;
assign addr[39504] = -306823237;
assign addr[39505] = -287884725;
assign addr[39506] = -268923386;
assign addr[39507] = -249940723;
assign addr[39508] = -230938242;
assign addr[39509] = -211917448;
assign addr[39510] = -192879850;
assign addr[39511] = -173826959;
assign addr[39512] = -154760284;
assign addr[39513] = -135681337;
assign addr[39514] = -116591632;
assign addr[39515] = -97492681;
assign addr[39516] = -78386000;
assign addr[39517] = -59273104;
assign addr[39518] = -40155507;
assign addr[39519] = -21034727;
assign addr[39520] = -1912278;
assign addr[39521] = 17210322;
assign addr[39522] = 36331557;
assign addr[39523] = 55449912;
assign addr[39524] = 74563870;
assign addr[39525] = 93671915;
assign addr[39526] = 112772533;
assign addr[39527] = 131864208;
assign addr[39528] = 150945428;
assign addr[39529] = 170014678;
assign addr[39530] = 189070447;
assign addr[39531] = 208111224;
assign addr[39532] = 227135500;
assign addr[39533] = 246141764;
assign addr[39534] = 265128512;
assign addr[39535] = 284094236;
assign addr[39536] = 303037433;
assign addr[39537] = 321956601;
assign addr[39538] = 340850240;
assign addr[39539] = 359716852;
assign addr[39540] = 378554940;
assign addr[39541] = 397363011;
assign addr[39542] = 416139574;
assign addr[39543] = 434883140;
assign addr[39544] = 453592221;
assign addr[39545] = 472265336;
assign addr[39546] = 490901003;
assign addr[39547] = 509497745;
assign addr[39548] = 528054086;
assign addr[39549] = 546568556;
assign addr[39550] = 565039687;
assign addr[39551] = 583466013;
assign addr[39552] = 601846074;
assign addr[39553] = 620178412;
assign addr[39554] = 638461574;
assign addr[39555] = 656694110;
assign addr[39556] = 674874574;
assign addr[39557] = 693001525;
assign addr[39558] = 711073524;
assign addr[39559] = 729089140;
assign addr[39560] = 747046944;
assign addr[39561] = 764945512;
assign addr[39562] = 782783424;
assign addr[39563] = 800559266;
assign addr[39564] = 818271628;
assign addr[39565] = 835919107;
assign addr[39566] = 853500302;
assign addr[39567] = 871013820;
assign addr[39568] = 888458272;
assign addr[39569] = 905832274;
assign addr[39570] = 923134450;
assign addr[39571] = 940363427;
assign addr[39572] = 957517838;
assign addr[39573] = 974596324;
assign addr[39574] = 991597531;
assign addr[39575] = 1008520110;
assign addr[39576] = 1025362720;
assign addr[39577] = 1042124025;
assign addr[39578] = 1058802695;
assign addr[39579] = 1075397409;
assign addr[39580] = 1091906851;
assign addr[39581] = 1108329711;
assign addr[39582] = 1124664687;
assign addr[39583] = 1140910484;
assign addr[39584] = 1157065814;
assign addr[39585] = 1173129396;
assign addr[39586] = 1189099956;
assign addr[39587] = 1204976227;
assign addr[39588] = 1220756951;
assign addr[39589] = 1236440877;
assign addr[39590] = 1252026760;
assign addr[39591] = 1267513365;
assign addr[39592] = 1282899464;
assign addr[39593] = 1298183838;
assign addr[39594] = 1313365273;
assign addr[39595] = 1328442566;
assign addr[39596] = 1343414522;
assign addr[39597] = 1358279953;
assign addr[39598] = 1373037681;
assign addr[39599] = 1387686535;
assign addr[39600] = 1402225355;
assign addr[39601] = 1416652986;
assign addr[39602] = 1430968286;
assign addr[39603] = 1445170118;
assign addr[39604] = 1459257358;
assign addr[39605] = 1473228887;
assign addr[39606] = 1487083598;
assign addr[39607] = 1500820393;
assign addr[39608] = 1514438181;
assign addr[39609] = 1527935884;
assign addr[39610] = 1541312431;
assign addr[39611] = 1554566762;
assign addr[39612] = 1567697824;
assign addr[39613] = 1580704578;
assign addr[39614] = 1593585992;
assign addr[39615] = 1606341043;
assign addr[39616] = 1618968722;
assign addr[39617] = 1631468027;
assign addr[39618] = 1643837966;
assign addr[39619] = 1656077559;
assign addr[39620] = 1668185835;
assign addr[39621] = 1680161834;
assign addr[39622] = 1692004606;
assign addr[39623] = 1703713213;
assign addr[39624] = 1715286726;
assign addr[39625] = 1726724227;
assign addr[39626] = 1738024810;
assign addr[39627] = 1749187577;
assign addr[39628] = 1760211645;
assign addr[39629] = 1771096139;
assign addr[39630] = 1781840195;
assign addr[39631] = 1792442963;
assign addr[39632] = 1802903601;
assign addr[39633] = 1813221279;
assign addr[39634] = 1823395180;
assign addr[39635] = 1833424497;
assign addr[39636] = 1843308435;
assign addr[39637] = 1853046210;
assign addr[39638] = 1862637049;
assign addr[39639] = 1872080193;
assign addr[39640] = 1881374892;
assign addr[39641] = 1890520410;
assign addr[39642] = 1899516021;
assign addr[39643] = 1908361011;
assign addr[39644] = 1917054681;
assign addr[39645] = 1925596340;
assign addr[39646] = 1933985310;
assign addr[39647] = 1942220928;
assign addr[39648] = 1950302539;
assign addr[39649] = 1958229503;
assign addr[39650] = 1966001192;
assign addr[39651] = 1973616989;
assign addr[39652] = 1981076290;
assign addr[39653] = 1988378503;
assign addr[39654] = 1995523051;
assign addr[39655] = 2002509365;
assign addr[39656] = 2009336893;
assign addr[39657] = 2016005093;
assign addr[39658] = 2022513436;
assign addr[39659] = 2028861406;
assign addr[39660] = 2035048499;
assign addr[39661] = 2041074226;
assign addr[39662] = 2046938108;
assign addr[39663] = 2052639680;
assign addr[39664] = 2058178491;
assign addr[39665] = 2063554100;
assign addr[39666] = 2068766083;
assign addr[39667] = 2073814024;
assign addr[39668] = 2078697525;
assign addr[39669] = 2083416198;
assign addr[39670] = 2087969669;
assign addr[39671] = 2092357577;
assign addr[39672] = 2096579573;
assign addr[39673] = 2100635323;
assign addr[39674] = 2104524506;
assign addr[39675] = 2108246813;
assign addr[39676] = 2111801949;
assign addr[39677] = 2115189632;
assign addr[39678] = 2118409593;
assign addr[39679] = 2121461578;
assign addr[39680] = 2124345343;
assign addr[39681] = 2127060661;
assign addr[39682] = 2129607316;
assign addr[39683] = 2131985106;
assign addr[39684] = 2134193842;
assign addr[39685] = 2136233350;
assign addr[39686] = 2138103468;
assign addr[39687] = 2139804048;
assign addr[39688] = 2141334954;
assign addr[39689] = 2142696065;
assign addr[39690] = 2143887273;
assign addr[39691] = 2144908484;
assign addr[39692] = 2145759618;
assign addr[39693] = 2146440605;
assign addr[39694] = 2146951393;
assign addr[39695] = 2147291941;
assign addr[39696] = 2147462221;
assign addr[39697] = 2147462221;
assign addr[39698] = 2147291941;
assign addr[39699] = 2146951393;
assign addr[39700] = 2146440605;
assign addr[39701] = 2145759618;
assign addr[39702] = 2144908484;
assign addr[39703] = 2143887273;
assign addr[39704] = 2142696065;
assign addr[39705] = 2141334954;
assign addr[39706] = 2139804048;
assign addr[39707] = 2138103468;
assign addr[39708] = 2136233350;
assign addr[39709] = 2134193842;
assign addr[39710] = 2131985106;
assign addr[39711] = 2129607316;
assign addr[39712] = 2127060661;
assign addr[39713] = 2124345343;
assign addr[39714] = 2121461578;
assign addr[39715] = 2118409593;
assign addr[39716] = 2115189632;
assign addr[39717] = 2111801949;
assign addr[39718] = 2108246813;
assign addr[39719] = 2104524506;
assign addr[39720] = 2100635323;
assign addr[39721] = 2096579573;
assign addr[39722] = 2092357577;
assign addr[39723] = 2087969669;
assign addr[39724] = 2083416198;
assign addr[39725] = 2078697525;
assign addr[39726] = 2073814024;
assign addr[39727] = 2068766083;
assign addr[39728] = 2063554100;
assign addr[39729] = 2058178491;
assign addr[39730] = 2052639680;
assign addr[39731] = 2046938108;
assign addr[39732] = 2041074226;
assign addr[39733] = 2035048499;
assign addr[39734] = 2028861406;
assign addr[39735] = 2022513436;
assign addr[39736] = 2016005093;
assign addr[39737] = 2009336893;
assign addr[39738] = 2002509365;
assign addr[39739] = 1995523051;
assign addr[39740] = 1988378503;
assign addr[39741] = 1981076290;
assign addr[39742] = 1973616989;
assign addr[39743] = 1966001192;
assign addr[39744] = 1958229503;
assign addr[39745] = 1950302539;
assign addr[39746] = 1942220928;
assign addr[39747] = 1933985310;
assign addr[39748] = 1925596340;
assign addr[39749] = 1917054681;
assign addr[39750] = 1908361011;
assign addr[39751] = 1899516021;
assign addr[39752] = 1890520410;
assign addr[39753] = 1881374892;
assign addr[39754] = 1872080193;
assign addr[39755] = 1862637049;
assign addr[39756] = 1853046210;
assign addr[39757] = 1843308435;
assign addr[39758] = 1833424497;
assign addr[39759] = 1823395180;
assign addr[39760] = 1813221279;
assign addr[39761] = 1802903601;
assign addr[39762] = 1792442963;
assign addr[39763] = 1781840195;
assign addr[39764] = 1771096139;
assign addr[39765] = 1760211645;
assign addr[39766] = 1749187577;
assign addr[39767] = 1738024810;
assign addr[39768] = 1726724227;
assign addr[39769] = 1715286726;
assign addr[39770] = 1703713213;
assign addr[39771] = 1692004606;
assign addr[39772] = 1680161834;
assign addr[39773] = 1668185835;
assign addr[39774] = 1656077559;
assign addr[39775] = 1643837966;
assign addr[39776] = 1631468027;
assign addr[39777] = 1618968722;
assign addr[39778] = 1606341043;
assign addr[39779] = 1593585992;
assign addr[39780] = 1580704578;
assign addr[39781] = 1567697824;
assign addr[39782] = 1554566762;
assign addr[39783] = 1541312431;
assign addr[39784] = 1527935884;
assign addr[39785] = 1514438181;
assign addr[39786] = 1500820393;
assign addr[39787] = 1487083598;
assign addr[39788] = 1473228887;
assign addr[39789] = 1459257358;
assign addr[39790] = 1445170118;
assign addr[39791] = 1430968286;
assign addr[39792] = 1416652986;
assign addr[39793] = 1402225355;
assign addr[39794] = 1387686535;
assign addr[39795] = 1373037681;
assign addr[39796] = 1358279953;
assign addr[39797] = 1343414522;
assign addr[39798] = 1328442566;
assign addr[39799] = 1313365273;
assign addr[39800] = 1298183838;
assign addr[39801] = 1282899464;
assign addr[39802] = 1267513365;
assign addr[39803] = 1252026760;
assign addr[39804] = 1236440877;
assign addr[39805] = 1220756951;
assign addr[39806] = 1204976227;
assign addr[39807] = 1189099956;
assign addr[39808] = 1173129396;
assign addr[39809] = 1157065814;
assign addr[39810] = 1140910484;
assign addr[39811] = 1124664687;
assign addr[39812] = 1108329711;
assign addr[39813] = 1091906851;
assign addr[39814] = 1075397409;
assign addr[39815] = 1058802695;
assign addr[39816] = 1042124025;
assign addr[39817] = 1025362720;
assign addr[39818] = 1008520110;
assign addr[39819] = 991597531;
assign addr[39820] = 974596324;
assign addr[39821] = 957517838;
assign addr[39822] = 940363427;
assign addr[39823] = 923134450;
assign addr[39824] = 905832274;
assign addr[39825] = 888458272;
assign addr[39826] = 871013820;
assign addr[39827] = 853500302;
assign addr[39828] = 835919107;
assign addr[39829] = 818271628;
assign addr[39830] = 800559266;
assign addr[39831] = 782783424;
assign addr[39832] = 764945512;
assign addr[39833] = 747046944;
assign addr[39834] = 729089140;
assign addr[39835] = 711073524;
assign addr[39836] = 693001525;
assign addr[39837] = 674874574;
assign addr[39838] = 656694110;
assign addr[39839] = 638461574;
assign addr[39840] = 620178412;
assign addr[39841] = 601846074;
assign addr[39842] = 583466013;
assign addr[39843] = 565039687;
assign addr[39844] = 546568556;
assign addr[39845] = 528054086;
assign addr[39846] = 509497745;
assign addr[39847] = 490901003;
assign addr[39848] = 472265336;
assign addr[39849] = 453592221;
assign addr[39850] = 434883140;
assign addr[39851] = 416139574;
assign addr[39852] = 397363011;
assign addr[39853] = 378554940;
assign addr[39854] = 359716852;
assign addr[39855] = 340850240;
assign addr[39856] = 321956601;
assign addr[39857] = 303037433;
assign addr[39858] = 284094236;
assign addr[39859] = 265128512;
assign addr[39860] = 246141764;
assign addr[39861] = 227135500;
assign addr[39862] = 208111224;
assign addr[39863] = 189070447;
assign addr[39864] = 170014678;
assign addr[39865] = 150945428;
assign addr[39866] = 131864208;
assign addr[39867] = 112772533;
assign addr[39868] = 93671915;
assign addr[39869] = 74563870;
assign addr[39870] = 55449912;
assign addr[39871] = 36331557;
assign addr[39872] = 17210322;
assign addr[39873] = -1912278;
assign addr[39874] = -21034727;
assign addr[39875] = -40155507;
assign addr[39876] = -59273104;
assign addr[39877] = -78386000;
assign addr[39878] = -97492681;
assign addr[39879] = -116591632;
assign addr[39880] = -135681337;
assign addr[39881] = -154760284;
assign addr[39882] = -173826959;
assign addr[39883] = -192879850;
assign addr[39884] = -211917448;
assign addr[39885] = -230938242;
assign addr[39886] = -249940723;
assign addr[39887] = -268923386;
assign addr[39888] = -287884725;
assign addr[39889] = -306823237;
assign addr[39890] = -325737419;
assign addr[39891] = -344625773;
assign addr[39892] = -363486799;
assign addr[39893] = -382319004;
assign addr[39894] = -401120892;
assign addr[39895] = -419890975;
assign addr[39896] = -438627762;
assign addr[39897] = -457329769;
assign addr[39898] = -475995513;
assign addr[39899] = -494623513;
assign addr[39900] = -513212292;
assign addr[39901] = -531760377;
assign addr[39902] = -550266296;
assign addr[39903] = -568728583;
assign addr[39904] = -587145773;
assign addr[39905] = -605516406;
assign addr[39906] = -623839025;
assign addr[39907] = -642112178;
assign addr[39908] = -660334415;
assign addr[39909] = -678504291;
assign addr[39910] = -696620367;
assign addr[39911] = -714681204;
assign addr[39912] = -732685372;
assign addr[39913] = -750631442;
assign addr[39914] = -768517992;
assign addr[39915] = -786343603;
assign addr[39916] = -804106861;
assign addr[39917] = -821806359;
assign addr[39918] = -839440693;
assign addr[39919] = -857008464;
assign addr[39920] = -874508280;
assign addr[39921] = -891938752;
assign addr[39922] = -909298500;
assign addr[39923] = -926586145;
assign addr[39924] = -943800318;
assign addr[39925] = -960939653;
assign addr[39926] = -978002791;
assign addr[39927] = -994988380;
assign addr[39928] = -1011895073;
assign addr[39929] = -1028721528;
assign addr[39930] = -1045466412;
assign addr[39931] = -1062128397;
assign addr[39932] = -1078706161;
assign addr[39933] = -1095198391;
assign addr[39934] = -1111603778;
assign addr[39935] = -1127921022;
assign addr[39936] = -1144148829;
assign addr[39937] = -1160285911;
assign addr[39938] = -1176330990;
assign addr[39939] = -1192282793;
assign addr[39940] = -1208140056;
assign addr[39941] = -1223901520;
assign addr[39942] = -1239565936;
assign addr[39943] = -1255132063;
assign addr[39944] = -1270598665;
assign addr[39945] = -1285964516;
assign addr[39946] = -1301228398;
assign addr[39947] = -1316389101;
assign addr[39948] = -1331445422;
assign addr[39949] = -1346396168;
assign addr[39950] = -1361240152;
assign addr[39951] = -1375976199;
assign addr[39952] = -1390603139;
assign addr[39953] = -1405119813;
assign addr[39954] = -1419525069;
assign addr[39955] = -1433817766;
assign addr[39956] = -1447996770;
assign addr[39957] = -1462060956;
assign addr[39958] = -1476009210;
assign addr[39959] = -1489840425;
assign addr[39960] = -1503553506;
assign addr[39961] = -1517147363;
assign addr[39962] = -1530620920;
assign addr[39963] = -1543973108;
assign addr[39964] = -1557202869;
assign addr[39965] = -1570309153;
assign addr[39966] = -1583290921;
assign addr[39967] = -1596147143;
assign addr[39968] = -1608876801;
assign addr[39969] = -1621478885;
assign addr[39970] = -1633952396;
assign addr[39971] = -1646296344;
assign addr[39972] = -1658509750;
assign addr[39973] = -1670591647;
assign addr[39974] = -1682541077;
assign addr[39975] = -1694357091;
assign addr[39976] = -1706038753;
assign addr[39977] = -1717585136;
assign addr[39978] = -1728995326;
assign addr[39979] = -1740268417;
assign addr[39980] = -1751403515;
assign addr[39981] = -1762399737;
assign addr[39982] = -1773256212;
assign addr[39983] = -1783972079;
assign addr[39984] = -1794546487;
assign addr[39985] = -1804978599;
assign addr[39986] = -1815267588;
assign addr[39987] = -1825412636;
assign addr[39988] = -1835412941;
assign addr[39989] = -1845267708;
assign addr[39990] = -1854976157;
assign addr[39991] = -1864537518;
assign addr[39992] = -1873951032;
assign addr[39993] = -1883215953;
assign addr[39994] = -1892331547;
assign addr[39995] = -1901297091;
assign addr[39996] = -1910111873;
assign addr[39997] = -1918775195;
assign addr[39998] = -1927286370;
assign addr[39999] = -1935644723;
assign addr[40000] = -1943849591;
assign addr[40001] = -1951900324;
assign addr[40002] = -1959796283;
assign addr[40003] = -1967536842;
assign addr[40004] = -1975121388;
assign addr[40005] = -1982549318;
assign addr[40006] = -1989820044;
assign addr[40007] = -1996932990;
assign addr[40008] = -2003887591;
assign addr[40009] = -2010683297;
assign addr[40010] = -2017319567;
assign addr[40011] = -2023795876;
assign addr[40012] = -2030111710;
assign addr[40013] = -2036266570;
assign addr[40014] = -2042259965;
assign addr[40015] = -2048091422;
assign addr[40016] = -2053760478;
assign addr[40017] = -2059266683;
assign addr[40018] = -2064609600;
assign addr[40019] = -2069788807;
assign addr[40020] = -2074803892;
assign addr[40021] = -2079654458;
assign addr[40022] = -2084340120;
assign addr[40023] = -2088860507;
assign addr[40024] = -2093215260;
assign addr[40025] = -2097404033;
assign addr[40026] = -2101426496;
assign addr[40027] = -2105282327;
assign addr[40028] = -2108971223;
assign addr[40029] = -2112492891;
assign addr[40030] = -2115847050;
assign addr[40031] = -2119033436;
assign addr[40032] = -2122051796;
assign addr[40033] = -2124901890;
assign addr[40034] = -2127583492;
assign addr[40035] = -2130096389;
assign addr[40036] = -2132440383;
assign addr[40037] = -2134615288;
assign addr[40038] = -2136620930;
assign addr[40039] = -2138457152;
assign addr[40040] = -2140123807;
assign addr[40041] = -2141620763;
assign addr[40042] = -2142947902;
assign addr[40043] = -2144105118;
assign addr[40044] = -2145092320;
assign addr[40045] = -2145909429;
assign addr[40046] = -2146556380;
assign addr[40047] = -2147033123;
assign addr[40048] = -2147339619;
assign addr[40049] = -2147475844;
assign addr[40050] = -2147441787;
assign addr[40051] = -2147237452;
assign addr[40052] = -2146862854;
assign addr[40053] = -2146318022;
assign addr[40054] = -2145603001;
assign addr[40055] = -2144717846;
assign addr[40056] = -2143662628;
assign addr[40057] = -2142437431;
assign addr[40058] = -2141042352;
assign addr[40059] = -2139477502;
assign addr[40060] = -2137743003;
assign addr[40061] = -2135838995;
assign addr[40062] = -2133765628;
assign addr[40063] = -2131523066;
assign addr[40064] = -2129111488;
assign addr[40065] = -2126531084;
assign addr[40066] = -2123782059;
assign addr[40067] = -2120864631;
assign addr[40068] = -2117779031;
assign addr[40069] = -2114525505;
assign addr[40070] = -2111104309;
assign addr[40071] = -2107515716;
assign addr[40072] = -2103760010;
assign addr[40073] = -2099837489;
assign addr[40074] = -2095748463;
assign addr[40075] = -2091493257;
assign addr[40076] = -2087072209;
assign addr[40077] = -2082485668;
assign addr[40078] = -2077733999;
assign addr[40079] = -2072817579;
assign addr[40080] = -2067736796;
assign addr[40081] = -2062492055;
assign addr[40082] = -2057083771;
assign addr[40083] = -2051512372;
assign addr[40084] = -2045778302;
assign addr[40085] = -2039882013;
assign addr[40086] = -2033823974;
assign addr[40087] = -2027604666;
assign addr[40088] = -2021224581;
assign addr[40089] = -2014684225;
assign addr[40090] = -2007984117;
assign addr[40091] = -2001124788;
assign addr[40092] = -1994106782;
assign addr[40093] = -1986930656;
assign addr[40094] = -1979596978;
assign addr[40095] = -1972106330;
assign addr[40096] = -1964459306;
assign addr[40097] = -1956656513;
assign addr[40098] = -1948698568;
assign addr[40099] = -1940586104;
assign addr[40100] = -1932319763;
assign addr[40101] = -1923900201;
assign addr[40102] = -1915328086;
assign addr[40103] = -1906604097;
assign addr[40104] = -1897728925;
assign addr[40105] = -1888703276;
assign addr[40106] = -1879527863;
assign addr[40107] = -1870203416;
assign addr[40108] = -1860730673;
assign addr[40109] = -1851110385;
assign addr[40110] = -1841343316;
assign addr[40111] = -1831430239;
assign addr[40112] = -1821371941;
assign addr[40113] = -1811169220;
assign addr[40114] = -1800822883;
assign addr[40115] = -1790333753;
assign addr[40116] = -1779702660;
assign addr[40117] = -1768930447;
assign addr[40118] = -1758017969;
assign addr[40119] = -1746966091;
assign addr[40120] = -1735775690;
assign addr[40121] = -1724447652;
assign addr[40122] = -1712982875;
assign addr[40123] = -1701382270;
assign addr[40124] = -1689646755;
assign addr[40125] = -1677777262;
assign addr[40126] = -1665774731;
assign addr[40127] = -1653640115;
assign addr[40128] = -1641374375;
assign addr[40129] = -1628978484;
assign addr[40130] = -1616453425;
assign addr[40131] = -1603800191;
assign addr[40132] = -1591019785;
assign addr[40133] = -1578113222;
assign addr[40134] = -1565081523;
assign addr[40135] = -1551925723;
assign addr[40136] = -1538646865;
assign addr[40137] = -1525246002;
assign addr[40138] = -1511724196;
assign addr[40139] = -1498082520;
assign addr[40140] = -1484322054;
assign addr[40141] = -1470443891;
assign addr[40142] = -1456449131;
assign addr[40143] = -1442338884;
assign addr[40144] = -1428114267;
assign addr[40145] = -1413776410;
assign addr[40146] = -1399326449;
assign addr[40147] = -1384765530;
assign addr[40148] = -1370094808;
assign addr[40149] = -1355315445;
assign addr[40150] = -1340428615;
assign addr[40151] = -1325435496;
assign addr[40152] = -1310337279;
assign addr[40153] = -1295135159;
assign addr[40154] = -1279830344;
assign addr[40155] = -1264424045;
assign addr[40156] = -1248917486;
assign addr[40157] = -1233311895;
assign addr[40158] = -1217608510;
assign addr[40159] = -1201808576;
assign addr[40160] = -1185913346;
assign addr[40161] = -1169924081;
assign addr[40162] = -1153842047;
assign addr[40163] = -1137668521;
assign addr[40164] = -1121404785;
assign addr[40165] = -1105052128;
assign addr[40166] = -1088611847;
assign addr[40167] = -1072085246;
assign addr[40168] = -1055473635;
assign addr[40169] = -1038778332;
assign addr[40170] = -1022000660;
assign addr[40171] = -1005141949;
assign addr[40172] = -988203537;
assign addr[40173] = -971186766;
assign addr[40174] = -954092986;
assign addr[40175] = -936923553;
assign addr[40176] = -919679827;
assign addr[40177] = -902363176;
assign addr[40178] = -884974973;
assign addr[40179] = -867516597;
assign addr[40180] = -849989433;
assign addr[40181] = -832394869;
assign addr[40182] = -814734301;
assign addr[40183] = -797009130;
assign addr[40184] = -779220762;
assign addr[40185] = -761370605;
assign addr[40186] = -743460077;
assign addr[40187] = -725490597;
assign addr[40188] = -707463589;
assign addr[40189] = -689380485;
assign addr[40190] = -671242716;
assign addr[40191] = -653051723;
assign addr[40192] = -634808946;
assign addr[40193] = -616515832;
assign addr[40194] = -598173833;
assign addr[40195] = -579784402;
assign addr[40196] = -561348998;
assign addr[40197] = -542869083;
assign addr[40198] = -524346121;
assign addr[40199] = -505781581;
assign addr[40200] = -487176937;
assign addr[40201] = -468533662;
assign addr[40202] = -449853235;
assign addr[40203] = -431137138;
assign addr[40204] = -412386854;
assign addr[40205] = -393603870;
assign addr[40206] = -374789676;
assign addr[40207] = -355945764;
assign addr[40208] = -337073627;
assign addr[40209] = -318174762;
assign addr[40210] = -299250668;
assign addr[40211] = -280302845;
assign addr[40212] = -261332796;
assign addr[40213] = -242342025;
assign addr[40214] = -223332037;
assign addr[40215] = -204304341;
assign addr[40216] = -185260444;
assign addr[40217] = -166201858;
assign addr[40218] = -147130093;
assign addr[40219] = -128046661;
assign addr[40220] = -108953076;
assign addr[40221] = -89850852;
assign addr[40222] = -70741503;
assign addr[40223] = -51626544;
assign addr[40224] = -32507492;
assign addr[40225] = -13385863;
assign addr[40226] = 5736829;
assign addr[40227] = 24859065;
assign addr[40228] = 43979330;
assign addr[40229] = 63096108;
assign addr[40230] = 82207882;
assign addr[40231] = 101313138;
assign addr[40232] = 120410361;
assign addr[40233] = 139498035;
assign addr[40234] = 158574649;
assign addr[40235] = 177638688;
assign addr[40236] = 196688642;
assign addr[40237] = 215722999;
assign addr[40238] = 234740251;
assign addr[40239] = 253738890;
assign addr[40240] = 272717408;
assign addr[40241] = 291674302;
assign addr[40242] = 310608068;
assign addr[40243] = 329517204;
assign addr[40244] = 348400212;
assign addr[40245] = 367255594;
assign addr[40246] = 386081854;
assign addr[40247] = 404877501;
assign addr[40248] = 423641043;
assign addr[40249] = 442370993;
assign addr[40250] = 461065866;
assign addr[40251] = 479724180;
assign addr[40252] = 498344454;
assign addr[40253] = 516925212;
assign addr[40254] = 535464981;
assign addr[40255] = 553962291;
assign addr[40256] = 572415676;
assign addr[40257] = 590823671;
assign addr[40258] = 609184818;
assign addr[40259] = 627497660;
assign addr[40260] = 645760745;
assign addr[40261] = 663972625;
assign addr[40262] = 682131857;
assign addr[40263] = 700236999;
assign addr[40264] = 718286617;
assign addr[40265] = 736279279;
assign addr[40266] = 754213559;
assign addr[40267] = 772088034;
assign addr[40268] = 789901288;
assign addr[40269] = 807651907;
assign addr[40270] = 825338484;
assign addr[40271] = 842959617;
assign addr[40272] = 860513908;
assign addr[40273] = 877999966;
assign addr[40274] = 895416404;
assign addr[40275] = 912761841;
assign addr[40276] = 930034901;
assign addr[40277] = 947234215;
assign addr[40278] = 964358420;
assign addr[40279] = 981406156;
assign addr[40280] = 998376073;
assign addr[40281] = 1015266825;
assign addr[40282] = 1032077073;
assign addr[40283] = 1048805483;
assign addr[40284] = 1065450729;
assign addr[40285] = 1082011492;
assign addr[40286] = 1098486458;
assign addr[40287] = 1114874320;
assign addr[40288] = 1131173780;
assign addr[40289] = 1147383544;
assign addr[40290] = 1163502328;
assign addr[40291] = 1179528853;
assign addr[40292] = 1195461849;
assign addr[40293] = 1211300053;
assign addr[40294] = 1227042207;
assign addr[40295] = 1242687064;
assign addr[40296] = 1258233384;
assign addr[40297] = 1273679934;
assign addr[40298] = 1289025489;
assign addr[40299] = 1304268832;
assign addr[40300] = 1319408754;
assign addr[40301] = 1334444055;
assign addr[40302] = 1349373543;
assign addr[40303] = 1364196034;
assign addr[40304] = 1378910353;
assign addr[40305] = 1393515332;
assign addr[40306] = 1408009814;
assign addr[40307] = 1422392650;
assign addr[40308] = 1436662698;
assign addr[40309] = 1450818828;
assign addr[40310] = 1464859917;
assign addr[40311] = 1478784851;
assign addr[40312] = 1492592527;
assign addr[40313] = 1506281850;
assign addr[40314] = 1519851733;
assign addr[40315] = 1533301101;
assign addr[40316] = 1546628888;
assign addr[40317] = 1559834037;
assign addr[40318] = 1572915501;
assign addr[40319] = 1585872242;
assign addr[40320] = 1598703233;
assign addr[40321] = 1611407456;
assign addr[40322] = 1623983905;
assign addr[40323] = 1636431582;
assign addr[40324] = 1648749499;
assign addr[40325] = 1660936681;
assign addr[40326] = 1672992161;
assign addr[40327] = 1684914983;
assign addr[40328] = 1696704201;
assign addr[40329] = 1708358881;
assign addr[40330] = 1719878099;
assign addr[40331] = 1731260941;
assign addr[40332] = 1742506504;
assign addr[40333] = 1753613897;
assign addr[40334] = 1764582240;
assign addr[40335] = 1775410662;
assign addr[40336] = 1786098304;
assign addr[40337] = 1796644320;
assign addr[40338] = 1807047873;
assign addr[40339] = 1817308138;
assign addr[40340] = 1827424302;
assign addr[40341] = 1837395562;
assign addr[40342] = 1847221128;
assign addr[40343] = 1856900221;
assign addr[40344] = 1866432072;
assign addr[40345] = 1875815927;
assign addr[40346] = 1885051042;
assign addr[40347] = 1894136683;
assign addr[40348] = 1903072131;
assign addr[40349] = 1911856677;
assign addr[40350] = 1920489624;
assign addr[40351] = 1928970288;
assign addr[40352] = 1937297997;
assign addr[40353] = 1945472089;
assign addr[40354] = 1953491918;
assign addr[40355] = 1961356847;
assign addr[40356] = 1969066252;
assign addr[40357] = 1976619522;
assign addr[40358] = 1984016058;
assign addr[40359] = 1991255274;
assign addr[40360] = 1998336596;
assign addr[40361] = 2005259462;
assign addr[40362] = 2012023322;
assign addr[40363] = 2018627642;
assign addr[40364] = 2025071897;
assign addr[40365] = 2031355576;
assign addr[40366] = 2037478181;
assign addr[40367] = 2043439226;
assign addr[40368] = 2049238240;
assign addr[40369] = 2054874761;
assign addr[40370] = 2060348343;
assign addr[40371] = 2065658552;
assign addr[40372] = 2070804967;
assign addr[40373] = 2075787180;
assign addr[40374] = 2080604795;
assign addr[40375] = 2085257431;
assign addr[40376] = 2089744719;
assign addr[40377] = 2094066304;
assign addr[40378] = 2098221841;
assign addr[40379] = 2102211002;
assign addr[40380] = 2106033471;
assign addr[40381] = 2109688944;
assign addr[40382] = 2113177132;
assign addr[40383] = 2116497758;
assign addr[40384] = 2119650558;
assign addr[40385] = 2122635283;
assign addr[40386] = 2125451696;
assign addr[40387] = 2128099574;
assign addr[40388] = 2130578706;
assign addr[40389] = 2132888897;
assign addr[40390] = 2135029962;
assign addr[40391] = 2137001733;
assign addr[40392] = 2138804053;
assign addr[40393] = 2140436778;
assign addr[40394] = 2141899780;
assign addr[40395] = 2143192942;
assign addr[40396] = 2144316162;
assign addr[40397] = 2145269351;
assign addr[40398] = 2146052433;
assign addr[40399] = 2146665347;
assign addr[40400] = 2147108043;
assign addr[40401] = 2147380486;
assign addr[40402] = 2147482655;
assign addr[40403] = 2147414542;
assign addr[40404] = 2147176152;
assign addr[40405] = 2146767505;
assign addr[40406] = 2146188631;
assign addr[40407] = 2145439578;
assign addr[40408] = 2144520405;
assign addr[40409] = 2143431184;
assign addr[40410] = 2142172003;
assign addr[40411] = 2140742960;
assign addr[40412] = 2139144169;
assign addr[40413] = 2137375758;
assign addr[40414] = 2135437865;
assign addr[40415] = 2133330646;
assign addr[40416] = 2131054266;
assign addr[40417] = 2128608907;
assign addr[40418] = 2125994762;
assign addr[40419] = 2123212038;
assign addr[40420] = 2120260957;
assign addr[40421] = 2117141752;
assign addr[40422] = 2113854671;
assign addr[40423] = 2110399974;
assign addr[40424] = 2106777935;
assign addr[40425] = 2102988841;
assign addr[40426] = 2099032994;
assign addr[40427] = 2094910706;
assign addr[40428] = 2090622304;
assign addr[40429] = 2086168128;
assign addr[40430] = 2081548533;
assign addr[40431] = 2076763883;
assign addr[40432] = 2071814558;
assign addr[40433] = 2066700952;
assign addr[40434] = 2061423468;
assign addr[40435] = 2055982526;
assign addr[40436] = 2050378558;
assign addr[40437] = 2044612007;
assign addr[40438] = 2038683330;
assign addr[40439] = 2032592999;
assign addr[40440] = 2026341495;
assign addr[40441] = 2019929315;
assign addr[40442] = 2013356967;
assign addr[40443] = 2006624971;
assign addr[40444] = 1999733863;
assign addr[40445] = 1992684188;
assign addr[40446] = 1985476506;
assign addr[40447] = 1978111387;
assign addr[40448] = 1970589416;
assign addr[40449] = 1962911189;
assign addr[40450] = 1955077316;
assign addr[40451] = 1947088417;
assign addr[40452] = 1938945125;
assign addr[40453] = 1930648088;
assign addr[40454] = 1922197961;
assign addr[40455] = 1913595416;
assign addr[40456] = 1904841135;
assign addr[40457] = 1895935811;
assign addr[40458] = 1886880151;
assign addr[40459] = 1877674873;
assign addr[40460] = 1868320707;
assign addr[40461] = 1858818395;
assign addr[40462] = 1849168689;
assign addr[40463] = 1839372356;
assign addr[40464] = 1829430172;
assign addr[40465] = 1819342925;
assign addr[40466] = 1809111415;
assign addr[40467] = 1798736454;
assign addr[40468] = 1788218865;
assign addr[40469] = 1777559480;
assign addr[40470] = 1766759146;
assign addr[40471] = 1755818718;
assign addr[40472] = 1744739065;
assign addr[40473] = 1733521064;
assign addr[40474] = 1722165606;
assign addr[40475] = 1710673591;
assign addr[40476] = 1699045930;
assign addr[40477] = 1687283545;
assign addr[40478] = 1675387369;
assign addr[40479] = 1663358344;
assign addr[40480] = 1651197426;
assign addr[40481] = 1638905577;
assign addr[40482] = 1626483774;
assign addr[40483] = 1613933000;
assign addr[40484] = 1601254251;
assign addr[40485] = 1588448533;
assign addr[40486] = 1575516860;
assign addr[40487] = 1562460258;
assign addr[40488] = 1549279763;
assign addr[40489] = 1535976419;
assign addr[40490] = 1522551282;
assign addr[40491] = 1509005416;
assign addr[40492] = 1495339895;
assign addr[40493] = 1481555802;
assign addr[40494] = 1467654232;
assign addr[40495] = 1453636285;
assign addr[40496] = 1439503074;
assign addr[40497] = 1425255719;
assign addr[40498] = 1410895350;
assign addr[40499] = 1396423105;
assign addr[40500] = 1381840133;
assign addr[40501] = 1367147589;
assign addr[40502] = 1352346639;
assign addr[40503] = 1337438456;
assign addr[40504] = 1322424222;
assign addr[40505] = 1307305128;
assign addr[40506] = 1292082373;
assign addr[40507] = 1276757164;
assign addr[40508] = 1261330715;
assign addr[40509] = 1245804251;
assign addr[40510] = 1230179002;
assign addr[40511] = 1214456207;
assign addr[40512] = 1198637114;
assign addr[40513] = 1182722976;
assign addr[40514] = 1166715055;
assign addr[40515] = 1150614620;
assign addr[40516] = 1134422949;
assign addr[40517] = 1118141326;
assign addr[40518] = 1101771040;
assign addr[40519] = 1085313391;
assign addr[40520] = 1068769683;
assign addr[40521] = 1052141228;
assign addr[40522] = 1035429345;
assign addr[40523] = 1018635358;
assign addr[40524] = 1001760600;
assign addr[40525] = 984806408;
assign addr[40526] = 967774128;
assign addr[40527] = 950665109;
assign addr[40528] = 933480707;
assign addr[40529] = 916222287;
assign addr[40530] = 898891215;
assign addr[40531] = 881488868;
assign addr[40532] = 864016623;
assign addr[40533] = 846475867;
assign addr[40534] = 828867991;
assign addr[40535] = 811194391;
assign addr[40536] = 793456467;
assign addr[40537] = 775655628;
assign addr[40538] = 757793284;
assign addr[40539] = 739870851;
assign addr[40540] = 721889752;
assign addr[40541] = 703851410;
assign addr[40542] = 685757258;
assign addr[40543] = 667608730;
assign addr[40544] = 649407264;
assign addr[40545] = 631154304;
assign addr[40546] = 612851297;
assign addr[40547] = 594499695;
assign addr[40548] = 576100953;
assign addr[40549] = 557656529;
assign addr[40550] = 539167887;
assign addr[40551] = 520636492;
assign addr[40552] = 502063814;
assign addr[40553] = 483451325;
assign addr[40554] = 464800501;
assign addr[40555] = 446112822;
assign addr[40556] = 427389768;
assign addr[40557] = 408632825;
assign addr[40558] = 389843480;
assign addr[40559] = 371023223;
assign addr[40560] = 352173546;
assign addr[40561] = 333295944;
assign addr[40562] = 314391913;
assign addr[40563] = 295462954;
assign addr[40564] = 276510565;
assign addr[40565] = 257536251;
assign addr[40566] = 238541516;
assign addr[40567] = 219527866;
assign addr[40568] = 200496809;
assign addr[40569] = 181449854;
assign addr[40570] = 162388511;
assign addr[40571] = 143314291;
assign addr[40572] = 124228708;
assign addr[40573] = 105133274;
assign addr[40574] = 86029503;
assign addr[40575] = 66918911;
assign addr[40576] = 47803013;
assign addr[40577] = 28683324;
assign addr[40578] = 9561361;
assign addr[40579] = -9561361;
assign addr[40580] = -28683324;
assign addr[40581] = -47803013;
assign addr[40582] = -66918911;
assign addr[40583] = -86029503;
assign addr[40584] = -105133274;
assign addr[40585] = -124228708;
assign addr[40586] = -143314291;
assign addr[40587] = -162388511;
assign addr[40588] = -181449854;
assign addr[40589] = -200496809;
assign addr[40590] = -219527866;
assign addr[40591] = -238541516;
assign addr[40592] = -257536251;
assign addr[40593] = -276510565;
assign addr[40594] = -295462953;
assign addr[40595] = -314391913;
assign addr[40596] = -333295944;
assign addr[40597] = -352173546;
assign addr[40598] = -371023223;
assign addr[40599] = -389843480;
assign addr[40600] = -408632825;
assign addr[40601] = -427389768;
assign addr[40602] = -446112822;
assign addr[40603] = -464800501;
assign addr[40604] = -483451325;
assign addr[40605] = -502063814;
assign addr[40606] = -520636492;
assign addr[40607] = -539167887;
assign addr[40608] = -557656529;
assign addr[40609] = -576100953;
assign addr[40610] = -594499695;
assign addr[40611] = -612851297;
assign addr[40612] = -631154304;
assign addr[40613] = -649407264;
assign addr[40614] = -667608730;
assign addr[40615] = -685757258;
assign addr[40616] = -703851410;
assign addr[40617] = -721889752;
assign addr[40618] = -739870851;
assign addr[40619] = -757793284;
assign addr[40620] = -775655628;
assign addr[40621] = -793456467;
assign addr[40622] = -811194391;
assign addr[40623] = -828867991;
assign addr[40624] = -846475867;
assign addr[40625] = -864016623;
assign addr[40626] = -881488868;
assign addr[40627] = -898891215;
assign addr[40628] = -916222287;
assign addr[40629] = -933480707;
assign addr[40630] = -950665109;
assign addr[40631] = -967774128;
assign addr[40632] = -984806408;
assign addr[40633] = -1001760600;
assign addr[40634] = -1018635358;
assign addr[40635] = -1035429345;
assign addr[40636] = -1052141228;
assign addr[40637] = -1068769683;
assign addr[40638] = -1085313391;
assign addr[40639] = -1101771040;
assign addr[40640] = -1118141326;
assign addr[40641] = -1134422949;
assign addr[40642] = -1150614620;
assign addr[40643] = -1166715055;
assign addr[40644] = -1182722976;
assign addr[40645] = -1198637114;
assign addr[40646] = -1214456207;
assign addr[40647] = -1230179002;
assign addr[40648] = -1245804251;
assign addr[40649] = -1261330715;
assign addr[40650] = -1276757164;
assign addr[40651] = -1292082373;
assign addr[40652] = -1307305128;
assign addr[40653] = -1322424222;
assign addr[40654] = -1337438456;
assign addr[40655] = -1352346639;
assign addr[40656] = -1367147589;
assign addr[40657] = -1381840133;
assign addr[40658] = -1396423105;
assign addr[40659] = -1410895350;
assign addr[40660] = -1425255719;
assign addr[40661] = -1439503074;
assign addr[40662] = -1453636285;
assign addr[40663] = -1467654232;
assign addr[40664] = -1481555802;
assign addr[40665] = -1495339895;
assign addr[40666] = -1509005416;
assign addr[40667] = -1522551282;
assign addr[40668] = -1535976419;
assign addr[40669] = -1549279763;
assign addr[40670] = -1562460258;
assign addr[40671] = -1575516860;
assign addr[40672] = -1588448533;
assign addr[40673] = -1601254251;
assign addr[40674] = -1613933000;
assign addr[40675] = -1626483774;
assign addr[40676] = -1638905577;
assign addr[40677] = -1651197426;
assign addr[40678] = -1663358344;
assign addr[40679] = -1675387369;
assign addr[40680] = -1687283545;
assign addr[40681] = -1699045930;
assign addr[40682] = -1710673591;
assign addr[40683] = -1722165606;
assign addr[40684] = -1733521064;
assign addr[40685] = -1744739065;
assign addr[40686] = -1755818718;
assign addr[40687] = -1766759146;
assign addr[40688] = -1777559480;
assign addr[40689] = -1788218865;
assign addr[40690] = -1798736454;
assign addr[40691] = -1809111415;
assign addr[40692] = -1819342925;
assign addr[40693] = -1829430172;
assign addr[40694] = -1839372356;
assign addr[40695] = -1849168689;
assign addr[40696] = -1858818395;
assign addr[40697] = -1868320707;
assign addr[40698] = -1877674873;
assign addr[40699] = -1886880151;
assign addr[40700] = -1895935811;
assign addr[40701] = -1904841135;
assign addr[40702] = -1913595416;
assign addr[40703] = -1922197961;
assign addr[40704] = -1930648088;
assign addr[40705] = -1938945125;
assign addr[40706] = -1947088417;
assign addr[40707] = -1955077316;
assign addr[40708] = -1962911189;
assign addr[40709] = -1970589416;
assign addr[40710] = -1978111387;
assign addr[40711] = -1985476506;
assign addr[40712] = -1992684188;
assign addr[40713] = -1999733863;
assign addr[40714] = -2006624971;
assign addr[40715] = -2013356967;
assign addr[40716] = -2019929315;
assign addr[40717] = -2026341495;
assign addr[40718] = -2032592999;
assign addr[40719] = -2038683330;
assign addr[40720] = -2044612007;
assign addr[40721] = -2050378558;
assign addr[40722] = -2055982526;
assign addr[40723] = -2061423468;
assign addr[40724] = -2066700952;
assign addr[40725] = -2071814558;
assign addr[40726] = -2076763883;
assign addr[40727] = -2081548533;
assign addr[40728] = -2086168128;
assign addr[40729] = -2090622304;
assign addr[40730] = -2094910706;
assign addr[40731] = -2099032994;
assign addr[40732] = -2102988841;
assign addr[40733] = -2106777935;
assign addr[40734] = -2110399974;
assign addr[40735] = -2113854671;
assign addr[40736] = -2117141752;
assign addr[40737] = -2120260957;
assign addr[40738] = -2123212038;
assign addr[40739] = -2125994762;
assign addr[40740] = -2128608907;
assign addr[40741] = -2131054266;
assign addr[40742] = -2133330646;
assign addr[40743] = -2135437865;
assign addr[40744] = -2137375758;
assign addr[40745] = -2139144169;
assign addr[40746] = -2140742960;
assign addr[40747] = -2142172003;
assign addr[40748] = -2143431184;
assign addr[40749] = -2144520405;
assign addr[40750] = -2145439578;
assign addr[40751] = -2146188631;
assign addr[40752] = -2146767505;
assign addr[40753] = -2147176152;
assign addr[40754] = -2147414542;
assign addr[40755] = -2147482655;
assign addr[40756] = -2147380486;
assign addr[40757] = -2147108043;
assign addr[40758] = -2146665347;
assign addr[40759] = -2146052433;
assign addr[40760] = -2145269351;
assign addr[40761] = -2144316162;
assign addr[40762] = -2143192942;
assign addr[40763] = -2141899780;
assign addr[40764] = -2140436778;
assign addr[40765] = -2138804053;
assign addr[40766] = -2137001733;
assign addr[40767] = -2135029962;
assign addr[40768] = -2132888897;
assign addr[40769] = -2130578706;
assign addr[40770] = -2128099574;
assign addr[40771] = -2125451696;
assign addr[40772] = -2122635283;
assign addr[40773] = -2119650558;
assign addr[40774] = -2116497758;
assign addr[40775] = -2113177132;
assign addr[40776] = -2109688944;
assign addr[40777] = -2106033471;
assign addr[40778] = -2102211002;
assign addr[40779] = -2098221841;
assign addr[40780] = -2094066304;
assign addr[40781] = -2089744719;
assign addr[40782] = -2085257431;
assign addr[40783] = -2080604795;
assign addr[40784] = -2075787180;
assign addr[40785] = -2070804967;
assign addr[40786] = -2065658552;
assign addr[40787] = -2060348343;
assign addr[40788] = -2054874761;
assign addr[40789] = -2049238240;
assign addr[40790] = -2043439226;
assign addr[40791] = -2037478181;
assign addr[40792] = -2031355576;
assign addr[40793] = -2025071897;
assign addr[40794] = -2018627642;
assign addr[40795] = -2012023322;
assign addr[40796] = -2005259462;
assign addr[40797] = -1998336596;
assign addr[40798] = -1991255274;
assign addr[40799] = -1984016058;
assign addr[40800] = -1976619522;
assign addr[40801] = -1969066252;
assign addr[40802] = -1961356847;
assign addr[40803] = -1953491918;
assign addr[40804] = -1945472089;
assign addr[40805] = -1937297997;
assign addr[40806] = -1928970288;
assign addr[40807] = -1920489624;
assign addr[40808] = -1911856677;
assign addr[40809] = -1903072131;
assign addr[40810] = -1894136683;
assign addr[40811] = -1885051042;
assign addr[40812] = -1875815927;
assign addr[40813] = -1866432072;
assign addr[40814] = -1856900221;
assign addr[40815] = -1847221128;
assign addr[40816] = -1837395562;
assign addr[40817] = -1827424302;
assign addr[40818] = -1817308138;
assign addr[40819] = -1807047873;
assign addr[40820] = -1796644320;
assign addr[40821] = -1786098304;
assign addr[40822] = -1775410662;
assign addr[40823] = -1764582240;
assign addr[40824] = -1753613897;
assign addr[40825] = -1742506504;
assign addr[40826] = -1731260941;
assign addr[40827] = -1719878099;
assign addr[40828] = -1708358881;
assign addr[40829] = -1696704201;
assign addr[40830] = -1684914983;
assign addr[40831] = -1672992161;
assign addr[40832] = -1660936681;
assign addr[40833] = -1648749499;
assign addr[40834] = -1636431582;
assign addr[40835] = -1623983905;
assign addr[40836] = -1611407456;
assign addr[40837] = -1598703233;
assign addr[40838] = -1585872242;
assign addr[40839] = -1572915501;
assign addr[40840] = -1559834037;
assign addr[40841] = -1546628888;
assign addr[40842] = -1533301101;
assign addr[40843] = -1519851733;
assign addr[40844] = -1506281850;
assign addr[40845] = -1492592527;
assign addr[40846] = -1478784851;
assign addr[40847] = -1464859917;
assign addr[40848] = -1450818828;
assign addr[40849] = -1436662698;
assign addr[40850] = -1422392650;
assign addr[40851] = -1408009814;
assign addr[40852] = -1393515332;
assign addr[40853] = -1378910353;
assign addr[40854] = -1364196034;
assign addr[40855] = -1349373543;
assign addr[40856] = -1334444055;
assign addr[40857] = -1319408754;
assign addr[40858] = -1304268832;
assign addr[40859] = -1289025489;
assign addr[40860] = -1273679934;
assign addr[40861] = -1258233384;
assign addr[40862] = -1242687064;
assign addr[40863] = -1227042207;
assign addr[40864] = -1211300053;
assign addr[40865] = -1195461849;
assign addr[40866] = -1179528853;
assign addr[40867] = -1163502328;
assign addr[40868] = -1147383544;
assign addr[40869] = -1131173780;
assign addr[40870] = -1114874320;
assign addr[40871] = -1098486458;
assign addr[40872] = -1082011492;
assign addr[40873] = -1065450729;
assign addr[40874] = -1048805483;
assign addr[40875] = -1032077073;
assign addr[40876] = -1015266825;
assign addr[40877] = -998376073;
assign addr[40878] = -981406156;
assign addr[40879] = -964358420;
assign addr[40880] = -947234215;
assign addr[40881] = -930034901;
assign addr[40882] = -912761841;
assign addr[40883] = -895416404;
assign addr[40884] = -877999966;
assign addr[40885] = -860513908;
assign addr[40886] = -842959617;
assign addr[40887] = -825338484;
assign addr[40888] = -807651907;
assign addr[40889] = -789901288;
assign addr[40890] = -772088034;
assign addr[40891] = -754213559;
assign addr[40892] = -736279279;
assign addr[40893] = -718286617;
assign addr[40894] = -700236999;
assign addr[40895] = -682131857;
assign addr[40896] = -663972625;
assign addr[40897] = -645760745;
assign addr[40898] = -627497660;
assign addr[40899] = -609184818;
assign addr[40900] = -590823671;
assign addr[40901] = -572415676;
assign addr[40902] = -553962291;
assign addr[40903] = -535464981;
assign addr[40904] = -516925212;
assign addr[40905] = -498344454;
assign addr[40906] = -479724180;
assign addr[40907] = -461065866;
assign addr[40908] = -442370993;
assign addr[40909] = -423641043;
assign addr[40910] = -404877501;
assign addr[40911] = -386081854;
assign addr[40912] = -367255594;
assign addr[40913] = -348400212;
assign addr[40914] = -329517204;
assign addr[40915] = -310608068;
assign addr[40916] = -291674302;
assign addr[40917] = -272717408;
assign addr[40918] = -253738890;
assign addr[40919] = -234740251;
assign addr[40920] = -215722999;
assign addr[40921] = -196688642;
assign addr[40922] = -177638688;
assign addr[40923] = -158574649;
assign addr[40924] = -139498035;
assign addr[40925] = -120410361;
assign addr[40926] = -101313138;
assign addr[40927] = -82207882;
assign addr[40928] = -63096108;
assign addr[40929] = -43979330;
assign addr[40930] = -24859065;
assign addr[40931] = -5736829;
assign addr[40932] = 13385863;
assign addr[40933] = 32507492;
assign addr[40934] = 51626544;
assign addr[40935] = 70741503;
assign addr[40936] = 89850852;
assign addr[40937] = 108953076;
assign addr[40938] = 128046661;
assign addr[40939] = 147130093;
assign addr[40940] = 166201858;
assign addr[40941] = 185260444;
assign addr[40942] = 204304341;
assign addr[40943] = 223332037;
assign addr[40944] = 242342025;
assign addr[40945] = 261332796;
assign addr[40946] = 280302845;
assign addr[40947] = 299250668;
assign addr[40948] = 318174762;
assign addr[40949] = 337073627;
assign addr[40950] = 355945764;
assign addr[40951] = 374789676;
assign addr[40952] = 393603870;
assign addr[40953] = 412386854;
assign addr[40954] = 431137138;
assign addr[40955] = 449853235;
assign addr[40956] = 468533662;
assign addr[40957] = 487176937;
assign addr[40958] = 505781581;
assign addr[40959] = 524346121;
assign addr[40960] = 542869083;
assign addr[40961] = 561348998;
assign addr[40962] = 579784402;
assign addr[40963] = 598173833;
assign addr[40964] = 616515832;
assign addr[40965] = 634808946;
assign addr[40966] = 653051723;
assign addr[40967] = 671242716;
assign addr[40968] = 689380485;
assign addr[40969] = 707463589;
assign addr[40970] = 725490597;
assign addr[40971] = 743460077;
assign addr[40972] = 761370605;
assign addr[40973] = 779220762;
assign addr[40974] = 797009130;
assign addr[40975] = 814734301;
assign addr[40976] = 832394869;
assign addr[40977] = 849989433;
assign addr[40978] = 867516597;
assign addr[40979] = 884974973;
assign addr[40980] = 902363176;
assign addr[40981] = 919679827;
assign addr[40982] = 936923553;
assign addr[40983] = 954092986;
assign addr[40984] = 971186766;
assign addr[40985] = 988203537;
assign addr[40986] = 1005141949;
assign addr[40987] = 1022000660;
assign addr[40988] = 1038778332;
assign addr[40989] = 1055473635;
assign addr[40990] = 1072085246;
assign addr[40991] = 1088611847;
assign addr[40992] = 1105052128;
assign addr[40993] = 1121404785;
assign addr[40994] = 1137668521;
assign addr[40995] = 1153842047;
assign addr[40996] = 1169924081;
assign addr[40997] = 1185913346;
assign addr[40998] = 1201808576;
assign addr[40999] = 1217608510;
assign addr[41000] = 1233311895;
assign addr[41001] = 1248917486;
assign addr[41002] = 1264424045;
assign addr[41003] = 1279830344;
assign addr[41004] = 1295135159;
assign addr[41005] = 1310337279;
assign addr[41006] = 1325435496;
assign addr[41007] = 1340428615;
assign addr[41008] = 1355315445;
assign addr[41009] = 1370094808;
assign addr[41010] = 1384765530;
assign addr[41011] = 1399326449;
assign addr[41012] = 1413776410;
assign addr[41013] = 1428114267;
assign addr[41014] = 1442338884;
assign addr[41015] = 1456449131;
assign addr[41016] = 1470443891;
assign addr[41017] = 1484322054;
assign addr[41018] = 1498082520;
assign addr[41019] = 1511724196;
assign addr[41020] = 1525246002;
assign addr[41021] = 1538646865;
assign addr[41022] = 1551925723;
assign addr[41023] = 1565081523;
assign addr[41024] = 1578113222;
assign addr[41025] = 1591019785;
assign addr[41026] = 1603800191;
assign addr[41027] = 1616453425;
assign addr[41028] = 1628978484;
assign addr[41029] = 1641374375;
assign addr[41030] = 1653640115;
assign addr[41031] = 1665774731;
assign addr[41032] = 1677777262;
assign addr[41033] = 1689646755;
assign addr[41034] = 1701382270;
assign addr[41035] = 1712982875;
assign addr[41036] = 1724447652;
assign addr[41037] = 1735775690;
assign addr[41038] = 1746966091;
assign addr[41039] = 1758017969;
assign addr[41040] = 1768930447;
assign addr[41041] = 1779702660;
assign addr[41042] = 1790333753;
assign addr[41043] = 1800822883;
assign addr[41044] = 1811169220;
assign addr[41045] = 1821371941;
assign addr[41046] = 1831430239;
assign addr[41047] = 1841343316;
assign addr[41048] = 1851110385;
assign addr[41049] = 1860730673;
assign addr[41050] = 1870203416;
assign addr[41051] = 1879527863;
assign addr[41052] = 1888703276;
assign addr[41053] = 1897728925;
assign addr[41054] = 1906604097;
assign addr[41055] = 1915328086;
assign addr[41056] = 1923900201;
assign addr[41057] = 1932319763;
assign addr[41058] = 1940586104;
assign addr[41059] = 1948698568;
assign addr[41060] = 1956656513;
assign addr[41061] = 1964459306;
assign addr[41062] = 1972106330;
assign addr[41063] = 1979596978;
assign addr[41064] = 1986930656;
assign addr[41065] = 1994106782;
assign addr[41066] = 2001124788;
assign addr[41067] = 2007984117;
assign addr[41068] = 2014684225;
assign addr[41069] = 2021224581;
assign addr[41070] = 2027604666;
assign addr[41071] = 2033823974;
assign addr[41072] = 2039882013;
assign addr[41073] = 2045778302;
assign addr[41074] = 2051512372;
assign addr[41075] = 2057083771;
assign addr[41076] = 2062492055;
assign addr[41077] = 2067736796;
assign addr[41078] = 2072817579;
assign addr[41079] = 2077733999;
assign addr[41080] = 2082485668;
assign addr[41081] = 2087072209;
assign addr[41082] = 2091493257;
assign addr[41083] = 2095748463;
assign addr[41084] = 2099837489;
assign addr[41085] = 2103760010;
assign addr[41086] = 2107515716;
assign addr[41087] = 2111104309;
assign addr[41088] = 2114525505;
assign addr[41089] = 2117779031;
assign addr[41090] = 2120864631;
assign addr[41091] = 2123782059;
assign addr[41092] = 2126531084;
assign addr[41093] = 2129111488;
assign addr[41094] = 2131523066;
assign addr[41095] = 2133765628;
assign addr[41096] = 2135838995;
assign addr[41097] = 2137743003;
assign addr[41098] = 2139477502;
assign addr[41099] = 2141042352;
assign addr[41100] = 2142437431;
assign addr[41101] = 2143662628;
assign addr[41102] = 2144717846;
assign addr[41103] = 2145603001;
assign addr[41104] = 2146318022;
assign addr[41105] = 2146862854;
assign addr[41106] = 2147237452;
assign addr[41107] = 2147441787;
assign addr[41108] = 2147475844;
assign addr[41109] = 2147339619;
assign addr[41110] = 2147033123;
assign addr[41111] = 2146556380;
assign addr[41112] = 2145909429;
assign addr[41113] = 2145092320;
assign addr[41114] = 2144105118;
assign addr[41115] = 2142947902;
assign addr[41116] = 2141620763;
assign addr[41117] = 2140123807;
assign addr[41118] = 2138457152;
assign addr[41119] = 2136620930;
assign addr[41120] = 2134615288;
assign addr[41121] = 2132440383;
assign addr[41122] = 2130096389;
assign addr[41123] = 2127583492;
assign addr[41124] = 2124901890;
assign addr[41125] = 2122051796;
assign addr[41126] = 2119033436;
assign addr[41127] = 2115847050;
assign addr[41128] = 2112492891;
assign addr[41129] = 2108971223;
assign addr[41130] = 2105282327;
assign addr[41131] = 2101426496;
assign addr[41132] = 2097404033;
assign addr[41133] = 2093215260;
assign addr[41134] = 2088860507;
assign addr[41135] = 2084340120;
assign addr[41136] = 2079654458;
assign addr[41137] = 2074803892;
assign addr[41138] = 2069788807;
assign addr[41139] = 2064609600;
assign addr[41140] = 2059266683;
assign addr[41141] = 2053760478;
assign addr[41142] = 2048091422;
assign addr[41143] = 2042259965;
assign addr[41144] = 2036266570;
assign addr[41145] = 2030111710;
assign addr[41146] = 2023795876;
assign addr[41147] = 2017319567;
assign addr[41148] = 2010683297;
assign addr[41149] = 2003887591;
assign addr[41150] = 1996932990;
assign addr[41151] = 1989820044;
assign addr[41152] = 1982549318;
assign addr[41153] = 1975121388;
assign addr[41154] = 1967536842;
assign addr[41155] = 1959796283;
assign addr[41156] = 1951900324;
assign addr[41157] = 1943849591;
assign addr[41158] = 1935644723;
assign addr[41159] = 1927286370;
assign addr[41160] = 1918775195;
assign addr[41161] = 1910111873;
assign addr[41162] = 1901297091;
assign addr[41163] = 1892331547;
assign addr[41164] = 1883215953;
assign addr[41165] = 1873951032;
assign addr[41166] = 1864537518;
assign addr[41167] = 1854976157;
assign addr[41168] = 1845267708;
assign addr[41169] = 1835412941;
assign addr[41170] = 1825412636;
assign addr[41171] = 1815267588;
assign addr[41172] = 1804978599;
assign addr[41173] = 1794546487;
assign addr[41174] = 1783972079;
assign addr[41175] = 1773256212;
assign addr[41176] = 1762399737;
assign addr[41177] = 1751403515;
assign addr[41178] = 1740268417;
assign addr[41179] = 1728995326;
assign addr[41180] = 1717585136;
assign addr[41181] = 1706038753;
assign addr[41182] = 1694357091;
assign addr[41183] = 1682541077;
assign addr[41184] = 1670591647;
assign addr[41185] = 1658509750;
assign addr[41186] = 1646296344;
assign addr[41187] = 1633952396;
assign addr[41188] = 1621478885;
assign addr[41189] = 1608876801;
assign addr[41190] = 1596147143;
assign addr[41191] = 1583290921;
assign addr[41192] = 1570309153;
assign addr[41193] = 1557202869;
assign addr[41194] = 1543973108;
assign addr[41195] = 1530620920;
assign addr[41196] = 1517147363;
assign addr[41197] = 1503553506;
assign addr[41198] = 1489840425;
assign addr[41199] = 1476009210;
assign addr[41200] = 1462060956;
assign addr[41201] = 1447996770;
assign addr[41202] = 1433817766;
assign addr[41203] = 1419525069;
assign addr[41204] = 1405119813;
assign addr[41205] = 1390603139;
assign addr[41206] = 1375976199;
assign addr[41207] = 1361240152;
assign addr[41208] = 1346396168;
assign addr[41209] = 1331445422;
assign addr[41210] = 1316389101;
assign addr[41211] = 1301228398;
assign addr[41212] = 1285964516;
assign addr[41213] = 1270598665;
assign addr[41214] = 1255132063;
assign addr[41215] = 1239565936;
assign addr[41216] = 1223901520;
assign addr[41217] = 1208140056;
assign addr[41218] = 1192282793;
assign addr[41219] = 1176330990;
assign addr[41220] = 1160285911;
assign addr[41221] = 1144148829;
assign addr[41222] = 1127921022;
assign addr[41223] = 1111603778;
assign addr[41224] = 1095198391;
assign addr[41225] = 1078706161;
assign addr[41226] = 1062128397;
assign addr[41227] = 1045466412;
assign addr[41228] = 1028721528;
assign addr[41229] = 1011895073;
assign addr[41230] = 994988380;
assign addr[41231] = 978002791;
assign addr[41232] = 960939653;
assign addr[41233] = 943800318;
assign addr[41234] = 926586145;
assign addr[41235] = 909298500;
assign addr[41236] = 891938752;
assign addr[41237] = 874508280;
assign addr[41238] = 857008464;
assign addr[41239] = 839440693;
assign addr[41240] = 821806359;
assign addr[41241] = 804106861;
assign addr[41242] = 786343603;
assign addr[41243] = 768517992;
assign addr[41244] = 750631442;
assign addr[41245] = 732685372;
assign addr[41246] = 714681204;
assign addr[41247] = 696620367;
assign addr[41248] = 678504291;
assign addr[41249] = 660334415;
assign addr[41250] = 642112178;
assign addr[41251] = 623839025;
assign addr[41252] = 605516406;
assign addr[41253] = 587145773;
assign addr[41254] = 568728583;
assign addr[41255] = 550266296;
assign addr[41256] = 531760377;
assign addr[41257] = 513212292;
assign addr[41258] = 494623513;
assign addr[41259] = 475995513;
assign addr[41260] = 457329769;
assign addr[41261] = 438627762;
assign addr[41262] = 419890975;
assign addr[41263] = 401120892;
assign addr[41264] = 382319004;
assign addr[41265] = 363486799;
assign addr[41266] = 344625773;
assign addr[41267] = 325737419;
assign addr[41268] = 306823237;
assign addr[41269] = 287884725;
assign addr[41270] = 268923386;
assign addr[41271] = 249940723;
assign addr[41272] = 230938242;
assign addr[41273] = 211917448;
assign addr[41274] = 192879850;
assign addr[41275] = 173826959;
assign addr[41276] = 154760284;
assign addr[41277] = 135681337;
assign addr[41278] = 116591632;
assign addr[41279] = 97492681;
assign addr[41280] = 78386000;
assign addr[41281] = 59273104;
assign addr[41282] = 40155507;
assign addr[41283] = 21034727;
assign addr[41284] = 1912278;
assign addr[41285] = -17210322;
assign addr[41286] = -36331557;
assign addr[41287] = -55449912;
assign addr[41288] = -74563870;
assign addr[41289] = -93671915;
assign addr[41290] = -112772533;
assign addr[41291] = -131864208;
assign addr[41292] = -150945428;
assign addr[41293] = -170014678;
assign addr[41294] = -189070447;
assign addr[41295] = -208111224;
assign addr[41296] = -227135500;
assign addr[41297] = -246141764;
assign addr[41298] = -265128512;
assign addr[41299] = -284094236;
assign addr[41300] = -303037433;
assign addr[41301] = -321956601;
assign addr[41302] = -340850240;
assign addr[41303] = -359716852;
assign addr[41304] = -378554940;
assign addr[41305] = -397363011;
assign addr[41306] = -416139574;
assign addr[41307] = -434883140;
assign addr[41308] = -453592221;
assign addr[41309] = -472265336;
assign addr[41310] = -490901003;
assign addr[41311] = -509497745;
assign addr[41312] = -528054086;
assign addr[41313] = -546568556;
assign addr[41314] = -565039687;
assign addr[41315] = -583466013;
assign addr[41316] = -601846074;
assign addr[41317] = -620178412;
assign addr[41318] = -638461574;
assign addr[41319] = -656694110;
assign addr[41320] = -674874574;
assign addr[41321] = -693001525;
assign addr[41322] = -711073524;
assign addr[41323] = -729089140;
assign addr[41324] = -747046944;
assign addr[41325] = -764945512;
assign addr[41326] = -782783424;
assign addr[41327] = -800559266;
assign addr[41328] = -818271628;
assign addr[41329] = -835919107;
assign addr[41330] = -853500302;
assign addr[41331] = -871013820;
assign addr[41332] = -888458272;
assign addr[41333] = -905832274;
assign addr[41334] = -923134450;
assign addr[41335] = -940363427;
assign addr[41336] = -957517838;
assign addr[41337] = -974596324;
assign addr[41338] = -991597531;
assign addr[41339] = -1008520110;
assign addr[41340] = -1025362720;
assign addr[41341] = -1042124025;
assign addr[41342] = -1058802695;
assign addr[41343] = -1075397409;
assign addr[41344] = -1091906851;
assign addr[41345] = -1108329711;
assign addr[41346] = -1124664687;
assign addr[41347] = -1140910484;
assign addr[41348] = -1157065814;
assign addr[41349] = -1173129396;
assign addr[41350] = -1189099956;
assign addr[41351] = -1204976227;
assign addr[41352] = -1220756951;
assign addr[41353] = -1236440877;
assign addr[41354] = -1252026760;
assign addr[41355] = -1267513365;
assign addr[41356] = -1282899464;
assign addr[41357] = -1298183838;
assign addr[41358] = -1313365273;
assign addr[41359] = -1328442566;
assign addr[41360] = -1343414522;
assign addr[41361] = -1358279953;
assign addr[41362] = -1373037681;
assign addr[41363] = -1387686535;
assign addr[41364] = -1402225355;
assign addr[41365] = -1416652986;
assign addr[41366] = -1430968286;
assign addr[41367] = -1445170118;
assign addr[41368] = -1459257358;
assign addr[41369] = -1473228887;
assign addr[41370] = -1487083598;
assign addr[41371] = -1500820393;
assign addr[41372] = -1514438181;
assign addr[41373] = -1527935884;
assign addr[41374] = -1541312431;
assign addr[41375] = -1554566762;
assign addr[41376] = -1567697824;
assign addr[41377] = -1580704578;
assign addr[41378] = -1593585992;
assign addr[41379] = -1606341043;
assign addr[41380] = -1618968722;
assign addr[41381] = -1631468027;
assign addr[41382] = -1643837966;
assign addr[41383] = -1656077559;
assign addr[41384] = -1668185835;
assign addr[41385] = -1680161834;
assign addr[41386] = -1692004606;
assign addr[41387] = -1703713213;
assign addr[41388] = -1715286726;
assign addr[41389] = -1726724227;
assign addr[41390] = -1738024810;
assign addr[41391] = -1749187577;
assign addr[41392] = -1760211645;
assign addr[41393] = -1771096139;
assign addr[41394] = -1781840195;
assign addr[41395] = -1792442963;
assign addr[41396] = -1802903601;
assign addr[41397] = -1813221279;
assign addr[41398] = -1823395180;
assign addr[41399] = -1833424497;
assign addr[41400] = -1843308435;
assign addr[41401] = -1853046210;
assign addr[41402] = -1862637049;
assign addr[41403] = -1872080193;
assign addr[41404] = -1881374892;
assign addr[41405] = -1890520410;
assign addr[41406] = -1899516021;
assign addr[41407] = -1908361011;
assign addr[41408] = -1917054681;
assign addr[41409] = -1925596340;
assign addr[41410] = -1933985310;
assign addr[41411] = -1942220928;
assign addr[41412] = -1950302539;
assign addr[41413] = -1958229503;
assign addr[41414] = -1966001192;
assign addr[41415] = -1973616989;
assign addr[41416] = -1981076290;
assign addr[41417] = -1988378503;
assign addr[41418] = -1995523051;
assign addr[41419] = -2002509365;
assign addr[41420] = -2009336893;
assign addr[41421] = -2016005093;
assign addr[41422] = -2022513436;
assign addr[41423] = -2028861406;
assign addr[41424] = -2035048499;
assign addr[41425] = -2041074226;
assign addr[41426] = -2046938108;
assign addr[41427] = -2052639680;
assign addr[41428] = -2058178491;
assign addr[41429] = -2063554100;
assign addr[41430] = -2068766083;
assign addr[41431] = -2073814024;
assign addr[41432] = -2078697525;
assign addr[41433] = -2083416198;
assign addr[41434] = -2087969669;
assign addr[41435] = -2092357577;
assign addr[41436] = -2096579573;
assign addr[41437] = -2100635323;
assign addr[41438] = -2104524506;
assign addr[41439] = -2108246813;
assign addr[41440] = -2111801949;
assign addr[41441] = -2115189632;
assign addr[41442] = -2118409593;
assign addr[41443] = -2121461578;
assign addr[41444] = -2124345343;
assign addr[41445] = -2127060661;
assign addr[41446] = -2129607316;
assign addr[41447] = -2131985106;
assign addr[41448] = -2134193842;
assign addr[41449] = -2136233350;
assign addr[41450] = -2138103468;
assign addr[41451] = -2139804048;
assign addr[41452] = -2141334954;
assign addr[41453] = -2142696065;
assign addr[41454] = -2143887273;
assign addr[41455] = -2144908484;
assign addr[41456] = -2145759618;
assign addr[41457] = -2146440605;
assign addr[41458] = -2146951393;
assign addr[41459] = -2147291941;
assign addr[41460] = -2147462221;
assign addr[41461] = -2147462221;
assign addr[41462] = -2147291941;
assign addr[41463] = -2146951393;
assign addr[41464] = -2146440605;
assign addr[41465] = -2145759618;
assign addr[41466] = -2144908484;
assign addr[41467] = -2143887273;
assign addr[41468] = -2142696065;
assign addr[41469] = -2141334954;
assign addr[41470] = -2139804048;
assign addr[41471] = -2138103468;
assign addr[41472] = -2136233350;
assign addr[41473] = -2134193842;
assign addr[41474] = -2131985106;
assign addr[41475] = -2129607316;
assign addr[41476] = -2127060661;
assign addr[41477] = -2124345343;
assign addr[41478] = -2121461578;
assign addr[41479] = -2118409593;
assign addr[41480] = -2115189632;
assign addr[41481] = -2111801949;
assign addr[41482] = -2108246813;
assign addr[41483] = -2104524506;
assign addr[41484] = -2100635323;
assign addr[41485] = -2096579573;
assign addr[41486] = -2092357577;
assign addr[41487] = -2087969669;
assign addr[41488] = -2083416198;
assign addr[41489] = -2078697525;
assign addr[41490] = -2073814024;
assign addr[41491] = -2068766083;
assign addr[41492] = -2063554100;
assign addr[41493] = -2058178491;
assign addr[41494] = -2052639680;
assign addr[41495] = -2046938108;
assign addr[41496] = -2041074226;
assign addr[41497] = -2035048499;
assign addr[41498] = -2028861406;
assign addr[41499] = -2022513436;
assign addr[41500] = -2016005093;
assign addr[41501] = -2009336893;
assign addr[41502] = -2002509365;
assign addr[41503] = -1995523051;
assign addr[41504] = -1988378503;
assign addr[41505] = -1981076290;
assign addr[41506] = -1973616989;
assign addr[41507] = -1966001192;
assign addr[41508] = -1958229503;
assign addr[41509] = -1950302539;
assign addr[41510] = -1942220928;
assign addr[41511] = -1933985310;
assign addr[41512] = -1925596340;
assign addr[41513] = -1917054681;
assign addr[41514] = -1908361011;
assign addr[41515] = -1899516021;
assign addr[41516] = -1890520410;
assign addr[41517] = -1881374892;
assign addr[41518] = -1872080193;
assign addr[41519] = -1862637049;
assign addr[41520] = -1853046210;
assign addr[41521] = -1843308435;
assign addr[41522] = -1833424497;
assign addr[41523] = -1823395180;
assign addr[41524] = -1813221279;
assign addr[41525] = -1802903601;
assign addr[41526] = -1792442963;
assign addr[41527] = -1781840195;
assign addr[41528] = -1771096139;
assign addr[41529] = -1760211645;
assign addr[41530] = -1749187577;
assign addr[41531] = -1738024810;
assign addr[41532] = -1726724227;
assign addr[41533] = -1715286726;
assign addr[41534] = -1703713213;
assign addr[41535] = -1692004606;
assign addr[41536] = -1680161834;
assign addr[41537] = -1668185835;
assign addr[41538] = -1656077559;
assign addr[41539] = -1643837966;
assign addr[41540] = -1631468027;
assign addr[41541] = -1618968722;
assign addr[41542] = -1606341043;
assign addr[41543] = -1593585992;
assign addr[41544] = -1580704578;
assign addr[41545] = -1567697824;
assign addr[41546] = -1554566762;
assign addr[41547] = -1541312431;
assign addr[41548] = -1527935884;
assign addr[41549] = -1514438181;
assign addr[41550] = -1500820393;
assign addr[41551] = -1487083598;
assign addr[41552] = -1473228887;
assign addr[41553] = -1459257358;
assign addr[41554] = -1445170118;
assign addr[41555] = -1430968286;
assign addr[41556] = -1416652986;
assign addr[41557] = -1402225355;
assign addr[41558] = -1387686535;
assign addr[41559] = -1373037681;
assign addr[41560] = -1358279953;
assign addr[41561] = -1343414522;
assign addr[41562] = -1328442566;
assign addr[41563] = -1313365273;
assign addr[41564] = -1298183838;
assign addr[41565] = -1282899464;
assign addr[41566] = -1267513365;
assign addr[41567] = -1252026760;
assign addr[41568] = -1236440877;
assign addr[41569] = -1220756951;
assign addr[41570] = -1204976227;
assign addr[41571] = -1189099956;
assign addr[41572] = -1173129396;
assign addr[41573] = -1157065814;
assign addr[41574] = -1140910484;
assign addr[41575] = -1124664687;
assign addr[41576] = -1108329711;
assign addr[41577] = -1091906851;
assign addr[41578] = -1075397409;
assign addr[41579] = -1058802695;
assign addr[41580] = -1042124025;
assign addr[41581] = -1025362720;
assign addr[41582] = -1008520110;
assign addr[41583] = -991597531;
assign addr[41584] = -974596324;
assign addr[41585] = -957517838;
assign addr[41586] = -940363427;
assign addr[41587] = -923134450;
assign addr[41588] = -905832274;
assign addr[41589] = -888458272;
assign addr[41590] = -871013820;
assign addr[41591] = -853500302;
assign addr[41592] = -835919107;
assign addr[41593] = -818271628;
assign addr[41594] = -800559266;
assign addr[41595] = -782783424;
assign addr[41596] = -764945512;
assign addr[41597] = -747046944;
assign addr[41598] = -729089140;
assign addr[41599] = -711073524;
assign addr[41600] = -693001525;
assign addr[41601] = -674874574;
assign addr[41602] = -656694110;
assign addr[41603] = -638461574;
assign addr[41604] = -620178412;
assign addr[41605] = -601846074;
assign addr[41606] = -583466013;
assign addr[41607] = -565039687;
assign addr[41608] = -546568556;
assign addr[41609] = -528054086;
assign addr[41610] = -509497745;
assign addr[41611] = -490901003;
assign addr[41612] = -472265336;
assign addr[41613] = -453592221;
assign addr[41614] = -434883140;
assign addr[41615] = -416139574;
assign addr[41616] = -397363011;
assign addr[41617] = -378554940;
assign addr[41618] = -359716852;
assign addr[41619] = -340850240;
assign addr[41620] = -321956601;
assign addr[41621] = -303037433;
assign addr[41622] = -284094236;
assign addr[41623] = -265128512;
assign addr[41624] = -246141764;
assign addr[41625] = -227135500;
assign addr[41626] = -208111224;
assign addr[41627] = -189070447;
assign addr[41628] = -170014678;
assign addr[41629] = -150945428;
assign addr[41630] = -131864208;
assign addr[41631] = -112772533;
assign addr[41632] = -93671915;
assign addr[41633] = -74563870;
assign addr[41634] = -55449912;
assign addr[41635] = -36331557;
assign addr[41636] = -17210322;
assign addr[41637] = 1912278;
assign addr[41638] = 21034727;
assign addr[41639] = 40155507;
assign addr[41640] = 59273104;
assign addr[41641] = 78386000;
assign addr[41642] = 97492681;
assign addr[41643] = 116591632;
assign addr[41644] = 135681337;
assign addr[41645] = 154760284;
assign addr[41646] = 173826959;
assign addr[41647] = 192879850;
assign addr[41648] = 211917448;
assign addr[41649] = 230938242;
assign addr[41650] = 249940723;
assign addr[41651] = 268923386;
assign addr[41652] = 287884725;
assign addr[41653] = 306823237;
assign addr[41654] = 325737419;
assign addr[41655] = 344625773;
assign addr[41656] = 363486799;
assign addr[41657] = 382319004;
assign addr[41658] = 401120892;
assign addr[41659] = 419890975;
assign addr[41660] = 438627762;
assign addr[41661] = 457329769;
assign addr[41662] = 475995513;
assign addr[41663] = 494623513;
assign addr[41664] = 513212292;
assign addr[41665] = 531760377;
assign addr[41666] = 550266296;
assign addr[41667] = 568728583;
assign addr[41668] = 587145773;
assign addr[41669] = 605516406;
assign addr[41670] = 623839025;
assign addr[41671] = 642112178;
assign addr[41672] = 660334415;
assign addr[41673] = 678504291;
assign addr[41674] = 696620367;
assign addr[41675] = 714681204;
assign addr[41676] = 732685372;
assign addr[41677] = 750631442;
assign addr[41678] = 768517992;
assign addr[41679] = 786343603;
assign addr[41680] = 804106861;
assign addr[41681] = 821806359;
assign addr[41682] = 839440693;
assign addr[41683] = 857008464;
assign addr[41684] = 874508280;
assign addr[41685] = 891938752;
assign addr[41686] = 909298500;
assign addr[41687] = 926586145;
assign addr[41688] = 943800318;
assign addr[41689] = 960939653;
assign addr[41690] = 978002791;
assign addr[41691] = 994988380;
assign addr[41692] = 1011895073;
assign addr[41693] = 1028721528;
assign addr[41694] = 1045466412;
assign addr[41695] = 1062128397;
assign addr[41696] = 1078706161;
assign addr[41697] = 1095198391;
assign addr[41698] = 1111603778;
assign addr[41699] = 1127921022;
assign addr[41700] = 1144148829;
assign addr[41701] = 1160285911;
assign addr[41702] = 1176330990;
assign addr[41703] = 1192282793;
assign addr[41704] = 1208140056;
assign addr[41705] = 1223901520;
assign addr[41706] = 1239565936;
assign addr[41707] = 1255132063;
assign addr[41708] = 1270598665;
assign addr[41709] = 1285964516;
assign addr[41710] = 1301228398;
assign addr[41711] = 1316389101;
assign addr[41712] = 1331445422;
assign addr[41713] = 1346396168;
assign addr[41714] = 1361240152;
assign addr[41715] = 1375976199;
assign addr[41716] = 1390603139;
assign addr[41717] = 1405119813;
assign addr[41718] = 1419525069;
assign addr[41719] = 1433817766;
assign addr[41720] = 1447996770;
assign addr[41721] = 1462060956;
assign addr[41722] = 1476009210;
assign addr[41723] = 1489840425;
assign addr[41724] = 1503553506;
assign addr[41725] = 1517147363;
assign addr[41726] = 1530620920;
assign addr[41727] = 1543973108;
assign addr[41728] = 1557202869;
assign addr[41729] = 1570309153;
assign addr[41730] = 1583290921;
assign addr[41731] = 1596147143;
assign addr[41732] = 1608876801;
assign addr[41733] = 1621478885;
assign addr[41734] = 1633952396;
assign addr[41735] = 1646296344;
assign addr[41736] = 1658509750;
assign addr[41737] = 1670591647;
assign addr[41738] = 1682541077;
assign addr[41739] = 1694357091;
assign addr[41740] = 1706038753;
assign addr[41741] = 1717585136;
assign addr[41742] = 1728995326;
assign addr[41743] = 1740268417;
assign addr[41744] = 1751403515;
assign addr[41745] = 1762399737;
assign addr[41746] = 1773256212;
assign addr[41747] = 1783972079;
assign addr[41748] = 1794546487;
assign addr[41749] = 1804978599;
assign addr[41750] = 1815267588;
assign addr[41751] = 1825412636;
assign addr[41752] = 1835412941;
assign addr[41753] = 1845267708;
assign addr[41754] = 1854976157;
assign addr[41755] = 1864537518;
assign addr[41756] = 1873951032;
assign addr[41757] = 1883215953;
assign addr[41758] = 1892331547;
assign addr[41759] = 1901297091;
assign addr[41760] = 1910111873;
assign addr[41761] = 1918775195;
assign addr[41762] = 1927286370;
assign addr[41763] = 1935644723;
assign addr[41764] = 1943849591;
assign addr[41765] = 1951900324;
assign addr[41766] = 1959796283;
assign addr[41767] = 1967536842;
assign addr[41768] = 1975121388;
assign addr[41769] = 1982549318;
assign addr[41770] = 1989820044;
assign addr[41771] = 1996932990;
assign addr[41772] = 2003887591;
assign addr[41773] = 2010683297;
assign addr[41774] = 2017319567;
assign addr[41775] = 2023795876;
assign addr[41776] = 2030111710;
assign addr[41777] = 2036266570;
assign addr[41778] = 2042259965;
assign addr[41779] = 2048091422;
assign addr[41780] = 2053760478;
assign addr[41781] = 2059266683;
assign addr[41782] = 2064609600;
assign addr[41783] = 2069788807;
assign addr[41784] = 2074803892;
assign addr[41785] = 2079654458;
assign addr[41786] = 2084340120;
assign addr[41787] = 2088860507;
assign addr[41788] = 2093215260;
assign addr[41789] = 2097404033;
assign addr[41790] = 2101426496;
assign addr[41791] = 2105282327;
assign addr[41792] = 2108971223;
assign addr[41793] = 2112492891;
assign addr[41794] = 2115847050;
assign addr[41795] = 2119033436;
assign addr[41796] = 2122051796;
assign addr[41797] = 2124901890;
assign addr[41798] = 2127583492;
assign addr[41799] = 2130096389;
assign addr[41800] = 2132440383;
assign addr[41801] = 2134615288;
assign addr[41802] = 2136620930;
assign addr[41803] = 2138457152;
assign addr[41804] = 2140123807;
assign addr[41805] = 2141620763;
assign addr[41806] = 2142947902;
assign addr[41807] = 2144105118;
assign addr[41808] = 2145092320;
assign addr[41809] = 2145909429;
assign addr[41810] = 2146556380;
assign addr[41811] = 2147033123;
assign addr[41812] = 2147339619;
assign addr[41813] = 2147475844;
assign addr[41814] = 2147441787;
assign addr[41815] = 2147237452;
assign addr[41816] = 2146862854;
assign addr[41817] = 2146318022;
assign addr[41818] = 2145603001;
assign addr[41819] = 2144717846;
assign addr[41820] = 2143662628;
assign addr[41821] = 2142437431;
assign addr[41822] = 2141042352;
assign addr[41823] = 2139477502;
assign addr[41824] = 2137743003;
assign addr[41825] = 2135838995;
assign addr[41826] = 2133765628;
assign addr[41827] = 2131523066;
assign addr[41828] = 2129111488;
assign addr[41829] = 2126531084;
assign addr[41830] = 2123782059;
assign addr[41831] = 2120864631;
assign addr[41832] = 2117779031;
assign addr[41833] = 2114525505;
assign addr[41834] = 2111104309;
assign addr[41835] = 2107515716;
assign addr[41836] = 2103760010;
assign addr[41837] = 2099837489;
assign addr[41838] = 2095748463;
assign addr[41839] = 2091493257;
assign addr[41840] = 2087072209;
assign addr[41841] = 2082485668;
assign addr[41842] = 2077733999;
assign addr[41843] = 2072817579;
assign addr[41844] = 2067736796;
assign addr[41845] = 2062492055;
assign addr[41846] = 2057083771;
assign addr[41847] = 2051512372;
assign addr[41848] = 2045778302;
assign addr[41849] = 2039882013;
assign addr[41850] = 2033823974;
assign addr[41851] = 2027604666;
assign addr[41852] = 2021224581;
assign addr[41853] = 2014684225;
assign addr[41854] = 2007984117;
assign addr[41855] = 2001124788;
assign addr[41856] = 1994106782;
assign addr[41857] = 1986930656;
assign addr[41858] = 1979596978;
assign addr[41859] = 1972106330;
assign addr[41860] = 1964459306;
assign addr[41861] = 1956656513;
assign addr[41862] = 1948698568;
assign addr[41863] = 1940586104;
assign addr[41864] = 1932319763;
assign addr[41865] = 1923900201;
assign addr[41866] = 1915328086;
assign addr[41867] = 1906604097;
assign addr[41868] = 1897728925;
assign addr[41869] = 1888703276;
assign addr[41870] = 1879527863;
assign addr[41871] = 1870203416;
assign addr[41872] = 1860730673;
assign addr[41873] = 1851110385;
assign addr[41874] = 1841343316;
assign addr[41875] = 1831430239;
assign addr[41876] = 1821371941;
assign addr[41877] = 1811169220;
assign addr[41878] = 1800822883;
assign addr[41879] = 1790333753;
assign addr[41880] = 1779702660;
assign addr[41881] = 1768930447;
assign addr[41882] = 1758017969;
assign addr[41883] = 1746966091;
assign addr[41884] = 1735775690;
assign addr[41885] = 1724447652;
assign addr[41886] = 1712982875;
assign addr[41887] = 1701382270;
assign addr[41888] = 1689646755;
assign addr[41889] = 1677777262;
assign addr[41890] = 1665774731;
assign addr[41891] = 1653640115;
assign addr[41892] = 1641374375;
assign addr[41893] = 1628978484;
assign addr[41894] = 1616453425;
assign addr[41895] = 1603800191;
assign addr[41896] = 1591019785;
assign addr[41897] = 1578113222;
assign addr[41898] = 1565081523;
assign addr[41899] = 1551925723;
assign addr[41900] = 1538646865;
assign addr[41901] = 1525246002;
assign addr[41902] = 1511724196;
assign addr[41903] = 1498082520;
assign addr[41904] = 1484322054;
assign addr[41905] = 1470443891;
assign addr[41906] = 1456449131;
assign addr[41907] = 1442338884;
assign addr[41908] = 1428114267;
assign addr[41909] = 1413776410;
assign addr[41910] = 1399326449;
assign addr[41911] = 1384765530;
assign addr[41912] = 1370094808;
assign addr[41913] = 1355315445;
assign addr[41914] = 1340428615;
assign addr[41915] = 1325435496;
assign addr[41916] = 1310337279;
assign addr[41917] = 1295135159;
assign addr[41918] = 1279830344;
assign addr[41919] = 1264424045;
assign addr[41920] = 1248917486;
assign addr[41921] = 1233311895;
assign addr[41922] = 1217608510;
assign addr[41923] = 1201808576;
assign addr[41924] = 1185913346;
assign addr[41925] = 1169924081;
assign addr[41926] = 1153842047;
assign addr[41927] = 1137668521;
assign addr[41928] = 1121404785;
assign addr[41929] = 1105052128;
assign addr[41930] = 1088611847;
assign addr[41931] = 1072085246;
assign addr[41932] = 1055473635;
assign addr[41933] = 1038778332;
assign addr[41934] = 1022000660;
assign addr[41935] = 1005141949;
assign addr[41936] = 988203537;
assign addr[41937] = 971186766;
assign addr[41938] = 954092986;
assign addr[41939] = 936923553;
assign addr[41940] = 919679827;
assign addr[41941] = 902363176;
assign addr[41942] = 884974973;
assign addr[41943] = 867516597;
assign addr[41944] = 849989433;
assign addr[41945] = 832394869;
assign addr[41946] = 814734301;
assign addr[41947] = 797009130;
assign addr[41948] = 779220762;
assign addr[41949] = 761370605;
assign addr[41950] = 743460077;
assign addr[41951] = 725490597;
assign addr[41952] = 707463589;
assign addr[41953] = 689380485;
assign addr[41954] = 671242716;
assign addr[41955] = 653051723;
assign addr[41956] = 634808946;
assign addr[41957] = 616515832;
assign addr[41958] = 598173833;
assign addr[41959] = 579784402;
assign addr[41960] = 561348998;
assign addr[41961] = 542869083;
assign addr[41962] = 524346121;
assign addr[41963] = 505781581;
assign addr[41964] = 487176937;
assign addr[41965] = 468533662;
assign addr[41966] = 449853235;
assign addr[41967] = 431137138;
assign addr[41968] = 412386854;
assign addr[41969] = 393603870;
assign addr[41970] = 374789676;
assign addr[41971] = 355945764;
assign addr[41972] = 337073627;
assign addr[41973] = 318174762;
assign addr[41974] = 299250668;
assign addr[41975] = 280302845;
assign addr[41976] = 261332796;
assign addr[41977] = 242342025;
assign addr[41978] = 223332037;
assign addr[41979] = 204304341;
assign addr[41980] = 185260444;
assign addr[41981] = 166201858;
assign addr[41982] = 147130093;
assign addr[41983] = 128046661;
assign addr[41984] = 108953076;
assign addr[41985] = 89850852;
assign addr[41986] = 70741503;
assign addr[41987] = 51626544;
assign addr[41988] = 32507492;
assign addr[41989] = 13385863;
assign addr[41990] = -5736829;
assign addr[41991] = -24859065;
assign addr[41992] = -43979330;
assign addr[41993] = -63096108;
assign addr[41994] = -82207882;
assign addr[41995] = -101313138;
assign addr[41996] = -120410361;
assign addr[41997] = -139498035;
assign addr[41998] = -158574649;
assign addr[41999] = -177638688;
assign addr[42000] = -196688642;
assign addr[42001] = -215722999;
assign addr[42002] = -234740251;
assign addr[42003] = -253738890;
assign addr[42004] = -272717408;
assign addr[42005] = -291674302;
assign addr[42006] = -310608068;
assign addr[42007] = -329517204;
assign addr[42008] = -348400212;
assign addr[42009] = -367255594;
assign addr[42010] = -386081854;
assign addr[42011] = -404877501;
assign addr[42012] = -423641043;
assign addr[42013] = -442370993;
assign addr[42014] = -461065866;
assign addr[42015] = -479724180;
assign addr[42016] = -498344454;
assign addr[42017] = -516925212;
assign addr[42018] = -535464981;
assign addr[42019] = -553962291;
assign addr[42020] = -572415676;
assign addr[42021] = -590823671;
assign addr[42022] = -609184818;
assign addr[42023] = -627497660;
assign addr[42024] = -645760745;
assign addr[42025] = -663972625;
assign addr[42026] = -682131857;
assign addr[42027] = -700236999;
assign addr[42028] = -718286617;
assign addr[42029] = -736279279;
assign addr[42030] = -754213559;
assign addr[42031] = -772088034;
assign addr[42032] = -789901288;
assign addr[42033] = -807651907;
assign addr[42034] = -825338484;
assign addr[42035] = -842959617;
assign addr[42036] = -860513908;
assign addr[42037] = -877999966;
assign addr[42038] = -895416404;
assign addr[42039] = -912761841;
assign addr[42040] = -930034901;
assign addr[42041] = -947234215;
assign addr[42042] = -964358420;
assign addr[42043] = -981406156;
assign addr[42044] = -998376073;
assign addr[42045] = -1015266825;
assign addr[42046] = -1032077073;
assign addr[42047] = -1048805483;
assign addr[42048] = -1065450729;
assign addr[42049] = -1082011492;
assign addr[42050] = -1098486458;
assign addr[42051] = -1114874320;
assign addr[42052] = -1131173780;
assign addr[42053] = -1147383544;
assign addr[42054] = -1163502328;
assign addr[42055] = -1179528853;
assign addr[42056] = -1195461849;
assign addr[42057] = -1211300053;
assign addr[42058] = -1227042207;
assign addr[42059] = -1242687064;
assign addr[42060] = -1258233384;
assign addr[42061] = -1273679934;
assign addr[42062] = -1289025489;
assign addr[42063] = -1304268832;
assign addr[42064] = -1319408754;
assign addr[42065] = -1334444055;
assign addr[42066] = -1349373543;
assign addr[42067] = -1364196034;
assign addr[42068] = -1378910353;
assign addr[42069] = -1393515332;
assign addr[42070] = -1408009814;
assign addr[42071] = -1422392650;
assign addr[42072] = -1436662698;
assign addr[42073] = -1450818828;
assign addr[42074] = -1464859917;
assign addr[42075] = -1478784851;
assign addr[42076] = -1492592527;
assign addr[42077] = -1506281850;
assign addr[42078] = -1519851733;
assign addr[42079] = -1533301101;
assign addr[42080] = -1546628888;
assign addr[42081] = -1559834037;
assign addr[42082] = -1572915501;
assign addr[42083] = -1585872242;
assign addr[42084] = -1598703233;
assign addr[42085] = -1611407456;
assign addr[42086] = -1623983905;
assign addr[42087] = -1636431582;
assign addr[42088] = -1648749499;
assign addr[42089] = -1660936681;
assign addr[42090] = -1672992161;
assign addr[42091] = -1684914983;
assign addr[42092] = -1696704201;
assign addr[42093] = -1708358881;
assign addr[42094] = -1719878099;
assign addr[42095] = -1731260941;
assign addr[42096] = -1742506504;
assign addr[42097] = -1753613897;
assign addr[42098] = -1764582240;
assign addr[42099] = -1775410662;
assign addr[42100] = -1786098304;
assign addr[42101] = -1796644320;
assign addr[42102] = -1807047873;
assign addr[42103] = -1817308138;
assign addr[42104] = -1827424302;
assign addr[42105] = -1837395562;
assign addr[42106] = -1847221128;
assign addr[42107] = -1856900221;
assign addr[42108] = -1866432072;
assign addr[42109] = -1875815927;
assign addr[42110] = -1885051042;
assign addr[42111] = -1894136683;
assign addr[42112] = -1903072131;
assign addr[42113] = -1911856677;
assign addr[42114] = -1920489624;
assign addr[42115] = -1928970288;
assign addr[42116] = -1937297997;
assign addr[42117] = -1945472089;
assign addr[42118] = -1953491918;
assign addr[42119] = -1961356847;
assign addr[42120] = -1969066252;
assign addr[42121] = -1976619522;
assign addr[42122] = -1984016058;
assign addr[42123] = -1991255274;
assign addr[42124] = -1998336596;
assign addr[42125] = -2005259462;
assign addr[42126] = -2012023322;
assign addr[42127] = -2018627642;
assign addr[42128] = -2025071897;
assign addr[42129] = -2031355576;
assign addr[42130] = -2037478181;
assign addr[42131] = -2043439226;
assign addr[42132] = -2049238240;
assign addr[42133] = -2054874761;
assign addr[42134] = -2060348343;
assign addr[42135] = -2065658552;
assign addr[42136] = -2070804967;
assign addr[42137] = -2075787180;
assign addr[42138] = -2080604795;
assign addr[42139] = -2085257431;
assign addr[42140] = -2089744719;
assign addr[42141] = -2094066304;
assign addr[42142] = -2098221841;
assign addr[42143] = -2102211002;
assign addr[42144] = -2106033471;
assign addr[42145] = -2109688944;
assign addr[42146] = -2113177132;
assign addr[42147] = -2116497758;
assign addr[42148] = -2119650558;
assign addr[42149] = -2122635283;
assign addr[42150] = -2125451696;
assign addr[42151] = -2128099574;
assign addr[42152] = -2130578706;
assign addr[42153] = -2132888897;
assign addr[42154] = -2135029962;
assign addr[42155] = -2137001733;
assign addr[42156] = -2138804053;
assign addr[42157] = -2140436778;
assign addr[42158] = -2141899780;
assign addr[42159] = -2143192942;
assign addr[42160] = -2144316162;
assign addr[42161] = -2145269351;
assign addr[42162] = -2146052433;
assign addr[42163] = -2146665347;
assign addr[42164] = -2147108043;
assign addr[42165] = -2147380486;
assign addr[42166] = -2147482655;
assign addr[42167] = -2147414542;
assign addr[42168] = -2147176152;
assign addr[42169] = -2146767505;
assign addr[42170] = -2146188631;
assign addr[42171] = -2145439578;
assign addr[42172] = -2144520405;
assign addr[42173] = -2143431184;
assign addr[42174] = -2142172003;
assign addr[42175] = -2140742960;
assign addr[42176] = -2139144169;
assign addr[42177] = -2137375758;
assign addr[42178] = -2135437865;
assign addr[42179] = -2133330646;
assign addr[42180] = -2131054266;
assign addr[42181] = -2128608907;
assign addr[42182] = -2125994762;
assign addr[42183] = -2123212038;
assign addr[42184] = -2120260957;
assign addr[42185] = -2117141752;
assign addr[42186] = -2113854671;
assign addr[42187] = -2110399974;
assign addr[42188] = -2106777935;
assign addr[42189] = -2102988841;
assign addr[42190] = -2099032994;
assign addr[42191] = -2094910706;
assign addr[42192] = -2090622304;
assign addr[42193] = -2086168128;
assign addr[42194] = -2081548533;
assign addr[42195] = -2076763883;
assign addr[42196] = -2071814558;
assign addr[42197] = -2066700952;
assign addr[42198] = -2061423468;
assign addr[42199] = -2055982526;
assign addr[42200] = -2050378558;
assign addr[42201] = -2044612007;
assign addr[42202] = -2038683330;
assign addr[42203] = -2032592999;
assign addr[42204] = -2026341495;
assign addr[42205] = -2019929315;
assign addr[42206] = -2013356967;
assign addr[42207] = -2006624971;
assign addr[42208] = -1999733863;
assign addr[42209] = -1992684188;
assign addr[42210] = -1985476506;
assign addr[42211] = -1978111387;
assign addr[42212] = -1970589416;
assign addr[42213] = -1962911189;
assign addr[42214] = -1955077316;
assign addr[42215] = -1947088417;
assign addr[42216] = -1938945125;
assign addr[42217] = -1930648088;
assign addr[42218] = -1922197961;
assign addr[42219] = -1913595416;
assign addr[42220] = -1904841135;
assign addr[42221] = -1895935811;
assign addr[42222] = -1886880151;
assign addr[42223] = -1877674873;
assign addr[42224] = -1868320707;
assign addr[42225] = -1858818395;
assign addr[42226] = -1849168689;
assign addr[42227] = -1839372356;
assign addr[42228] = -1829430172;
assign addr[42229] = -1819342925;
assign addr[42230] = -1809111415;
assign addr[42231] = -1798736454;
assign addr[42232] = -1788218865;
assign addr[42233] = -1777559480;
assign addr[42234] = -1766759146;
assign addr[42235] = -1755818718;
assign addr[42236] = -1744739065;
assign addr[42237] = -1733521064;
assign addr[42238] = -1722165606;
assign addr[42239] = -1710673591;
assign addr[42240] = -1699045930;
assign addr[42241] = -1687283545;
assign addr[42242] = -1675387369;
assign addr[42243] = -1663358344;
assign addr[42244] = -1651197426;
assign addr[42245] = -1638905577;
assign addr[42246] = -1626483774;
assign addr[42247] = -1613933000;
assign addr[42248] = -1601254251;
assign addr[42249] = -1588448533;
assign addr[42250] = -1575516860;
assign addr[42251] = -1562460258;
assign addr[42252] = -1549279763;
assign addr[42253] = -1535976419;
assign addr[42254] = -1522551282;
assign addr[42255] = -1509005416;
assign addr[42256] = -1495339895;
assign addr[42257] = -1481555802;
assign addr[42258] = -1467654232;
assign addr[42259] = -1453636285;
assign addr[42260] = -1439503074;
assign addr[42261] = -1425255719;
assign addr[42262] = -1410895350;
assign addr[42263] = -1396423105;
assign addr[42264] = -1381840133;
assign addr[42265] = -1367147589;
assign addr[42266] = -1352346639;
assign addr[42267] = -1337438456;
assign addr[42268] = -1322424222;
assign addr[42269] = -1307305128;
assign addr[42270] = -1292082373;
assign addr[42271] = -1276757164;
assign addr[42272] = -1261330715;
assign addr[42273] = -1245804251;
assign addr[42274] = -1230179002;
assign addr[42275] = -1214456207;
assign addr[42276] = -1198637114;
assign addr[42277] = -1182722976;
assign addr[42278] = -1166715055;
assign addr[42279] = -1150614620;
assign addr[42280] = -1134422949;
assign addr[42281] = -1118141326;
assign addr[42282] = -1101771040;
assign addr[42283] = -1085313391;
assign addr[42284] = -1068769683;
assign addr[42285] = -1052141228;
assign addr[42286] = -1035429345;
assign addr[42287] = -1018635358;
assign addr[42288] = -1001760600;
assign addr[42289] = -984806408;
assign addr[42290] = -967774128;
assign addr[42291] = -950665109;
assign addr[42292] = -933480707;
assign addr[42293] = -916222287;
assign addr[42294] = -898891215;
assign addr[42295] = -881488868;
assign addr[42296] = -864016623;
assign addr[42297] = -846475867;
assign addr[42298] = -828867991;
assign addr[42299] = -811194391;
assign addr[42300] = -793456467;
assign addr[42301] = -775655628;
assign addr[42302] = -757793284;
assign addr[42303] = -739870851;
assign addr[42304] = -721889752;
assign addr[42305] = -703851410;
assign addr[42306] = -685757258;
assign addr[42307] = -667608730;
assign addr[42308] = -649407264;
assign addr[42309] = -631154304;
assign addr[42310] = -612851297;
assign addr[42311] = -594499695;
assign addr[42312] = -576100953;
assign addr[42313] = -557656529;
assign addr[42314] = -539167887;
assign addr[42315] = -520636492;
assign addr[42316] = -502063814;
assign addr[42317] = -483451325;
assign addr[42318] = -464800501;
assign addr[42319] = -446112822;
assign addr[42320] = -427389768;
assign addr[42321] = -408632825;
assign addr[42322] = -389843480;
assign addr[42323] = -371023223;
assign addr[42324] = -352173546;
assign addr[42325] = -333295944;
assign addr[42326] = -314391913;
assign addr[42327] = -295462954;
assign addr[42328] = -276510565;
assign addr[42329] = -257536251;
assign addr[42330] = -238541516;
assign addr[42331] = -219527866;
assign addr[42332] = -200496809;
assign addr[42333] = -181449854;
assign addr[42334] = -162388511;
assign addr[42335] = -143314291;
assign addr[42336] = -124228708;
assign addr[42337] = -105133274;
assign addr[42338] = -86029503;
assign addr[42339] = -66918911;
assign addr[42340] = -47803013;
assign addr[42341] = -28683324;
assign addr[42342] = -9561361;
assign addr[42343] = 9561361;
assign addr[42344] = 28683324;
assign addr[42345] = 47803013;
assign addr[42346] = 66918911;
assign addr[42347] = 86029503;
assign addr[42348] = 105133274;
assign addr[42349] = 124228708;
assign addr[42350] = 143314291;
assign addr[42351] = 162388511;
assign addr[42352] = 181449854;
assign addr[42353] = 200496809;
assign addr[42354] = 219527866;
assign addr[42355] = 238541516;
assign addr[42356] = 257536251;
assign addr[42357] = 276510565;
assign addr[42358] = 295462953;
assign addr[42359] = 314391913;
assign addr[42360] = 333295944;
assign addr[42361] = 352173546;
assign addr[42362] = 371023223;
assign addr[42363] = 389843480;
assign addr[42364] = 408632825;
assign addr[42365] = 427389768;
assign addr[42366] = 446112822;
assign addr[42367] = 464800501;
assign addr[42368] = 483451325;
assign addr[42369] = 502063814;
assign addr[42370] = 520636492;
assign addr[42371] = 539167887;
assign addr[42372] = 557656529;
assign addr[42373] = 576100953;
assign addr[42374] = 594499695;
assign addr[42375] = 612851297;
assign addr[42376] = 631154304;
assign addr[42377] = 649407264;
assign addr[42378] = 667608730;
assign addr[42379] = 685757258;
assign addr[42380] = 703851410;
assign addr[42381] = 721889752;
assign addr[42382] = 739870851;
assign addr[42383] = 757793284;
assign addr[42384] = 775655628;
assign addr[42385] = 793456467;
assign addr[42386] = 811194391;
assign addr[42387] = 828867991;
assign addr[42388] = 846475867;
assign addr[42389] = 864016623;
assign addr[42390] = 881488868;
assign addr[42391] = 898891215;
assign addr[42392] = 916222287;
assign addr[42393] = 933480707;
assign addr[42394] = 950665109;
assign addr[42395] = 967774128;
assign addr[42396] = 984806408;
assign addr[42397] = 1001760600;
assign addr[42398] = 1018635358;
assign addr[42399] = 1035429345;
assign addr[42400] = 1052141228;
assign addr[42401] = 1068769683;
assign addr[42402] = 1085313391;
assign addr[42403] = 1101771040;
assign addr[42404] = 1118141326;
assign addr[42405] = 1134422949;
assign addr[42406] = 1150614620;
assign addr[42407] = 1166715055;
assign addr[42408] = 1182722976;
assign addr[42409] = 1198637114;
assign addr[42410] = 1214456207;
assign addr[42411] = 1230179002;
assign addr[42412] = 1245804251;
assign addr[42413] = 1261330715;
assign addr[42414] = 1276757164;
assign addr[42415] = 1292082373;
assign addr[42416] = 1307305128;
assign addr[42417] = 1322424222;
assign addr[42418] = 1337438456;
assign addr[42419] = 1352346639;
assign addr[42420] = 1367147589;
assign addr[42421] = 1381840133;
assign addr[42422] = 1396423105;
assign addr[42423] = 1410895350;
assign addr[42424] = 1425255719;
assign addr[42425] = 1439503074;
assign addr[42426] = 1453636285;
assign addr[42427] = 1467654232;
assign addr[42428] = 1481555802;
assign addr[42429] = 1495339895;
assign addr[42430] = 1509005416;
assign addr[42431] = 1522551282;
assign addr[42432] = 1535976419;
assign addr[42433] = 1549279763;
assign addr[42434] = 1562460258;
assign addr[42435] = 1575516860;
assign addr[42436] = 1588448533;
assign addr[42437] = 1601254251;
assign addr[42438] = 1613933000;
assign addr[42439] = 1626483774;
assign addr[42440] = 1638905577;
assign addr[42441] = 1651197426;
assign addr[42442] = 1663358344;
assign addr[42443] = 1675387369;
assign addr[42444] = 1687283545;
assign addr[42445] = 1699045930;
assign addr[42446] = 1710673591;
assign addr[42447] = 1722165606;
assign addr[42448] = 1733521064;
assign addr[42449] = 1744739065;
assign addr[42450] = 1755818718;
assign addr[42451] = 1766759146;
assign addr[42452] = 1777559480;
assign addr[42453] = 1788218865;
assign addr[42454] = 1798736454;
assign addr[42455] = 1809111415;
assign addr[42456] = 1819342925;
assign addr[42457] = 1829430172;
assign addr[42458] = 1839372356;
assign addr[42459] = 1849168689;
assign addr[42460] = 1858818395;
assign addr[42461] = 1868320707;
assign addr[42462] = 1877674873;
assign addr[42463] = 1886880151;
assign addr[42464] = 1895935811;
assign addr[42465] = 1904841135;
assign addr[42466] = 1913595416;
assign addr[42467] = 1922197961;
assign addr[42468] = 1930648088;
assign addr[42469] = 1938945125;
assign addr[42470] = 1947088417;
assign addr[42471] = 1955077316;
assign addr[42472] = 1962911189;
assign addr[42473] = 1970589416;
assign addr[42474] = 1978111387;
assign addr[42475] = 1985476506;
assign addr[42476] = 1992684188;
assign addr[42477] = 1999733863;
assign addr[42478] = 2006624971;
assign addr[42479] = 2013356967;
assign addr[42480] = 2019929315;
assign addr[42481] = 2026341495;
assign addr[42482] = 2032592999;
assign addr[42483] = 2038683330;
assign addr[42484] = 2044612007;
assign addr[42485] = 2050378558;
assign addr[42486] = 2055982526;
assign addr[42487] = 2061423468;
assign addr[42488] = 2066700952;
assign addr[42489] = 2071814558;
assign addr[42490] = 2076763883;
assign addr[42491] = 2081548533;
assign addr[42492] = 2086168128;
assign addr[42493] = 2090622304;
assign addr[42494] = 2094910706;
assign addr[42495] = 2099032994;
assign addr[42496] = 2102988841;
assign addr[42497] = 2106777935;
assign addr[42498] = 2110399974;
assign addr[42499] = 2113854671;
assign addr[42500] = 2117141752;
assign addr[42501] = 2120260957;
assign addr[42502] = 2123212038;
assign addr[42503] = 2125994762;
assign addr[42504] = 2128608907;
assign addr[42505] = 2131054266;
assign addr[42506] = 2133330646;
assign addr[42507] = 2135437865;
assign addr[42508] = 2137375758;
assign addr[42509] = 2139144169;
assign addr[42510] = 2140742960;
assign addr[42511] = 2142172003;
assign addr[42512] = 2143431184;
assign addr[42513] = 2144520405;
assign addr[42514] = 2145439578;
assign addr[42515] = 2146188631;
assign addr[42516] = 2146767505;
assign addr[42517] = 2147176152;
assign addr[42518] = 2147414542;
assign addr[42519] = 2147482655;
assign addr[42520] = 2147380486;
assign addr[42521] = 2147108043;
assign addr[42522] = 2146665347;
assign addr[42523] = 2146052433;
assign addr[42524] = 2145269351;
assign addr[42525] = 2144316162;
assign addr[42526] = 2143192942;
assign addr[42527] = 2141899780;
assign addr[42528] = 2140436778;
assign addr[42529] = 2138804053;
assign addr[42530] = 2137001733;
assign addr[42531] = 2135029962;
assign addr[42532] = 2132888897;
assign addr[42533] = 2130578706;
assign addr[42534] = 2128099574;
assign addr[42535] = 2125451696;
assign addr[42536] = 2122635283;
assign addr[42537] = 2119650558;
assign addr[42538] = 2116497758;
assign addr[42539] = 2113177132;
assign addr[42540] = 2109688944;
assign addr[42541] = 2106033471;
assign addr[42542] = 2102211002;
assign addr[42543] = 2098221841;
assign addr[42544] = 2094066304;
assign addr[42545] = 2089744719;
assign addr[42546] = 2085257431;
assign addr[42547] = 2080604795;
assign addr[42548] = 2075787180;
assign addr[42549] = 2070804967;
assign addr[42550] = 2065658552;
assign addr[42551] = 2060348343;
assign addr[42552] = 2054874761;
assign addr[42553] = 2049238240;
assign addr[42554] = 2043439226;
assign addr[42555] = 2037478181;
assign addr[42556] = 2031355576;
assign addr[42557] = 2025071897;
assign addr[42558] = 2018627642;
assign addr[42559] = 2012023322;
assign addr[42560] = 2005259462;
assign addr[42561] = 1998336596;
assign addr[42562] = 1991255274;
assign addr[42563] = 1984016058;
assign addr[42564] = 1976619522;
assign addr[42565] = 1969066252;
assign addr[42566] = 1961356847;
assign addr[42567] = 1953491918;
assign addr[42568] = 1945472089;
assign addr[42569] = 1937297997;
assign addr[42570] = 1928970288;
assign addr[42571] = 1920489624;
assign addr[42572] = 1911856677;
assign addr[42573] = 1903072131;
assign addr[42574] = 1894136683;
assign addr[42575] = 1885051042;
assign addr[42576] = 1875815927;
assign addr[42577] = 1866432072;
assign addr[42578] = 1856900221;
assign addr[42579] = 1847221128;
assign addr[42580] = 1837395562;
assign addr[42581] = 1827424302;
assign addr[42582] = 1817308138;
assign addr[42583] = 1807047873;
assign addr[42584] = 1796644320;
assign addr[42585] = 1786098304;
assign addr[42586] = 1775410662;
assign addr[42587] = 1764582240;
assign addr[42588] = 1753613897;
assign addr[42589] = 1742506504;
assign addr[42590] = 1731260941;
assign addr[42591] = 1719878099;
assign addr[42592] = 1708358881;
assign addr[42593] = 1696704201;
assign addr[42594] = 1684914983;
assign addr[42595] = 1672992161;
assign addr[42596] = 1660936681;
assign addr[42597] = 1648749499;
assign addr[42598] = 1636431582;
assign addr[42599] = 1623983905;
assign addr[42600] = 1611407456;
assign addr[42601] = 1598703233;
assign addr[42602] = 1585872242;
assign addr[42603] = 1572915501;
assign addr[42604] = 1559834037;
assign addr[42605] = 1546628888;
assign addr[42606] = 1533301101;
assign addr[42607] = 1519851733;
assign addr[42608] = 1506281850;
assign addr[42609] = 1492592527;
assign addr[42610] = 1478784851;
assign addr[42611] = 1464859917;
assign addr[42612] = 1450818828;
assign addr[42613] = 1436662698;
assign addr[42614] = 1422392650;
assign addr[42615] = 1408009814;
assign addr[42616] = 1393515332;
assign addr[42617] = 1378910353;
assign addr[42618] = 1364196034;
assign addr[42619] = 1349373543;
assign addr[42620] = 1334444055;
assign addr[42621] = 1319408754;
assign addr[42622] = 1304268832;
assign addr[42623] = 1289025489;
assign addr[42624] = 1273679934;
assign addr[42625] = 1258233384;
assign addr[42626] = 1242687064;
assign addr[42627] = 1227042207;
assign addr[42628] = 1211300053;
assign addr[42629] = 1195461849;
assign addr[42630] = 1179528853;
assign addr[42631] = 1163502328;
assign addr[42632] = 1147383544;
assign addr[42633] = 1131173780;
assign addr[42634] = 1114874320;
assign addr[42635] = 1098486458;
assign addr[42636] = 1082011492;
assign addr[42637] = 1065450729;
assign addr[42638] = 1048805483;
assign addr[42639] = 1032077073;
assign addr[42640] = 1015266825;
assign addr[42641] = 998376073;
assign addr[42642] = 981406156;
assign addr[42643] = 964358420;
assign addr[42644] = 947234215;
assign addr[42645] = 930034901;
assign addr[42646] = 912761841;
assign addr[42647] = 895416404;
assign addr[42648] = 877999966;
assign addr[42649] = 860513908;
assign addr[42650] = 842959617;
assign addr[42651] = 825338484;
assign addr[42652] = 807651907;
assign addr[42653] = 789901288;
assign addr[42654] = 772088034;
assign addr[42655] = 754213559;
assign addr[42656] = 736279279;
assign addr[42657] = 718286617;
assign addr[42658] = 700236999;
assign addr[42659] = 682131857;
assign addr[42660] = 663972625;
assign addr[42661] = 645760745;
assign addr[42662] = 627497660;
assign addr[42663] = 609184818;
assign addr[42664] = 590823671;
assign addr[42665] = 572415676;
assign addr[42666] = 553962291;
assign addr[42667] = 535464981;
assign addr[42668] = 516925212;
assign addr[42669] = 498344454;
assign addr[42670] = 479724180;
assign addr[42671] = 461065866;
assign addr[42672] = 442370993;
assign addr[42673] = 423641043;
assign addr[42674] = 404877501;
assign addr[42675] = 386081854;
assign addr[42676] = 367255594;
assign addr[42677] = 348400212;
assign addr[42678] = 329517204;
assign addr[42679] = 310608068;
assign addr[42680] = 291674302;
assign addr[42681] = 272717408;
assign addr[42682] = 253738890;
assign addr[42683] = 234740251;
assign addr[42684] = 215722999;
assign addr[42685] = 196688642;
assign addr[42686] = 177638688;
assign addr[42687] = 158574649;
assign addr[42688] = 139498035;
assign addr[42689] = 120410361;
assign addr[42690] = 101313138;
assign addr[42691] = 82207882;
assign addr[42692] = 63096108;
assign addr[42693] = 43979330;
assign addr[42694] = 24859065;
assign addr[42695] = 5736829;
assign addr[42696] = -13385863;
assign addr[42697] = -32507492;
assign addr[42698] = -51626544;
assign addr[42699] = -70741503;
assign addr[42700] = -89850852;
assign addr[42701] = -108953076;
assign addr[42702] = -128046661;
assign addr[42703] = -147130093;
assign addr[42704] = -166201858;
assign addr[42705] = -185260444;
assign addr[42706] = -204304341;
assign addr[42707] = -223332037;
assign addr[42708] = -242342025;
assign addr[42709] = -261332796;
assign addr[42710] = -280302845;
assign addr[42711] = -299250668;
assign addr[42712] = -318174762;
assign addr[42713] = -337073627;
assign addr[42714] = -355945764;
assign addr[42715] = -374789676;
assign addr[42716] = -393603870;
assign addr[42717] = -412386854;
assign addr[42718] = -431137138;
assign addr[42719] = -449853235;
assign addr[42720] = -468533662;
assign addr[42721] = -487176937;
assign addr[42722] = -505781581;
assign addr[42723] = -524346121;
assign addr[42724] = -542869083;
assign addr[42725] = -561348998;
assign addr[42726] = -579784402;
assign addr[42727] = -598173833;
assign addr[42728] = -616515832;
assign addr[42729] = -634808946;
assign addr[42730] = -653051723;
assign addr[42731] = -671242716;
assign addr[42732] = -689380485;
assign addr[42733] = -707463589;
assign addr[42734] = -725490597;
assign addr[42735] = -743460077;
assign addr[42736] = -761370605;
assign addr[42737] = -779220762;
assign addr[42738] = -797009130;
assign addr[42739] = -814734301;
assign addr[42740] = -832394869;
assign addr[42741] = -849989433;
assign addr[42742] = -867516597;
assign addr[42743] = -884974973;
assign addr[42744] = -902363176;
assign addr[42745] = -919679827;
assign addr[42746] = -936923553;
assign addr[42747] = -954092986;
assign addr[42748] = -971186766;
assign addr[42749] = -988203537;
assign addr[42750] = -1005141949;
assign addr[42751] = -1022000660;
assign addr[42752] = -1038778332;
assign addr[42753] = -1055473635;
assign addr[42754] = -1072085246;
assign addr[42755] = -1088611847;
assign addr[42756] = -1105052128;
assign addr[42757] = -1121404785;
assign addr[42758] = -1137668521;
assign addr[42759] = -1153842047;
assign addr[42760] = -1169924081;
assign addr[42761] = -1185913346;
assign addr[42762] = -1201808576;
assign addr[42763] = -1217608510;
assign addr[42764] = -1233311895;
assign addr[42765] = -1248917486;
assign addr[42766] = -1264424045;
assign addr[42767] = -1279830344;
assign addr[42768] = -1295135159;
assign addr[42769] = -1310337279;
assign addr[42770] = -1325435496;
assign addr[42771] = -1340428615;
assign addr[42772] = -1355315445;
assign addr[42773] = -1370094808;
assign addr[42774] = -1384765530;
assign addr[42775] = -1399326449;
assign addr[42776] = -1413776410;
assign addr[42777] = -1428114267;
assign addr[42778] = -1442338884;
assign addr[42779] = -1456449131;
assign addr[42780] = -1470443891;
assign addr[42781] = -1484322054;
assign addr[42782] = -1498082520;
assign addr[42783] = -1511724196;
assign addr[42784] = -1525246002;
assign addr[42785] = -1538646865;
assign addr[42786] = -1551925723;
assign addr[42787] = -1565081523;
assign addr[42788] = -1578113222;
assign addr[42789] = -1591019785;
assign addr[42790] = -1603800191;
assign addr[42791] = -1616453425;
assign addr[42792] = -1628978484;
assign addr[42793] = -1641374375;
assign addr[42794] = -1653640115;
assign addr[42795] = -1665774731;
assign addr[42796] = -1677777262;
assign addr[42797] = -1689646755;
assign addr[42798] = -1701382270;
assign addr[42799] = -1712982875;
assign addr[42800] = -1724447652;
assign addr[42801] = -1735775690;
assign addr[42802] = -1746966091;
assign addr[42803] = -1758017969;
assign addr[42804] = -1768930447;
assign addr[42805] = -1779702660;
assign addr[42806] = -1790333753;
assign addr[42807] = -1800822883;
assign addr[42808] = -1811169220;
assign addr[42809] = -1821371941;
assign addr[42810] = -1831430239;
assign addr[42811] = -1841343316;
assign addr[42812] = -1851110385;
assign addr[42813] = -1860730673;
assign addr[42814] = -1870203416;
assign addr[42815] = -1879527863;
assign addr[42816] = -1888703276;
assign addr[42817] = -1897728925;
assign addr[42818] = -1906604097;
assign addr[42819] = -1915328086;
assign addr[42820] = -1923900201;
assign addr[42821] = -1932319763;
assign addr[42822] = -1940586104;
assign addr[42823] = -1948698568;
assign addr[42824] = -1956656513;
assign addr[42825] = -1964459306;
assign addr[42826] = -1972106330;
assign addr[42827] = -1979596978;
assign addr[42828] = -1986930656;
assign addr[42829] = -1994106782;
assign addr[42830] = -2001124788;
assign addr[42831] = -2007984117;
assign addr[42832] = -2014684225;
assign addr[42833] = -2021224581;
assign addr[42834] = -2027604666;
assign addr[42835] = -2033823974;
assign addr[42836] = -2039882013;
assign addr[42837] = -2045778302;
assign addr[42838] = -2051512372;
assign addr[42839] = -2057083771;
assign addr[42840] = -2062492055;
assign addr[42841] = -2067736796;
assign addr[42842] = -2072817579;
assign addr[42843] = -2077733999;
assign addr[42844] = -2082485668;
assign addr[42845] = -2087072209;
assign addr[42846] = -2091493257;
assign addr[42847] = -2095748463;
assign addr[42848] = -2099837489;
assign addr[42849] = -2103760010;
assign addr[42850] = -2107515716;
assign addr[42851] = -2111104309;
assign addr[42852] = -2114525505;
assign addr[42853] = -2117779031;
assign addr[42854] = -2120864631;
assign addr[42855] = -2123782059;
assign addr[42856] = -2126531084;
assign addr[42857] = -2129111488;
assign addr[42858] = -2131523066;
assign addr[42859] = -2133765628;
assign addr[42860] = -2135838995;
assign addr[42861] = -2137743003;
assign addr[42862] = -2139477502;
assign addr[42863] = -2141042352;
assign addr[42864] = -2142437431;
assign addr[42865] = -2143662628;
assign addr[42866] = -2144717846;
assign addr[42867] = -2145603001;
assign addr[42868] = -2146318022;
assign addr[42869] = -2146862854;
assign addr[42870] = -2147237452;
assign addr[42871] = -2147441787;
assign addr[42872] = -2147475844;
assign addr[42873] = -2147339619;
assign addr[42874] = -2147033123;
assign addr[42875] = -2146556380;
assign addr[42876] = -2145909429;
assign addr[42877] = -2145092320;
assign addr[42878] = -2144105118;
assign addr[42879] = -2142947902;
assign addr[42880] = -2141620763;
assign addr[42881] = -2140123807;
assign addr[42882] = -2138457152;
assign addr[42883] = -2136620930;
assign addr[42884] = -2134615288;
assign addr[42885] = -2132440383;
assign addr[42886] = -2130096389;
assign addr[42887] = -2127583492;
assign addr[42888] = -2124901890;
assign addr[42889] = -2122051796;
assign addr[42890] = -2119033436;
assign addr[42891] = -2115847050;
assign addr[42892] = -2112492891;
assign addr[42893] = -2108971223;
assign addr[42894] = -2105282327;
assign addr[42895] = -2101426496;
assign addr[42896] = -2097404033;
assign addr[42897] = -2093215260;
assign addr[42898] = -2088860507;
assign addr[42899] = -2084340120;
assign addr[42900] = -2079654458;
assign addr[42901] = -2074803892;
assign addr[42902] = -2069788807;
assign addr[42903] = -2064609600;
assign addr[42904] = -2059266683;
assign addr[42905] = -2053760478;
assign addr[42906] = -2048091422;
assign addr[42907] = -2042259965;
assign addr[42908] = -2036266570;
assign addr[42909] = -2030111710;
assign addr[42910] = -2023795876;
assign addr[42911] = -2017319567;
assign addr[42912] = -2010683297;
assign addr[42913] = -2003887591;
assign addr[42914] = -1996932990;
assign addr[42915] = -1989820044;
assign addr[42916] = -1982549318;
assign addr[42917] = -1975121388;
assign addr[42918] = -1967536842;
assign addr[42919] = -1959796283;
assign addr[42920] = -1951900324;
assign addr[42921] = -1943849591;
assign addr[42922] = -1935644723;
assign addr[42923] = -1927286370;
assign addr[42924] = -1918775195;
assign addr[42925] = -1910111873;
assign addr[42926] = -1901297091;
assign addr[42927] = -1892331547;
assign addr[42928] = -1883215953;
assign addr[42929] = -1873951032;
assign addr[42930] = -1864537518;
assign addr[42931] = -1854976157;
assign addr[42932] = -1845267708;
assign addr[42933] = -1835412941;
assign addr[42934] = -1825412636;
assign addr[42935] = -1815267588;
assign addr[42936] = -1804978599;
assign addr[42937] = -1794546487;
assign addr[42938] = -1783972079;
assign addr[42939] = -1773256212;
assign addr[42940] = -1762399737;
assign addr[42941] = -1751403515;
assign addr[42942] = -1740268417;
assign addr[42943] = -1728995326;
assign addr[42944] = -1717585136;
assign addr[42945] = -1706038753;
assign addr[42946] = -1694357091;
assign addr[42947] = -1682541077;
assign addr[42948] = -1670591647;
assign addr[42949] = -1658509750;
assign addr[42950] = -1646296344;
assign addr[42951] = -1633952396;
assign addr[42952] = -1621478885;
assign addr[42953] = -1608876801;
assign addr[42954] = -1596147143;
assign addr[42955] = -1583290921;
assign addr[42956] = -1570309153;
assign addr[42957] = -1557202869;
assign addr[42958] = -1543973108;
assign addr[42959] = -1530620920;
assign addr[42960] = -1517147363;
assign addr[42961] = -1503553506;
assign addr[42962] = -1489840425;
assign addr[42963] = -1476009210;
assign addr[42964] = -1462060956;
assign addr[42965] = -1447996770;
assign addr[42966] = -1433817766;
assign addr[42967] = -1419525069;
assign addr[42968] = -1405119813;
assign addr[42969] = -1390603139;
assign addr[42970] = -1375976199;
assign addr[42971] = -1361240152;
assign addr[42972] = -1346396168;
assign addr[42973] = -1331445422;
assign addr[42974] = -1316389101;
assign addr[42975] = -1301228398;
assign addr[42976] = -1285964516;
assign addr[42977] = -1270598665;
assign addr[42978] = -1255132063;
assign addr[42979] = -1239565936;
assign addr[42980] = -1223901520;
assign addr[42981] = -1208140056;
assign addr[42982] = -1192282793;
assign addr[42983] = -1176330990;
assign addr[42984] = -1160285911;
assign addr[42985] = -1144148829;
assign addr[42986] = -1127921022;
assign addr[42987] = -1111603778;
assign addr[42988] = -1095198391;
assign addr[42989] = -1078706161;
assign addr[42990] = -1062128397;
assign addr[42991] = -1045466412;
assign addr[42992] = -1028721528;
assign addr[42993] = -1011895073;
assign addr[42994] = -994988380;
assign addr[42995] = -978002791;
assign addr[42996] = -960939653;
assign addr[42997] = -943800318;
assign addr[42998] = -926586145;
assign addr[42999] = -909298500;
assign addr[43000] = -891938752;
assign addr[43001] = -874508280;
assign addr[43002] = -857008464;
assign addr[43003] = -839440693;
assign addr[43004] = -821806359;
assign addr[43005] = -804106861;
assign addr[43006] = -786343603;
assign addr[43007] = -768517992;
assign addr[43008] = -750631442;
assign addr[43009] = -732685372;
assign addr[43010] = -714681204;
assign addr[43011] = -696620367;
assign addr[43012] = -678504291;
assign addr[43013] = -660334415;
assign addr[43014] = -642112178;
assign addr[43015] = -623839025;
assign addr[43016] = -605516406;
assign addr[43017] = -587145773;
assign addr[43018] = -568728583;
assign addr[43019] = -550266296;
assign addr[43020] = -531760377;
assign addr[43021] = -513212292;
assign addr[43022] = -494623513;
assign addr[43023] = -475995513;
assign addr[43024] = -457329769;
assign addr[43025] = -438627762;
assign addr[43026] = -419890975;
assign addr[43027] = -401120892;
assign addr[43028] = -382319004;
assign addr[43029] = -363486799;
assign addr[43030] = -344625773;
assign addr[43031] = -325737419;
assign addr[43032] = -306823237;
assign addr[43033] = -287884725;
assign addr[43034] = -268923386;
assign addr[43035] = -249940723;
assign addr[43036] = -230938242;
assign addr[43037] = -211917448;
assign addr[43038] = -192879850;
assign addr[43039] = -173826959;
assign addr[43040] = -154760284;
assign addr[43041] = -135681337;
assign addr[43042] = -116591632;
assign addr[43043] = -97492681;
assign addr[43044] = -78386000;
assign addr[43045] = -59273104;
assign addr[43046] = -40155507;
assign addr[43047] = -21034727;
assign addr[43048] = -1912278;
assign addr[43049] = 17210322;
assign addr[43050] = 36331557;
assign addr[43051] = 55449912;
assign addr[43052] = 74563870;
assign addr[43053] = 93671915;
assign addr[43054] = 112772533;
assign addr[43055] = 131864208;
assign addr[43056] = 150945428;
assign addr[43057] = 170014678;
assign addr[43058] = 189070447;
assign addr[43059] = 208111224;
assign addr[43060] = 227135500;
assign addr[43061] = 246141764;
assign addr[43062] = 265128512;
assign addr[43063] = 284094236;
assign addr[43064] = 303037433;
assign addr[43065] = 321956601;
assign addr[43066] = 340850240;
assign addr[43067] = 359716852;
assign addr[43068] = 378554940;
assign addr[43069] = 397363011;
assign addr[43070] = 416139574;
assign addr[43071] = 434883140;
assign addr[43072] = 453592221;
assign addr[43073] = 472265336;
assign addr[43074] = 490901003;
assign addr[43075] = 509497745;
assign addr[43076] = 528054086;
assign addr[43077] = 546568556;
assign addr[43078] = 565039687;
assign addr[43079] = 583466013;
assign addr[43080] = 601846074;
assign addr[43081] = 620178412;
assign addr[43082] = 638461574;
assign addr[43083] = 656694110;
assign addr[43084] = 674874574;
assign addr[43085] = 693001525;
assign addr[43086] = 711073524;
assign addr[43087] = 729089140;
assign addr[43088] = 747046944;
assign addr[43089] = 764945512;
assign addr[43090] = 782783424;
assign addr[43091] = 800559266;
assign addr[43092] = 818271628;
assign addr[43093] = 835919107;
assign addr[43094] = 853500302;
assign addr[43095] = 871013820;
assign addr[43096] = 888458272;
assign addr[43097] = 905832274;
assign addr[43098] = 923134450;
assign addr[43099] = 940363427;
assign addr[43100] = 957517838;
assign addr[43101] = 974596324;
assign addr[43102] = 991597531;
assign addr[43103] = 1008520110;
assign addr[43104] = 1025362720;
assign addr[43105] = 1042124025;
assign addr[43106] = 1058802695;
assign addr[43107] = 1075397409;
assign addr[43108] = 1091906851;
assign addr[43109] = 1108329711;
assign addr[43110] = 1124664687;
assign addr[43111] = 1140910484;
assign addr[43112] = 1157065814;
assign addr[43113] = 1173129396;
assign addr[43114] = 1189099956;
assign addr[43115] = 1204976227;
assign addr[43116] = 1220756951;
assign addr[43117] = 1236440877;
assign addr[43118] = 1252026760;
assign addr[43119] = 1267513365;
assign addr[43120] = 1282899464;
assign addr[43121] = 1298183838;
assign addr[43122] = 1313365273;
assign addr[43123] = 1328442566;
assign addr[43124] = 1343414522;
assign addr[43125] = 1358279953;
assign addr[43126] = 1373037681;
assign addr[43127] = 1387686535;
assign addr[43128] = 1402225355;
assign addr[43129] = 1416652986;
assign addr[43130] = 1430968286;
assign addr[43131] = 1445170118;
assign addr[43132] = 1459257358;
assign addr[43133] = 1473228887;
assign addr[43134] = 1487083598;
assign addr[43135] = 1500820393;
assign addr[43136] = 1514438181;
assign addr[43137] = 1527935884;
assign addr[43138] = 1541312431;
assign addr[43139] = 1554566762;
assign addr[43140] = 1567697824;
assign addr[43141] = 1580704578;
assign addr[43142] = 1593585992;
assign addr[43143] = 1606341043;
assign addr[43144] = 1618968722;
assign addr[43145] = 1631468027;
assign addr[43146] = 1643837966;
assign addr[43147] = 1656077559;
assign addr[43148] = 1668185835;
assign addr[43149] = 1680161834;
assign addr[43150] = 1692004606;
assign addr[43151] = 1703713213;
assign addr[43152] = 1715286726;
assign addr[43153] = 1726724227;
assign addr[43154] = 1738024810;
assign addr[43155] = 1749187577;
assign addr[43156] = 1760211645;
assign addr[43157] = 1771096139;
assign addr[43158] = 1781840195;
assign addr[43159] = 1792442963;
assign addr[43160] = 1802903601;
assign addr[43161] = 1813221279;
assign addr[43162] = 1823395180;
assign addr[43163] = 1833424497;
assign addr[43164] = 1843308435;
assign addr[43165] = 1853046210;
assign addr[43166] = 1862637049;
assign addr[43167] = 1872080193;
assign addr[43168] = 1881374892;
assign addr[43169] = 1890520410;
assign addr[43170] = 1899516021;
assign addr[43171] = 1908361011;
assign addr[43172] = 1917054681;
assign addr[43173] = 1925596340;
assign addr[43174] = 1933985310;
assign addr[43175] = 1942220928;
assign addr[43176] = 1950302539;
assign addr[43177] = 1958229503;
assign addr[43178] = 1966001192;
assign addr[43179] = 1973616989;
assign addr[43180] = 1981076290;
assign addr[43181] = 1988378503;
assign addr[43182] = 1995523051;
assign addr[43183] = 2002509365;
assign addr[43184] = 2009336893;
assign addr[43185] = 2016005093;
assign addr[43186] = 2022513436;
assign addr[43187] = 2028861406;
assign addr[43188] = 2035048499;
assign addr[43189] = 2041074226;
assign addr[43190] = 2046938108;
assign addr[43191] = 2052639680;
assign addr[43192] = 2058178491;
assign addr[43193] = 2063554100;
assign addr[43194] = 2068766083;
assign addr[43195] = 2073814024;
assign addr[43196] = 2078697525;
assign addr[43197] = 2083416198;
assign addr[43198] = 2087969669;
assign addr[43199] = 2092357577;
assign addr[43200] = 2096579573;
assign addr[43201] = 2100635323;
assign addr[43202] = 2104524506;
assign addr[43203] = 2108246813;
assign addr[43204] = 2111801949;
assign addr[43205] = 2115189632;
assign addr[43206] = 2118409593;
assign addr[43207] = 2121461578;
assign addr[43208] = 2124345343;
assign addr[43209] = 2127060661;
assign addr[43210] = 2129607316;
assign addr[43211] = 2131985106;
assign addr[43212] = 2134193842;
assign addr[43213] = 2136233350;
assign addr[43214] = 2138103468;
assign addr[43215] = 2139804048;
assign addr[43216] = 2141334954;
assign addr[43217] = 2142696065;
assign addr[43218] = 2143887273;
assign addr[43219] = 2144908484;
assign addr[43220] = 2145759618;
assign addr[43221] = 2146440605;
assign addr[43222] = 2146951393;
assign addr[43223] = 2147291941;
assign addr[43224] = 2147462221;
assign addr[43225] = 2147462221;
assign addr[43226] = 2147291941;
assign addr[43227] = 2146951393;
assign addr[43228] = 2146440605;
assign addr[43229] = 2145759618;
assign addr[43230] = 2144908484;
assign addr[43231] = 2143887273;
assign addr[43232] = 2142696065;
assign addr[43233] = 2141334954;
assign addr[43234] = 2139804048;
assign addr[43235] = 2138103468;
assign addr[43236] = 2136233350;
assign addr[43237] = 2134193842;
assign addr[43238] = 2131985106;
assign addr[43239] = 2129607316;
assign addr[43240] = 2127060661;
assign addr[43241] = 2124345343;
assign addr[43242] = 2121461578;
assign addr[43243] = 2118409593;
assign addr[43244] = 2115189632;
assign addr[43245] = 2111801949;
assign addr[43246] = 2108246813;
assign addr[43247] = 2104524506;
assign addr[43248] = 2100635323;
assign addr[43249] = 2096579573;
assign addr[43250] = 2092357577;
assign addr[43251] = 2087969669;
assign addr[43252] = 2083416198;
assign addr[43253] = 2078697525;
assign addr[43254] = 2073814024;
assign addr[43255] = 2068766083;
assign addr[43256] = 2063554100;
assign addr[43257] = 2058178491;
assign addr[43258] = 2052639680;
assign addr[43259] = 2046938108;
assign addr[43260] = 2041074226;
assign addr[43261] = 2035048499;
assign addr[43262] = 2028861406;
assign addr[43263] = 2022513436;
assign addr[43264] = 2016005093;
assign addr[43265] = 2009336893;
assign addr[43266] = 2002509365;
assign addr[43267] = 1995523051;
assign addr[43268] = 1988378503;
assign addr[43269] = 1981076290;
assign addr[43270] = 1973616989;
assign addr[43271] = 1966001192;
assign addr[43272] = 1958229503;
assign addr[43273] = 1950302539;
assign addr[43274] = 1942220928;
assign addr[43275] = 1933985310;
assign addr[43276] = 1925596340;
assign addr[43277] = 1917054681;
assign addr[43278] = 1908361011;
assign addr[43279] = 1899516021;
assign addr[43280] = 1890520410;
assign addr[43281] = 1881374892;
assign addr[43282] = 1872080193;
assign addr[43283] = 1862637049;
assign addr[43284] = 1853046210;
assign addr[43285] = 1843308435;
assign addr[43286] = 1833424497;
assign addr[43287] = 1823395180;
assign addr[43288] = 1813221279;
assign addr[43289] = 1802903601;
assign addr[43290] = 1792442963;
assign addr[43291] = 1781840195;
assign addr[43292] = 1771096139;
assign addr[43293] = 1760211645;
assign addr[43294] = 1749187577;
assign addr[43295] = 1738024810;
assign addr[43296] = 1726724227;
assign addr[43297] = 1715286726;
assign addr[43298] = 1703713213;
assign addr[43299] = 1692004606;
assign addr[43300] = 1680161834;
assign addr[43301] = 1668185835;
assign addr[43302] = 1656077559;
assign addr[43303] = 1643837966;
assign addr[43304] = 1631468027;
assign addr[43305] = 1618968722;
assign addr[43306] = 1606341043;
assign addr[43307] = 1593585992;
assign addr[43308] = 1580704578;
assign addr[43309] = 1567697824;
assign addr[43310] = 1554566762;
assign addr[43311] = 1541312431;
assign addr[43312] = 1527935884;
assign addr[43313] = 1514438181;
assign addr[43314] = 1500820393;
assign addr[43315] = 1487083598;
assign addr[43316] = 1473228887;
assign addr[43317] = 1459257358;
assign addr[43318] = 1445170118;
assign addr[43319] = 1430968286;
assign addr[43320] = 1416652986;
assign addr[43321] = 1402225355;
assign addr[43322] = 1387686535;
assign addr[43323] = 1373037681;
assign addr[43324] = 1358279953;
assign addr[43325] = 1343414522;
assign addr[43326] = 1328442566;
assign addr[43327] = 1313365273;
assign addr[43328] = 1298183838;
assign addr[43329] = 1282899464;
assign addr[43330] = 1267513365;
assign addr[43331] = 1252026760;
assign addr[43332] = 1236440877;
assign addr[43333] = 1220756951;
assign addr[43334] = 1204976227;
assign addr[43335] = 1189099956;
assign addr[43336] = 1173129396;
assign addr[43337] = 1157065814;
assign addr[43338] = 1140910484;
assign addr[43339] = 1124664687;
assign addr[43340] = 1108329711;
assign addr[43341] = 1091906851;
assign addr[43342] = 1075397409;
assign addr[43343] = 1058802695;
assign addr[43344] = 1042124025;
assign addr[43345] = 1025362720;
assign addr[43346] = 1008520110;
assign addr[43347] = 991597531;
assign addr[43348] = 974596324;
assign addr[43349] = 957517838;
assign addr[43350] = 940363427;
assign addr[43351] = 923134450;
assign addr[43352] = 905832274;
assign addr[43353] = 888458272;
assign addr[43354] = 871013820;
assign addr[43355] = 853500302;
assign addr[43356] = 835919107;
assign addr[43357] = 818271628;
assign addr[43358] = 800559266;
assign addr[43359] = 782783424;
assign addr[43360] = 764945512;
assign addr[43361] = 747046944;
assign addr[43362] = 729089140;
assign addr[43363] = 711073524;
assign addr[43364] = 693001525;
assign addr[43365] = 674874574;
assign addr[43366] = 656694110;
assign addr[43367] = 638461574;
assign addr[43368] = 620178412;
assign addr[43369] = 601846074;
assign addr[43370] = 583466013;
assign addr[43371] = 565039687;
assign addr[43372] = 546568556;
assign addr[43373] = 528054086;
assign addr[43374] = 509497745;
assign addr[43375] = 490901003;
assign addr[43376] = 472265336;
assign addr[43377] = 453592221;
assign addr[43378] = 434883140;
assign addr[43379] = 416139574;
assign addr[43380] = 397363011;
assign addr[43381] = 378554940;
assign addr[43382] = 359716852;
assign addr[43383] = 340850240;
assign addr[43384] = 321956601;
assign addr[43385] = 303037433;
assign addr[43386] = 284094236;
assign addr[43387] = 265128512;
assign addr[43388] = 246141764;
assign addr[43389] = 227135500;
assign addr[43390] = 208111224;
assign addr[43391] = 189070447;
assign addr[43392] = 170014678;
assign addr[43393] = 150945428;
assign addr[43394] = 131864208;
assign addr[43395] = 112772533;
assign addr[43396] = 93671915;
assign addr[43397] = 74563870;
assign addr[43398] = 55449912;
assign addr[43399] = 36331557;
assign addr[43400] = 17210322;
assign addr[43401] = -1912278;
assign addr[43402] = -21034727;
assign addr[43403] = -40155507;
assign addr[43404] = -59273104;
assign addr[43405] = -78386000;
assign addr[43406] = -97492681;
assign addr[43407] = -116591632;
assign addr[43408] = -135681337;
assign addr[43409] = -154760284;
assign addr[43410] = -173826959;
assign addr[43411] = -192879850;
assign addr[43412] = -211917448;
assign addr[43413] = -230938242;
assign addr[43414] = -249940723;
assign addr[43415] = -268923386;
assign addr[43416] = -287884725;
assign addr[43417] = -306823237;
assign addr[43418] = -325737419;
assign addr[43419] = -344625773;
assign addr[43420] = -363486799;
assign addr[43421] = -382319004;
assign addr[43422] = -401120892;
assign addr[43423] = -419890975;
assign addr[43424] = -438627762;
assign addr[43425] = -457329769;
assign addr[43426] = -475995513;
assign addr[43427] = -494623513;
assign addr[43428] = -513212292;
assign addr[43429] = -531760377;
assign addr[43430] = -550266296;
assign addr[43431] = -568728583;
assign addr[43432] = -587145773;
assign addr[43433] = -605516406;
assign addr[43434] = -623839025;
assign addr[43435] = -642112178;
assign addr[43436] = -660334415;
assign addr[43437] = -678504291;
assign addr[43438] = -696620367;
assign addr[43439] = -714681204;
assign addr[43440] = -732685372;
assign addr[43441] = -750631442;
assign addr[43442] = -768517992;
assign addr[43443] = -786343603;
assign addr[43444] = -804106861;
assign addr[43445] = -821806359;
assign addr[43446] = -839440693;
assign addr[43447] = -857008464;
assign addr[43448] = -874508280;
assign addr[43449] = -891938752;
assign addr[43450] = -909298500;
assign addr[43451] = -926586145;
assign addr[43452] = -943800318;
assign addr[43453] = -960939653;
assign addr[43454] = -978002791;
assign addr[43455] = -994988380;
assign addr[43456] = -1011895073;
assign addr[43457] = -1028721528;
assign addr[43458] = -1045466412;
assign addr[43459] = -1062128397;
assign addr[43460] = -1078706161;
assign addr[43461] = -1095198391;
assign addr[43462] = -1111603778;
assign addr[43463] = -1127921022;
assign addr[43464] = -1144148829;
assign addr[43465] = -1160285911;
assign addr[43466] = -1176330990;
assign addr[43467] = -1192282793;
assign addr[43468] = -1208140056;
assign addr[43469] = -1223901520;
assign addr[43470] = -1239565936;
assign addr[43471] = -1255132063;
assign addr[43472] = -1270598665;
assign addr[43473] = -1285964516;
assign addr[43474] = -1301228398;
assign addr[43475] = -1316389101;
assign addr[43476] = -1331445422;
assign addr[43477] = -1346396168;
assign addr[43478] = -1361240152;
assign addr[43479] = -1375976199;
assign addr[43480] = -1390603139;
assign addr[43481] = -1405119813;
assign addr[43482] = -1419525069;
assign addr[43483] = -1433817766;
assign addr[43484] = -1447996770;
assign addr[43485] = -1462060956;
assign addr[43486] = -1476009210;
assign addr[43487] = -1489840425;
assign addr[43488] = -1503553506;
assign addr[43489] = -1517147363;
assign addr[43490] = -1530620920;
assign addr[43491] = -1543973108;
assign addr[43492] = -1557202869;
assign addr[43493] = -1570309153;
assign addr[43494] = -1583290921;
assign addr[43495] = -1596147143;
assign addr[43496] = -1608876801;
assign addr[43497] = -1621478885;
assign addr[43498] = -1633952396;
assign addr[43499] = -1646296344;
assign addr[43500] = -1658509750;
assign addr[43501] = -1670591647;
assign addr[43502] = -1682541077;
assign addr[43503] = -1694357091;
assign addr[43504] = -1706038753;
assign addr[43505] = -1717585136;
assign addr[43506] = -1728995326;
assign addr[43507] = -1740268417;
assign addr[43508] = -1751403515;
assign addr[43509] = -1762399737;
assign addr[43510] = -1773256212;
assign addr[43511] = -1783972079;
assign addr[43512] = -1794546487;
assign addr[43513] = -1804978599;
assign addr[43514] = -1815267588;
assign addr[43515] = -1825412636;
assign addr[43516] = -1835412941;
assign addr[43517] = -1845267708;
assign addr[43518] = -1854976157;
assign addr[43519] = -1864537518;
assign addr[43520] = -1873951032;
assign addr[43521] = -1883215953;
assign addr[43522] = -1892331547;
assign addr[43523] = -1901297091;
assign addr[43524] = -1910111873;
assign addr[43525] = -1918775195;
assign addr[43526] = -1927286370;
assign addr[43527] = -1935644723;
assign addr[43528] = -1943849591;
assign addr[43529] = -1951900324;
assign addr[43530] = -1959796283;
assign addr[43531] = -1967536842;
assign addr[43532] = -1975121388;
assign addr[43533] = -1982549318;
assign addr[43534] = -1989820044;
assign addr[43535] = -1996932990;
assign addr[43536] = -2003887591;
assign addr[43537] = -2010683297;
assign addr[43538] = -2017319567;
assign addr[43539] = -2023795876;
assign addr[43540] = -2030111710;
assign addr[43541] = -2036266570;
assign addr[43542] = -2042259965;
assign addr[43543] = -2048091422;
assign addr[43544] = -2053760478;
assign addr[43545] = -2059266683;
assign addr[43546] = -2064609600;
assign addr[43547] = -2069788807;
assign addr[43548] = -2074803892;
assign addr[43549] = -2079654458;
assign addr[43550] = -2084340120;
assign addr[43551] = -2088860507;
assign addr[43552] = -2093215260;
assign addr[43553] = -2097404033;
assign addr[43554] = -2101426496;
assign addr[43555] = -2105282327;
assign addr[43556] = -2108971223;
assign addr[43557] = -2112492891;
assign addr[43558] = -2115847050;
assign addr[43559] = -2119033436;
assign addr[43560] = -2122051796;
assign addr[43561] = -2124901890;
assign addr[43562] = -2127583492;
assign addr[43563] = -2130096389;
assign addr[43564] = -2132440383;
assign addr[43565] = -2134615288;
assign addr[43566] = -2136620930;
assign addr[43567] = -2138457152;
assign addr[43568] = -2140123807;
assign addr[43569] = -2141620763;
assign addr[43570] = -2142947902;
assign addr[43571] = -2144105118;
assign addr[43572] = -2145092320;
assign addr[43573] = -2145909429;
assign addr[43574] = -2146556380;
assign addr[43575] = -2147033123;
assign addr[43576] = -2147339619;
assign addr[43577] = -2147475844;
assign addr[43578] = -2147441787;
assign addr[43579] = -2147237452;
assign addr[43580] = -2146862854;
assign addr[43581] = -2146318022;
assign addr[43582] = -2145603001;
assign addr[43583] = -2144717846;
assign addr[43584] = -2143662628;
assign addr[43585] = -2142437431;
assign addr[43586] = -2141042352;
assign addr[43587] = -2139477502;
assign addr[43588] = -2137743003;
assign addr[43589] = -2135838995;
assign addr[43590] = -2133765628;
assign addr[43591] = -2131523066;
assign addr[43592] = -2129111488;
assign addr[43593] = -2126531084;
assign addr[43594] = -2123782059;
assign addr[43595] = -2120864631;
assign addr[43596] = -2117779031;
assign addr[43597] = -2114525505;
assign addr[43598] = -2111104309;
assign addr[43599] = -2107515716;
assign addr[43600] = -2103760010;
assign addr[43601] = -2099837489;
assign addr[43602] = -2095748463;
assign addr[43603] = -2091493257;
assign addr[43604] = -2087072209;
assign addr[43605] = -2082485668;
assign addr[43606] = -2077733999;
assign addr[43607] = -2072817579;
assign addr[43608] = -2067736796;
assign addr[43609] = -2062492055;
assign addr[43610] = -2057083771;
assign addr[43611] = -2051512372;
assign addr[43612] = -2045778302;
assign addr[43613] = -2039882013;
assign addr[43614] = -2033823974;
assign addr[43615] = -2027604666;
assign addr[43616] = -2021224581;
assign addr[43617] = -2014684225;
assign addr[43618] = -2007984117;
assign addr[43619] = -2001124788;
assign addr[43620] = -1994106782;
assign addr[43621] = -1986930656;
assign addr[43622] = -1979596978;
assign addr[43623] = -1972106330;
assign addr[43624] = -1964459306;
assign addr[43625] = -1956656513;
assign addr[43626] = -1948698568;
assign addr[43627] = -1940586104;
assign addr[43628] = -1932319763;
assign addr[43629] = -1923900201;
assign addr[43630] = -1915328086;
assign addr[43631] = -1906604097;
assign addr[43632] = -1897728925;
assign addr[43633] = -1888703276;
assign addr[43634] = -1879527863;
assign addr[43635] = -1870203416;
assign addr[43636] = -1860730673;
assign addr[43637] = -1851110385;
assign addr[43638] = -1841343316;
assign addr[43639] = -1831430239;
assign addr[43640] = -1821371941;
assign addr[43641] = -1811169220;
assign addr[43642] = -1800822883;
assign addr[43643] = -1790333753;
assign addr[43644] = -1779702660;
assign addr[43645] = -1768930447;
assign addr[43646] = -1758017969;
assign addr[43647] = -1746966091;
assign addr[43648] = -1735775690;
assign addr[43649] = -1724447652;
assign addr[43650] = -1712982875;
assign addr[43651] = -1701382270;
assign addr[43652] = -1689646755;
assign addr[43653] = -1677777262;
assign addr[43654] = -1665774731;
assign addr[43655] = -1653640115;
assign addr[43656] = -1641374375;
assign addr[43657] = -1628978484;
assign addr[43658] = -1616453425;
assign addr[43659] = -1603800191;
assign addr[43660] = -1591019785;
assign addr[43661] = -1578113222;
assign addr[43662] = -1565081523;
assign addr[43663] = -1551925723;
assign addr[43664] = -1538646865;
assign addr[43665] = -1525246002;
assign addr[43666] = -1511724196;
assign addr[43667] = -1498082520;
assign addr[43668] = -1484322054;
assign addr[43669] = -1470443891;
assign addr[43670] = -1456449131;
assign addr[43671] = -1442338884;
assign addr[43672] = -1428114267;
assign addr[43673] = -1413776410;
assign addr[43674] = -1399326449;
assign addr[43675] = -1384765530;
assign addr[43676] = -1370094808;
assign addr[43677] = -1355315445;
assign addr[43678] = -1340428615;
assign addr[43679] = -1325435496;
assign addr[43680] = -1310337279;
assign addr[43681] = -1295135159;
assign addr[43682] = -1279830344;
assign addr[43683] = -1264424045;
assign addr[43684] = -1248917486;
assign addr[43685] = -1233311895;
assign addr[43686] = -1217608510;
assign addr[43687] = -1201808576;
assign addr[43688] = -1185913346;
assign addr[43689] = -1169924081;
assign addr[43690] = -1153842047;
assign addr[43691] = -1137668521;
assign addr[43692] = -1121404785;
assign addr[43693] = -1105052128;
assign addr[43694] = -1088611847;
assign addr[43695] = -1072085246;
assign addr[43696] = -1055473635;
assign addr[43697] = -1038778332;
assign addr[43698] = -1022000660;
assign addr[43699] = -1005141949;
assign addr[43700] = -988203537;
assign addr[43701] = -971186766;
assign addr[43702] = -954092986;
assign addr[43703] = -936923553;
assign addr[43704] = -919679827;
assign addr[43705] = -902363176;
assign addr[43706] = -884974973;
assign addr[43707] = -867516597;
assign addr[43708] = -849989433;
assign addr[43709] = -832394869;
assign addr[43710] = -814734301;
assign addr[43711] = -797009130;
assign addr[43712] = -779220762;
assign addr[43713] = -761370605;
assign addr[43714] = -743460077;
assign addr[43715] = -725490597;
assign addr[43716] = -707463589;
assign addr[43717] = -689380485;
assign addr[43718] = -671242716;
assign addr[43719] = -653051723;
assign addr[43720] = -634808946;
assign addr[43721] = -616515832;
assign addr[43722] = -598173833;
assign addr[43723] = -579784402;
assign addr[43724] = -561348998;
assign addr[43725] = -542869083;
assign addr[43726] = -524346121;
assign addr[43727] = -505781581;
assign addr[43728] = -487176937;
assign addr[43729] = -468533662;
assign addr[43730] = -449853235;
assign addr[43731] = -431137138;
assign addr[43732] = -412386854;
assign addr[43733] = -393603870;
assign addr[43734] = -374789676;
assign addr[43735] = -355945764;
assign addr[43736] = -337073627;
assign addr[43737] = -318174762;
assign addr[43738] = -299250668;
assign addr[43739] = -280302845;
assign addr[43740] = -261332796;
assign addr[43741] = -242342025;
assign addr[43742] = -223332037;
assign addr[43743] = -204304341;
assign addr[43744] = -185260444;
assign addr[43745] = -166201858;
assign addr[43746] = -147130093;
assign addr[43747] = -128046661;
assign addr[43748] = -108953076;
assign addr[43749] = -89850852;
assign addr[43750] = -70741503;
assign addr[43751] = -51626544;
assign addr[43752] = -32507492;
assign addr[43753] = -13385863;
assign addr[43754] = 5736829;
assign addr[43755] = 24859065;
assign addr[43756] = 43979330;
assign addr[43757] = 63096108;
assign addr[43758] = 82207882;
assign addr[43759] = 101313138;
assign addr[43760] = 120410361;
assign addr[43761] = 139498035;
assign addr[43762] = 158574649;
assign addr[43763] = 177638688;
assign addr[43764] = 196688642;
assign addr[43765] = 215722999;
assign addr[43766] = 234740251;
assign addr[43767] = 253738890;
assign addr[43768] = 272717408;
assign addr[43769] = 291674302;
assign addr[43770] = 310608068;
assign addr[43771] = 329517204;
assign addr[43772] = 348400212;
assign addr[43773] = 367255594;
assign addr[43774] = 386081854;
assign addr[43775] = 404877501;
assign addr[43776] = 423641043;
assign addr[43777] = 442370993;
assign addr[43778] = 461065866;
assign addr[43779] = 479724180;
assign addr[43780] = 498344454;
assign addr[43781] = 516925212;
assign addr[43782] = 535464981;
assign addr[43783] = 553962291;
assign addr[43784] = 572415676;
assign addr[43785] = 590823671;
assign addr[43786] = 609184818;
assign addr[43787] = 627497660;
assign addr[43788] = 645760745;
assign addr[43789] = 663972625;
assign addr[43790] = 682131857;
assign addr[43791] = 700236999;
assign addr[43792] = 718286617;
assign addr[43793] = 736279279;
assign addr[43794] = 754213559;
assign addr[43795] = 772088034;
assign addr[43796] = 789901288;
assign addr[43797] = 807651907;
assign addr[43798] = 825338484;
assign addr[43799] = 842959617;
assign addr[43800] = 860513908;
assign addr[43801] = 877999966;
assign addr[43802] = 895416404;
assign addr[43803] = 912761841;
assign addr[43804] = 930034901;
assign addr[43805] = 947234215;
assign addr[43806] = 964358420;
assign addr[43807] = 981406156;
assign addr[43808] = 998376073;
assign addr[43809] = 1015266825;
assign addr[43810] = 1032077073;
assign addr[43811] = 1048805483;
assign addr[43812] = 1065450729;
assign addr[43813] = 1082011492;
assign addr[43814] = 1098486458;
assign addr[43815] = 1114874320;
assign addr[43816] = 1131173780;
assign addr[43817] = 1147383544;
assign addr[43818] = 1163502328;
assign addr[43819] = 1179528853;
assign addr[43820] = 1195461849;
assign addr[43821] = 1211300053;
assign addr[43822] = 1227042207;
assign addr[43823] = 1242687064;
assign addr[43824] = 1258233384;
assign addr[43825] = 1273679934;
assign addr[43826] = 1289025489;
assign addr[43827] = 1304268832;
assign addr[43828] = 1319408754;
assign addr[43829] = 1334444055;
assign addr[43830] = 1349373543;
assign addr[43831] = 1364196034;
assign addr[43832] = 1378910353;
assign addr[43833] = 1393515332;
assign addr[43834] = 1408009814;
assign addr[43835] = 1422392650;
assign addr[43836] = 1436662698;
assign addr[43837] = 1450818828;
assign addr[43838] = 1464859917;
assign addr[43839] = 1478784851;
assign addr[43840] = 1492592527;
assign addr[43841] = 1506281850;
assign addr[43842] = 1519851733;
assign addr[43843] = 1533301101;
assign addr[43844] = 1546628888;
assign addr[43845] = 1559834037;
assign addr[43846] = 1572915501;
assign addr[43847] = 1585872242;
assign addr[43848] = 1598703233;
assign addr[43849] = 1611407456;
assign addr[43850] = 1623983905;
assign addr[43851] = 1636431582;
assign addr[43852] = 1648749499;
assign addr[43853] = 1660936681;
assign addr[43854] = 1672992161;
assign addr[43855] = 1684914983;
assign addr[43856] = 1696704201;
assign addr[43857] = 1708358881;
assign addr[43858] = 1719878099;
assign addr[43859] = 1731260941;
assign addr[43860] = 1742506504;
assign addr[43861] = 1753613897;
assign addr[43862] = 1764582240;
assign addr[43863] = 1775410662;
assign addr[43864] = 1786098304;
assign addr[43865] = 1796644320;
assign addr[43866] = 1807047873;
assign addr[43867] = 1817308138;
assign addr[43868] = 1827424302;
assign addr[43869] = 1837395562;
assign addr[43870] = 1847221128;
assign addr[43871] = 1856900221;
assign addr[43872] = 1866432072;
assign addr[43873] = 1875815927;
assign addr[43874] = 1885051042;
assign addr[43875] = 1894136683;
assign addr[43876] = 1903072131;
assign addr[43877] = 1911856677;
assign addr[43878] = 1920489624;
assign addr[43879] = 1928970288;
assign addr[43880] = 1937297997;
assign addr[43881] = 1945472089;
assign addr[43882] = 1953491918;
assign addr[43883] = 1961356847;
assign addr[43884] = 1969066252;
assign addr[43885] = 1976619522;
assign addr[43886] = 1984016058;
assign addr[43887] = 1991255274;
assign addr[43888] = 1998336596;
assign addr[43889] = 2005259462;
assign addr[43890] = 2012023322;
assign addr[43891] = 2018627642;
assign addr[43892] = 2025071897;
assign addr[43893] = 2031355576;
assign addr[43894] = 2037478181;
assign addr[43895] = 2043439226;
assign addr[43896] = 2049238240;
assign addr[43897] = 2054874761;
assign addr[43898] = 2060348343;
assign addr[43899] = 2065658552;
assign addr[43900] = 2070804967;
assign addr[43901] = 2075787180;
assign addr[43902] = 2080604795;
assign addr[43903] = 2085257431;
assign addr[43904] = 2089744719;
assign addr[43905] = 2094066304;
assign addr[43906] = 2098221841;
assign addr[43907] = 2102211002;
assign addr[43908] = 2106033471;
assign addr[43909] = 2109688944;
assign addr[43910] = 2113177132;
assign addr[43911] = 2116497758;
assign addr[43912] = 2119650558;
assign addr[43913] = 2122635283;
assign addr[43914] = 2125451696;
assign addr[43915] = 2128099574;
assign addr[43916] = 2130578706;
assign addr[43917] = 2132888897;
assign addr[43918] = 2135029962;
assign addr[43919] = 2137001733;
assign addr[43920] = 2138804053;
assign addr[43921] = 2140436778;
assign addr[43922] = 2141899780;
assign addr[43923] = 2143192942;
assign addr[43924] = 2144316162;
assign addr[43925] = 2145269351;
assign addr[43926] = 2146052433;
assign addr[43927] = 2146665347;
assign addr[43928] = 2147108043;
assign addr[43929] = 2147380486;
assign addr[43930] = 2147482655;
assign addr[43931] = 2147414542;
assign addr[43932] = 2147176152;
assign addr[43933] = 2146767505;
assign addr[43934] = 2146188631;
assign addr[43935] = 2145439578;
assign addr[43936] = 2144520405;
assign addr[43937] = 2143431184;
assign addr[43938] = 2142172003;
assign addr[43939] = 2140742960;
assign addr[43940] = 2139144169;
assign addr[43941] = 2137375758;
assign addr[43942] = 2135437865;
assign addr[43943] = 2133330646;
assign addr[43944] = 2131054266;
assign addr[43945] = 2128608907;
assign addr[43946] = 2125994762;
assign addr[43947] = 2123212038;
assign addr[43948] = 2120260957;
assign addr[43949] = 2117141752;
assign addr[43950] = 2113854671;
assign addr[43951] = 2110399974;
assign addr[43952] = 2106777935;
assign addr[43953] = 2102988841;
assign addr[43954] = 2099032994;
assign addr[43955] = 2094910706;
assign addr[43956] = 2090622304;
assign addr[43957] = 2086168128;
assign addr[43958] = 2081548533;
assign addr[43959] = 2076763883;
assign addr[43960] = 2071814558;
assign addr[43961] = 2066700952;
assign addr[43962] = 2061423468;
assign addr[43963] = 2055982526;
assign addr[43964] = 2050378558;
assign addr[43965] = 2044612007;
assign addr[43966] = 2038683330;
assign addr[43967] = 2032592999;
assign addr[43968] = 2026341495;
assign addr[43969] = 2019929315;
assign addr[43970] = 2013356967;
assign addr[43971] = 2006624971;
assign addr[43972] = 1999733863;
assign addr[43973] = 1992684188;
assign addr[43974] = 1985476506;
assign addr[43975] = 1978111387;
assign addr[43976] = 1970589416;
assign addr[43977] = 1962911189;
assign addr[43978] = 1955077316;
assign addr[43979] = 1947088417;
assign addr[43980] = 1938945125;
assign addr[43981] = 1930648088;
assign addr[43982] = 1922197961;
assign addr[43983] = 1913595416;
assign addr[43984] = 1904841135;
assign addr[43985] = 1895935811;
assign addr[43986] = 1886880151;
assign addr[43987] = 1877674873;
assign addr[43988] = 1868320707;
assign addr[43989] = 1858818395;
assign addr[43990] = 1849168689;
assign addr[43991] = 1839372356;
assign addr[43992] = 1829430172;
assign addr[43993] = 1819342925;
assign addr[43994] = 1809111415;
assign addr[43995] = 1798736454;
assign addr[43996] = 1788218865;
assign addr[43997] = 1777559480;
assign addr[43998] = 1766759146;
assign addr[43999] = 1755818718;
assign addr[44000] = 1744739065;
assign addr[44001] = 1733521064;
assign addr[44002] = 1722165606;
assign addr[44003] = 1710673591;
assign addr[44004] = 1699045930;
assign addr[44005] = 1687283545;
assign addr[44006] = 1675387369;
assign addr[44007] = 1663358344;
assign addr[44008] = 1651197426;
assign addr[44009] = 1638905577;
assign addr[44010] = 1626483774;
assign addr[44011] = 1613933000;
assign addr[44012] = 1601254251;
assign addr[44013] = 1588448533;
assign addr[44014] = 1575516860;
assign addr[44015] = 1562460258;
assign addr[44016] = 1549279763;
assign addr[44017] = 1535976419;
assign addr[44018] = 1522551282;
assign addr[44019] = 1509005416;
assign addr[44020] = 1495339895;
assign addr[44021] = 1481555802;
assign addr[44022] = 1467654232;
assign addr[44023] = 1453636285;
assign addr[44024] = 1439503074;
assign addr[44025] = 1425255719;
assign addr[44026] = 1410895350;
assign addr[44027] = 1396423105;
assign addr[44028] = 1381840133;
assign addr[44029] = 1367147589;
assign addr[44030] = 1352346639;
assign addr[44031] = 1337438456;
assign addr[44032] = 1322424222;
assign addr[44033] = 1307305128;
assign addr[44034] = 1292082373;
assign addr[44035] = 1276757164;
assign addr[44036] = 1261330715;
assign addr[44037] = 1245804251;
assign addr[44038] = 1230179002;
assign addr[44039] = 1214456207;
assign addr[44040] = 1198637114;
assign addr[44041] = 1182722976;
assign addr[44042] = 1166715055;
assign addr[44043] = 1150614620;
assign addr[44044] = 1134422949;
assign addr[44045] = 1118141326;
assign addr[44046] = 1101771040;
assign addr[44047] = 1085313391;
assign addr[44048] = 1068769683;
assign addr[44049] = 1052141228;
assign addr[44050] = 1035429345;
assign addr[44051] = 1018635358;
assign addr[44052] = 1001760600;
assign addr[44053] = 984806408;
assign addr[44054] = 967774128;
assign addr[44055] = 950665109;
assign addr[44056] = 933480707;
assign addr[44057] = 916222287;
assign addr[44058] = 898891215;
assign addr[44059] = 881488868;
assign addr[44060] = 864016623;
assign addr[44061] = 846475867;
assign addr[44062] = 828867991;
assign addr[44063] = 811194391;
assign addr[44064] = 793456467;
assign addr[44065] = 775655628;
assign addr[44066] = 757793284;
assign addr[44067] = 739870851;
assign addr[44068] = 721889752;
assign addr[44069] = 703851410;
assign addr[44070] = 685757258;
assign addr[44071] = 667608730;
assign addr[44072] = 649407264;
assign addr[44073] = 631154304;
assign addr[44074] = 612851297;
assign addr[44075] = 594499695;
assign addr[44076] = 576100953;
assign addr[44077] = 557656529;
assign addr[44078] = 539167887;
assign addr[44079] = 520636492;
assign addr[44080] = 502063814;
assign addr[44081] = 483451325;
assign addr[44082] = 464800501;
assign addr[44083] = 446112822;
assign addr[44084] = 427389768;
assign addr[44085] = 408632825;
assign addr[44086] = 389843480;
assign addr[44087] = 371023223;
assign addr[44088] = 352173546;
assign addr[44089] = 333295944;
assign addr[44090] = 314391913;
assign addr[44091] = 295462954;
assign addr[44092] = 276510565;
assign addr[44093] = 257536251;
assign addr[44094] = 238541516;
assign addr[44095] = 219527866;
assign addr[44096] = 200496809;
assign addr[44097] = 181449854;
assign addr[44098] = 162388511;
assign addr[44099] = 143314291;
assign addr[44100] = 124228708;
assign addr[44101] = 105133274;
assign addr[44102] = 86029503;
assign addr[44103] = 66918911;
assign addr[44104] = 47803013;
assign addr[44105] = 28683324;
assign addr[44106] = 9561361;
assign addr[44107] = -9561361;
assign addr[44108] = -28683324;
assign addr[44109] = -47803013;
assign addr[44110] = -66918911;
assign addr[44111] = -86029503;
assign addr[44112] = -105133274;
assign addr[44113] = -124228708;
assign addr[44114] = -143314291;
assign addr[44115] = -162388511;
assign addr[44116] = -181449854;
assign addr[44117] = -200496809;
assign addr[44118] = -219527866;
assign addr[44119] = -238541516;
assign addr[44120] = -257536251;
assign addr[44121] = -276510565;
assign addr[44122] = -295462953;
assign addr[44123] = -314391913;
assign addr[44124] = -333295944;
assign addr[44125] = -352173546;
assign addr[44126] = -371023223;
assign addr[44127] = -389843480;
assign addr[44128] = -408632825;
assign addr[44129] = -427389768;
assign addr[44130] = -446112822;
assign addr[44131] = -464800501;
assign addr[44132] = -483451325;
assign addr[44133] = -502063814;
assign addr[44134] = -520636492;
assign addr[44135] = -539167887;
assign addr[44136] = -557656529;
assign addr[44137] = -576100953;
assign addr[44138] = -594499695;
assign addr[44139] = -612851297;
assign addr[44140] = -631154304;
assign addr[44141] = -649407264;
assign addr[44142] = -667608730;
assign addr[44143] = -685757258;
assign addr[44144] = -703851410;
assign addr[44145] = -721889752;
assign addr[44146] = -739870851;
assign addr[44147] = -757793284;
assign addr[44148] = -775655628;
assign addr[44149] = -793456467;
assign addr[44150] = -811194391;
assign addr[44151] = -828867991;
assign addr[44152] = -846475867;
assign addr[44153] = -864016623;
assign addr[44154] = -881488868;
assign addr[44155] = -898891215;
assign addr[44156] = -916222287;
assign addr[44157] = -933480707;
assign addr[44158] = -950665109;
assign addr[44159] = -967774128;
assign addr[44160] = -984806408;
assign addr[44161] = -1001760600;
assign addr[44162] = -1018635358;
assign addr[44163] = -1035429345;
assign addr[44164] = -1052141228;
assign addr[44165] = -1068769683;
assign addr[44166] = -1085313391;
assign addr[44167] = -1101771040;
assign addr[44168] = -1118141326;
assign addr[44169] = -1134422949;
assign addr[44170] = -1150614620;
assign addr[44171] = -1166715055;
assign addr[44172] = -1182722976;
assign addr[44173] = -1198637114;
assign addr[44174] = -1214456207;
assign addr[44175] = -1230179002;
assign addr[44176] = -1245804251;
assign addr[44177] = -1261330715;
assign addr[44178] = -1276757164;
assign addr[44179] = -1292082373;
assign addr[44180] = -1307305128;
assign addr[44181] = -1322424222;
assign addr[44182] = -1337438456;
assign addr[44183] = -1352346639;
assign addr[44184] = -1367147589;
assign addr[44185] = -1381840133;
assign addr[44186] = -1396423105;
assign addr[44187] = -1410895350;
assign addr[44188] = -1425255719;
assign addr[44189] = -1439503074;
assign addr[44190] = -1453636285;
assign addr[44191] = -1467654232;
assign addr[44192] = -1481555802;
assign addr[44193] = -1495339895;
assign addr[44194] = -1509005416;
assign addr[44195] = -1522551282;
assign addr[44196] = -1535976419;
assign addr[44197] = -1549279763;
assign addr[44198] = -1562460258;
assign addr[44199] = -1575516860;
assign addr[44200] = -1588448533;
assign addr[44201] = -1601254251;
assign addr[44202] = -1613933000;
assign addr[44203] = -1626483774;
assign addr[44204] = -1638905577;
assign addr[44205] = -1651197426;
assign addr[44206] = -1663358344;
assign addr[44207] = -1675387369;
assign addr[44208] = -1687283545;
assign addr[44209] = -1699045930;
assign addr[44210] = -1710673591;
assign addr[44211] = -1722165606;
assign addr[44212] = -1733521064;
assign addr[44213] = -1744739065;
assign addr[44214] = -1755818718;
assign addr[44215] = -1766759146;
assign addr[44216] = -1777559480;
assign addr[44217] = -1788218865;
assign addr[44218] = -1798736454;
assign addr[44219] = -1809111415;
assign addr[44220] = -1819342925;
assign addr[44221] = -1829430172;
assign addr[44222] = -1839372356;
assign addr[44223] = -1849168689;
assign addr[44224] = -1858818395;
assign addr[44225] = -1868320707;
assign addr[44226] = -1877674873;
assign addr[44227] = -1886880151;
assign addr[44228] = -1895935811;
assign addr[44229] = -1904841135;
assign addr[44230] = -1913595416;
assign addr[44231] = -1922197961;
assign addr[44232] = -1930648088;
assign addr[44233] = -1938945125;
assign addr[44234] = -1947088417;
assign addr[44235] = -1955077316;
assign addr[44236] = -1962911189;
assign addr[44237] = -1970589416;
assign addr[44238] = -1978111387;
assign addr[44239] = -1985476506;
assign addr[44240] = -1992684188;
assign addr[44241] = -1999733863;
assign addr[44242] = -2006624971;
assign addr[44243] = -2013356967;
assign addr[44244] = -2019929315;
assign addr[44245] = -2026341495;
assign addr[44246] = -2032592999;
assign addr[44247] = -2038683330;
assign addr[44248] = -2044612007;
assign addr[44249] = -2050378558;
assign addr[44250] = -2055982526;
assign addr[44251] = -2061423468;
assign addr[44252] = -2066700952;
assign addr[44253] = -2071814558;
assign addr[44254] = -2076763883;
assign addr[44255] = -2081548533;
assign addr[44256] = -2086168128;
assign addr[44257] = -2090622304;
assign addr[44258] = -2094910706;
assign addr[44259] = -2099032994;
assign addr[44260] = -2102988841;
assign addr[44261] = -2106777935;
assign addr[44262] = -2110399974;
assign addr[44263] = -2113854671;
assign addr[44264] = -2117141752;
assign addr[44265] = -2120260957;
assign addr[44266] = -2123212038;
assign addr[44267] = -2125994762;
assign addr[44268] = -2128608907;
assign addr[44269] = -2131054266;
assign addr[44270] = -2133330646;
assign addr[44271] = -2135437865;
assign addr[44272] = -2137375758;
assign addr[44273] = -2139144169;
assign addr[44274] = -2140742960;
assign addr[44275] = -2142172003;
assign addr[44276] = -2143431184;
assign addr[44277] = -2144520405;
assign addr[44278] = -2145439578;
assign addr[44279] = -2146188631;
assign addr[44280] = -2146767505;
assign addr[44281] = -2147176152;
assign addr[44282] = -2147414542;
assign addr[44283] = -2147482655;
assign addr[44284] = -2147380486;
assign addr[44285] = -2147108043;
assign addr[44286] = -2146665347;
assign addr[44287] = -2146052433;
assign addr[44288] = -2145269351;
assign addr[44289] = -2144316162;
assign addr[44290] = -2143192942;
assign addr[44291] = -2141899780;
assign addr[44292] = -2140436778;
assign addr[44293] = -2138804053;
assign addr[44294] = -2137001733;
assign addr[44295] = -2135029962;
assign addr[44296] = -2132888897;
assign addr[44297] = -2130578706;
assign addr[44298] = -2128099574;
assign addr[44299] = -2125451696;
assign addr[44300] = -2122635283;
assign addr[44301] = -2119650558;
assign addr[44302] = -2116497758;
assign addr[44303] = -2113177132;
assign addr[44304] = -2109688944;
assign addr[44305] = -2106033471;
assign addr[44306] = -2102211002;
assign addr[44307] = -2098221841;
assign addr[44308] = -2094066304;
assign addr[44309] = -2089744719;
assign addr[44310] = -2085257431;
assign addr[44311] = -2080604795;
assign addr[44312] = -2075787180;
assign addr[44313] = -2070804967;
assign addr[44314] = -2065658552;
assign addr[44315] = -2060348343;
assign addr[44316] = -2054874761;
assign addr[44317] = -2049238240;
assign addr[44318] = -2043439226;
assign addr[44319] = -2037478181;
assign addr[44320] = -2031355576;
assign addr[44321] = -2025071897;
assign addr[44322] = -2018627642;
assign addr[44323] = -2012023322;
assign addr[44324] = -2005259462;
assign addr[44325] = -1998336596;
assign addr[44326] = -1991255274;
assign addr[44327] = -1984016058;
assign addr[44328] = -1976619522;
assign addr[44329] = -1969066252;
assign addr[44330] = -1961356847;
assign addr[44331] = -1953491918;
assign addr[44332] = -1945472089;
assign addr[44333] = -1937297997;
assign addr[44334] = -1928970288;
assign addr[44335] = -1920489624;
assign addr[44336] = -1911856677;
assign addr[44337] = -1903072131;
assign addr[44338] = -1894136683;
assign addr[44339] = -1885051042;
assign addr[44340] = -1875815927;
assign addr[44341] = -1866432072;
assign addr[44342] = -1856900221;
assign addr[44343] = -1847221128;
assign addr[44344] = -1837395562;
assign addr[44345] = -1827424302;
assign addr[44346] = -1817308138;
assign addr[44347] = -1807047873;
assign addr[44348] = -1796644320;
assign addr[44349] = -1786098304;
assign addr[44350] = -1775410662;
assign addr[44351] = -1764582240;
assign addr[44352] = -1753613897;
assign addr[44353] = -1742506504;
assign addr[44354] = -1731260941;
assign addr[44355] = -1719878099;
assign addr[44356] = -1708358881;
assign addr[44357] = -1696704201;
assign addr[44358] = -1684914983;
assign addr[44359] = -1672992161;
assign addr[44360] = -1660936681;
assign addr[44361] = -1648749499;
assign addr[44362] = -1636431582;
assign addr[44363] = -1623983905;
assign addr[44364] = -1611407456;
assign addr[44365] = -1598703233;
assign addr[44366] = -1585872242;
assign addr[44367] = -1572915501;
assign addr[44368] = -1559834037;
assign addr[44369] = -1546628888;
assign addr[44370] = -1533301101;
assign addr[44371] = -1519851733;
assign addr[44372] = -1506281850;
assign addr[44373] = -1492592527;
assign addr[44374] = -1478784851;
assign addr[44375] = -1464859917;
assign addr[44376] = -1450818828;
assign addr[44377] = -1436662698;
assign addr[44378] = -1422392650;
assign addr[44379] = -1408009814;
assign addr[44380] = -1393515332;
assign addr[44381] = -1378910353;
assign addr[44382] = -1364196034;
assign addr[44383] = -1349373543;
assign addr[44384] = -1334444055;
assign addr[44385] = -1319408754;
assign addr[44386] = -1304268832;
assign addr[44387] = -1289025489;
assign addr[44388] = -1273679934;
assign addr[44389] = -1258233384;
assign addr[44390] = -1242687064;
assign addr[44391] = -1227042207;
assign addr[44392] = -1211300053;
assign addr[44393] = -1195461849;
assign addr[44394] = -1179528853;
assign addr[44395] = -1163502328;
assign addr[44396] = -1147383544;
assign addr[44397] = -1131173780;
assign addr[44398] = -1114874320;
assign addr[44399] = -1098486458;
assign addr[44400] = -1082011492;
assign addr[44401] = -1065450729;
assign addr[44402] = -1048805483;
assign addr[44403] = -1032077073;
assign addr[44404] = -1015266825;
assign addr[44405] = -998376073;
assign addr[44406] = -981406156;
assign addr[44407] = -964358420;
assign addr[44408] = -947234215;
assign addr[44409] = -930034901;
assign addr[44410] = -912761841;
assign addr[44411] = -895416404;
assign addr[44412] = -877999966;
assign addr[44413] = -860513908;
assign addr[44414] = -842959617;
assign addr[44415] = -825338484;
assign addr[44416] = -807651907;
assign addr[44417] = -789901288;
assign addr[44418] = -772088034;
assign addr[44419] = -754213559;
assign addr[44420] = -736279279;
assign addr[44421] = -718286617;
assign addr[44422] = -700236999;
assign addr[44423] = -682131857;
assign addr[44424] = -663972625;
assign addr[44425] = -645760745;
assign addr[44426] = -627497660;
assign addr[44427] = -609184818;
assign addr[44428] = -590823671;
assign addr[44429] = -572415676;
assign addr[44430] = -553962291;
assign addr[44431] = -535464981;
assign addr[44432] = -516925212;
assign addr[44433] = -498344454;
assign addr[44434] = -479724180;
assign addr[44435] = -461065866;
assign addr[44436] = -442370993;
assign addr[44437] = -423641043;
assign addr[44438] = -404877501;
assign addr[44439] = -386081854;
assign addr[44440] = -367255594;
assign addr[44441] = -348400212;
assign addr[44442] = -329517204;
assign addr[44443] = -310608068;
assign addr[44444] = -291674302;
assign addr[44445] = -272717408;
assign addr[44446] = -253738890;
assign addr[44447] = -234740251;
assign addr[44448] = -215722999;
assign addr[44449] = -196688642;
assign addr[44450] = -177638688;
assign addr[44451] = -158574649;
assign addr[44452] = -139498035;
assign addr[44453] = -120410361;
assign addr[44454] = -101313138;
assign addr[44455] = -82207882;
assign addr[44456] = -63096108;
assign addr[44457] = -43979330;
assign addr[44458] = -24859065;
assign addr[44459] = -5736829;
assign addr[44460] = 13385863;
assign addr[44461] = 32507492;
assign addr[44462] = 51626544;
assign addr[44463] = 70741503;
assign addr[44464] = 89850852;
assign addr[44465] = 108953076;
assign addr[44466] = 128046661;
assign addr[44467] = 147130093;
assign addr[44468] = 166201858;
assign addr[44469] = 185260444;
assign addr[44470] = 204304341;
assign addr[44471] = 223332037;
assign addr[44472] = 242342025;
assign addr[44473] = 261332796;
assign addr[44474] = 280302845;
assign addr[44475] = 299250668;
assign addr[44476] = 318174762;
assign addr[44477] = 337073627;
assign addr[44478] = 355945764;
assign addr[44479] = 374789676;
assign addr[44480] = 393603870;
assign addr[44481] = 412386854;
assign addr[44482] = 431137138;
assign addr[44483] = 449853235;
assign addr[44484] = 468533662;
assign addr[44485] = 487176937;
assign addr[44486] = 505781581;
assign addr[44487] = 524346121;
assign addr[44488] = 542869083;
assign addr[44489] = 561348998;
assign addr[44490] = 579784402;
assign addr[44491] = 598173833;
assign addr[44492] = 616515832;
assign addr[44493] = 634808946;
assign addr[44494] = 653051723;
assign addr[44495] = 671242716;
assign addr[44496] = 689380485;
assign addr[44497] = 707463589;
assign addr[44498] = 725490597;
assign addr[44499] = 743460077;
assign addr[44500] = 761370605;
assign addr[44501] = 779220762;
assign addr[44502] = 797009130;
assign addr[44503] = 814734301;
assign addr[44504] = 832394869;
assign addr[44505] = 849989433;
assign addr[44506] = 867516597;
assign addr[44507] = 884974973;
assign addr[44508] = 902363176;
assign addr[44509] = 919679827;
assign addr[44510] = 936923553;
assign addr[44511] = 954092986;
assign addr[44512] = 971186766;
assign addr[44513] = 988203537;
assign addr[44514] = 1005141949;
assign addr[44515] = 1022000660;
assign addr[44516] = 1038778332;
assign addr[44517] = 1055473635;
assign addr[44518] = 1072085246;
assign addr[44519] = 1088611847;
assign addr[44520] = 1105052128;
assign addr[44521] = 1121404785;
assign addr[44522] = 1137668521;
assign addr[44523] = 1153842047;
assign addr[44524] = 1169924081;
assign addr[44525] = 1185913346;
assign addr[44526] = 1201808576;
assign addr[44527] = 1217608510;
assign addr[44528] = 1233311895;
assign addr[44529] = 1248917486;
assign addr[44530] = 1264424045;
assign addr[44531] = 1279830344;
assign addr[44532] = 1295135159;
assign addr[44533] = 1310337279;
assign addr[44534] = 1325435496;
assign addr[44535] = 1340428615;
assign addr[44536] = 1355315445;
assign addr[44537] = 1370094808;
assign addr[44538] = 1384765530;
assign addr[44539] = 1399326449;
assign addr[44540] = 1413776410;
assign addr[44541] = 1428114267;
assign addr[44542] = 1442338884;
assign addr[44543] = 1456449131;
assign addr[44544] = 1470443891;
assign addr[44545] = 1484322054;
assign addr[44546] = 1498082520;
assign addr[44547] = 1511724196;
assign addr[44548] = 1525246002;
assign addr[44549] = 1538646865;
assign addr[44550] = 1551925723;
assign addr[44551] = 1565081523;
assign addr[44552] = 1578113222;
assign addr[44553] = 1591019785;
assign addr[44554] = 1603800191;
assign addr[44555] = 1616453425;
assign addr[44556] = 1628978484;
assign addr[44557] = 1641374375;
assign addr[44558] = 1653640115;
assign addr[44559] = 1665774731;
assign addr[44560] = 1677777262;
assign addr[44561] = 1689646755;
assign addr[44562] = 1701382270;
assign addr[44563] = 1712982875;
assign addr[44564] = 1724447652;
assign addr[44565] = 1735775690;
assign addr[44566] = 1746966091;
assign addr[44567] = 1758017969;
assign addr[44568] = 1768930447;
assign addr[44569] = 1779702660;
assign addr[44570] = 1790333753;
assign addr[44571] = 1800822883;
assign addr[44572] = 1811169220;
assign addr[44573] = 1821371941;
assign addr[44574] = 1831430239;
assign addr[44575] = 1841343316;
assign addr[44576] = 1851110385;
assign addr[44577] = 1860730673;
assign addr[44578] = 1870203416;
assign addr[44579] = 1879527863;
assign addr[44580] = 1888703276;
assign addr[44581] = 1897728925;
assign addr[44582] = 1906604097;
assign addr[44583] = 1915328086;
assign addr[44584] = 1923900201;
assign addr[44585] = 1932319763;
assign addr[44586] = 1940586104;
assign addr[44587] = 1948698568;
assign addr[44588] = 1956656513;
assign addr[44589] = 1964459306;
assign addr[44590] = 1972106330;
assign addr[44591] = 1979596978;
assign addr[44592] = 1986930656;
assign addr[44593] = 1994106782;
assign addr[44594] = 2001124788;
assign addr[44595] = 2007984117;
assign addr[44596] = 2014684225;
assign addr[44597] = 2021224581;
assign addr[44598] = 2027604666;
assign addr[44599] = 2033823974;
assign addr[44600] = 2039882013;
assign addr[44601] = 2045778302;
assign addr[44602] = 2051512372;
assign addr[44603] = 2057083771;
assign addr[44604] = 2062492055;
assign addr[44605] = 2067736796;
assign addr[44606] = 2072817579;
assign addr[44607] = 2077733999;
assign addr[44608] = 2082485668;
assign addr[44609] = 2087072209;
assign addr[44610] = 2091493257;
assign addr[44611] = 2095748463;
assign addr[44612] = 2099837489;
assign addr[44613] = 2103760010;
assign addr[44614] = 2107515716;
assign addr[44615] = 2111104309;
assign addr[44616] = 2114525505;
assign addr[44617] = 2117779031;
assign addr[44618] = 2120864631;
assign addr[44619] = 2123782059;
assign addr[44620] = 2126531084;
assign addr[44621] = 2129111488;
assign addr[44622] = 2131523066;
assign addr[44623] = 2133765628;
assign addr[44624] = 2135838995;
assign addr[44625] = 2137743003;
assign addr[44626] = 2139477502;
assign addr[44627] = 2141042352;
assign addr[44628] = 2142437431;
assign addr[44629] = 2143662628;
assign addr[44630] = 2144717846;
assign addr[44631] = 2145603001;
assign addr[44632] = 2146318022;
assign addr[44633] = 2146862854;
assign addr[44634] = 2147237452;
assign addr[44635] = 2147441787;
assign addr[44636] = 2147475844;
assign addr[44637] = 2147339619;
assign addr[44638] = 2147033123;
assign addr[44639] = 2146556380;
assign addr[44640] = 2145909429;
assign addr[44641] = 2145092320;
assign addr[44642] = 2144105118;
assign addr[44643] = 2142947902;
assign addr[44644] = 2141620763;
assign addr[44645] = 2140123807;
assign addr[44646] = 2138457152;
assign addr[44647] = 2136620930;
assign addr[44648] = 2134615288;
assign addr[44649] = 2132440383;
assign addr[44650] = 2130096389;
assign addr[44651] = 2127583492;
assign addr[44652] = 2124901890;
assign addr[44653] = 2122051796;
assign addr[44654] = 2119033436;
assign addr[44655] = 2115847050;
assign addr[44656] = 2112492891;
assign addr[44657] = 2108971223;
assign addr[44658] = 2105282327;
assign addr[44659] = 2101426496;
assign addr[44660] = 2097404033;
assign addr[44661] = 2093215260;
assign addr[44662] = 2088860507;
assign addr[44663] = 2084340120;
assign addr[44664] = 2079654458;
assign addr[44665] = 2074803892;
assign addr[44666] = 2069788807;
assign addr[44667] = 2064609600;
assign addr[44668] = 2059266683;
assign addr[44669] = 2053760478;
assign addr[44670] = 2048091422;
assign addr[44671] = 2042259965;
assign addr[44672] = 2036266570;
assign addr[44673] = 2030111710;
assign addr[44674] = 2023795876;
assign addr[44675] = 2017319567;
assign addr[44676] = 2010683297;
assign addr[44677] = 2003887591;
assign addr[44678] = 1996932990;
assign addr[44679] = 1989820044;
assign addr[44680] = 1982549318;
assign addr[44681] = 1975121388;
assign addr[44682] = 1967536842;
assign addr[44683] = 1959796283;
assign addr[44684] = 1951900324;
assign addr[44685] = 1943849591;
assign addr[44686] = 1935644723;
assign addr[44687] = 1927286370;
assign addr[44688] = 1918775195;
assign addr[44689] = 1910111873;
assign addr[44690] = 1901297091;
assign addr[44691] = 1892331547;
assign addr[44692] = 1883215953;
assign addr[44693] = 1873951032;
assign addr[44694] = 1864537518;
assign addr[44695] = 1854976157;
assign addr[44696] = 1845267708;
assign addr[44697] = 1835412941;
assign addr[44698] = 1825412636;
assign addr[44699] = 1815267588;
assign addr[44700] = 1804978599;
assign addr[44701] = 1794546487;
assign addr[44702] = 1783972079;
assign addr[44703] = 1773256212;
assign addr[44704] = 1762399737;
assign addr[44705] = 1751403515;
assign addr[44706] = 1740268417;
assign addr[44707] = 1728995326;
assign addr[44708] = 1717585136;
assign addr[44709] = 1706038753;
assign addr[44710] = 1694357091;
assign addr[44711] = 1682541077;
assign addr[44712] = 1670591647;
assign addr[44713] = 1658509750;
assign addr[44714] = 1646296344;
assign addr[44715] = 1633952396;
assign addr[44716] = 1621478885;
assign addr[44717] = 1608876801;
assign addr[44718] = 1596147143;
assign addr[44719] = 1583290921;
assign addr[44720] = 1570309153;
assign addr[44721] = 1557202869;
assign addr[44722] = 1543973108;
assign addr[44723] = 1530620920;
assign addr[44724] = 1517147363;
assign addr[44725] = 1503553506;
assign addr[44726] = 1489840425;
assign addr[44727] = 1476009210;
assign addr[44728] = 1462060956;
assign addr[44729] = 1447996770;
assign addr[44730] = 1433817766;
assign addr[44731] = 1419525069;
assign addr[44732] = 1405119813;
assign addr[44733] = 1390603139;
assign addr[44734] = 1375976199;
assign addr[44735] = 1361240152;
assign addr[44736] = 1346396168;
assign addr[44737] = 1331445422;
assign addr[44738] = 1316389101;
assign addr[44739] = 1301228398;
assign addr[44740] = 1285964516;
assign addr[44741] = 1270598665;
assign addr[44742] = 1255132063;
assign addr[44743] = 1239565936;
assign addr[44744] = 1223901520;
assign addr[44745] = 1208140056;
assign addr[44746] = 1192282793;
assign addr[44747] = 1176330990;
assign addr[44748] = 1160285911;
assign addr[44749] = 1144148829;
assign addr[44750] = 1127921022;
assign addr[44751] = 1111603778;
assign addr[44752] = 1095198391;
assign addr[44753] = 1078706161;
assign addr[44754] = 1062128397;
assign addr[44755] = 1045466412;
assign addr[44756] = 1028721528;
assign addr[44757] = 1011895073;
assign addr[44758] = 994988380;
assign addr[44759] = 978002791;
assign addr[44760] = 960939653;
assign addr[44761] = 943800318;
assign addr[44762] = 926586145;
assign addr[44763] = 909298500;
assign addr[44764] = 891938752;
assign addr[44765] = 874508280;
assign addr[44766] = 857008464;
assign addr[44767] = 839440693;
assign addr[44768] = 821806359;
assign addr[44769] = 804106861;
assign addr[44770] = 786343603;
assign addr[44771] = 768517992;
assign addr[44772] = 750631442;
assign addr[44773] = 732685372;
assign addr[44774] = 714681204;
assign addr[44775] = 696620367;
assign addr[44776] = 678504291;
assign addr[44777] = 660334415;
assign addr[44778] = 642112178;
assign addr[44779] = 623839025;
assign addr[44780] = 605516406;
assign addr[44781] = 587145773;
assign addr[44782] = 568728583;
assign addr[44783] = 550266296;
assign addr[44784] = 531760377;
assign addr[44785] = 513212292;
assign addr[44786] = 494623513;
assign addr[44787] = 475995513;
assign addr[44788] = 457329769;
assign addr[44789] = 438627762;
assign addr[44790] = 419890975;
assign addr[44791] = 401120892;
assign addr[44792] = 382319004;
assign addr[44793] = 363486799;
assign addr[44794] = 344625773;
assign addr[44795] = 325737419;
assign addr[44796] = 306823237;
assign addr[44797] = 287884725;
assign addr[44798] = 268923386;
assign addr[44799] = 249940723;
assign addr[44800] = 230938242;
assign addr[44801] = 211917448;
assign addr[44802] = 192879850;
assign addr[44803] = 173826959;
assign addr[44804] = 154760284;
assign addr[44805] = 135681337;
assign addr[44806] = 116591632;
assign addr[44807] = 97492681;
assign addr[44808] = 78386000;
assign addr[44809] = 59273104;
assign addr[44810] = 40155507;
assign addr[44811] = 21034727;
assign addr[44812] = 1912278;
assign addr[44813] = -17210322;
assign addr[44814] = -36331557;
assign addr[44815] = -55449912;
assign addr[44816] = -74563870;
assign addr[44817] = -93671915;
assign addr[44818] = -112772533;
assign addr[44819] = -131864208;
assign addr[44820] = -150945428;
assign addr[44821] = -170014678;
assign addr[44822] = -189070447;
assign addr[44823] = -208111224;
assign addr[44824] = -227135500;
assign addr[44825] = -246141764;
assign addr[44826] = -265128512;
assign addr[44827] = -284094236;
assign addr[44828] = -303037433;
assign addr[44829] = -321956601;
assign addr[44830] = -340850240;
assign addr[44831] = -359716852;
assign addr[44832] = -378554940;
assign addr[44833] = -397363011;
assign addr[44834] = -416139574;
assign addr[44835] = -434883140;
assign addr[44836] = -453592221;
assign addr[44837] = -472265336;
assign addr[44838] = -490901003;
assign addr[44839] = -509497745;
assign addr[44840] = -528054086;
assign addr[44841] = -546568556;
assign addr[44842] = -565039687;
assign addr[44843] = -583466013;
assign addr[44844] = -601846074;
assign addr[44845] = -620178412;
assign addr[44846] = -638461574;
assign addr[44847] = -656694110;
assign addr[44848] = -674874574;
assign addr[44849] = -693001525;
assign addr[44850] = -711073524;
assign addr[44851] = -729089140;
assign addr[44852] = -747046944;
assign addr[44853] = -764945512;
assign addr[44854] = -782783424;
assign addr[44855] = -800559266;
assign addr[44856] = -818271628;
assign addr[44857] = -835919107;
assign addr[44858] = -853500302;
assign addr[44859] = -871013820;
assign addr[44860] = -888458272;
assign addr[44861] = -905832274;
assign addr[44862] = -923134450;
assign addr[44863] = -940363427;
assign addr[44864] = -957517838;
assign addr[44865] = -974596324;
assign addr[44866] = -991597531;
assign addr[44867] = -1008520110;
assign addr[44868] = -1025362720;
assign addr[44869] = -1042124025;
assign addr[44870] = -1058802695;
assign addr[44871] = -1075397409;
assign addr[44872] = -1091906851;
assign addr[44873] = -1108329711;
assign addr[44874] = -1124664687;
assign addr[44875] = -1140910484;
assign addr[44876] = -1157065814;
assign addr[44877] = -1173129396;
assign addr[44878] = -1189099956;
assign addr[44879] = -1204976227;
assign addr[44880] = -1220756951;
assign addr[44881] = -1236440877;
assign addr[44882] = -1252026760;
assign addr[44883] = -1267513365;
assign addr[44884] = -1282899464;
assign addr[44885] = -1298183838;
assign addr[44886] = -1313365273;
assign addr[44887] = -1328442566;
assign addr[44888] = -1343414522;
assign addr[44889] = -1358279953;
assign addr[44890] = -1373037681;
assign addr[44891] = -1387686535;
assign addr[44892] = -1402225355;
assign addr[44893] = -1416652986;
assign addr[44894] = -1430968286;
assign addr[44895] = -1445170118;
assign addr[44896] = -1459257358;
assign addr[44897] = -1473228887;
assign addr[44898] = -1487083598;
assign addr[44899] = -1500820393;
assign addr[44900] = -1514438181;
assign addr[44901] = -1527935884;
assign addr[44902] = -1541312431;
assign addr[44903] = -1554566762;
assign addr[44904] = -1567697824;
assign addr[44905] = -1580704578;
assign addr[44906] = -1593585992;
assign addr[44907] = -1606341043;
assign addr[44908] = -1618968722;
assign addr[44909] = -1631468027;
assign addr[44910] = -1643837966;
assign addr[44911] = -1656077559;
assign addr[44912] = -1668185835;
assign addr[44913] = -1680161834;
assign addr[44914] = -1692004606;
assign addr[44915] = -1703713213;
assign addr[44916] = -1715286726;
assign addr[44917] = -1726724227;
assign addr[44918] = -1738024810;
assign addr[44919] = -1749187577;
assign addr[44920] = -1760211645;
assign addr[44921] = -1771096139;
assign addr[44922] = -1781840195;
assign addr[44923] = -1792442963;
assign addr[44924] = -1802903601;
assign addr[44925] = -1813221279;
assign addr[44926] = -1823395180;
assign addr[44927] = -1833424497;
assign addr[44928] = -1843308435;
assign addr[44929] = -1853046210;
assign addr[44930] = -1862637049;
assign addr[44931] = -1872080193;
assign addr[44932] = -1881374892;
assign addr[44933] = -1890520410;
assign addr[44934] = -1899516021;
assign addr[44935] = -1908361011;
assign addr[44936] = -1917054681;
assign addr[44937] = -1925596340;
assign addr[44938] = -1933985310;
assign addr[44939] = -1942220928;
assign addr[44940] = -1950302539;
assign addr[44941] = -1958229503;
assign addr[44942] = -1966001192;
assign addr[44943] = -1973616989;
assign addr[44944] = -1981076290;
assign addr[44945] = -1988378503;
assign addr[44946] = -1995523051;
assign addr[44947] = -2002509365;
assign addr[44948] = -2009336893;
assign addr[44949] = -2016005093;
assign addr[44950] = -2022513436;
assign addr[44951] = -2028861406;
assign addr[44952] = -2035048499;
assign addr[44953] = -2041074226;
assign addr[44954] = -2046938108;
assign addr[44955] = -2052639680;
assign addr[44956] = -2058178491;
assign addr[44957] = -2063554100;
assign addr[44958] = -2068766083;
assign addr[44959] = -2073814024;
assign addr[44960] = -2078697525;
assign addr[44961] = -2083416198;
assign addr[44962] = -2087969669;
assign addr[44963] = -2092357577;
assign addr[44964] = -2096579573;
assign addr[44965] = -2100635323;
assign addr[44966] = -2104524506;
assign addr[44967] = -2108246813;
assign addr[44968] = -2111801949;
assign addr[44969] = -2115189632;
assign addr[44970] = -2118409593;
assign addr[44971] = -2121461578;
assign addr[44972] = -2124345343;
assign addr[44973] = -2127060661;
assign addr[44974] = -2129607316;
assign addr[44975] = -2131985106;
assign addr[44976] = -2134193842;
assign addr[44977] = -2136233350;
assign addr[44978] = -2138103468;
assign addr[44979] = -2139804048;
assign addr[44980] = -2141334954;
assign addr[44981] = -2142696065;
assign addr[44982] = -2143887273;
assign addr[44983] = -2144908484;
assign addr[44984] = -2145759618;
assign addr[44985] = -2146440605;
assign addr[44986] = -2146951393;
assign addr[44987] = -2147291941;
assign addr[44988] = -2147462221;
assign addr[44989] = -2147462221;
assign addr[44990] = -2147291941;
assign addr[44991] = -2146951393;
assign addr[44992] = -2146440605;
assign addr[44993] = -2145759618;
assign addr[44994] = -2144908484;
assign addr[44995] = -2143887273;
assign addr[44996] = -2142696065;
assign addr[44997] = -2141334954;
assign addr[44998] = -2139804048;
assign addr[44999] = -2138103468;
assign addr[45000] = -2136233350;
assign addr[45001] = -2134193842;
assign addr[45002] = -2131985106;
assign addr[45003] = -2129607316;
assign addr[45004] = -2127060661;
assign addr[45005] = -2124345343;
assign addr[45006] = -2121461578;
assign addr[45007] = -2118409593;
assign addr[45008] = -2115189632;
assign addr[45009] = -2111801949;
assign addr[45010] = -2108246813;
assign addr[45011] = -2104524506;
assign addr[45012] = -2100635323;
assign addr[45013] = -2096579573;
assign addr[45014] = -2092357577;
assign addr[45015] = -2087969669;
assign addr[45016] = -2083416198;
assign addr[45017] = -2078697525;
assign addr[45018] = -2073814024;
assign addr[45019] = -2068766083;
assign addr[45020] = -2063554100;
assign addr[45021] = -2058178491;
assign addr[45022] = -2052639680;
assign addr[45023] = -2046938108;
assign addr[45024] = -2041074226;
assign addr[45025] = -2035048499;
assign addr[45026] = -2028861406;
assign addr[45027] = -2022513436;
assign addr[45028] = -2016005093;
assign addr[45029] = -2009336893;
assign addr[45030] = -2002509365;
assign addr[45031] = -1995523051;
assign addr[45032] = -1988378503;
assign addr[45033] = -1981076290;
assign addr[45034] = -1973616989;
assign addr[45035] = -1966001192;
assign addr[45036] = -1958229503;
assign addr[45037] = -1950302539;
assign addr[45038] = -1942220928;
assign addr[45039] = -1933985310;
assign addr[45040] = -1925596340;
assign addr[45041] = -1917054681;
assign addr[45042] = -1908361011;
assign addr[45043] = -1899516021;
assign addr[45044] = -1890520410;
assign addr[45045] = -1881374892;
assign addr[45046] = -1872080193;
assign addr[45047] = -1862637049;
assign addr[45048] = -1853046210;
assign addr[45049] = -1843308435;
assign addr[45050] = -1833424497;
assign addr[45051] = -1823395180;
assign addr[45052] = -1813221279;
assign addr[45053] = -1802903601;
assign addr[45054] = -1792442963;
assign addr[45055] = -1781840195;
assign addr[45056] = -1771096139;
assign addr[45057] = -1760211645;
assign addr[45058] = -1749187577;
assign addr[45059] = -1738024810;
assign addr[45060] = -1726724227;
assign addr[45061] = -1715286726;
assign addr[45062] = -1703713213;
assign addr[45063] = -1692004606;
assign addr[45064] = -1680161834;
assign addr[45065] = -1668185835;
assign addr[45066] = -1656077559;
assign addr[45067] = -1643837966;
assign addr[45068] = -1631468027;
assign addr[45069] = -1618968722;
assign addr[45070] = -1606341043;
assign addr[45071] = -1593585992;
assign addr[45072] = -1580704578;
assign addr[45073] = -1567697824;
assign addr[45074] = -1554566762;
assign addr[45075] = -1541312431;
assign addr[45076] = -1527935884;
assign addr[45077] = -1514438181;
assign addr[45078] = -1500820393;
assign addr[45079] = -1487083598;
assign addr[45080] = -1473228887;
assign addr[45081] = -1459257358;
assign addr[45082] = -1445170118;
assign addr[45083] = -1430968286;
assign addr[45084] = -1416652986;
assign addr[45085] = -1402225355;
assign addr[45086] = -1387686535;
assign addr[45087] = -1373037681;
assign addr[45088] = -1358279953;
assign addr[45089] = -1343414522;
assign addr[45090] = -1328442566;
assign addr[45091] = -1313365273;
assign addr[45092] = -1298183838;
assign addr[45093] = -1282899464;
assign addr[45094] = -1267513365;
assign addr[45095] = -1252026760;
assign addr[45096] = -1236440877;
assign addr[45097] = -1220756951;
assign addr[45098] = -1204976227;
assign addr[45099] = -1189099956;
assign addr[45100] = -1173129396;
assign addr[45101] = -1157065814;
assign addr[45102] = -1140910484;
assign addr[45103] = -1124664687;
assign addr[45104] = -1108329711;
assign addr[45105] = -1091906851;
assign addr[45106] = -1075397409;
assign addr[45107] = -1058802695;
assign addr[45108] = -1042124025;
assign addr[45109] = -1025362720;
assign addr[45110] = -1008520110;
assign addr[45111] = -991597531;
assign addr[45112] = -974596324;
assign addr[45113] = -957517838;
assign addr[45114] = -940363427;
assign addr[45115] = -923134450;
assign addr[45116] = -905832274;
assign addr[45117] = -888458272;
assign addr[45118] = -871013820;
assign addr[45119] = -853500302;
assign addr[45120] = -835919107;
assign addr[45121] = -818271628;
assign addr[45122] = -800559266;
assign addr[45123] = -782783424;
assign addr[45124] = -764945512;
assign addr[45125] = -747046944;
assign addr[45126] = -729089140;
assign addr[45127] = -711073525;
assign addr[45128] = -693001525;
assign addr[45129] = -674874574;
assign addr[45130] = -656694110;
assign addr[45131] = -638461574;
assign addr[45132] = -620178412;
assign addr[45133] = -601846074;
assign addr[45134] = -583466013;
assign addr[45135] = -565039687;
assign addr[45136] = -546568556;
assign addr[45137] = -528054086;
assign addr[45138] = -509497745;
assign addr[45139] = -490901003;
assign addr[45140] = -472265336;
assign addr[45141] = -453592221;
assign addr[45142] = -434883140;
assign addr[45143] = -416139574;
assign addr[45144] = -397363011;
assign addr[45145] = -378554940;
assign addr[45146] = -359716852;
assign addr[45147] = -340850240;
assign addr[45148] = -321956601;
assign addr[45149] = -303037433;
assign addr[45150] = -284094236;
assign addr[45151] = -265128512;
assign addr[45152] = -246141764;
assign addr[45153] = -227135500;
assign addr[45154] = -208111224;
assign addr[45155] = -189070447;
assign addr[45156] = -170014678;
assign addr[45157] = -150945428;
assign addr[45158] = -131864208;
assign addr[45159] = -112772533;
assign addr[45160] = -93671915;
assign addr[45161] = -74563870;
assign addr[45162] = -55449912;
assign addr[45163] = -36331557;
assign addr[45164] = -17210322;
assign addr[45165] = 1912278;
assign addr[45166] = 21034727;
assign addr[45167] = 40155507;
assign addr[45168] = 59273104;
assign addr[45169] = 78386000;
assign addr[45170] = 97492681;
assign addr[45171] = 116591632;
assign addr[45172] = 135681337;
assign addr[45173] = 154760284;
assign addr[45174] = 173826959;
assign addr[45175] = 192879850;
assign addr[45176] = 211917448;
assign addr[45177] = 230938242;
assign addr[45178] = 249940723;
assign addr[45179] = 268923386;
assign addr[45180] = 287884725;
assign addr[45181] = 306823237;
assign addr[45182] = 325737419;
assign addr[45183] = 344625773;
assign addr[45184] = 363486799;
assign addr[45185] = 382319004;
assign addr[45186] = 401120892;
assign addr[45187] = 419890975;
assign addr[45188] = 438627762;
assign addr[45189] = 457329769;
assign addr[45190] = 475995513;
assign addr[45191] = 494623513;
assign addr[45192] = 513212292;
assign addr[45193] = 531760377;
assign addr[45194] = 550266296;
assign addr[45195] = 568728583;
assign addr[45196] = 587145773;
assign addr[45197] = 605516406;
assign addr[45198] = 623839025;
assign addr[45199] = 642112178;
assign addr[45200] = 660334415;
assign addr[45201] = 678504291;
assign addr[45202] = 696620367;
assign addr[45203] = 714681204;
assign addr[45204] = 732685372;
assign addr[45205] = 750631442;
assign addr[45206] = 768517992;
assign addr[45207] = 786343603;
assign addr[45208] = 804106861;
assign addr[45209] = 821806359;
assign addr[45210] = 839440693;
assign addr[45211] = 857008464;
assign addr[45212] = 874508280;
assign addr[45213] = 891938752;
assign addr[45214] = 909298500;
assign addr[45215] = 926586145;
assign addr[45216] = 943800318;
assign addr[45217] = 960939653;
assign addr[45218] = 978002791;
assign addr[45219] = 994988380;
assign addr[45220] = 1011895073;
assign addr[45221] = 1028721528;
assign addr[45222] = 1045466412;
assign addr[45223] = 1062128397;
assign addr[45224] = 1078706161;
assign addr[45225] = 1095198391;
assign addr[45226] = 1111603778;
assign addr[45227] = 1127921022;
assign addr[45228] = 1144148829;
assign addr[45229] = 1160285911;
assign addr[45230] = 1176330990;
assign addr[45231] = 1192282793;
assign addr[45232] = 1208140056;
assign addr[45233] = 1223901520;
assign addr[45234] = 1239565936;
assign addr[45235] = 1255132063;
assign addr[45236] = 1270598665;
assign addr[45237] = 1285964516;
assign addr[45238] = 1301228398;
assign addr[45239] = 1316389101;
assign addr[45240] = 1331445422;
assign addr[45241] = 1346396168;
assign addr[45242] = 1361240152;
assign addr[45243] = 1375976199;
assign addr[45244] = 1390603139;
assign addr[45245] = 1405119813;
assign addr[45246] = 1419525069;
assign addr[45247] = 1433817766;
assign addr[45248] = 1447996770;
assign addr[45249] = 1462060956;
assign addr[45250] = 1476009210;
assign addr[45251] = 1489840425;
assign addr[45252] = 1503553506;
assign addr[45253] = 1517147363;
assign addr[45254] = 1530620920;
assign addr[45255] = 1543973108;
assign addr[45256] = 1557202869;
assign addr[45257] = 1570309153;
assign addr[45258] = 1583290921;
assign addr[45259] = 1596147143;
assign addr[45260] = 1608876801;
assign addr[45261] = 1621478885;
assign addr[45262] = 1633952396;
assign addr[45263] = 1646296344;
assign addr[45264] = 1658509750;
assign addr[45265] = 1670591647;
assign addr[45266] = 1682541077;
assign addr[45267] = 1694357091;
assign addr[45268] = 1706038753;
assign addr[45269] = 1717585136;
assign addr[45270] = 1728995326;
assign addr[45271] = 1740268417;
assign addr[45272] = 1751403515;
assign addr[45273] = 1762399737;
assign addr[45274] = 1773256212;
assign addr[45275] = 1783972079;
assign addr[45276] = 1794546487;
assign addr[45277] = 1804978599;
assign addr[45278] = 1815267588;
assign addr[45279] = 1825412636;
assign addr[45280] = 1835412941;
assign addr[45281] = 1845267708;
assign addr[45282] = 1854976157;
assign addr[45283] = 1864537518;
assign addr[45284] = 1873951032;
assign addr[45285] = 1883215953;
assign addr[45286] = 1892331547;
assign addr[45287] = 1901297091;
assign addr[45288] = 1910111873;
assign addr[45289] = 1918775195;
assign addr[45290] = 1927286370;
assign addr[45291] = 1935644723;
assign addr[45292] = 1943849591;
assign addr[45293] = 1951900324;
assign addr[45294] = 1959796283;
assign addr[45295] = 1967536842;
assign addr[45296] = 1975121388;
assign addr[45297] = 1982549318;
assign addr[45298] = 1989820044;
assign addr[45299] = 1996932990;
assign addr[45300] = 2003887591;
assign addr[45301] = 2010683297;
assign addr[45302] = 2017319567;
assign addr[45303] = 2023795876;
assign addr[45304] = 2030111710;
assign addr[45305] = 2036266570;
assign addr[45306] = 2042259965;
assign addr[45307] = 2048091422;
assign addr[45308] = 2053760478;
assign addr[45309] = 2059266683;
assign addr[45310] = 2064609600;
assign addr[45311] = 2069788807;
assign addr[45312] = 2074803892;
assign addr[45313] = 2079654458;
assign addr[45314] = 2084340120;
assign addr[45315] = 2088860507;
assign addr[45316] = 2093215260;
assign addr[45317] = 2097404033;
assign addr[45318] = 2101426496;
assign addr[45319] = 2105282327;
assign addr[45320] = 2108971223;
assign addr[45321] = 2112492891;
assign addr[45322] = 2115847050;
assign addr[45323] = 2119033436;
assign addr[45324] = 2122051796;
assign addr[45325] = 2124901890;
assign addr[45326] = 2127583492;
assign addr[45327] = 2130096389;
assign addr[45328] = 2132440383;
assign addr[45329] = 2134615288;
assign addr[45330] = 2136620930;
assign addr[45331] = 2138457152;
assign addr[45332] = 2140123807;
assign addr[45333] = 2141620763;
assign addr[45334] = 2142947902;
assign addr[45335] = 2144105118;
assign addr[45336] = 2145092320;
assign addr[45337] = 2145909429;
assign addr[45338] = 2146556380;
assign addr[45339] = 2147033123;
assign addr[45340] = 2147339619;
assign addr[45341] = 2147475844;
assign addr[45342] = 2147441787;
assign addr[45343] = 2147237452;
assign addr[45344] = 2146862854;
assign addr[45345] = 2146318022;
assign addr[45346] = 2145603001;
assign addr[45347] = 2144717846;
assign addr[45348] = 2143662628;
assign addr[45349] = 2142437431;
assign addr[45350] = 2141042352;
assign addr[45351] = 2139477502;
assign addr[45352] = 2137743003;
assign addr[45353] = 2135838995;
assign addr[45354] = 2133765628;
assign addr[45355] = 2131523066;
assign addr[45356] = 2129111488;
assign addr[45357] = 2126531084;
assign addr[45358] = 2123782059;
assign addr[45359] = 2120864631;
assign addr[45360] = 2117779031;
assign addr[45361] = 2114525505;
assign addr[45362] = 2111104309;
assign addr[45363] = 2107515716;
assign addr[45364] = 2103760010;
assign addr[45365] = 2099837489;
assign addr[45366] = 2095748463;
assign addr[45367] = 2091493257;
assign addr[45368] = 2087072209;
assign addr[45369] = 2082485668;
assign addr[45370] = 2077733999;
assign addr[45371] = 2072817579;
assign addr[45372] = 2067736796;
assign addr[45373] = 2062492055;
assign addr[45374] = 2057083771;
assign addr[45375] = 2051512372;
assign addr[45376] = 2045778302;
assign addr[45377] = 2039882013;
assign addr[45378] = 2033823974;
assign addr[45379] = 2027604666;
assign addr[45380] = 2021224581;
assign addr[45381] = 2014684225;
assign addr[45382] = 2007984117;
assign addr[45383] = 2001124788;
assign addr[45384] = 1994106782;
assign addr[45385] = 1986930656;
assign addr[45386] = 1979596978;
assign addr[45387] = 1972106330;
assign addr[45388] = 1964459306;
assign addr[45389] = 1956656513;
assign addr[45390] = 1948698568;
assign addr[45391] = 1940586104;
assign addr[45392] = 1932319763;
assign addr[45393] = 1923900201;
assign addr[45394] = 1915328086;
assign addr[45395] = 1906604097;
assign addr[45396] = 1897728925;
assign addr[45397] = 1888703276;
assign addr[45398] = 1879527863;
assign addr[45399] = 1870203416;
assign addr[45400] = 1860730673;
assign addr[45401] = 1851110385;
assign addr[45402] = 1841343316;
assign addr[45403] = 1831430239;
assign addr[45404] = 1821371941;
assign addr[45405] = 1811169220;
assign addr[45406] = 1800822883;
assign addr[45407] = 1790333753;
assign addr[45408] = 1779702660;
assign addr[45409] = 1768930447;
assign addr[45410] = 1758017969;
assign addr[45411] = 1746966091;
assign addr[45412] = 1735775690;
assign addr[45413] = 1724447652;
assign addr[45414] = 1712982875;
assign addr[45415] = 1701382270;
assign addr[45416] = 1689646755;
assign addr[45417] = 1677777262;
assign addr[45418] = 1665774731;
assign addr[45419] = 1653640115;
assign addr[45420] = 1641374375;
assign addr[45421] = 1628978484;
assign addr[45422] = 1616453425;
assign addr[45423] = 1603800191;
assign addr[45424] = 1591019785;
assign addr[45425] = 1578113222;
assign addr[45426] = 1565081523;
assign addr[45427] = 1551925723;
assign addr[45428] = 1538646865;
assign addr[45429] = 1525246002;
assign addr[45430] = 1511724196;
assign addr[45431] = 1498082520;
assign addr[45432] = 1484322054;
assign addr[45433] = 1470443891;
assign addr[45434] = 1456449131;
assign addr[45435] = 1442338884;
assign addr[45436] = 1428114267;
assign addr[45437] = 1413776410;
assign addr[45438] = 1399326449;
assign addr[45439] = 1384765530;
assign addr[45440] = 1370094808;
assign addr[45441] = 1355315445;
assign addr[45442] = 1340428615;
assign addr[45443] = 1325435496;
assign addr[45444] = 1310337279;
assign addr[45445] = 1295135159;
assign addr[45446] = 1279830344;
assign addr[45447] = 1264424045;
assign addr[45448] = 1248917486;
assign addr[45449] = 1233311895;
assign addr[45450] = 1217608510;
assign addr[45451] = 1201808576;
assign addr[45452] = 1185913346;
assign addr[45453] = 1169924081;
assign addr[45454] = 1153842047;
assign addr[45455] = 1137668521;
assign addr[45456] = 1121404785;
assign addr[45457] = 1105052128;
assign addr[45458] = 1088611847;
assign addr[45459] = 1072085246;
assign addr[45460] = 1055473635;
assign addr[45461] = 1038778332;
assign addr[45462] = 1022000660;
assign addr[45463] = 1005141949;
assign addr[45464] = 988203537;
assign addr[45465] = 971186766;
assign addr[45466] = 954092986;
assign addr[45467] = 936923553;
assign addr[45468] = 919679827;
assign addr[45469] = 902363176;
assign addr[45470] = 884974973;
assign addr[45471] = 867516597;
assign addr[45472] = 849989433;
assign addr[45473] = 832394869;
assign addr[45474] = 814734301;
assign addr[45475] = 797009130;
assign addr[45476] = 779220762;
assign addr[45477] = 761370605;
assign addr[45478] = 743460077;
assign addr[45479] = 725490597;
assign addr[45480] = 707463589;
assign addr[45481] = 689380485;
assign addr[45482] = 671242716;
assign addr[45483] = 653051723;
assign addr[45484] = 634808946;
assign addr[45485] = 616515832;
assign addr[45486] = 598173833;
assign addr[45487] = 579784402;
assign addr[45488] = 561348998;
assign addr[45489] = 542869083;
assign addr[45490] = 524346121;
assign addr[45491] = 505781581;
assign addr[45492] = 487176937;
assign addr[45493] = 468533662;
assign addr[45494] = 449853235;
assign addr[45495] = 431137138;
assign addr[45496] = 412386854;
assign addr[45497] = 393603870;
assign addr[45498] = 374789676;
assign addr[45499] = 355945764;
assign addr[45500] = 337073627;
assign addr[45501] = 318174762;
assign addr[45502] = 299250668;
assign addr[45503] = 280302845;
assign addr[45504] = 261332796;
assign addr[45505] = 242342025;
assign addr[45506] = 223332037;
assign addr[45507] = 204304341;
assign addr[45508] = 185260444;
assign addr[45509] = 166201858;
assign addr[45510] = 147130093;
assign addr[45511] = 128046661;
assign addr[45512] = 108953076;
assign addr[45513] = 89850852;
assign addr[45514] = 70741503;
assign addr[45515] = 51626544;
assign addr[45516] = 32507492;
assign addr[45517] = 13385863;
assign addr[45518] = -5736829;
assign addr[45519] = -24859065;
assign addr[45520] = -43979330;
assign addr[45521] = -63096108;
assign addr[45522] = -82207882;
assign addr[45523] = -101313138;
assign addr[45524] = -120410361;
assign addr[45525] = -139498035;
assign addr[45526] = -158574649;
assign addr[45527] = -177638688;
assign addr[45528] = -196688642;
assign addr[45529] = -215722999;
assign addr[45530] = -234740251;
assign addr[45531] = -253738890;
assign addr[45532] = -272717408;
assign addr[45533] = -291674302;
assign addr[45534] = -310608068;
assign addr[45535] = -329517204;
assign addr[45536] = -348400212;
assign addr[45537] = -367255594;
assign addr[45538] = -386081854;
assign addr[45539] = -404877501;
assign addr[45540] = -423641043;
assign addr[45541] = -442370993;
assign addr[45542] = -461065866;
assign addr[45543] = -479724180;
assign addr[45544] = -498344454;
assign addr[45545] = -516925212;
assign addr[45546] = -535464981;
assign addr[45547] = -553962291;
assign addr[45548] = -572415676;
assign addr[45549] = -590823671;
assign addr[45550] = -609184818;
assign addr[45551] = -627497660;
assign addr[45552] = -645760745;
assign addr[45553] = -663972625;
assign addr[45554] = -682131857;
assign addr[45555] = -700236999;
assign addr[45556] = -718286617;
assign addr[45557] = -736279279;
assign addr[45558] = -754213559;
assign addr[45559] = -772088034;
assign addr[45560] = -789901288;
assign addr[45561] = -807651907;
assign addr[45562] = -825338484;
assign addr[45563] = -842959617;
assign addr[45564] = -860513908;
assign addr[45565] = -877999966;
assign addr[45566] = -895416404;
assign addr[45567] = -912761841;
assign addr[45568] = -930034901;
assign addr[45569] = -947234215;
assign addr[45570] = -964358420;
assign addr[45571] = -981406156;
assign addr[45572] = -998376073;
assign addr[45573] = -1015266825;
assign addr[45574] = -1032077073;
assign addr[45575] = -1048805483;
assign addr[45576] = -1065450729;
assign addr[45577] = -1082011492;
assign addr[45578] = -1098486458;
assign addr[45579] = -1114874320;
assign addr[45580] = -1131173780;
assign addr[45581] = -1147383544;
assign addr[45582] = -1163502328;
assign addr[45583] = -1179528853;
assign addr[45584] = -1195461849;
assign addr[45585] = -1211300053;
assign addr[45586] = -1227042207;
assign addr[45587] = -1242687064;
assign addr[45588] = -1258233384;
assign addr[45589] = -1273679934;
assign addr[45590] = -1289025489;
assign addr[45591] = -1304268832;
assign addr[45592] = -1319408754;
assign addr[45593] = -1334444055;
assign addr[45594] = -1349373543;
assign addr[45595] = -1364196034;
assign addr[45596] = -1378910353;
assign addr[45597] = -1393515332;
assign addr[45598] = -1408009814;
assign addr[45599] = -1422392650;
assign addr[45600] = -1436662698;
assign addr[45601] = -1450818828;
assign addr[45602] = -1464859917;
assign addr[45603] = -1478784851;
assign addr[45604] = -1492592527;
assign addr[45605] = -1506281850;
assign addr[45606] = -1519851733;
assign addr[45607] = -1533301101;
assign addr[45608] = -1546628888;
assign addr[45609] = -1559834037;
assign addr[45610] = -1572915501;
assign addr[45611] = -1585872242;
assign addr[45612] = -1598703233;
assign addr[45613] = -1611407456;
assign addr[45614] = -1623983905;
assign addr[45615] = -1636431582;
assign addr[45616] = -1648749499;
assign addr[45617] = -1660936681;
assign addr[45618] = -1672992161;
assign addr[45619] = -1684914983;
assign addr[45620] = -1696704201;
assign addr[45621] = -1708358881;
assign addr[45622] = -1719878099;
assign addr[45623] = -1731260941;
assign addr[45624] = -1742506504;
assign addr[45625] = -1753613897;
assign addr[45626] = -1764582240;
assign addr[45627] = -1775410662;
assign addr[45628] = -1786098304;
assign addr[45629] = -1796644320;
assign addr[45630] = -1807047873;
assign addr[45631] = -1817308138;
assign addr[45632] = -1827424302;
assign addr[45633] = -1837395562;
assign addr[45634] = -1847221128;
assign addr[45635] = -1856900221;
assign addr[45636] = -1866432072;
assign addr[45637] = -1875815927;
assign addr[45638] = -1885051042;
assign addr[45639] = -1894136683;
assign addr[45640] = -1903072131;
assign addr[45641] = -1911856677;
assign addr[45642] = -1920489624;
assign addr[45643] = -1928970288;
assign addr[45644] = -1937297997;
assign addr[45645] = -1945472089;
assign addr[45646] = -1953491918;
assign addr[45647] = -1961356847;
assign addr[45648] = -1969066252;
assign addr[45649] = -1976619522;
assign addr[45650] = -1984016058;
assign addr[45651] = -1991255274;
assign addr[45652] = -1998336596;
assign addr[45653] = -2005259462;
assign addr[45654] = -2012023322;
assign addr[45655] = -2018627642;
assign addr[45656] = -2025071897;
assign addr[45657] = -2031355576;
assign addr[45658] = -2037478181;
assign addr[45659] = -2043439226;
assign addr[45660] = -2049238240;
assign addr[45661] = -2054874761;
assign addr[45662] = -2060348343;
assign addr[45663] = -2065658552;
assign addr[45664] = -2070804967;
assign addr[45665] = -2075787180;
assign addr[45666] = -2080604795;
assign addr[45667] = -2085257431;
assign addr[45668] = -2089744719;
assign addr[45669] = -2094066304;
assign addr[45670] = -2098221841;
assign addr[45671] = -2102211002;
assign addr[45672] = -2106033471;
assign addr[45673] = -2109688944;
assign addr[45674] = -2113177132;
assign addr[45675] = -2116497758;
assign addr[45676] = -2119650558;
assign addr[45677] = -2122635283;
assign addr[45678] = -2125451696;
assign addr[45679] = -2128099574;
assign addr[45680] = -2130578706;
assign addr[45681] = -2132888897;
assign addr[45682] = -2135029962;
assign addr[45683] = -2137001733;
assign addr[45684] = -2138804053;
assign addr[45685] = -2140436778;
assign addr[45686] = -2141899780;
assign addr[45687] = -2143192942;
assign addr[45688] = -2144316162;
assign addr[45689] = -2145269351;
assign addr[45690] = -2146052433;
assign addr[45691] = -2146665347;
assign addr[45692] = -2147108043;
assign addr[45693] = -2147380486;
assign addr[45694] = -2147482655;
assign addr[45695] = -2147414542;
assign addr[45696] = -2147176152;
assign addr[45697] = -2146767505;
assign addr[45698] = -2146188631;
assign addr[45699] = -2145439578;
assign addr[45700] = -2144520405;
assign addr[45701] = -2143431184;
assign addr[45702] = -2142172003;
assign addr[45703] = -2140742960;
assign addr[45704] = -2139144169;
assign addr[45705] = -2137375758;
assign addr[45706] = -2135437865;
assign addr[45707] = -2133330646;
assign addr[45708] = -2131054266;
assign addr[45709] = -2128608907;
assign addr[45710] = -2125994762;
assign addr[45711] = -2123212038;
assign addr[45712] = -2120260957;
assign addr[45713] = -2117141752;
assign addr[45714] = -2113854671;
assign addr[45715] = -2110399974;
assign addr[45716] = -2106777935;
assign addr[45717] = -2102988841;
assign addr[45718] = -2099032994;
assign addr[45719] = -2094910706;
assign addr[45720] = -2090622304;
assign addr[45721] = -2086168128;
assign addr[45722] = -2081548533;
assign addr[45723] = -2076763883;
assign addr[45724] = -2071814558;
assign addr[45725] = -2066700952;
assign addr[45726] = -2061423468;
assign addr[45727] = -2055982526;
assign addr[45728] = -2050378558;
assign addr[45729] = -2044612007;
assign addr[45730] = -2038683330;
assign addr[45731] = -2032592999;
assign addr[45732] = -2026341495;
assign addr[45733] = -2019929315;
assign addr[45734] = -2013356967;
assign addr[45735] = -2006624971;
assign addr[45736] = -1999733863;
assign addr[45737] = -1992684188;
assign addr[45738] = -1985476506;
assign addr[45739] = -1978111387;
assign addr[45740] = -1970589416;
assign addr[45741] = -1962911189;
assign addr[45742] = -1955077316;
assign addr[45743] = -1947088417;
assign addr[45744] = -1938945125;
assign addr[45745] = -1930648088;
assign addr[45746] = -1922197961;
assign addr[45747] = -1913595416;
assign addr[45748] = -1904841135;
assign addr[45749] = -1895935811;
assign addr[45750] = -1886880151;
assign addr[45751] = -1877674873;
assign addr[45752] = -1868320707;
assign addr[45753] = -1858818395;
assign addr[45754] = -1849168689;
assign addr[45755] = -1839372356;
assign addr[45756] = -1829430172;
assign addr[45757] = -1819342925;
assign addr[45758] = -1809111415;
assign addr[45759] = -1798736454;
assign addr[45760] = -1788218865;
assign addr[45761] = -1777559480;
assign addr[45762] = -1766759146;
assign addr[45763] = -1755818718;
assign addr[45764] = -1744739065;
assign addr[45765] = -1733521064;
assign addr[45766] = -1722165606;
assign addr[45767] = -1710673591;
assign addr[45768] = -1699045930;
assign addr[45769] = -1687283545;
assign addr[45770] = -1675387369;
assign addr[45771] = -1663358344;
assign addr[45772] = -1651197426;
assign addr[45773] = -1638905577;
assign addr[45774] = -1626483774;
assign addr[45775] = -1613933000;
assign addr[45776] = -1601254251;
assign addr[45777] = -1588448533;
assign addr[45778] = -1575516860;
assign addr[45779] = -1562460258;
assign addr[45780] = -1549279763;
assign addr[45781] = -1535976419;
assign addr[45782] = -1522551282;
assign addr[45783] = -1509005416;
assign addr[45784] = -1495339895;
assign addr[45785] = -1481555802;
assign addr[45786] = -1467654232;
assign addr[45787] = -1453636285;
assign addr[45788] = -1439503074;
assign addr[45789] = -1425255719;
assign addr[45790] = -1410895350;
assign addr[45791] = -1396423105;
assign addr[45792] = -1381840133;
assign addr[45793] = -1367147589;
assign addr[45794] = -1352346639;
assign addr[45795] = -1337438456;
assign addr[45796] = -1322424222;
assign addr[45797] = -1307305128;
assign addr[45798] = -1292082373;
assign addr[45799] = -1276757164;
assign addr[45800] = -1261330715;
assign addr[45801] = -1245804251;
assign addr[45802] = -1230179002;
assign addr[45803] = -1214456207;
assign addr[45804] = -1198637114;
assign addr[45805] = -1182722976;
assign addr[45806] = -1166715055;
assign addr[45807] = -1150614620;
assign addr[45808] = -1134422949;
assign addr[45809] = -1118141326;
assign addr[45810] = -1101771040;
assign addr[45811] = -1085313391;
assign addr[45812] = -1068769683;
assign addr[45813] = -1052141228;
assign addr[45814] = -1035429345;
assign addr[45815] = -1018635358;
assign addr[45816] = -1001760600;
assign addr[45817] = -984806408;
assign addr[45818] = -967774128;
assign addr[45819] = -950665109;
assign addr[45820] = -933480707;
assign addr[45821] = -916222287;
assign addr[45822] = -898891215;
assign addr[45823] = -881488868;
assign addr[45824] = -864016623;
assign addr[45825] = -846475867;
assign addr[45826] = -828867991;
assign addr[45827] = -811194391;
assign addr[45828] = -793456467;
assign addr[45829] = -775655628;
assign addr[45830] = -757793284;
assign addr[45831] = -739870851;
assign addr[45832] = -721889752;
assign addr[45833] = -703851410;
assign addr[45834] = -685757258;
assign addr[45835] = -667608730;
assign addr[45836] = -649407264;
assign addr[45837] = -631154304;
assign addr[45838] = -612851297;
assign addr[45839] = -594499695;
assign addr[45840] = -576100953;
assign addr[45841] = -557656529;
assign addr[45842] = -539167887;
assign addr[45843] = -520636492;
assign addr[45844] = -502063814;
assign addr[45845] = -483451325;
assign addr[45846] = -464800501;
assign addr[45847] = -446112822;
assign addr[45848] = -427389768;
assign addr[45849] = -408632825;
assign addr[45850] = -389843480;
assign addr[45851] = -371023223;
assign addr[45852] = -352173546;
assign addr[45853] = -333295944;
assign addr[45854] = -314391913;
assign addr[45855] = -295462954;
assign addr[45856] = -276510565;
assign addr[45857] = -257536251;
assign addr[45858] = -238541516;
assign addr[45859] = -219527866;
assign addr[45860] = -200496809;
assign addr[45861] = -181449854;
assign addr[45862] = -162388511;
assign addr[45863] = -143314291;
assign addr[45864] = -124228708;
assign addr[45865] = -105133274;
assign addr[45866] = -86029503;
assign addr[45867] = -66918911;
assign addr[45868] = -47803013;
assign addr[45869] = -28683324;
assign addr[45870] = -9561361;
assign addr[45871] = 9561361;
assign addr[45872] = 28683324;
assign addr[45873] = 47803013;
assign addr[45874] = 66918911;
assign addr[45875] = 86029503;
assign addr[45876] = 105133274;
assign addr[45877] = 124228708;
assign addr[45878] = 143314291;
assign addr[45879] = 162388511;
assign addr[45880] = 181449854;
assign addr[45881] = 200496809;
assign addr[45882] = 219527866;
assign addr[45883] = 238541516;
assign addr[45884] = 257536251;
assign addr[45885] = 276510565;
assign addr[45886] = 295462953;
assign addr[45887] = 314391913;
assign addr[45888] = 333295944;
assign addr[45889] = 352173546;
assign addr[45890] = 371023223;
assign addr[45891] = 389843480;
assign addr[45892] = 408632825;
assign addr[45893] = 427389768;
assign addr[45894] = 446112822;
assign addr[45895] = 464800501;
assign addr[45896] = 483451325;
assign addr[45897] = 502063814;
assign addr[45898] = 520636492;
assign addr[45899] = 539167887;
assign addr[45900] = 557656529;
assign addr[45901] = 576100953;
assign addr[45902] = 594499695;
assign addr[45903] = 612851297;
assign addr[45904] = 631154304;
assign addr[45905] = 649407264;
assign addr[45906] = 667608730;
assign addr[45907] = 685757258;
assign addr[45908] = 703851410;
assign addr[45909] = 721889752;
assign addr[45910] = 739870851;
assign addr[45911] = 757793284;
assign addr[45912] = 775655628;
assign addr[45913] = 793456467;
assign addr[45914] = 811194391;
assign addr[45915] = 828867991;
assign addr[45916] = 846475867;
assign addr[45917] = 864016623;
assign addr[45918] = 881488868;
assign addr[45919] = 898891215;
assign addr[45920] = 916222287;
assign addr[45921] = 933480707;
assign addr[45922] = 950665109;
assign addr[45923] = 967774128;
assign addr[45924] = 984806408;
assign addr[45925] = 1001760600;
assign addr[45926] = 1018635358;
assign addr[45927] = 1035429345;
assign addr[45928] = 1052141228;
assign addr[45929] = 1068769683;
assign addr[45930] = 1085313391;
assign addr[45931] = 1101771040;
assign addr[45932] = 1118141326;
assign addr[45933] = 1134422949;
assign addr[45934] = 1150614620;
assign addr[45935] = 1166715055;
assign addr[45936] = 1182722976;
assign addr[45937] = 1198637114;
assign addr[45938] = 1214456207;
assign addr[45939] = 1230179002;
assign addr[45940] = 1245804251;
assign addr[45941] = 1261330715;
assign addr[45942] = 1276757164;
assign addr[45943] = 1292082373;
assign addr[45944] = 1307305128;
assign addr[45945] = 1322424222;
assign addr[45946] = 1337438456;
assign addr[45947] = 1352346639;
assign addr[45948] = 1367147589;
assign addr[45949] = 1381840133;
assign addr[45950] = 1396423105;
assign addr[45951] = 1410895350;
assign addr[45952] = 1425255719;
assign addr[45953] = 1439503074;
assign addr[45954] = 1453636285;
assign addr[45955] = 1467654232;
assign addr[45956] = 1481555802;
assign addr[45957] = 1495339895;
assign addr[45958] = 1509005416;
assign addr[45959] = 1522551282;
assign addr[45960] = 1535976419;
assign addr[45961] = 1549279763;
assign addr[45962] = 1562460258;
assign addr[45963] = 1575516860;
assign addr[45964] = 1588448533;
assign addr[45965] = 1601254251;
assign addr[45966] = 1613933000;
assign addr[45967] = 1626483774;
assign addr[45968] = 1638905577;
assign addr[45969] = 1651197426;
assign addr[45970] = 1663358344;
assign addr[45971] = 1675387369;
assign addr[45972] = 1687283545;
assign addr[45973] = 1699045930;
assign addr[45974] = 1710673591;
assign addr[45975] = 1722165606;
assign addr[45976] = 1733521064;
assign addr[45977] = 1744739065;
assign addr[45978] = 1755818718;
assign addr[45979] = 1766759146;
assign addr[45980] = 1777559480;
assign addr[45981] = 1788218865;
assign addr[45982] = 1798736454;
assign addr[45983] = 1809111415;
assign addr[45984] = 1819342925;
assign addr[45985] = 1829430172;
assign addr[45986] = 1839372356;
assign addr[45987] = 1849168689;
assign addr[45988] = 1858818395;
assign addr[45989] = 1868320707;
assign addr[45990] = 1877674873;
assign addr[45991] = 1886880151;
assign addr[45992] = 1895935811;
assign addr[45993] = 1904841135;
assign addr[45994] = 1913595416;
assign addr[45995] = 1922197961;
assign addr[45996] = 1930648088;
assign addr[45997] = 1938945125;
assign addr[45998] = 1947088417;
assign addr[45999] = 1955077316;
assign addr[46000] = 1962911189;
assign addr[46001] = 1970589416;
assign addr[46002] = 1978111387;
assign addr[46003] = 1985476506;
assign addr[46004] = 1992684188;
assign addr[46005] = 1999733863;
assign addr[46006] = 2006624971;
assign addr[46007] = 2013356967;
assign addr[46008] = 2019929315;
assign addr[46009] = 2026341495;
assign addr[46010] = 2032592999;
assign addr[46011] = 2038683330;
assign addr[46012] = 2044612007;
assign addr[46013] = 2050378558;
assign addr[46014] = 2055982526;
assign addr[46015] = 2061423468;
assign addr[46016] = 2066700952;
assign addr[46017] = 2071814558;
assign addr[46018] = 2076763883;
assign addr[46019] = 2081548533;
assign addr[46020] = 2086168128;
assign addr[46021] = 2090622304;
assign addr[46022] = 2094910706;
assign addr[46023] = 2099032994;
assign addr[46024] = 2102988841;
assign addr[46025] = 2106777935;
assign addr[46026] = 2110399974;
assign addr[46027] = 2113854671;
assign addr[46028] = 2117141752;
assign addr[46029] = 2120260957;
assign addr[46030] = 2123212038;
assign addr[46031] = 2125994762;
assign addr[46032] = 2128608907;
assign addr[46033] = 2131054266;
assign addr[46034] = 2133330646;
assign addr[46035] = 2135437865;
assign addr[46036] = 2137375758;
assign addr[46037] = 2139144169;
assign addr[46038] = 2140742960;
assign addr[46039] = 2142172003;
assign addr[46040] = 2143431184;
assign addr[46041] = 2144520405;
assign addr[46042] = 2145439578;
assign addr[46043] = 2146188631;
assign addr[46044] = 2146767505;
assign addr[46045] = 2147176152;
assign addr[46046] = 2147414542;
assign addr[46047] = 2147482655;
assign addr[46048] = 2147380486;
assign addr[46049] = 2147108043;
assign addr[46050] = 2146665347;
assign addr[46051] = 2146052433;
assign addr[46052] = 2145269351;
assign addr[46053] = 2144316162;
assign addr[46054] = 2143192942;
assign addr[46055] = 2141899780;
assign addr[46056] = 2140436778;
assign addr[46057] = 2138804053;
assign addr[46058] = 2137001733;
assign addr[46059] = 2135029962;
assign addr[46060] = 2132888897;
assign addr[46061] = 2130578706;
assign addr[46062] = 2128099574;
assign addr[46063] = 2125451696;
assign addr[46064] = 2122635283;
assign addr[46065] = 2119650558;
assign addr[46066] = 2116497758;
assign addr[46067] = 2113177132;
assign addr[46068] = 2109688944;
assign addr[46069] = 2106033471;
assign addr[46070] = 2102211002;
assign addr[46071] = 2098221841;
assign addr[46072] = 2094066304;
assign addr[46073] = 2089744719;
assign addr[46074] = 2085257431;
assign addr[46075] = 2080604795;
assign addr[46076] = 2075787180;
assign addr[46077] = 2070804967;
assign addr[46078] = 2065658552;
assign addr[46079] = 2060348343;
assign addr[46080] = 2054874761;
assign addr[46081] = 2049238240;
assign addr[46082] = 2043439226;
assign addr[46083] = 2037478181;
assign addr[46084] = 2031355576;
assign addr[46085] = 2025071897;
assign addr[46086] = 2018627642;
assign addr[46087] = 2012023322;
assign addr[46088] = 2005259462;
assign addr[46089] = 1998336596;
assign addr[46090] = 1991255274;
assign addr[46091] = 1984016058;
assign addr[46092] = 1976619522;
assign addr[46093] = 1969066252;
assign addr[46094] = 1961356847;
assign addr[46095] = 1953491918;
assign addr[46096] = 1945472089;
assign addr[46097] = 1937297997;
assign addr[46098] = 1928970288;
assign addr[46099] = 1920489624;
assign addr[46100] = 1911856677;
assign addr[46101] = 1903072131;
assign addr[46102] = 1894136683;
assign addr[46103] = 1885051042;
assign addr[46104] = 1875815927;
assign addr[46105] = 1866432072;
assign addr[46106] = 1856900221;
assign addr[46107] = 1847221128;
assign addr[46108] = 1837395562;
assign addr[46109] = 1827424302;
assign addr[46110] = 1817308138;
assign addr[46111] = 1807047873;
assign addr[46112] = 1796644320;
assign addr[46113] = 1786098304;
assign addr[46114] = 1775410662;
assign addr[46115] = 1764582240;
assign addr[46116] = 1753613897;
assign addr[46117] = 1742506504;
assign addr[46118] = 1731260941;
assign addr[46119] = 1719878099;
assign addr[46120] = 1708358881;
assign addr[46121] = 1696704201;
assign addr[46122] = 1684914983;
assign addr[46123] = 1672992161;
assign addr[46124] = 1660936681;
assign addr[46125] = 1648749499;
assign addr[46126] = 1636431582;
assign addr[46127] = 1623983905;
assign addr[46128] = 1611407456;
assign addr[46129] = 1598703233;
assign addr[46130] = 1585872242;
assign addr[46131] = 1572915501;
assign addr[46132] = 1559834037;
assign addr[46133] = 1546628888;
assign addr[46134] = 1533301101;
assign addr[46135] = 1519851733;
assign addr[46136] = 1506281850;
assign addr[46137] = 1492592527;
assign addr[46138] = 1478784851;
assign addr[46139] = 1464859917;
assign addr[46140] = 1450818828;
assign addr[46141] = 1436662698;
assign addr[46142] = 1422392650;
assign addr[46143] = 1408009814;
assign addr[46144] = 1393515332;
assign addr[46145] = 1378910353;
assign addr[46146] = 1364196034;
assign addr[46147] = 1349373543;
assign addr[46148] = 1334444055;
assign addr[46149] = 1319408754;
assign addr[46150] = 1304268832;
assign addr[46151] = 1289025489;
assign addr[46152] = 1273679934;
assign addr[46153] = 1258233384;
assign addr[46154] = 1242687064;
assign addr[46155] = 1227042207;
assign addr[46156] = 1211300053;
assign addr[46157] = 1195461849;
assign addr[46158] = 1179528853;
assign addr[46159] = 1163502328;
assign addr[46160] = 1147383544;
assign addr[46161] = 1131173780;
assign addr[46162] = 1114874320;
assign addr[46163] = 1098486458;
assign addr[46164] = 1082011492;
assign addr[46165] = 1065450729;
assign addr[46166] = 1048805483;
assign addr[46167] = 1032077073;
assign addr[46168] = 1015266825;
assign addr[46169] = 998376073;
assign addr[46170] = 981406156;
assign addr[46171] = 964358420;
assign addr[46172] = 947234215;
assign addr[46173] = 930034901;
assign addr[46174] = 912761841;
assign addr[46175] = 895416404;
assign addr[46176] = 877999966;
assign addr[46177] = 860513908;
assign addr[46178] = 842959617;
assign addr[46179] = 825338484;
assign addr[46180] = 807651907;
assign addr[46181] = 789901288;
assign addr[46182] = 772088034;
assign addr[46183] = 754213559;
assign addr[46184] = 736279279;
assign addr[46185] = 718286617;
assign addr[46186] = 700236999;
assign addr[46187] = 682131857;
assign addr[46188] = 663972625;
assign addr[46189] = 645760745;
assign addr[46190] = 627497660;
assign addr[46191] = 609184818;
assign addr[46192] = 590823671;
assign addr[46193] = 572415676;
assign addr[46194] = 553962291;
assign addr[46195] = 535464981;
assign addr[46196] = 516925212;
assign addr[46197] = 498344454;
assign addr[46198] = 479724180;
assign addr[46199] = 461065866;
assign addr[46200] = 442370993;
assign addr[46201] = 423641043;
assign addr[46202] = 404877501;
assign addr[46203] = 386081854;
assign addr[46204] = 367255594;
assign addr[46205] = 348400212;
assign addr[46206] = 329517204;
assign addr[46207] = 310608068;
assign addr[46208] = 291674302;
assign addr[46209] = 272717408;
assign addr[46210] = 253738890;
assign addr[46211] = 234740251;
assign addr[46212] = 215722999;
assign addr[46213] = 196688642;
assign addr[46214] = 177638688;
assign addr[46215] = 158574649;
assign addr[46216] = 139498035;
assign addr[46217] = 120410361;
assign addr[46218] = 101313138;
assign addr[46219] = 82207882;
assign addr[46220] = 63096108;
assign addr[46221] = 43979330;
assign addr[46222] = 24859065;
assign addr[46223] = 5736829;
assign addr[46224] = -13385863;
assign addr[46225] = -32507492;
assign addr[46226] = -51626544;
assign addr[46227] = -70741503;
assign addr[46228] = -89850852;
assign addr[46229] = -108953076;
assign addr[46230] = -128046661;
assign addr[46231] = -147130093;
assign addr[46232] = -166201858;
assign addr[46233] = -185260444;
assign addr[46234] = -204304341;
assign addr[46235] = -223332037;
assign addr[46236] = -242342025;
assign addr[46237] = -261332796;
assign addr[46238] = -280302845;
assign addr[46239] = -299250668;
assign addr[46240] = -318174762;
assign addr[46241] = -337073627;
assign addr[46242] = -355945764;
assign addr[46243] = -374789676;
assign addr[46244] = -393603870;
assign addr[46245] = -412386854;
assign addr[46246] = -431137138;
assign addr[46247] = -449853235;
assign addr[46248] = -468533662;
assign addr[46249] = -487176937;
assign addr[46250] = -505781581;
assign addr[46251] = -524346121;
assign addr[46252] = -542869083;
assign addr[46253] = -561348998;
assign addr[46254] = -579784402;
assign addr[46255] = -598173833;
assign addr[46256] = -616515832;
assign addr[46257] = -634808946;
assign addr[46258] = -653051723;
assign addr[46259] = -671242716;
assign addr[46260] = -689380485;
assign addr[46261] = -707463589;
assign addr[46262] = -725490597;
assign addr[46263] = -743460077;
assign addr[46264] = -761370605;
assign addr[46265] = -779220762;
assign addr[46266] = -797009130;
assign addr[46267] = -814734301;
assign addr[46268] = -832394869;
assign addr[46269] = -849989433;
assign addr[46270] = -867516597;
assign addr[46271] = -884974973;
assign addr[46272] = -902363176;
assign addr[46273] = -919679827;
assign addr[46274] = -936923553;
assign addr[46275] = -954092986;
assign addr[46276] = -971186766;
assign addr[46277] = -988203537;
assign addr[46278] = -1005141949;
assign addr[46279] = -1022000660;
assign addr[46280] = -1038778332;
assign addr[46281] = -1055473635;
assign addr[46282] = -1072085246;
assign addr[46283] = -1088611847;
assign addr[46284] = -1105052128;
assign addr[46285] = -1121404785;
assign addr[46286] = -1137668521;
assign addr[46287] = -1153842047;
assign addr[46288] = -1169924081;
assign addr[46289] = -1185913346;
assign addr[46290] = -1201808576;
assign addr[46291] = -1217608510;
assign addr[46292] = -1233311895;
assign addr[46293] = -1248917486;
assign addr[46294] = -1264424045;
assign addr[46295] = -1279830344;
assign addr[46296] = -1295135159;
assign addr[46297] = -1310337279;
assign addr[46298] = -1325435496;
assign addr[46299] = -1340428615;
assign addr[46300] = -1355315445;
assign addr[46301] = -1370094808;
assign addr[46302] = -1384765530;
assign addr[46303] = -1399326449;
assign addr[46304] = -1413776410;
assign addr[46305] = -1428114267;
assign addr[46306] = -1442338884;
assign addr[46307] = -1456449131;
assign addr[46308] = -1470443891;
assign addr[46309] = -1484322054;
assign addr[46310] = -1498082520;
assign addr[46311] = -1511724196;
assign addr[46312] = -1525246002;
assign addr[46313] = -1538646865;
assign addr[46314] = -1551925723;
assign addr[46315] = -1565081523;
assign addr[46316] = -1578113222;
assign addr[46317] = -1591019785;
assign addr[46318] = -1603800191;
assign addr[46319] = -1616453425;
assign addr[46320] = -1628978484;
assign addr[46321] = -1641374375;
assign addr[46322] = -1653640115;
assign addr[46323] = -1665774731;
assign addr[46324] = -1677777262;
assign addr[46325] = -1689646755;
assign addr[46326] = -1701382270;
assign addr[46327] = -1712982875;
assign addr[46328] = -1724447652;
assign addr[46329] = -1735775690;
assign addr[46330] = -1746966091;
assign addr[46331] = -1758017969;
assign addr[46332] = -1768930447;
assign addr[46333] = -1779702660;
assign addr[46334] = -1790333753;
assign addr[46335] = -1800822883;
assign addr[46336] = -1811169220;
assign addr[46337] = -1821371941;
assign addr[46338] = -1831430239;
assign addr[46339] = -1841343316;
assign addr[46340] = -1851110385;
assign addr[46341] = -1860730673;
assign addr[46342] = -1870203416;
assign addr[46343] = -1879527863;
assign addr[46344] = -1888703276;
assign addr[46345] = -1897728925;
assign addr[46346] = -1906604097;
assign addr[46347] = -1915328086;
assign addr[46348] = -1923900201;
assign addr[46349] = -1932319763;
assign addr[46350] = -1940586104;
assign addr[46351] = -1948698568;
assign addr[46352] = -1956656513;
assign addr[46353] = -1964459306;
assign addr[46354] = -1972106330;
assign addr[46355] = -1979596978;
assign addr[46356] = -1986930656;
assign addr[46357] = -1994106782;
assign addr[46358] = -2001124788;
assign addr[46359] = -2007984117;
assign addr[46360] = -2014684225;
assign addr[46361] = -2021224581;
assign addr[46362] = -2027604666;
assign addr[46363] = -2033823974;
assign addr[46364] = -2039882013;
assign addr[46365] = -2045778302;
assign addr[46366] = -2051512372;
assign addr[46367] = -2057083771;
assign addr[46368] = -2062492055;
assign addr[46369] = -2067736796;
assign addr[46370] = -2072817579;
assign addr[46371] = -2077733999;
assign addr[46372] = -2082485668;
assign addr[46373] = -2087072209;
assign addr[46374] = -2091493257;
assign addr[46375] = -2095748463;
assign addr[46376] = -2099837489;
assign addr[46377] = -2103760010;
assign addr[46378] = -2107515716;
assign addr[46379] = -2111104309;
assign addr[46380] = -2114525505;
assign addr[46381] = -2117779031;
assign addr[46382] = -2120864631;
assign addr[46383] = -2123782059;
assign addr[46384] = -2126531084;
assign addr[46385] = -2129111488;
assign addr[46386] = -2131523066;
assign addr[46387] = -2133765628;
assign addr[46388] = -2135838995;
assign addr[46389] = -2137743003;
assign addr[46390] = -2139477502;
assign addr[46391] = -2141042352;
assign addr[46392] = -2142437431;
assign addr[46393] = -2143662628;
assign addr[46394] = -2144717846;
assign addr[46395] = -2145603001;
assign addr[46396] = -2146318022;
assign addr[46397] = -2146862854;
assign addr[46398] = -2147237452;
assign addr[46399] = -2147441787;
assign addr[46400] = -2147475844;
assign addr[46401] = -2147339619;
assign addr[46402] = -2147033123;
assign addr[46403] = -2146556380;
assign addr[46404] = -2145909429;
assign addr[46405] = -2145092320;
assign addr[46406] = -2144105118;
assign addr[46407] = -2142947902;
assign addr[46408] = -2141620763;
assign addr[46409] = -2140123807;
assign addr[46410] = -2138457152;
assign addr[46411] = -2136620930;
assign addr[46412] = -2134615288;
assign addr[46413] = -2132440383;
assign addr[46414] = -2130096389;
assign addr[46415] = -2127583492;
assign addr[46416] = -2124901890;
assign addr[46417] = -2122051796;
assign addr[46418] = -2119033436;
assign addr[46419] = -2115847050;
assign addr[46420] = -2112492891;
assign addr[46421] = -2108971223;
assign addr[46422] = -2105282327;
assign addr[46423] = -2101426496;
assign addr[46424] = -2097404033;
assign addr[46425] = -2093215260;
assign addr[46426] = -2088860507;
assign addr[46427] = -2084340120;
assign addr[46428] = -2079654458;
assign addr[46429] = -2074803892;
assign addr[46430] = -2069788807;
assign addr[46431] = -2064609600;
assign addr[46432] = -2059266683;
assign addr[46433] = -2053760478;
assign addr[46434] = -2048091422;
assign addr[46435] = -2042259965;
assign addr[46436] = -2036266570;
assign addr[46437] = -2030111710;
assign addr[46438] = -2023795876;
assign addr[46439] = -2017319567;
assign addr[46440] = -2010683297;
assign addr[46441] = -2003887591;
assign addr[46442] = -1996932990;
assign addr[46443] = -1989820044;
assign addr[46444] = -1982549318;
assign addr[46445] = -1975121388;
assign addr[46446] = -1967536842;
assign addr[46447] = -1959796283;
assign addr[46448] = -1951900324;
assign addr[46449] = -1943849591;
assign addr[46450] = -1935644723;
assign addr[46451] = -1927286370;
assign addr[46452] = -1918775195;
assign addr[46453] = -1910111873;
assign addr[46454] = -1901297091;
assign addr[46455] = -1892331547;
assign addr[46456] = -1883215953;
assign addr[46457] = -1873951032;
assign addr[46458] = -1864537518;
assign addr[46459] = -1854976157;
assign addr[46460] = -1845267708;
assign addr[46461] = -1835412941;
assign addr[46462] = -1825412636;
assign addr[46463] = -1815267588;
assign addr[46464] = -1804978599;
assign addr[46465] = -1794546487;
assign addr[46466] = -1783972079;
assign addr[46467] = -1773256212;
assign addr[46468] = -1762399737;
assign addr[46469] = -1751403515;
assign addr[46470] = -1740268417;
assign addr[46471] = -1728995326;
assign addr[46472] = -1717585136;
assign addr[46473] = -1706038753;
assign addr[46474] = -1694357091;
assign addr[46475] = -1682541077;
assign addr[46476] = -1670591647;
assign addr[46477] = -1658509750;
assign addr[46478] = -1646296344;
assign addr[46479] = -1633952396;
assign addr[46480] = -1621478885;
assign addr[46481] = -1608876801;
assign addr[46482] = -1596147143;
assign addr[46483] = -1583290921;
assign addr[46484] = -1570309153;
assign addr[46485] = -1557202869;
assign addr[46486] = -1543973108;
assign addr[46487] = -1530620920;
assign addr[46488] = -1517147363;
assign addr[46489] = -1503553506;
assign addr[46490] = -1489840425;
assign addr[46491] = -1476009210;
assign addr[46492] = -1462060956;
assign addr[46493] = -1447996770;
assign addr[46494] = -1433817766;
assign addr[46495] = -1419525069;
assign addr[46496] = -1405119813;
assign addr[46497] = -1390603139;
assign addr[46498] = -1375976199;
assign addr[46499] = -1361240152;
assign addr[46500] = -1346396168;
assign addr[46501] = -1331445422;
assign addr[46502] = -1316389101;
assign addr[46503] = -1301228398;
assign addr[46504] = -1285964516;
assign addr[46505] = -1270598665;
assign addr[46506] = -1255132063;
assign addr[46507] = -1239565936;
assign addr[46508] = -1223901520;
assign addr[46509] = -1208140056;
assign addr[46510] = -1192282793;
assign addr[46511] = -1176330990;
assign addr[46512] = -1160285911;
assign addr[46513] = -1144148829;
assign addr[46514] = -1127921022;
assign addr[46515] = -1111603778;
assign addr[46516] = -1095198391;
assign addr[46517] = -1078706161;
assign addr[46518] = -1062128397;
assign addr[46519] = -1045466412;
assign addr[46520] = -1028721528;
assign addr[46521] = -1011895073;
assign addr[46522] = -994988380;
assign addr[46523] = -978002791;
assign addr[46524] = -960939653;
assign addr[46525] = -943800318;
assign addr[46526] = -926586145;
assign addr[46527] = -909298500;
assign addr[46528] = -891938752;
assign addr[46529] = -874508280;
assign addr[46530] = -857008464;
assign addr[46531] = -839440693;
assign addr[46532] = -821806359;
assign addr[46533] = -804106861;
assign addr[46534] = -786343603;
assign addr[46535] = -768517992;
assign addr[46536] = -750631442;
assign addr[46537] = -732685372;
assign addr[46538] = -714681204;
assign addr[46539] = -696620367;
assign addr[46540] = -678504291;
assign addr[46541] = -660334415;
assign addr[46542] = -642112178;
assign addr[46543] = -623839025;
assign addr[46544] = -605516406;
assign addr[46545] = -587145773;
assign addr[46546] = -568728583;
assign addr[46547] = -550266296;
assign addr[46548] = -531760377;
assign addr[46549] = -513212292;
assign addr[46550] = -494623513;
assign addr[46551] = -475995513;
assign addr[46552] = -457329769;
assign addr[46553] = -438627762;
assign addr[46554] = -419890975;
assign addr[46555] = -401120892;
assign addr[46556] = -382319004;
assign addr[46557] = -363486799;
assign addr[46558] = -344625773;
assign addr[46559] = -325737419;
assign addr[46560] = -306823237;
assign addr[46561] = -287884725;
assign addr[46562] = -268923386;
assign addr[46563] = -249940723;
assign addr[46564] = -230938242;
assign addr[46565] = -211917448;
assign addr[46566] = -192879850;
assign addr[46567] = -173826959;
assign addr[46568] = -154760284;
assign addr[46569] = -135681337;
assign addr[46570] = -116591632;
assign addr[46571] = -97492681;
assign addr[46572] = -78386000;
assign addr[46573] = -59273104;
assign addr[46574] = -40155507;
assign addr[46575] = -21034727;
assign addr[46576] = -1912278;
assign addr[46577] = 17210322;
assign addr[46578] = 36331557;
assign addr[46579] = 55449912;
assign addr[46580] = 74563870;
assign addr[46581] = 93671915;
assign addr[46582] = 112772533;
assign addr[46583] = 131864208;
assign addr[46584] = 150945428;
assign addr[46585] = 170014678;
assign addr[46586] = 189070447;
assign addr[46587] = 208111224;
assign addr[46588] = 227135500;
assign addr[46589] = 246141764;
assign addr[46590] = 265128512;
assign addr[46591] = 284094236;
assign addr[46592] = 303037433;
assign addr[46593] = 321956601;
assign addr[46594] = 340850240;
assign addr[46595] = 359716852;
assign addr[46596] = 378554940;
assign addr[46597] = 397363011;
assign addr[46598] = 416139574;
assign addr[46599] = 434883140;
assign addr[46600] = 453592221;
assign addr[46601] = 472265336;
assign addr[46602] = 490901003;
assign addr[46603] = 509497745;
assign addr[46604] = 528054086;
assign addr[46605] = 546568556;
assign addr[46606] = 565039687;
assign addr[46607] = 583466013;
assign addr[46608] = 601846074;
assign addr[46609] = 620178412;
assign addr[46610] = 638461574;
assign addr[46611] = 656694110;
assign addr[46612] = 674874574;
assign addr[46613] = 693001525;
assign addr[46614] = 711073524;
assign addr[46615] = 729089140;
assign addr[46616] = 747046944;
assign addr[46617] = 764945512;
assign addr[46618] = 782783424;
assign addr[46619] = 800559266;
assign addr[46620] = 818271628;
assign addr[46621] = 835919107;
assign addr[46622] = 853500302;
assign addr[46623] = 871013820;
assign addr[46624] = 888458272;
assign addr[46625] = 905832274;
assign addr[46626] = 923134450;
assign addr[46627] = 940363427;
assign addr[46628] = 957517838;
assign addr[46629] = 974596324;
assign addr[46630] = 991597531;
assign addr[46631] = 1008520110;
assign addr[46632] = 1025362720;
assign addr[46633] = 1042124025;
assign addr[46634] = 1058802695;
assign addr[46635] = 1075397409;
assign addr[46636] = 1091906851;
assign addr[46637] = 1108329711;
assign addr[46638] = 1124664687;
assign addr[46639] = 1140910484;
assign addr[46640] = 1157065814;
assign addr[46641] = 1173129396;
assign addr[46642] = 1189099956;
assign addr[46643] = 1204976227;
assign addr[46644] = 1220756951;
assign addr[46645] = 1236440877;
assign addr[46646] = 1252026760;
assign addr[46647] = 1267513365;
assign addr[46648] = 1282899464;
assign addr[46649] = 1298183838;
assign addr[46650] = 1313365273;
assign addr[46651] = 1328442566;
assign addr[46652] = 1343414522;
assign addr[46653] = 1358279953;
assign addr[46654] = 1373037681;
assign addr[46655] = 1387686535;
assign addr[46656] = 1402225355;
assign addr[46657] = 1416652986;
assign addr[46658] = 1430968286;
assign addr[46659] = 1445170118;
assign addr[46660] = 1459257358;
assign addr[46661] = 1473228887;
assign addr[46662] = 1487083598;
assign addr[46663] = 1500820393;
assign addr[46664] = 1514438181;
assign addr[46665] = 1527935884;
assign addr[46666] = 1541312431;
assign addr[46667] = 1554566762;
assign addr[46668] = 1567697824;
assign addr[46669] = 1580704578;
assign addr[46670] = 1593585992;
assign addr[46671] = 1606341043;
assign addr[46672] = 1618968722;
assign addr[46673] = 1631468027;
assign addr[46674] = 1643837966;
assign addr[46675] = 1656077559;
assign addr[46676] = 1668185835;
assign addr[46677] = 1680161834;
assign addr[46678] = 1692004606;
assign addr[46679] = 1703713213;
assign addr[46680] = 1715286726;
assign addr[46681] = 1726724227;
assign addr[46682] = 1738024810;
assign addr[46683] = 1749187577;
assign addr[46684] = 1760211645;
assign addr[46685] = 1771096139;
assign addr[46686] = 1781840195;
assign addr[46687] = 1792442963;
assign addr[46688] = 1802903601;
assign addr[46689] = 1813221279;
assign addr[46690] = 1823395180;
assign addr[46691] = 1833424497;
assign addr[46692] = 1843308435;
assign addr[46693] = 1853046210;
assign addr[46694] = 1862637049;
assign addr[46695] = 1872080193;
assign addr[46696] = 1881374892;
assign addr[46697] = 1890520410;
assign addr[46698] = 1899516021;
assign addr[46699] = 1908361011;
assign addr[46700] = 1917054681;
assign addr[46701] = 1925596340;
assign addr[46702] = 1933985310;
assign addr[46703] = 1942220928;
assign addr[46704] = 1950302539;
assign addr[46705] = 1958229503;
assign addr[46706] = 1966001192;
assign addr[46707] = 1973616989;
assign addr[46708] = 1981076290;
assign addr[46709] = 1988378503;
assign addr[46710] = 1995523051;
assign addr[46711] = 2002509365;
assign addr[46712] = 2009336893;
assign addr[46713] = 2016005093;
assign addr[46714] = 2022513436;
assign addr[46715] = 2028861406;
assign addr[46716] = 2035048499;
assign addr[46717] = 2041074226;
assign addr[46718] = 2046938108;
assign addr[46719] = 2052639680;
assign addr[46720] = 2058178491;
assign addr[46721] = 2063554100;
assign addr[46722] = 2068766083;
assign addr[46723] = 2073814024;
assign addr[46724] = 2078697525;
assign addr[46725] = 2083416198;
assign addr[46726] = 2087969669;
assign addr[46727] = 2092357577;
assign addr[46728] = 2096579573;
assign addr[46729] = 2100635323;
assign addr[46730] = 2104524506;
assign addr[46731] = 2108246813;
assign addr[46732] = 2111801949;
assign addr[46733] = 2115189632;
assign addr[46734] = 2118409593;
assign addr[46735] = 2121461578;
assign addr[46736] = 2124345343;
assign addr[46737] = 2127060661;
assign addr[46738] = 2129607316;
assign addr[46739] = 2131985106;
assign addr[46740] = 2134193842;
assign addr[46741] = 2136233350;
assign addr[46742] = 2138103468;
assign addr[46743] = 2139804048;
assign addr[46744] = 2141334954;
assign addr[46745] = 2142696065;
assign addr[46746] = 2143887273;
assign addr[46747] = 2144908484;
assign addr[46748] = 2145759618;
assign addr[46749] = 2146440605;
assign addr[46750] = 2146951393;
assign addr[46751] = 2147291941;
assign addr[46752] = 2147462221;
assign addr[46753] = 2147462221;
assign addr[46754] = 2147291941;
assign addr[46755] = 2146951393;
assign addr[46756] = 2146440605;
assign addr[46757] = 2145759618;
assign addr[46758] = 2144908484;
assign addr[46759] = 2143887273;
assign addr[46760] = 2142696065;
assign addr[46761] = 2141334954;
assign addr[46762] = 2139804048;
assign addr[46763] = 2138103468;
assign addr[46764] = 2136233350;
assign addr[46765] = 2134193842;
assign addr[46766] = 2131985106;
assign addr[46767] = 2129607316;
assign addr[46768] = 2127060661;
assign addr[46769] = 2124345343;
assign addr[46770] = 2121461578;
assign addr[46771] = 2118409593;
assign addr[46772] = 2115189632;
assign addr[46773] = 2111801949;
assign addr[46774] = 2108246813;
assign addr[46775] = 2104524506;
assign addr[46776] = 2100635323;
assign addr[46777] = 2096579573;
assign addr[46778] = 2092357577;
assign addr[46779] = 2087969669;
assign addr[46780] = 2083416198;
assign addr[46781] = 2078697525;
assign addr[46782] = 2073814024;
assign addr[46783] = 2068766083;
assign addr[46784] = 2063554100;
assign addr[46785] = 2058178491;
assign addr[46786] = 2052639680;
assign addr[46787] = 2046938108;
assign addr[46788] = 2041074226;
assign addr[46789] = 2035048499;
assign addr[46790] = 2028861406;
assign addr[46791] = 2022513436;
assign addr[46792] = 2016005093;
assign addr[46793] = 2009336893;
assign addr[46794] = 2002509365;
assign addr[46795] = 1995523051;
assign addr[46796] = 1988378503;
assign addr[46797] = 1981076290;
assign addr[46798] = 1973616989;
assign addr[46799] = 1966001192;
assign addr[46800] = 1958229503;
assign addr[46801] = 1950302539;
assign addr[46802] = 1942220928;
assign addr[46803] = 1933985310;
assign addr[46804] = 1925596340;
assign addr[46805] = 1917054681;
assign addr[46806] = 1908361011;
assign addr[46807] = 1899516021;
assign addr[46808] = 1890520410;
assign addr[46809] = 1881374892;
assign addr[46810] = 1872080193;
assign addr[46811] = 1862637049;
assign addr[46812] = 1853046210;
assign addr[46813] = 1843308435;
assign addr[46814] = 1833424497;
assign addr[46815] = 1823395180;
assign addr[46816] = 1813221279;
assign addr[46817] = 1802903601;
assign addr[46818] = 1792442963;
assign addr[46819] = 1781840195;
assign addr[46820] = 1771096139;
assign addr[46821] = 1760211645;
assign addr[46822] = 1749187577;
assign addr[46823] = 1738024810;
assign addr[46824] = 1726724227;
assign addr[46825] = 1715286726;
assign addr[46826] = 1703713213;
assign addr[46827] = 1692004606;
assign addr[46828] = 1680161834;
assign addr[46829] = 1668185835;
assign addr[46830] = 1656077559;
assign addr[46831] = 1643837966;
assign addr[46832] = 1631468027;
assign addr[46833] = 1618968722;
assign addr[46834] = 1606341043;
assign addr[46835] = 1593585992;
assign addr[46836] = 1580704578;
assign addr[46837] = 1567697824;
assign addr[46838] = 1554566762;
assign addr[46839] = 1541312431;
assign addr[46840] = 1527935884;
assign addr[46841] = 1514438181;
assign addr[46842] = 1500820393;
assign addr[46843] = 1487083598;
assign addr[46844] = 1473228887;
assign addr[46845] = 1459257358;
assign addr[46846] = 1445170118;
assign addr[46847] = 1430968286;
assign addr[46848] = 1416652986;
assign addr[46849] = 1402225355;
assign addr[46850] = 1387686535;
assign addr[46851] = 1373037681;
assign addr[46852] = 1358279953;
assign addr[46853] = 1343414522;
assign addr[46854] = 1328442566;
assign addr[46855] = 1313365273;
assign addr[46856] = 1298183838;
assign addr[46857] = 1282899464;
assign addr[46858] = 1267513365;
assign addr[46859] = 1252026760;
assign addr[46860] = 1236440877;
assign addr[46861] = 1220756951;
assign addr[46862] = 1204976227;
assign addr[46863] = 1189099956;
assign addr[46864] = 1173129396;
assign addr[46865] = 1157065814;
assign addr[46866] = 1140910484;
assign addr[46867] = 1124664687;
assign addr[46868] = 1108329711;
assign addr[46869] = 1091906851;
assign addr[46870] = 1075397409;
assign addr[46871] = 1058802695;
assign addr[46872] = 1042124025;
assign addr[46873] = 1025362720;
assign addr[46874] = 1008520110;
assign addr[46875] = 991597531;
assign addr[46876] = 974596324;
assign addr[46877] = 957517838;
assign addr[46878] = 940363427;
assign addr[46879] = 923134450;
assign addr[46880] = 905832274;
assign addr[46881] = 888458272;
assign addr[46882] = 871013820;
assign addr[46883] = 853500302;
assign addr[46884] = 835919107;
assign addr[46885] = 818271628;
assign addr[46886] = 800559266;
assign addr[46887] = 782783424;
assign addr[46888] = 764945512;
assign addr[46889] = 747046944;
assign addr[46890] = 729089140;
assign addr[46891] = 711073525;
assign addr[46892] = 693001525;
assign addr[46893] = 674874574;
assign addr[46894] = 656694110;
assign addr[46895] = 638461574;
assign addr[46896] = 620178412;
assign addr[46897] = 601846074;
assign addr[46898] = 583466013;
assign addr[46899] = 565039687;
assign addr[46900] = 546568556;
assign addr[46901] = 528054086;
assign addr[46902] = 509497745;
assign addr[46903] = 490901003;
assign addr[46904] = 472265336;
assign addr[46905] = 453592221;
assign addr[46906] = 434883140;
assign addr[46907] = 416139574;
assign addr[46908] = 397363011;
assign addr[46909] = 378554940;
assign addr[46910] = 359716852;
assign addr[46911] = 340850240;
assign addr[46912] = 321956601;
assign addr[46913] = 303037433;
assign addr[46914] = 284094236;
assign addr[46915] = 265128512;
assign addr[46916] = 246141764;
assign addr[46917] = 227135500;
assign addr[46918] = 208111224;
assign addr[46919] = 189070447;
assign addr[46920] = 170014678;
assign addr[46921] = 150945428;
assign addr[46922] = 131864208;
assign addr[46923] = 112772533;
assign addr[46924] = 93671915;
assign addr[46925] = 74563870;
assign addr[46926] = 55449912;
assign addr[46927] = 36331557;
assign addr[46928] = 17210322;
assign addr[46929] = -1912278;
assign addr[46930] = -21034727;
assign addr[46931] = -40155507;
assign addr[46932] = -59273104;
assign addr[46933] = -78386000;
assign addr[46934] = -97492681;
assign addr[46935] = -116591632;
assign addr[46936] = -135681337;
assign addr[46937] = -154760284;
assign addr[46938] = -173826959;
assign addr[46939] = -192879850;
assign addr[46940] = -211917448;
assign addr[46941] = -230938242;
assign addr[46942] = -249940723;
assign addr[46943] = -268923386;
assign addr[46944] = -287884725;
assign addr[46945] = -306823237;
assign addr[46946] = -325737419;
assign addr[46947] = -344625773;
assign addr[46948] = -363486799;
assign addr[46949] = -382319004;
assign addr[46950] = -401120892;
assign addr[46951] = -419890975;
assign addr[46952] = -438627762;
assign addr[46953] = -457329769;
assign addr[46954] = -475995513;
assign addr[46955] = -494623513;
assign addr[46956] = -513212292;
assign addr[46957] = -531760377;
assign addr[46958] = -550266296;
assign addr[46959] = -568728583;
assign addr[46960] = -587145773;
assign addr[46961] = -605516406;
assign addr[46962] = -623839025;
assign addr[46963] = -642112178;
assign addr[46964] = -660334415;
assign addr[46965] = -678504291;
assign addr[46966] = -696620367;
assign addr[46967] = -714681204;
assign addr[46968] = -732685372;
assign addr[46969] = -750631442;
assign addr[46970] = -768517992;
assign addr[46971] = -786343603;
assign addr[46972] = -804106861;
assign addr[46973] = -821806359;
assign addr[46974] = -839440693;
assign addr[46975] = -857008464;
assign addr[46976] = -874508280;
assign addr[46977] = -891938752;
assign addr[46978] = -909298500;
assign addr[46979] = -926586145;
assign addr[46980] = -943800318;
assign addr[46981] = -960939653;
assign addr[46982] = -978002791;
assign addr[46983] = -994988380;
assign addr[46984] = -1011895073;
assign addr[46985] = -1028721528;
assign addr[46986] = -1045466412;
assign addr[46987] = -1062128397;
assign addr[46988] = -1078706161;
assign addr[46989] = -1095198391;
assign addr[46990] = -1111603778;
assign addr[46991] = -1127921022;
assign addr[46992] = -1144148829;
assign addr[46993] = -1160285911;
assign addr[46994] = -1176330990;
assign addr[46995] = -1192282793;
assign addr[46996] = -1208140056;
assign addr[46997] = -1223901520;
assign addr[46998] = -1239565936;
assign addr[46999] = -1255132063;
assign addr[47000] = -1270598665;
assign addr[47001] = -1285964516;
assign addr[47002] = -1301228398;
assign addr[47003] = -1316389101;
assign addr[47004] = -1331445422;
assign addr[47005] = -1346396168;
assign addr[47006] = -1361240152;
assign addr[47007] = -1375976199;
assign addr[47008] = -1390603139;
assign addr[47009] = -1405119813;
assign addr[47010] = -1419525069;
assign addr[47011] = -1433817766;
assign addr[47012] = -1447996770;
assign addr[47013] = -1462060956;
assign addr[47014] = -1476009210;
assign addr[47015] = -1489840425;
assign addr[47016] = -1503553506;
assign addr[47017] = -1517147363;
assign addr[47018] = -1530620920;
assign addr[47019] = -1543973108;
assign addr[47020] = -1557202869;
assign addr[47021] = -1570309153;
assign addr[47022] = -1583290921;
assign addr[47023] = -1596147143;
assign addr[47024] = -1608876801;
assign addr[47025] = -1621478885;
assign addr[47026] = -1633952396;
assign addr[47027] = -1646296344;
assign addr[47028] = -1658509750;
assign addr[47029] = -1670591647;
assign addr[47030] = -1682541077;
assign addr[47031] = -1694357091;
assign addr[47032] = -1706038753;
assign addr[47033] = -1717585136;
assign addr[47034] = -1728995326;
assign addr[47035] = -1740268417;
assign addr[47036] = -1751403515;
assign addr[47037] = -1762399737;
assign addr[47038] = -1773256212;
assign addr[47039] = -1783972079;
assign addr[47040] = -1794546487;
assign addr[47041] = -1804978599;
assign addr[47042] = -1815267588;
assign addr[47043] = -1825412636;
assign addr[47044] = -1835412941;
assign addr[47045] = -1845267708;
assign addr[47046] = -1854976157;
assign addr[47047] = -1864537518;
assign addr[47048] = -1873951032;
assign addr[47049] = -1883215953;
assign addr[47050] = -1892331547;
assign addr[47051] = -1901297091;
assign addr[47052] = -1910111873;
assign addr[47053] = -1918775195;
assign addr[47054] = -1927286370;
assign addr[47055] = -1935644723;
assign addr[47056] = -1943849591;
assign addr[47057] = -1951900324;
assign addr[47058] = -1959796283;
assign addr[47059] = -1967536842;
assign addr[47060] = -1975121388;
assign addr[47061] = -1982549318;
assign addr[47062] = -1989820044;
assign addr[47063] = -1996932990;
assign addr[47064] = -2003887591;
assign addr[47065] = -2010683297;
assign addr[47066] = -2017319567;
assign addr[47067] = -2023795876;
assign addr[47068] = -2030111710;
assign addr[47069] = -2036266570;
assign addr[47070] = -2042259965;
assign addr[47071] = -2048091422;
assign addr[47072] = -2053760478;
assign addr[47073] = -2059266683;
assign addr[47074] = -2064609600;
assign addr[47075] = -2069788807;
assign addr[47076] = -2074803892;
assign addr[47077] = -2079654458;
assign addr[47078] = -2084340120;
assign addr[47079] = -2088860507;
assign addr[47080] = -2093215260;
assign addr[47081] = -2097404033;
assign addr[47082] = -2101426496;
assign addr[47083] = -2105282327;
assign addr[47084] = -2108971223;
assign addr[47085] = -2112492891;
assign addr[47086] = -2115847050;
assign addr[47087] = -2119033436;
assign addr[47088] = -2122051796;
assign addr[47089] = -2124901890;
assign addr[47090] = -2127583492;
assign addr[47091] = -2130096389;
assign addr[47092] = -2132440383;
assign addr[47093] = -2134615288;
assign addr[47094] = -2136620930;
assign addr[47095] = -2138457152;
assign addr[47096] = -2140123807;
assign addr[47097] = -2141620763;
assign addr[47098] = -2142947902;
assign addr[47099] = -2144105118;
assign addr[47100] = -2145092320;
assign addr[47101] = -2145909429;
assign addr[47102] = -2146556380;
assign addr[47103] = -2147033123;
assign addr[47104] = -2147339619;
assign addr[47105] = -2147475844;
assign addr[47106] = -2147441787;
assign addr[47107] = -2147237452;
assign addr[47108] = -2146862854;
assign addr[47109] = -2146318022;
assign addr[47110] = -2145603001;
assign addr[47111] = -2144717846;
assign addr[47112] = -2143662628;
assign addr[47113] = -2142437431;
assign addr[47114] = -2141042352;
assign addr[47115] = -2139477502;
assign addr[47116] = -2137743003;
assign addr[47117] = -2135838995;
assign addr[47118] = -2133765628;
assign addr[47119] = -2131523066;
assign addr[47120] = -2129111488;
assign addr[47121] = -2126531084;
assign addr[47122] = -2123782059;
assign addr[47123] = -2120864631;
assign addr[47124] = -2117779031;
assign addr[47125] = -2114525505;
assign addr[47126] = -2111104309;
assign addr[47127] = -2107515716;
assign addr[47128] = -2103760010;
assign addr[47129] = -2099837489;
assign addr[47130] = -2095748463;
assign addr[47131] = -2091493257;
assign addr[47132] = -2087072209;
assign addr[47133] = -2082485668;
assign addr[47134] = -2077733999;
assign addr[47135] = -2072817579;
assign addr[47136] = -2067736796;
assign addr[47137] = -2062492055;
assign addr[47138] = -2057083771;
assign addr[47139] = -2051512372;
assign addr[47140] = -2045778302;
assign addr[47141] = -2039882013;
assign addr[47142] = -2033823974;
assign addr[47143] = -2027604666;
assign addr[47144] = -2021224581;
assign addr[47145] = -2014684225;
assign addr[47146] = -2007984117;
assign addr[47147] = -2001124788;
assign addr[47148] = -1994106782;
assign addr[47149] = -1986930656;
assign addr[47150] = -1979596978;
assign addr[47151] = -1972106330;
assign addr[47152] = -1964459306;
assign addr[47153] = -1956656513;
assign addr[47154] = -1948698568;
assign addr[47155] = -1940586104;
assign addr[47156] = -1932319763;
assign addr[47157] = -1923900201;
assign addr[47158] = -1915328086;
assign addr[47159] = -1906604097;
assign addr[47160] = -1897728925;
assign addr[47161] = -1888703276;
assign addr[47162] = -1879527863;
assign addr[47163] = -1870203416;
assign addr[47164] = -1860730673;
assign addr[47165] = -1851110385;
assign addr[47166] = -1841343316;
assign addr[47167] = -1831430239;
assign addr[47168] = -1821371941;
assign addr[47169] = -1811169220;
assign addr[47170] = -1800822883;
assign addr[47171] = -1790333753;
assign addr[47172] = -1779702660;
assign addr[47173] = -1768930447;
assign addr[47174] = -1758017969;
assign addr[47175] = -1746966091;
assign addr[47176] = -1735775690;
assign addr[47177] = -1724447652;
assign addr[47178] = -1712982875;
assign addr[47179] = -1701382270;
assign addr[47180] = -1689646755;
assign addr[47181] = -1677777262;
assign addr[47182] = -1665774731;
assign addr[47183] = -1653640115;
assign addr[47184] = -1641374375;
assign addr[47185] = -1628978484;
assign addr[47186] = -1616453425;
assign addr[47187] = -1603800191;
assign addr[47188] = -1591019785;
assign addr[47189] = -1578113222;
assign addr[47190] = -1565081523;
assign addr[47191] = -1551925723;
assign addr[47192] = -1538646865;
assign addr[47193] = -1525246002;
assign addr[47194] = -1511724196;
assign addr[47195] = -1498082520;
assign addr[47196] = -1484322054;
assign addr[47197] = -1470443891;
assign addr[47198] = -1456449131;
assign addr[47199] = -1442338884;
assign addr[47200] = -1428114267;
assign addr[47201] = -1413776410;
assign addr[47202] = -1399326449;
assign addr[47203] = -1384765530;
assign addr[47204] = -1370094808;
assign addr[47205] = -1355315445;
assign addr[47206] = -1340428615;
assign addr[47207] = -1325435496;
assign addr[47208] = -1310337279;
assign addr[47209] = -1295135159;
assign addr[47210] = -1279830344;
assign addr[47211] = -1264424045;
assign addr[47212] = -1248917486;
assign addr[47213] = -1233311895;
assign addr[47214] = -1217608510;
assign addr[47215] = -1201808576;
assign addr[47216] = -1185913346;
assign addr[47217] = -1169924081;
assign addr[47218] = -1153842047;
assign addr[47219] = -1137668521;
assign addr[47220] = -1121404785;
assign addr[47221] = -1105052128;
assign addr[47222] = -1088611847;
assign addr[47223] = -1072085246;
assign addr[47224] = -1055473635;
assign addr[47225] = -1038778332;
assign addr[47226] = -1022000660;
assign addr[47227] = -1005141949;
assign addr[47228] = -988203537;
assign addr[47229] = -971186766;
assign addr[47230] = -954092986;
assign addr[47231] = -936923553;
assign addr[47232] = -919679827;
assign addr[47233] = -902363176;
assign addr[47234] = -884974973;
assign addr[47235] = -867516597;
assign addr[47236] = -849989433;
assign addr[47237] = -832394869;
assign addr[47238] = -814734301;
assign addr[47239] = -797009130;
assign addr[47240] = -779220762;
assign addr[47241] = -761370605;
assign addr[47242] = -743460077;
assign addr[47243] = -725490597;
assign addr[47244] = -707463589;
assign addr[47245] = -689380485;
assign addr[47246] = -671242716;
assign addr[47247] = -653051723;
assign addr[47248] = -634808946;
assign addr[47249] = -616515832;
assign addr[47250] = -598173833;
assign addr[47251] = -579784402;
assign addr[47252] = -561348998;
assign addr[47253] = -542869083;
assign addr[47254] = -524346121;
assign addr[47255] = -505781581;
assign addr[47256] = -487176937;
assign addr[47257] = -468533662;
assign addr[47258] = -449853235;
assign addr[47259] = -431137138;
assign addr[47260] = -412386854;
assign addr[47261] = -393603870;
assign addr[47262] = -374789676;
assign addr[47263] = -355945764;
assign addr[47264] = -337073627;
assign addr[47265] = -318174762;
assign addr[47266] = -299250668;
assign addr[47267] = -280302845;
assign addr[47268] = -261332796;
assign addr[47269] = -242342025;
assign addr[47270] = -223332037;
assign addr[47271] = -204304341;
assign addr[47272] = -185260444;
assign addr[47273] = -166201858;
assign addr[47274] = -147130093;
assign addr[47275] = -128046661;
assign addr[47276] = -108953076;
assign addr[47277] = -89850852;
assign addr[47278] = -70741503;
assign addr[47279] = -51626544;
assign addr[47280] = -32507492;
assign addr[47281] = -13385863;
assign addr[47282] = 5736829;
assign addr[47283] = 24859065;
assign addr[47284] = 43979330;
assign addr[47285] = 63096108;
assign addr[47286] = 82207882;
assign addr[47287] = 101313138;
assign addr[47288] = 120410361;
assign addr[47289] = 139498035;
assign addr[47290] = 158574649;
assign addr[47291] = 177638688;
assign addr[47292] = 196688642;
assign addr[47293] = 215722999;
assign addr[47294] = 234740251;
assign addr[47295] = 253738890;
assign addr[47296] = 272717408;
assign addr[47297] = 291674302;
assign addr[47298] = 310608068;
assign addr[47299] = 329517204;
assign addr[47300] = 348400212;
assign addr[47301] = 367255594;
assign addr[47302] = 386081854;
assign addr[47303] = 404877501;
assign addr[47304] = 423641043;
assign addr[47305] = 442370993;
assign addr[47306] = 461065866;
assign addr[47307] = 479724180;
assign addr[47308] = 498344454;
assign addr[47309] = 516925212;
assign addr[47310] = 535464981;
assign addr[47311] = 553962291;
assign addr[47312] = 572415676;
assign addr[47313] = 590823671;
assign addr[47314] = 609184818;
assign addr[47315] = 627497660;
assign addr[47316] = 645760745;
assign addr[47317] = 663972625;
assign addr[47318] = 682131857;
assign addr[47319] = 700236999;
assign addr[47320] = 718286617;
assign addr[47321] = 736279279;
assign addr[47322] = 754213559;
assign addr[47323] = 772088034;
assign addr[47324] = 789901288;
assign addr[47325] = 807651907;
assign addr[47326] = 825338484;
assign addr[47327] = 842959617;
assign addr[47328] = 860513908;
assign addr[47329] = 877999966;
assign addr[47330] = 895416404;
assign addr[47331] = 912761841;
assign addr[47332] = 930034901;
assign addr[47333] = 947234215;
assign addr[47334] = 964358420;
assign addr[47335] = 981406156;
assign addr[47336] = 998376073;
assign addr[47337] = 1015266825;
assign addr[47338] = 1032077073;
assign addr[47339] = 1048805483;
assign addr[47340] = 1065450729;
assign addr[47341] = 1082011492;
assign addr[47342] = 1098486458;
assign addr[47343] = 1114874320;
assign addr[47344] = 1131173780;
assign addr[47345] = 1147383544;
assign addr[47346] = 1163502328;
assign addr[47347] = 1179528853;
assign addr[47348] = 1195461849;
assign addr[47349] = 1211300053;
assign addr[47350] = 1227042207;
assign addr[47351] = 1242687064;
assign addr[47352] = 1258233384;
assign addr[47353] = 1273679934;
assign addr[47354] = 1289025489;
assign addr[47355] = 1304268832;
assign addr[47356] = 1319408754;
assign addr[47357] = 1334444055;
assign addr[47358] = 1349373543;
assign addr[47359] = 1364196034;
assign addr[47360] = 1378910353;
assign addr[47361] = 1393515332;
assign addr[47362] = 1408009814;
assign addr[47363] = 1422392650;
assign addr[47364] = 1436662698;
assign addr[47365] = 1450818828;
assign addr[47366] = 1464859917;
assign addr[47367] = 1478784851;
assign addr[47368] = 1492592527;
assign addr[47369] = 1506281850;
assign addr[47370] = 1519851733;
assign addr[47371] = 1533301101;
assign addr[47372] = 1546628888;
assign addr[47373] = 1559834037;
assign addr[47374] = 1572915501;
assign addr[47375] = 1585872242;
assign addr[47376] = 1598703233;
assign addr[47377] = 1611407456;
assign addr[47378] = 1623983905;
assign addr[47379] = 1636431582;
assign addr[47380] = 1648749499;
assign addr[47381] = 1660936681;
assign addr[47382] = 1672992161;
assign addr[47383] = 1684914983;
assign addr[47384] = 1696704201;
assign addr[47385] = 1708358881;
assign addr[47386] = 1719878099;
assign addr[47387] = 1731260941;
assign addr[47388] = 1742506504;
assign addr[47389] = 1753613897;
assign addr[47390] = 1764582240;
assign addr[47391] = 1775410662;
assign addr[47392] = 1786098304;
assign addr[47393] = 1796644320;
assign addr[47394] = 1807047873;
assign addr[47395] = 1817308138;
assign addr[47396] = 1827424302;
assign addr[47397] = 1837395562;
assign addr[47398] = 1847221128;
assign addr[47399] = 1856900221;
assign addr[47400] = 1866432072;
assign addr[47401] = 1875815927;
assign addr[47402] = 1885051042;
assign addr[47403] = 1894136683;
assign addr[47404] = 1903072131;
assign addr[47405] = 1911856677;
assign addr[47406] = 1920489624;
assign addr[47407] = 1928970288;
assign addr[47408] = 1937297997;
assign addr[47409] = 1945472089;
assign addr[47410] = 1953491918;
assign addr[47411] = 1961356847;
assign addr[47412] = 1969066252;
assign addr[47413] = 1976619522;
assign addr[47414] = 1984016058;
assign addr[47415] = 1991255274;
assign addr[47416] = 1998336596;
assign addr[47417] = 2005259462;
assign addr[47418] = 2012023322;
assign addr[47419] = 2018627642;
assign addr[47420] = 2025071897;
assign addr[47421] = 2031355576;
assign addr[47422] = 2037478181;
assign addr[47423] = 2043439226;
assign addr[47424] = 2049238240;
assign addr[47425] = 2054874761;
assign addr[47426] = 2060348343;
assign addr[47427] = 2065658552;
assign addr[47428] = 2070804967;
assign addr[47429] = 2075787180;
assign addr[47430] = 2080604795;
assign addr[47431] = 2085257431;
assign addr[47432] = 2089744719;
assign addr[47433] = 2094066304;
assign addr[47434] = 2098221841;
assign addr[47435] = 2102211002;
assign addr[47436] = 2106033471;
assign addr[47437] = 2109688944;
assign addr[47438] = 2113177132;
assign addr[47439] = 2116497758;
assign addr[47440] = 2119650558;
assign addr[47441] = 2122635283;
assign addr[47442] = 2125451696;
assign addr[47443] = 2128099574;
assign addr[47444] = 2130578706;
assign addr[47445] = 2132888897;
assign addr[47446] = 2135029962;
assign addr[47447] = 2137001733;
assign addr[47448] = 2138804053;
assign addr[47449] = 2140436778;
assign addr[47450] = 2141899780;
assign addr[47451] = 2143192942;
assign addr[47452] = 2144316162;
assign addr[47453] = 2145269351;
assign addr[47454] = 2146052433;
assign addr[47455] = 2146665347;
assign addr[47456] = 2147108043;
assign addr[47457] = 2147380486;
assign addr[47458] = 2147482655;
assign addr[47459] = 2147414542;
assign addr[47460] = 2147176152;
assign addr[47461] = 2146767505;
assign addr[47462] = 2146188631;
assign addr[47463] = 2145439578;
assign addr[47464] = 2144520405;
assign addr[47465] = 2143431184;
assign addr[47466] = 2142172003;
assign addr[47467] = 2140742960;
assign addr[47468] = 2139144169;
assign addr[47469] = 2137375758;
assign addr[47470] = 2135437865;
assign addr[47471] = 2133330646;
assign addr[47472] = 2131054266;
assign addr[47473] = 2128608907;
assign addr[47474] = 2125994762;
assign addr[47475] = 2123212038;
assign addr[47476] = 2120260957;
assign addr[47477] = 2117141752;
assign addr[47478] = 2113854671;
assign addr[47479] = 2110399974;
assign addr[47480] = 2106777935;
assign addr[47481] = 2102988841;
assign addr[47482] = 2099032994;
assign addr[47483] = 2094910706;
assign addr[47484] = 2090622304;
assign addr[47485] = 2086168128;
assign addr[47486] = 2081548533;
assign addr[47487] = 2076763883;
assign addr[47488] = 2071814558;
assign addr[47489] = 2066700952;
assign addr[47490] = 2061423468;
assign addr[47491] = 2055982526;
assign addr[47492] = 2050378558;
assign addr[47493] = 2044612007;
assign addr[47494] = 2038683330;
assign addr[47495] = 2032592999;
assign addr[47496] = 2026341495;
assign addr[47497] = 2019929315;
assign addr[47498] = 2013356967;
assign addr[47499] = 2006624971;
assign addr[47500] = 1999733863;
assign addr[47501] = 1992684188;
assign addr[47502] = 1985476506;
assign addr[47503] = 1978111387;
assign addr[47504] = 1970589416;
assign addr[47505] = 1962911189;
assign addr[47506] = 1955077316;
assign addr[47507] = 1947088417;
assign addr[47508] = 1938945125;
assign addr[47509] = 1930648088;
assign addr[47510] = 1922197961;
assign addr[47511] = 1913595416;
assign addr[47512] = 1904841135;
assign addr[47513] = 1895935811;
assign addr[47514] = 1886880151;
assign addr[47515] = 1877674873;
assign addr[47516] = 1868320707;
assign addr[47517] = 1858818395;
assign addr[47518] = 1849168689;
assign addr[47519] = 1839372356;
assign addr[47520] = 1829430172;
assign addr[47521] = 1819342925;
assign addr[47522] = 1809111415;
assign addr[47523] = 1798736454;
assign addr[47524] = 1788218865;
assign addr[47525] = 1777559480;
assign addr[47526] = 1766759146;
assign addr[47527] = 1755818718;
assign addr[47528] = 1744739065;
assign addr[47529] = 1733521064;
assign addr[47530] = 1722165606;
assign addr[47531] = 1710673591;
assign addr[47532] = 1699045930;
assign addr[47533] = 1687283545;
assign addr[47534] = 1675387369;
assign addr[47535] = 1663358344;
assign addr[47536] = 1651197426;
assign addr[47537] = 1638905577;
assign addr[47538] = 1626483774;
assign addr[47539] = 1613933000;
assign addr[47540] = 1601254251;
assign addr[47541] = 1588448533;
assign addr[47542] = 1575516860;
assign addr[47543] = 1562460258;
assign addr[47544] = 1549279763;
assign addr[47545] = 1535976419;
assign addr[47546] = 1522551282;
assign addr[47547] = 1509005416;
assign addr[47548] = 1495339895;
assign addr[47549] = 1481555802;
assign addr[47550] = 1467654232;
assign addr[47551] = 1453636285;
assign addr[47552] = 1439503074;
assign addr[47553] = 1425255719;
assign addr[47554] = 1410895350;
assign addr[47555] = 1396423105;
assign addr[47556] = 1381840133;
assign addr[47557] = 1367147589;
assign addr[47558] = 1352346639;
assign addr[47559] = 1337438456;
assign addr[47560] = 1322424222;
assign addr[47561] = 1307305128;
assign addr[47562] = 1292082373;
assign addr[47563] = 1276757164;
assign addr[47564] = 1261330715;
assign addr[47565] = 1245804251;
assign addr[47566] = 1230179002;
assign addr[47567] = 1214456207;
assign addr[47568] = 1198637114;
assign addr[47569] = 1182722976;
assign addr[47570] = 1166715055;
assign addr[47571] = 1150614620;
assign addr[47572] = 1134422949;
assign addr[47573] = 1118141326;
assign addr[47574] = 1101771040;
assign addr[47575] = 1085313391;
assign addr[47576] = 1068769683;
assign addr[47577] = 1052141228;
assign addr[47578] = 1035429345;
assign addr[47579] = 1018635358;
assign addr[47580] = 1001760600;
assign addr[47581] = 984806408;
assign addr[47582] = 967774128;
assign addr[47583] = 950665109;
assign addr[47584] = 933480707;
assign addr[47585] = 916222287;
assign addr[47586] = 898891215;
assign addr[47587] = 881488868;
assign addr[47588] = 864016623;
assign addr[47589] = 846475867;
assign addr[47590] = 828867991;
assign addr[47591] = 811194391;
assign addr[47592] = 793456467;
assign addr[47593] = 775655628;
assign addr[47594] = 757793284;
assign addr[47595] = 739870851;
assign addr[47596] = 721889752;
assign addr[47597] = 703851410;
assign addr[47598] = 685757258;
assign addr[47599] = 667608730;
assign addr[47600] = 649407264;
assign addr[47601] = 631154304;
assign addr[47602] = 612851297;
assign addr[47603] = 594499695;
assign addr[47604] = 576100953;
assign addr[47605] = 557656529;
assign addr[47606] = 539167887;
assign addr[47607] = 520636492;
assign addr[47608] = 502063814;
assign addr[47609] = 483451325;
assign addr[47610] = 464800501;
assign addr[47611] = 446112822;
assign addr[47612] = 427389768;
assign addr[47613] = 408632825;
assign addr[47614] = 389843480;
assign addr[47615] = 371023223;
assign addr[47616] = 352173546;
assign addr[47617] = 333295944;
assign addr[47618] = 314391913;
assign addr[47619] = 295462954;
assign addr[47620] = 276510565;
assign addr[47621] = 257536251;
assign addr[47622] = 238541516;
assign addr[47623] = 219527866;
assign addr[47624] = 200496809;
assign addr[47625] = 181449854;
assign addr[47626] = 162388511;
assign addr[47627] = 143314291;
assign addr[47628] = 124228708;
assign addr[47629] = 105133274;
assign addr[47630] = 86029503;
assign addr[47631] = 66918911;
assign addr[47632] = 47803013;
assign addr[47633] = 28683324;
assign addr[47634] = 9561361;
assign addr[47635] = -9561361;
assign addr[47636] = -28683324;
assign addr[47637] = -47803013;
assign addr[47638] = -66918911;
assign addr[47639] = -86029503;
assign addr[47640] = -105133274;
assign addr[47641] = -124228708;
assign addr[47642] = -143314291;
assign addr[47643] = -162388511;
assign addr[47644] = -181449854;
assign addr[47645] = -200496809;
assign addr[47646] = -219527866;
assign addr[47647] = -238541516;
assign addr[47648] = -257536251;
assign addr[47649] = -276510565;
assign addr[47650] = -295462953;
assign addr[47651] = -314391913;
assign addr[47652] = -333295944;
assign addr[47653] = -352173546;
assign addr[47654] = -371023223;
assign addr[47655] = -389843480;
assign addr[47656] = -408632825;
assign addr[47657] = -427389768;
assign addr[47658] = -446112822;
assign addr[47659] = -464800501;
assign addr[47660] = -483451325;
assign addr[47661] = -502063814;
assign addr[47662] = -520636492;
assign addr[47663] = -539167887;
assign addr[47664] = -557656529;
assign addr[47665] = -576100953;
assign addr[47666] = -594499695;
assign addr[47667] = -612851297;
assign addr[47668] = -631154304;
assign addr[47669] = -649407264;
assign addr[47670] = -667608730;
assign addr[47671] = -685757258;
assign addr[47672] = -703851410;
assign addr[47673] = -721889752;
assign addr[47674] = -739870851;
assign addr[47675] = -757793284;
assign addr[47676] = -775655628;
assign addr[47677] = -793456467;
assign addr[47678] = -811194391;
assign addr[47679] = -828867991;
assign addr[47680] = -846475867;
assign addr[47681] = -864016623;
assign addr[47682] = -881488868;
assign addr[47683] = -898891215;
assign addr[47684] = -916222287;
assign addr[47685] = -933480707;
assign addr[47686] = -950665109;
assign addr[47687] = -967774128;
assign addr[47688] = -984806408;
assign addr[47689] = -1001760600;
assign addr[47690] = -1018635358;
assign addr[47691] = -1035429345;
assign addr[47692] = -1052141228;
assign addr[47693] = -1068769683;
assign addr[47694] = -1085313391;
assign addr[47695] = -1101771040;
assign addr[47696] = -1118141326;
assign addr[47697] = -1134422949;
assign addr[47698] = -1150614620;
assign addr[47699] = -1166715055;
assign addr[47700] = -1182722976;
assign addr[47701] = -1198637114;
assign addr[47702] = -1214456207;
assign addr[47703] = -1230179002;
assign addr[47704] = -1245804251;
assign addr[47705] = -1261330715;
assign addr[47706] = -1276757164;
assign addr[47707] = -1292082373;
assign addr[47708] = -1307305128;
assign addr[47709] = -1322424222;
assign addr[47710] = -1337438456;
assign addr[47711] = -1352346639;
assign addr[47712] = -1367147589;
assign addr[47713] = -1381840133;
assign addr[47714] = -1396423105;
assign addr[47715] = -1410895350;
assign addr[47716] = -1425255719;
assign addr[47717] = -1439503074;
assign addr[47718] = -1453636285;
assign addr[47719] = -1467654232;
assign addr[47720] = -1481555802;
assign addr[47721] = -1495339895;
assign addr[47722] = -1509005416;
assign addr[47723] = -1522551282;
assign addr[47724] = -1535976419;
assign addr[47725] = -1549279763;
assign addr[47726] = -1562460258;
assign addr[47727] = -1575516860;
assign addr[47728] = -1588448533;
assign addr[47729] = -1601254251;
assign addr[47730] = -1613933000;
assign addr[47731] = -1626483774;
assign addr[47732] = -1638905577;
assign addr[47733] = -1651197426;
assign addr[47734] = -1663358344;
assign addr[47735] = -1675387369;
assign addr[47736] = -1687283545;
assign addr[47737] = -1699045930;
assign addr[47738] = -1710673591;
assign addr[47739] = -1722165606;
assign addr[47740] = -1733521064;
assign addr[47741] = -1744739065;
assign addr[47742] = -1755818718;
assign addr[47743] = -1766759146;
assign addr[47744] = -1777559480;
assign addr[47745] = -1788218865;
assign addr[47746] = -1798736454;
assign addr[47747] = -1809111415;
assign addr[47748] = -1819342925;
assign addr[47749] = -1829430172;
assign addr[47750] = -1839372356;
assign addr[47751] = -1849168689;
assign addr[47752] = -1858818395;
assign addr[47753] = -1868320707;
assign addr[47754] = -1877674873;
assign addr[47755] = -1886880151;
assign addr[47756] = -1895935811;
assign addr[47757] = -1904841135;
assign addr[47758] = -1913595416;
assign addr[47759] = -1922197961;
assign addr[47760] = -1930648088;
assign addr[47761] = -1938945125;
assign addr[47762] = -1947088417;
assign addr[47763] = -1955077316;
assign addr[47764] = -1962911189;
assign addr[47765] = -1970589416;
assign addr[47766] = -1978111387;
assign addr[47767] = -1985476506;
assign addr[47768] = -1992684188;
assign addr[47769] = -1999733863;
assign addr[47770] = -2006624971;
assign addr[47771] = -2013356967;
assign addr[47772] = -2019929315;
assign addr[47773] = -2026341495;
assign addr[47774] = -2032592999;
assign addr[47775] = -2038683330;
assign addr[47776] = -2044612007;
assign addr[47777] = -2050378558;
assign addr[47778] = -2055982526;
assign addr[47779] = -2061423468;
assign addr[47780] = -2066700952;
assign addr[47781] = -2071814558;
assign addr[47782] = -2076763883;
assign addr[47783] = -2081548533;
assign addr[47784] = -2086168128;
assign addr[47785] = -2090622304;
assign addr[47786] = -2094910706;
assign addr[47787] = -2099032994;
assign addr[47788] = -2102988841;
assign addr[47789] = -2106777935;
assign addr[47790] = -2110399974;
assign addr[47791] = -2113854671;
assign addr[47792] = -2117141752;
assign addr[47793] = -2120260957;
assign addr[47794] = -2123212038;
assign addr[47795] = -2125994762;
assign addr[47796] = -2128608907;
assign addr[47797] = -2131054266;
assign addr[47798] = -2133330646;
assign addr[47799] = -2135437865;
assign addr[47800] = -2137375758;
assign addr[47801] = -2139144169;
assign addr[47802] = -2140742960;
assign addr[47803] = -2142172003;
assign addr[47804] = -2143431184;
assign addr[47805] = -2144520405;
assign addr[47806] = -2145439578;
assign addr[47807] = -2146188631;
assign addr[47808] = -2146767505;
assign addr[47809] = -2147176152;
assign addr[47810] = -2147414542;
assign addr[47811] = -2147482655;
assign addr[47812] = -2147380486;
assign addr[47813] = -2147108043;
assign addr[47814] = -2146665347;
assign addr[47815] = -2146052433;
assign addr[47816] = -2145269351;
assign addr[47817] = -2144316162;
assign addr[47818] = -2143192942;
assign addr[47819] = -2141899780;
assign addr[47820] = -2140436778;
assign addr[47821] = -2138804053;
assign addr[47822] = -2137001733;
assign addr[47823] = -2135029962;
assign addr[47824] = -2132888897;
assign addr[47825] = -2130578706;
assign addr[47826] = -2128099574;
assign addr[47827] = -2125451696;
assign addr[47828] = -2122635283;
assign addr[47829] = -2119650558;
assign addr[47830] = -2116497758;
assign addr[47831] = -2113177132;
assign addr[47832] = -2109688944;
assign addr[47833] = -2106033471;
assign addr[47834] = -2102211002;
assign addr[47835] = -2098221841;
assign addr[47836] = -2094066304;
assign addr[47837] = -2089744719;
assign addr[47838] = -2085257431;
assign addr[47839] = -2080604795;
assign addr[47840] = -2075787180;
assign addr[47841] = -2070804967;
assign addr[47842] = -2065658552;
assign addr[47843] = -2060348343;
assign addr[47844] = -2054874761;
assign addr[47845] = -2049238240;
assign addr[47846] = -2043439226;
assign addr[47847] = -2037478181;
assign addr[47848] = -2031355576;
assign addr[47849] = -2025071897;
assign addr[47850] = -2018627642;
assign addr[47851] = -2012023322;
assign addr[47852] = -2005259462;
assign addr[47853] = -1998336596;
assign addr[47854] = -1991255274;
assign addr[47855] = -1984016058;
assign addr[47856] = -1976619522;
assign addr[47857] = -1969066252;
assign addr[47858] = -1961356847;
assign addr[47859] = -1953491918;
assign addr[47860] = -1945472089;
assign addr[47861] = -1937297997;
assign addr[47862] = -1928970288;
assign addr[47863] = -1920489624;
assign addr[47864] = -1911856677;
assign addr[47865] = -1903072131;
assign addr[47866] = -1894136683;
assign addr[47867] = -1885051042;
assign addr[47868] = -1875815927;
assign addr[47869] = -1866432072;
assign addr[47870] = -1856900221;
assign addr[47871] = -1847221128;
assign addr[47872] = -1837395562;
assign addr[47873] = -1827424302;
assign addr[47874] = -1817308138;
assign addr[47875] = -1807047873;
assign addr[47876] = -1796644320;
assign addr[47877] = -1786098304;
assign addr[47878] = -1775410662;
assign addr[47879] = -1764582240;
assign addr[47880] = -1753613897;
assign addr[47881] = -1742506504;
assign addr[47882] = -1731260941;
assign addr[47883] = -1719878099;
assign addr[47884] = -1708358881;
assign addr[47885] = -1696704201;
assign addr[47886] = -1684914983;
assign addr[47887] = -1672992161;
assign addr[47888] = -1660936681;
assign addr[47889] = -1648749499;
assign addr[47890] = -1636431582;
assign addr[47891] = -1623983905;
assign addr[47892] = -1611407456;
assign addr[47893] = -1598703233;
assign addr[47894] = -1585872242;
assign addr[47895] = -1572915501;
assign addr[47896] = -1559834037;
assign addr[47897] = -1546628888;
assign addr[47898] = -1533301101;
assign addr[47899] = -1519851733;
assign addr[47900] = -1506281850;
assign addr[47901] = -1492592527;
assign addr[47902] = -1478784851;
assign addr[47903] = -1464859917;
assign addr[47904] = -1450818828;
assign addr[47905] = -1436662698;
assign addr[47906] = -1422392650;
assign addr[47907] = -1408009814;
assign addr[47908] = -1393515332;
assign addr[47909] = -1378910353;
assign addr[47910] = -1364196034;
assign addr[47911] = -1349373543;
assign addr[47912] = -1334444055;
assign addr[47913] = -1319408754;
assign addr[47914] = -1304268832;
assign addr[47915] = -1289025489;
assign addr[47916] = -1273679934;
assign addr[47917] = -1258233384;
assign addr[47918] = -1242687064;
assign addr[47919] = -1227042207;
assign addr[47920] = -1211300053;
assign addr[47921] = -1195461849;
assign addr[47922] = -1179528853;
assign addr[47923] = -1163502328;
assign addr[47924] = -1147383544;
assign addr[47925] = -1131173780;
assign addr[47926] = -1114874320;
assign addr[47927] = -1098486458;
assign addr[47928] = -1082011492;
assign addr[47929] = -1065450729;
assign addr[47930] = -1048805483;
assign addr[47931] = -1032077073;
assign addr[47932] = -1015266825;
assign addr[47933] = -998376073;
assign addr[47934] = -981406156;
assign addr[47935] = -964358420;
assign addr[47936] = -947234215;
assign addr[47937] = -930034901;
assign addr[47938] = -912761841;
assign addr[47939] = -895416404;
assign addr[47940] = -877999966;
assign addr[47941] = -860513908;
assign addr[47942] = -842959617;
assign addr[47943] = -825338484;
assign addr[47944] = -807651907;
assign addr[47945] = -789901288;
assign addr[47946] = -772088034;
assign addr[47947] = -754213559;
assign addr[47948] = -736279279;
assign addr[47949] = -718286617;
assign addr[47950] = -700236999;
assign addr[47951] = -682131857;
assign addr[47952] = -663972625;
assign addr[47953] = -645760745;
assign addr[47954] = -627497660;
assign addr[47955] = -609184818;
assign addr[47956] = -590823671;
assign addr[47957] = -572415676;
assign addr[47958] = -553962291;
assign addr[47959] = -535464981;
assign addr[47960] = -516925212;
assign addr[47961] = -498344454;
assign addr[47962] = -479724180;
assign addr[47963] = -461065866;
assign addr[47964] = -442370993;
assign addr[47965] = -423641043;
assign addr[47966] = -404877501;
assign addr[47967] = -386081854;
assign addr[47968] = -367255594;
assign addr[47969] = -348400212;
assign addr[47970] = -329517204;
assign addr[47971] = -310608068;
assign addr[47972] = -291674302;
assign addr[47973] = -272717408;
assign addr[47974] = -253738890;
assign addr[47975] = -234740251;
assign addr[47976] = -215722999;
assign addr[47977] = -196688642;
assign addr[47978] = -177638688;
assign addr[47979] = -158574649;
assign addr[47980] = -139498035;
assign addr[47981] = -120410361;
assign addr[47982] = -101313138;
assign addr[47983] = -82207882;
assign addr[47984] = -63096108;
assign addr[47985] = -43979330;
assign addr[47986] = -24859065;
assign addr[47987] = -5736829;
assign addr[47988] = 13385863;
assign addr[47989] = 32507492;
assign addr[47990] = 51626544;
assign addr[47991] = 70741503;
assign addr[47992] = 89850852;
assign addr[47993] = 108953076;
assign addr[47994] = 128046661;
assign addr[47995] = 147130093;
assign addr[47996] = 166201858;
assign addr[47997] = 185260444;
assign addr[47998] = 204304341;
assign addr[47999] = 223332037;
assign addr[48000] = 242342025;
assign addr[48001] = 261332796;
assign addr[48002] = 280302845;
assign addr[48003] = 299250668;
assign addr[48004] = 318174762;
assign addr[48005] = 337073627;
assign addr[48006] = 355945764;
assign addr[48007] = 374789676;
assign addr[48008] = 393603870;
assign addr[48009] = 412386854;
assign addr[48010] = 431137138;
assign addr[48011] = 449853235;
assign addr[48012] = 468533662;
assign addr[48013] = 487176937;
assign addr[48014] = 505781581;
assign addr[48015] = 524346121;
assign addr[48016] = 542869083;
assign addr[48017] = 561348998;
assign addr[48018] = 579784402;
assign addr[48019] = 598173833;
assign addr[48020] = 616515832;
assign addr[48021] = 634808946;
assign addr[48022] = 653051723;
assign addr[48023] = 671242716;
assign addr[48024] = 689380485;
assign addr[48025] = 707463589;
assign addr[48026] = 725490597;
assign addr[48027] = 743460077;
assign addr[48028] = 761370605;
assign addr[48029] = 779220762;
assign addr[48030] = 797009130;
assign addr[48031] = 814734301;
assign addr[48032] = 832394869;
assign addr[48033] = 849989433;
assign addr[48034] = 867516597;
assign addr[48035] = 884974973;
assign addr[48036] = 902363176;
assign addr[48037] = 919679827;
assign addr[48038] = 936923553;
assign addr[48039] = 954092986;
assign addr[48040] = 971186766;
assign addr[48041] = 988203537;
assign addr[48042] = 1005141949;
assign addr[48043] = 1022000660;
assign addr[48044] = 1038778332;
assign addr[48045] = 1055473635;
assign addr[48046] = 1072085246;
assign addr[48047] = 1088611847;
assign addr[48048] = 1105052128;
assign addr[48049] = 1121404785;
assign addr[48050] = 1137668521;
assign addr[48051] = 1153842047;
assign addr[48052] = 1169924081;
assign addr[48053] = 1185913346;
assign addr[48054] = 1201808576;
assign addr[48055] = 1217608510;
assign addr[48056] = 1233311895;
assign addr[48057] = 1248917486;
assign addr[48058] = 1264424045;
assign addr[48059] = 1279830344;
assign addr[48060] = 1295135159;
assign addr[48061] = 1310337279;
assign addr[48062] = 1325435496;
assign addr[48063] = 1340428615;
assign addr[48064] = 1355315445;
assign addr[48065] = 1370094808;
assign addr[48066] = 1384765530;
assign addr[48067] = 1399326449;
assign addr[48068] = 1413776410;
assign addr[48069] = 1428114267;
assign addr[48070] = 1442338884;
assign addr[48071] = 1456449131;
assign addr[48072] = 1470443891;
assign addr[48073] = 1484322054;
assign addr[48074] = 1498082520;
assign addr[48075] = 1511724196;
assign addr[48076] = 1525246002;
assign addr[48077] = 1538646865;
assign addr[48078] = 1551925723;
assign addr[48079] = 1565081523;
assign addr[48080] = 1578113222;
assign addr[48081] = 1591019785;
assign addr[48082] = 1603800191;
assign addr[48083] = 1616453425;
assign addr[48084] = 1628978484;
assign addr[48085] = 1641374375;
assign addr[48086] = 1653640115;
assign addr[48087] = 1665774731;
assign addr[48088] = 1677777262;
assign addr[48089] = 1689646755;
assign addr[48090] = 1701382270;
assign addr[48091] = 1712982875;
assign addr[48092] = 1724447652;
assign addr[48093] = 1735775690;
assign addr[48094] = 1746966091;
assign addr[48095] = 1758017969;
assign addr[48096] = 1768930447;
assign addr[48097] = 1779702660;
assign addr[48098] = 1790333753;
assign addr[48099] = 1800822883;
assign addr[48100] = 1811169220;
assign addr[48101] = 1821371941;
assign addr[48102] = 1831430239;
assign addr[48103] = 1841343316;
assign addr[48104] = 1851110385;
assign addr[48105] = 1860730673;
assign addr[48106] = 1870203416;
assign addr[48107] = 1879527863;
assign addr[48108] = 1888703276;
assign addr[48109] = 1897728925;
assign addr[48110] = 1906604097;
assign addr[48111] = 1915328086;
assign addr[48112] = 1923900201;
assign addr[48113] = 1932319763;
assign addr[48114] = 1940586104;
assign addr[48115] = 1948698568;
assign addr[48116] = 1956656513;
assign addr[48117] = 1964459306;
assign addr[48118] = 1972106330;
assign addr[48119] = 1979596978;
assign addr[48120] = 1986930656;
assign addr[48121] = 1994106782;
assign addr[48122] = 2001124788;
assign addr[48123] = 2007984117;
assign addr[48124] = 2014684225;
assign addr[48125] = 2021224581;
assign addr[48126] = 2027604666;
assign addr[48127] = 2033823974;
assign addr[48128] = 2039882013;
assign addr[48129] = 2045778302;
assign addr[48130] = 2051512372;
assign addr[48131] = 2057083771;
assign addr[48132] = 2062492055;
assign addr[48133] = 2067736796;
assign addr[48134] = 2072817579;
assign addr[48135] = 2077733999;
assign addr[48136] = 2082485668;
assign addr[48137] = 2087072209;
assign addr[48138] = 2091493257;
assign addr[48139] = 2095748463;
assign addr[48140] = 2099837489;
assign addr[48141] = 2103760010;
assign addr[48142] = 2107515716;
assign addr[48143] = 2111104309;
assign addr[48144] = 2114525505;
assign addr[48145] = 2117779031;
assign addr[48146] = 2120864631;
assign addr[48147] = 2123782059;
assign addr[48148] = 2126531084;
assign addr[48149] = 2129111488;
assign addr[48150] = 2131523066;
assign addr[48151] = 2133765628;
assign addr[48152] = 2135838995;
assign addr[48153] = 2137743003;
assign addr[48154] = 2139477502;
assign addr[48155] = 2141042352;
assign addr[48156] = 2142437431;
assign addr[48157] = 2143662628;
assign addr[48158] = 2144717846;
assign addr[48159] = 2145603001;
assign addr[48160] = 2146318022;
assign addr[48161] = 2146862854;
assign addr[48162] = 2147237452;
assign addr[48163] = 2147441787;
assign addr[48164] = 2147475844;
assign addr[48165] = 2147339619;
assign addr[48166] = 2147033123;
assign addr[48167] = 2146556380;
assign addr[48168] = 2145909429;
assign addr[48169] = 2145092320;
assign addr[48170] = 2144105118;
assign addr[48171] = 2142947902;
assign addr[48172] = 2141620763;
assign addr[48173] = 2140123807;
assign addr[48174] = 2138457152;
assign addr[48175] = 2136620930;
assign addr[48176] = 2134615288;
assign addr[48177] = 2132440383;
assign addr[48178] = 2130096389;
assign addr[48179] = 2127583492;
assign addr[48180] = 2124901890;
assign addr[48181] = 2122051796;
assign addr[48182] = 2119033436;
assign addr[48183] = 2115847050;
assign addr[48184] = 2112492891;
assign addr[48185] = 2108971223;
assign addr[48186] = 2105282327;
assign addr[48187] = 2101426496;
assign addr[48188] = 2097404033;
assign addr[48189] = 2093215260;
assign addr[48190] = 2088860507;
assign addr[48191] = 2084340120;
assign addr[48192] = 2079654458;
assign addr[48193] = 2074803892;
assign addr[48194] = 2069788807;
assign addr[48195] = 2064609600;
assign addr[48196] = 2059266683;
assign addr[48197] = 2053760478;
assign addr[48198] = 2048091422;
assign addr[48199] = 2042259965;
assign addr[48200] = 2036266570;
assign addr[48201] = 2030111710;
assign addr[48202] = 2023795876;
assign addr[48203] = 2017319567;
assign addr[48204] = 2010683297;
assign addr[48205] = 2003887591;
assign addr[48206] = 1996932990;
assign addr[48207] = 1989820044;
assign addr[48208] = 1982549318;
assign addr[48209] = 1975121388;
assign addr[48210] = 1967536842;
assign addr[48211] = 1959796283;
assign addr[48212] = 1951900324;
assign addr[48213] = 1943849591;
assign addr[48214] = 1935644723;
assign addr[48215] = 1927286370;
assign addr[48216] = 1918775195;
assign addr[48217] = 1910111873;
assign addr[48218] = 1901297091;
assign addr[48219] = 1892331547;
assign addr[48220] = 1883215953;
assign addr[48221] = 1873951032;
assign addr[48222] = 1864537518;
assign addr[48223] = 1854976157;
assign addr[48224] = 1845267708;
assign addr[48225] = 1835412941;
assign addr[48226] = 1825412636;
assign addr[48227] = 1815267588;
assign addr[48228] = 1804978599;
assign addr[48229] = 1794546487;
assign addr[48230] = 1783972079;
assign addr[48231] = 1773256212;
assign addr[48232] = 1762399737;
assign addr[48233] = 1751403515;
assign addr[48234] = 1740268417;
assign addr[48235] = 1728995326;
assign addr[48236] = 1717585136;
assign addr[48237] = 1706038753;
assign addr[48238] = 1694357091;
assign addr[48239] = 1682541077;
assign addr[48240] = 1670591647;
assign addr[48241] = 1658509750;
assign addr[48242] = 1646296344;
assign addr[48243] = 1633952396;
assign addr[48244] = 1621478885;
assign addr[48245] = 1608876801;
assign addr[48246] = 1596147143;
assign addr[48247] = 1583290921;
assign addr[48248] = 1570309153;
assign addr[48249] = 1557202869;
assign addr[48250] = 1543973108;
assign addr[48251] = 1530620920;
assign addr[48252] = 1517147363;
assign addr[48253] = 1503553506;
assign addr[48254] = 1489840425;
assign addr[48255] = 1476009210;
assign addr[48256] = 1462060956;
assign addr[48257] = 1447996770;
assign addr[48258] = 1433817766;
assign addr[48259] = 1419525069;
assign addr[48260] = 1405119813;
assign addr[48261] = 1390603139;
assign addr[48262] = 1375976199;
assign addr[48263] = 1361240152;
assign addr[48264] = 1346396168;
assign addr[48265] = 1331445422;
assign addr[48266] = 1316389101;
assign addr[48267] = 1301228398;
assign addr[48268] = 1285964516;
assign addr[48269] = 1270598665;
assign addr[48270] = 1255132063;
assign addr[48271] = 1239565936;
assign addr[48272] = 1223901520;
assign addr[48273] = 1208140056;
assign addr[48274] = 1192282793;
assign addr[48275] = 1176330990;
assign addr[48276] = 1160285911;
assign addr[48277] = 1144148829;
assign addr[48278] = 1127921022;
assign addr[48279] = 1111603778;
assign addr[48280] = 1095198391;
assign addr[48281] = 1078706161;
assign addr[48282] = 1062128397;
assign addr[48283] = 1045466412;
assign addr[48284] = 1028721528;
assign addr[48285] = 1011895073;
assign addr[48286] = 994988380;
assign addr[48287] = 978002791;
assign addr[48288] = 960939653;
assign addr[48289] = 943800318;
assign addr[48290] = 926586145;
assign addr[48291] = 909298500;
assign addr[48292] = 891938752;
assign addr[48293] = 874508280;
assign addr[48294] = 857008464;
assign addr[48295] = 839440693;
assign addr[48296] = 821806359;
assign addr[48297] = 804106861;
assign addr[48298] = 786343603;
assign addr[48299] = 768517992;
assign addr[48300] = 750631442;
assign addr[48301] = 732685372;
assign addr[48302] = 714681204;
assign addr[48303] = 696620367;
assign addr[48304] = 678504291;
assign addr[48305] = 660334415;
assign addr[48306] = 642112178;
assign addr[48307] = 623839025;
assign addr[48308] = 605516406;
assign addr[48309] = 587145773;
assign addr[48310] = 568728583;
assign addr[48311] = 550266296;
assign addr[48312] = 531760377;
assign addr[48313] = 513212292;
assign addr[48314] = 494623513;
assign addr[48315] = 475995513;
assign addr[48316] = 457329769;
assign addr[48317] = 438627762;
assign addr[48318] = 419890975;
assign addr[48319] = 401120892;
assign addr[48320] = 382319004;
assign addr[48321] = 363486799;
assign addr[48322] = 344625773;
assign addr[48323] = 325737419;
assign addr[48324] = 306823237;
assign addr[48325] = 287884725;
assign addr[48326] = 268923386;
assign addr[48327] = 249940723;
assign addr[48328] = 230938242;
assign addr[48329] = 211917448;
assign addr[48330] = 192879850;
assign addr[48331] = 173826959;
assign addr[48332] = 154760284;
assign addr[48333] = 135681337;
assign addr[48334] = 116591632;
assign addr[48335] = 97492681;
assign addr[48336] = 78386000;
assign addr[48337] = 59273104;
assign addr[48338] = 40155507;
assign addr[48339] = 21034727;
assign addr[48340] = 1912278;
assign addr[48341] = -17210322;
assign addr[48342] = -36331557;
assign addr[48343] = -55449912;
assign addr[48344] = -74563870;
assign addr[48345] = -93671915;
assign addr[48346] = -112772533;
assign addr[48347] = -131864208;
assign addr[48348] = -150945428;
assign addr[48349] = -170014678;
assign addr[48350] = -189070447;
assign addr[48351] = -208111224;
assign addr[48352] = -227135500;
assign addr[48353] = -246141764;
assign addr[48354] = -265128512;
assign addr[48355] = -284094236;
assign addr[48356] = -303037433;
assign addr[48357] = -321956601;
assign addr[48358] = -340850240;
assign addr[48359] = -359716852;
assign addr[48360] = -378554940;
assign addr[48361] = -397363011;
assign addr[48362] = -416139574;
assign addr[48363] = -434883140;
assign addr[48364] = -453592221;
assign addr[48365] = -472265336;
assign addr[48366] = -490901003;
assign addr[48367] = -509497745;
assign addr[48368] = -528054086;
assign addr[48369] = -546568556;
assign addr[48370] = -565039687;
assign addr[48371] = -583466013;
assign addr[48372] = -601846074;
assign addr[48373] = -620178412;
assign addr[48374] = -638461574;
assign addr[48375] = -656694110;
assign addr[48376] = -674874574;
assign addr[48377] = -693001525;
assign addr[48378] = -711073524;
assign addr[48379] = -729089140;
assign addr[48380] = -747046944;
assign addr[48381] = -764945512;
assign addr[48382] = -782783424;
assign addr[48383] = -800559266;
assign addr[48384] = -818271628;
assign addr[48385] = -835919107;
assign addr[48386] = -853500302;
assign addr[48387] = -871013820;
assign addr[48388] = -888458272;
assign addr[48389] = -905832274;
assign addr[48390] = -923134450;
assign addr[48391] = -940363427;
assign addr[48392] = -957517838;
assign addr[48393] = -974596324;
assign addr[48394] = -991597531;
assign addr[48395] = -1008520110;
assign addr[48396] = -1025362720;
assign addr[48397] = -1042124025;
assign addr[48398] = -1058802695;
assign addr[48399] = -1075397409;
assign addr[48400] = -1091906851;
assign addr[48401] = -1108329711;
assign addr[48402] = -1124664687;
assign addr[48403] = -1140910484;
assign addr[48404] = -1157065814;
assign addr[48405] = -1173129396;
assign addr[48406] = -1189099956;
assign addr[48407] = -1204976227;
assign addr[48408] = -1220756951;
assign addr[48409] = -1236440877;
assign addr[48410] = -1252026760;
assign addr[48411] = -1267513365;
assign addr[48412] = -1282899464;
assign addr[48413] = -1298183838;
assign addr[48414] = -1313365273;
assign addr[48415] = -1328442566;
assign addr[48416] = -1343414522;
assign addr[48417] = -1358279953;
assign addr[48418] = -1373037681;
assign addr[48419] = -1387686535;
assign addr[48420] = -1402225355;
assign addr[48421] = -1416652986;
assign addr[48422] = -1430968286;
assign addr[48423] = -1445170118;
assign addr[48424] = -1459257358;
assign addr[48425] = -1473228887;
assign addr[48426] = -1487083598;
assign addr[48427] = -1500820393;
assign addr[48428] = -1514438181;
assign addr[48429] = -1527935884;
assign addr[48430] = -1541312431;
assign addr[48431] = -1554566762;
assign addr[48432] = -1567697824;
assign addr[48433] = -1580704578;
assign addr[48434] = -1593585992;
assign addr[48435] = -1606341043;
assign addr[48436] = -1618968722;
assign addr[48437] = -1631468027;
assign addr[48438] = -1643837966;
assign addr[48439] = -1656077559;
assign addr[48440] = -1668185835;
assign addr[48441] = -1680161834;
assign addr[48442] = -1692004606;
assign addr[48443] = -1703713213;
assign addr[48444] = -1715286726;
assign addr[48445] = -1726724227;
assign addr[48446] = -1738024810;
assign addr[48447] = -1749187577;
assign addr[48448] = -1760211645;
assign addr[48449] = -1771096139;
assign addr[48450] = -1781840195;
assign addr[48451] = -1792442963;
assign addr[48452] = -1802903601;
assign addr[48453] = -1813221279;
assign addr[48454] = -1823395180;
assign addr[48455] = -1833424497;
assign addr[48456] = -1843308435;
assign addr[48457] = -1853046210;
assign addr[48458] = -1862637049;
assign addr[48459] = -1872080193;
assign addr[48460] = -1881374892;
assign addr[48461] = -1890520410;
assign addr[48462] = -1899516021;
assign addr[48463] = -1908361011;
assign addr[48464] = -1917054681;
assign addr[48465] = -1925596340;
assign addr[48466] = -1933985310;
assign addr[48467] = -1942220928;
assign addr[48468] = -1950302539;
assign addr[48469] = -1958229503;
assign addr[48470] = -1966001192;
assign addr[48471] = -1973616989;
assign addr[48472] = -1981076290;
assign addr[48473] = -1988378503;
assign addr[48474] = -1995523051;
assign addr[48475] = -2002509365;
assign addr[48476] = -2009336893;
assign addr[48477] = -2016005093;
assign addr[48478] = -2022513436;
assign addr[48479] = -2028861406;
assign addr[48480] = -2035048499;
assign addr[48481] = -2041074226;
assign addr[48482] = -2046938108;
assign addr[48483] = -2052639680;
assign addr[48484] = -2058178491;
assign addr[48485] = -2063554100;
assign addr[48486] = -2068766083;
assign addr[48487] = -2073814024;
assign addr[48488] = -2078697525;
assign addr[48489] = -2083416198;
assign addr[48490] = -2087969669;
assign addr[48491] = -2092357577;
assign addr[48492] = -2096579573;
assign addr[48493] = -2100635323;
assign addr[48494] = -2104524506;
assign addr[48495] = -2108246813;
assign addr[48496] = -2111801949;
assign addr[48497] = -2115189632;
assign addr[48498] = -2118409593;
assign addr[48499] = -2121461578;
assign addr[48500] = -2124345343;
assign addr[48501] = -2127060661;
assign addr[48502] = -2129607316;
assign addr[48503] = -2131985106;
assign addr[48504] = -2134193842;
assign addr[48505] = -2136233350;
assign addr[48506] = -2138103468;
assign addr[48507] = -2139804048;
assign addr[48508] = -2141334954;
assign addr[48509] = -2142696065;
assign addr[48510] = -2143887273;
assign addr[48511] = -2144908484;
assign addr[48512] = -2145759618;
assign addr[48513] = -2146440605;
assign addr[48514] = -2146951393;
assign addr[48515] = -2147291941;
assign addr[48516] = -2147462221;
assign addr[48517] = -2147462221;
assign addr[48518] = -2147291941;
assign addr[48519] = -2146951393;
assign addr[48520] = -2146440605;
assign addr[48521] = -2145759618;
assign addr[48522] = -2144908484;
assign addr[48523] = -2143887273;
assign addr[48524] = -2142696065;
assign addr[48525] = -2141334954;
assign addr[48526] = -2139804048;
assign addr[48527] = -2138103468;
assign addr[48528] = -2136233350;
assign addr[48529] = -2134193842;
assign addr[48530] = -2131985106;
assign addr[48531] = -2129607316;
assign addr[48532] = -2127060661;
assign addr[48533] = -2124345343;
assign addr[48534] = -2121461578;
assign addr[48535] = -2118409593;
assign addr[48536] = -2115189632;
assign addr[48537] = -2111801949;
assign addr[48538] = -2108246813;
assign addr[48539] = -2104524506;
assign addr[48540] = -2100635323;
assign addr[48541] = -2096579573;
assign addr[48542] = -2092357577;
assign addr[48543] = -2087969669;
assign addr[48544] = -2083416198;
assign addr[48545] = -2078697525;
assign addr[48546] = -2073814024;
assign addr[48547] = -2068766083;
assign addr[48548] = -2063554100;
assign addr[48549] = -2058178491;
assign addr[48550] = -2052639680;
assign addr[48551] = -2046938108;
assign addr[48552] = -2041074226;
assign addr[48553] = -2035048499;
assign addr[48554] = -2028861406;
assign addr[48555] = -2022513436;
assign addr[48556] = -2016005093;
assign addr[48557] = -2009336893;
assign addr[48558] = -2002509365;
assign addr[48559] = -1995523051;
assign addr[48560] = -1988378503;
assign addr[48561] = -1981076290;
assign addr[48562] = -1973616989;
assign addr[48563] = -1966001192;
assign addr[48564] = -1958229503;
assign addr[48565] = -1950302539;
assign addr[48566] = -1942220928;
assign addr[48567] = -1933985310;
assign addr[48568] = -1925596340;
assign addr[48569] = -1917054681;
assign addr[48570] = -1908361011;
assign addr[48571] = -1899516021;
assign addr[48572] = -1890520410;
assign addr[48573] = -1881374892;
assign addr[48574] = -1872080193;
assign addr[48575] = -1862637049;
assign addr[48576] = -1853046210;
assign addr[48577] = -1843308435;
assign addr[48578] = -1833424497;
assign addr[48579] = -1823395180;
assign addr[48580] = -1813221279;
assign addr[48581] = -1802903601;
assign addr[48582] = -1792442963;
assign addr[48583] = -1781840195;
assign addr[48584] = -1771096139;
assign addr[48585] = -1760211645;
assign addr[48586] = -1749187577;
assign addr[48587] = -1738024810;
assign addr[48588] = -1726724227;
assign addr[48589] = -1715286726;
assign addr[48590] = -1703713213;
assign addr[48591] = -1692004606;
assign addr[48592] = -1680161834;
assign addr[48593] = -1668185835;
assign addr[48594] = -1656077559;
assign addr[48595] = -1643837966;
assign addr[48596] = -1631468027;
assign addr[48597] = -1618968722;
assign addr[48598] = -1606341043;
assign addr[48599] = -1593585992;
assign addr[48600] = -1580704578;
assign addr[48601] = -1567697824;
assign addr[48602] = -1554566762;
assign addr[48603] = -1541312431;
assign addr[48604] = -1527935884;
assign addr[48605] = -1514438181;
assign addr[48606] = -1500820393;
assign addr[48607] = -1487083598;
assign addr[48608] = -1473228887;
assign addr[48609] = -1459257358;
assign addr[48610] = -1445170118;
assign addr[48611] = -1430968286;
assign addr[48612] = -1416652986;
assign addr[48613] = -1402225355;
assign addr[48614] = -1387686535;
assign addr[48615] = -1373037681;
assign addr[48616] = -1358279953;
assign addr[48617] = -1343414522;
assign addr[48618] = -1328442566;
assign addr[48619] = -1313365273;
assign addr[48620] = -1298183838;
assign addr[48621] = -1282899464;
assign addr[48622] = -1267513365;
assign addr[48623] = -1252026760;
assign addr[48624] = -1236440877;
assign addr[48625] = -1220756951;
assign addr[48626] = -1204976227;
assign addr[48627] = -1189099956;
assign addr[48628] = -1173129396;
assign addr[48629] = -1157065814;
assign addr[48630] = -1140910484;
assign addr[48631] = -1124664687;
assign addr[48632] = -1108329711;
assign addr[48633] = -1091906851;
assign addr[48634] = -1075397409;
assign addr[48635] = -1058802695;
assign addr[48636] = -1042124025;
assign addr[48637] = -1025362720;
assign addr[48638] = -1008520110;
assign addr[48639] = -991597531;
assign addr[48640] = -974596324;
assign addr[48641] = -957517838;
assign addr[48642] = -940363427;
assign addr[48643] = -923134450;
assign addr[48644] = -905832274;
assign addr[48645] = -888458272;
assign addr[48646] = -871013820;
assign addr[48647] = -853500302;
assign addr[48648] = -835919107;
assign addr[48649] = -818271628;
assign addr[48650] = -800559266;
assign addr[48651] = -782783424;
assign addr[48652] = -764945512;
assign addr[48653] = -747046944;
assign addr[48654] = -729089140;
assign addr[48655] = -711073524;
assign addr[48656] = -693001525;
assign addr[48657] = -674874574;
assign addr[48658] = -656694110;
assign addr[48659] = -638461574;
assign addr[48660] = -620178412;
assign addr[48661] = -601846074;
assign addr[48662] = -583466013;
assign addr[48663] = -565039687;
assign addr[48664] = -546568556;
assign addr[48665] = -528054086;
assign addr[48666] = -509497745;
assign addr[48667] = -490901003;
assign addr[48668] = -472265336;
assign addr[48669] = -453592221;
assign addr[48670] = -434883140;
assign addr[48671] = -416139574;
assign addr[48672] = -397363011;
assign addr[48673] = -378554940;
assign addr[48674] = -359716852;
assign addr[48675] = -340850240;
assign addr[48676] = -321956601;
assign addr[48677] = -303037433;
assign addr[48678] = -284094236;
assign addr[48679] = -265128512;
assign addr[48680] = -246141764;
assign addr[48681] = -227135500;
assign addr[48682] = -208111224;
assign addr[48683] = -189070447;
assign addr[48684] = -170014678;
assign addr[48685] = -150945428;
assign addr[48686] = -131864208;
assign addr[48687] = -112772533;
assign addr[48688] = -93671915;
assign addr[48689] = -74563870;
assign addr[48690] = -55449912;
assign addr[48691] = -36331557;
assign addr[48692] = -17210322;
assign addr[48693] = 1912278;
assign addr[48694] = 21034727;
assign addr[48695] = 40155507;
assign addr[48696] = 59273104;
assign addr[48697] = 78386000;
assign addr[48698] = 97492681;
assign addr[48699] = 116591632;
assign addr[48700] = 135681337;
assign addr[48701] = 154760284;
assign addr[48702] = 173826959;
assign addr[48703] = 192879850;
assign addr[48704] = 211917448;
assign addr[48705] = 230938242;
assign addr[48706] = 249940723;
assign addr[48707] = 268923386;
assign addr[48708] = 287884725;
assign addr[48709] = 306823237;
assign addr[48710] = 325737419;
assign addr[48711] = 344625773;
assign addr[48712] = 363486799;
assign addr[48713] = 382319004;
assign addr[48714] = 401120892;
assign addr[48715] = 419890975;
assign addr[48716] = 438627762;
assign addr[48717] = 457329769;
assign addr[48718] = 475995513;
assign addr[48719] = 494623513;
assign addr[48720] = 513212292;
assign addr[48721] = 531760377;
assign addr[48722] = 550266296;
assign addr[48723] = 568728583;
assign addr[48724] = 587145773;
assign addr[48725] = 605516406;
assign addr[48726] = 623839025;
assign addr[48727] = 642112178;
assign addr[48728] = 660334415;
assign addr[48729] = 678504291;
assign addr[48730] = 696620367;
assign addr[48731] = 714681204;
assign addr[48732] = 732685372;
assign addr[48733] = 750631442;
assign addr[48734] = 768517992;
assign addr[48735] = 786343603;
assign addr[48736] = 804106861;
assign addr[48737] = 821806359;
assign addr[48738] = 839440693;
assign addr[48739] = 857008464;
assign addr[48740] = 874508280;
assign addr[48741] = 891938752;
assign addr[48742] = 909298500;
assign addr[48743] = 926586145;
assign addr[48744] = 943800318;
assign addr[48745] = 960939653;
assign addr[48746] = 978002791;
assign addr[48747] = 994988380;
assign addr[48748] = 1011895073;
assign addr[48749] = 1028721528;
assign addr[48750] = 1045466412;
assign addr[48751] = 1062128397;
assign addr[48752] = 1078706161;
assign addr[48753] = 1095198391;
assign addr[48754] = 1111603778;
assign addr[48755] = 1127921022;
assign addr[48756] = 1144148829;
assign addr[48757] = 1160285911;
assign addr[48758] = 1176330990;
assign addr[48759] = 1192282793;
assign addr[48760] = 1208140056;
assign addr[48761] = 1223901520;
assign addr[48762] = 1239565936;
assign addr[48763] = 1255132063;
assign addr[48764] = 1270598665;
assign addr[48765] = 1285964516;
assign addr[48766] = 1301228398;
assign addr[48767] = 1316389101;
assign addr[48768] = 1331445422;
assign addr[48769] = 1346396168;
assign addr[48770] = 1361240152;
assign addr[48771] = 1375976199;
assign addr[48772] = 1390603139;
assign addr[48773] = 1405119813;
assign addr[48774] = 1419525069;
assign addr[48775] = 1433817766;
assign addr[48776] = 1447996770;
assign addr[48777] = 1462060956;
assign addr[48778] = 1476009210;
assign addr[48779] = 1489840425;
assign addr[48780] = 1503553506;
assign addr[48781] = 1517147363;
assign addr[48782] = 1530620920;
assign addr[48783] = 1543973108;
assign addr[48784] = 1557202869;
assign addr[48785] = 1570309153;
assign addr[48786] = 1583290921;
assign addr[48787] = 1596147143;
assign addr[48788] = 1608876801;
assign addr[48789] = 1621478885;
assign addr[48790] = 1633952396;
assign addr[48791] = 1646296344;
assign addr[48792] = 1658509750;
assign addr[48793] = 1670591647;
assign addr[48794] = 1682541077;
assign addr[48795] = 1694357091;
assign addr[48796] = 1706038753;
assign addr[48797] = 1717585136;
assign addr[48798] = 1728995326;
assign addr[48799] = 1740268417;
assign addr[48800] = 1751403515;
assign addr[48801] = 1762399737;
assign addr[48802] = 1773256212;
assign addr[48803] = 1783972079;
assign addr[48804] = 1794546487;
assign addr[48805] = 1804978599;
assign addr[48806] = 1815267588;
assign addr[48807] = 1825412636;
assign addr[48808] = 1835412941;
assign addr[48809] = 1845267708;
assign addr[48810] = 1854976157;
assign addr[48811] = 1864537518;
assign addr[48812] = 1873951032;
assign addr[48813] = 1883215953;
assign addr[48814] = 1892331547;
assign addr[48815] = 1901297091;
assign addr[48816] = 1910111873;
assign addr[48817] = 1918775195;
assign addr[48818] = 1927286370;
assign addr[48819] = 1935644723;
assign addr[48820] = 1943849591;
assign addr[48821] = 1951900324;
assign addr[48822] = 1959796283;
assign addr[48823] = 1967536842;
assign addr[48824] = 1975121388;
assign addr[48825] = 1982549318;
assign addr[48826] = 1989820044;
assign addr[48827] = 1996932990;
assign addr[48828] = 2003887591;
assign addr[48829] = 2010683297;
assign addr[48830] = 2017319567;
assign addr[48831] = 2023795876;
assign addr[48832] = 2030111710;
assign addr[48833] = 2036266570;
assign addr[48834] = 2042259965;
assign addr[48835] = 2048091422;
assign addr[48836] = 2053760478;
assign addr[48837] = 2059266683;
assign addr[48838] = 2064609600;
assign addr[48839] = 2069788807;
assign addr[48840] = 2074803892;
assign addr[48841] = 2079654458;
assign addr[48842] = 2084340120;
assign addr[48843] = 2088860507;
assign addr[48844] = 2093215260;
assign addr[48845] = 2097404033;
assign addr[48846] = 2101426496;
assign addr[48847] = 2105282327;
assign addr[48848] = 2108971223;
assign addr[48849] = 2112492891;
assign addr[48850] = 2115847050;
assign addr[48851] = 2119033436;
assign addr[48852] = 2122051796;
assign addr[48853] = 2124901890;
assign addr[48854] = 2127583492;
assign addr[48855] = 2130096389;
assign addr[48856] = 2132440383;
assign addr[48857] = 2134615288;
assign addr[48858] = 2136620930;
assign addr[48859] = 2138457152;
assign addr[48860] = 2140123807;
assign addr[48861] = 2141620763;
assign addr[48862] = 2142947902;
assign addr[48863] = 2144105118;
assign addr[48864] = 2145092320;
assign addr[48865] = 2145909429;
assign addr[48866] = 2146556380;
assign addr[48867] = 2147033123;
assign addr[48868] = 2147339619;
assign addr[48869] = 2147475844;
assign addr[48870] = 2147441787;
assign addr[48871] = 2147237452;
assign addr[48872] = 2146862854;
assign addr[48873] = 2146318022;
assign addr[48874] = 2145603001;
assign addr[48875] = 2144717846;
assign addr[48876] = 2143662628;
assign addr[48877] = 2142437431;
assign addr[48878] = 2141042352;
assign addr[48879] = 2139477502;
assign addr[48880] = 2137743003;
assign addr[48881] = 2135838995;
assign addr[48882] = 2133765628;
assign addr[48883] = 2131523066;
assign addr[48884] = 2129111488;
assign addr[48885] = 2126531084;
assign addr[48886] = 2123782059;
assign addr[48887] = 2120864631;
assign addr[48888] = 2117779031;
assign addr[48889] = 2114525505;
assign addr[48890] = 2111104309;
assign addr[48891] = 2107515716;
assign addr[48892] = 2103760010;
assign addr[48893] = 2099837489;
assign addr[48894] = 2095748463;
assign addr[48895] = 2091493257;
assign addr[48896] = 2087072209;
assign addr[48897] = 2082485668;
assign addr[48898] = 2077733999;
assign addr[48899] = 2072817579;
assign addr[48900] = 2067736796;
assign addr[48901] = 2062492055;
assign addr[48902] = 2057083771;
assign addr[48903] = 2051512372;
assign addr[48904] = 2045778302;
assign addr[48905] = 2039882013;
assign addr[48906] = 2033823974;
assign addr[48907] = 2027604666;
assign addr[48908] = 2021224581;
assign addr[48909] = 2014684225;
assign addr[48910] = 2007984117;
assign addr[48911] = 2001124788;
assign addr[48912] = 1994106782;
assign addr[48913] = 1986930656;
assign addr[48914] = 1979596978;
assign addr[48915] = 1972106330;
assign addr[48916] = 1964459306;
assign addr[48917] = 1956656513;
assign addr[48918] = 1948698568;
assign addr[48919] = 1940586104;
assign addr[48920] = 1932319763;
assign addr[48921] = 1923900201;
assign addr[48922] = 1915328086;
assign addr[48923] = 1906604097;
assign addr[48924] = 1897728925;
assign addr[48925] = 1888703276;
assign addr[48926] = 1879527863;
assign addr[48927] = 1870203416;
assign addr[48928] = 1860730673;
assign addr[48929] = 1851110385;
assign addr[48930] = 1841343316;
assign addr[48931] = 1831430239;
assign addr[48932] = 1821371941;
assign addr[48933] = 1811169220;
assign addr[48934] = 1800822883;
assign addr[48935] = 1790333753;
assign addr[48936] = 1779702660;
assign addr[48937] = 1768930447;
assign addr[48938] = 1758017969;
assign addr[48939] = 1746966091;
assign addr[48940] = 1735775690;
assign addr[48941] = 1724447652;
assign addr[48942] = 1712982875;
assign addr[48943] = 1701382270;
assign addr[48944] = 1689646755;
assign addr[48945] = 1677777262;
assign addr[48946] = 1665774731;
assign addr[48947] = 1653640115;
assign addr[48948] = 1641374375;
assign addr[48949] = 1628978484;
assign addr[48950] = 1616453425;
assign addr[48951] = 1603800191;
assign addr[48952] = 1591019785;
assign addr[48953] = 1578113222;
assign addr[48954] = 1565081523;
assign addr[48955] = 1551925723;
assign addr[48956] = 1538646865;
assign addr[48957] = 1525246002;
assign addr[48958] = 1511724196;
assign addr[48959] = 1498082520;
assign addr[48960] = 1484322054;
assign addr[48961] = 1470443891;
assign addr[48962] = 1456449131;
assign addr[48963] = 1442338884;
assign addr[48964] = 1428114267;
assign addr[48965] = 1413776410;
assign addr[48966] = 1399326449;
assign addr[48967] = 1384765530;
assign addr[48968] = 1370094808;
assign addr[48969] = 1355315445;
assign addr[48970] = 1340428615;
assign addr[48971] = 1325435496;
assign addr[48972] = 1310337279;
assign addr[48973] = 1295135159;
assign addr[48974] = 1279830344;
assign addr[48975] = 1264424045;
assign addr[48976] = 1248917486;
assign addr[48977] = 1233311895;
assign addr[48978] = 1217608510;
assign addr[48979] = 1201808576;
assign addr[48980] = 1185913346;
assign addr[48981] = 1169924081;
assign addr[48982] = 1153842047;
assign addr[48983] = 1137668521;
assign addr[48984] = 1121404785;
assign addr[48985] = 1105052128;
assign addr[48986] = 1088611847;
assign addr[48987] = 1072085246;
assign addr[48988] = 1055473635;
assign addr[48989] = 1038778332;
assign addr[48990] = 1022000660;
assign addr[48991] = 1005141949;
assign addr[48992] = 988203537;
assign addr[48993] = 971186766;
assign addr[48994] = 954092986;
assign addr[48995] = 936923553;
assign addr[48996] = 919679827;
assign addr[48997] = 902363176;
assign addr[48998] = 884974973;
assign addr[48999] = 867516597;
assign addr[49000] = 849989433;
assign addr[49001] = 832394869;
assign addr[49002] = 814734301;
assign addr[49003] = 797009130;
assign addr[49004] = 779220762;
assign addr[49005] = 761370605;
assign addr[49006] = 743460077;
assign addr[49007] = 725490597;
assign addr[49008] = 707463589;
assign addr[49009] = 689380485;
assign addr[49010] = 671242716;
assign addr[49011] = 653051723;
assign addr[49012] = 634808946;
assign addr[49013] = 616515832;
assign addr[49014] = 598173833;
assign addr[49015] = 579784402;
assign addr[49016] = 561348998;
assign addr[49017] = 542869083;
assign addr[49018] = 524346121;
assign addr[49019] = 505781581;
assign addr[49020] = 487176937;
assign addr[49021] = 468533662;
assign addr[49022] = 449853235;
assign addr[49023] = 431137138;
assign addr[49024] = 412386854;
assign addr[49025] = 393603870;
assign addr[49026] = 374789676;
assign addr[49027] = 355945764;
assign addr[49028] = 337073627;
assign addr[49029] = 318174762;
assign addr[49030] = 299250668;
assign addr[49031] = 280302845;
assign addr[49032] = 261332796;
assign addr[49033] = 242342025;
assign addr[49034] = 223332037;
assign addr[49035] = 204304341;
assign addr[49036] = 185260444;
assign addr[49037] = 166201858;
assign addr[49038] = 147130093;
assign addr[49039] = 128046661;
assign addr[49040] = 108953076;
assign addr[49041] = 89850852;
assign addr[49042] = 70741503;
assign addr[49043] = 51626544;
assign addr[49044] = 32507492;
assign addr[49045] = 13385863;
assign addr[49046] = -5736829;
assign addr[49047] = -24859065;
assign addr[49048] = -43979330;
assign addr[49049] = -63096108;
assign addr[49050] = -82207882;
assign addr[49051] = -101313138;
assign addr[49052] = -120410361;
assign addr[49053] = -139498035;
assign addr[49054] = -158574649;
assign addr[49055] = -177638688;
assign addr[49056] = -196688642;
assign addr[49057] = -215722999;
assign addr[49058] = -234740251;
assign addr[49059] = -253738890;
assign addr[49060] = -272717408;
assign addr[49061] = -291674302;
assign addr[49062] = -310608068;
assign addr[49063] = -329517204;
assign addr[49064] = -348400212;
assign addr[49065] = -367255594;
assign addr[49066] = -386081854;
assign addr[49067] = -404877501;
assign addr[49068] = -423641043;
assign addr[49069] = -442370993;
assign addr[49070] = -461065866;
assign addr[49071] = -479724180;
assign addr[49072] = -498344454;
assign addr[49073] = -516925212;
assign addr[49074] = -535464981;
assign addr[49075] = -553962291;
assign addr[49076] = -572415676;
assign addr[49077] = -590823671;
assign addr[49078] = -609184818;
assign addr[49079] = -627497660;
assign addr[49080] = -645760745;
assign addr[49081] = -663972625;
assign addr[49082] = -682131857;
assign addr[49083] = -700236999;
assign addr[49084] = -718286617;
assign addr[49085] = -736279279;
assign addr[49086] = -754213559;
assign addr[49087] = -772088034;
assign addr[49088] = -789901288;
assign addr[49089] = -807651907;
assign addr[49090] = -825338484;
assign addr[49091] = -842959617;
assign addr[49092] = -860513908;
assign addr[49093] = -877999966;
assign addr[49094] = -895416404;
assign addr[49095] = -912761841;
assign addr[49096] = -930034901;
assign addr[49097] = -947234215;
assign addr[49098] = -964358420;
assign addr[49099] = -981406156;
assign addr[49100] = -998376073;
assign addr[49101] = -1015266825;
assign addr[49102] = -1032077073;
assign addr[49103] = -1048805483;
assign addr[49104] = -1065450729;
assign addr[49105] = -1082011492;
assign addr[49106] = -1098486458;
assign addr[49107] = -1114874320;
assign addr[49108] = -1131173780;
assign addr[49109] = -1147383544;
assign addr[49110] = -1163502328;
assign addr[49111] = -1179528853;
assign addr[49112] = -1195461849;
assign addr[49113] = -1211300053;
assign addr[49114] = -1227042207;
assign addr[49115] = -1242687064;
assign addr[49116] = -1258233384;
assign addr[49117] = -1273679934;
assign addr[49118] = -1289025489;
assign addr[49119] = -1304268832;
assign addr[49120] = -1319408754;
assign addr[49121] = -1334444055;
assign addr[49122] = -1349373543;
assign addr[49123] = -1364196034;
assign addr[49124] = -1378910353;
assign addr[49125] = -1393515332;
assign addr[49126] = -1408009814;
assign addr[49127] = -1422392650;
assign addr[49128] = -1436662698;
assign addr[49129] = -1450818828;
assign addr[49130] = -1464859917;
assign addr[49131] = -1478784851;
assign addr[49132] = -1492592527;
assign addr[49133] = -1506281850;
assign addr[49134] = -1519851733;
assign addr[49135] = -1533301101;
assign addr[49136] = -1546628888;
assign addr[49137] = -1559834037;
assign addr[49138] = -1572915501;
assign addr[49139] = -1585872242;
assign addr[49140] = -1598703233;
assign addr[49141] = -1611407456;
assign addr[49142] = -1623983905;
assign addr[49143] = -1636431582;
assign addr[49144] = -1648749499;
assign addr[49145] = -1660936681;
assign addr[49146] = -1672992161;
assign addr[49147] = -1684914983;
assign addr[49148] = -1696704201;
assign addr[49149] = -1708358881;
assign addr[49150] = -1719878099;
assign addr[49151] = -1731260941;
assign addr[49152] = -1742506504;
assign addr[49153] = -1753613897;
assign addr[49154] = -1764582240;
assign addr[49155] = -1775410662;
assign addr[49156] = -1786098304;
assign addr[49157] = -1796644320;
assign addr[49158] = -1807047873;
assign addr[49159] = -1817308138;
assign addr[49160] = -1827424302;
assign addr[49161] = -1837395562;
assign addr[49162] = -1847221128;
assign addr[49163] = -1856900221;
assign addr[49164] = -1866432072;
assign addr[49165] = -1875815927;
assign addr[49166] = -1885051042;
assign addr[49167] = -1894136683;
assign addr[49168] = -1903072131;
assign addr[49169] = -1911856677;
assign addr[49170] = -1920489624;
assign addr[49171] = -1928970288;
assign addr[49172] = -1937297997;
assign addr[49173] = -1945472089;
assign addr[49174] = -1953491918;
assign addr[49175] = -1961356847;
assign addr[49176] = -1969066252;
assign addr[49177] = -1976619522;
assign addr[49178] = -1984016058;
assign addr[49179] = -1991255274;
assign addr[49180] = -1998336596;
assign addr[49181] = -2005259462;
assign addr[49182] = -2012023322;
assign addr[49183] = -2018627642;
assign addr[49184] = -2025071897;
assign addr[49185] = -2031355576;
assign addr[49186] = -2037478181;
assign addr[49187] = -2043439226;
assign addr[49188] = -2049238240;
assign addr[49189] = -2054874761;
assign addr[49190] = -2060348343;
assign addr[49191] = -2065658552;
assign addr[49192] = -2070804967;
assign addr[49193] = -2075787180;
assign addr[49194] = -2080604795;
assign addr[49195] = -2085257431;
assign addr[49196] = -2089744719;
assign addr[49197] = -2094066304;
assign addr[49198] = -2098221841;
assign addr[49199] = -2102211002;
assign addr[49200] = -2106033471;
assign addr[49201] = -2109688944;
assign addr[49202] = -2113177132;
assign addr[49203] = -2116497758;
assign addr[49204] = -2119650558;
assign addr[49205] = -2122635283;
assign addr[49206] = -2125451696;
assign addr[49207] = -2128099574;
assign addr[49208] = -2130578706;
assign addr[49209] = -2132888897;
assign addr[49210] = -2135029962;
assign addr[49211] = -2137001733;
assign addr[49212] = -2138804053;
assign addr[49213] = -2140436778;
assign addr[49214] = -2141899780;
assign addr[49215] = -2143192942;
assign addr[49216] = -2144316162;
assign addr[49217] = -2145269351;
assign addr[49218] = -2146052433;
assign addr[49219] = -2146665347;
assign addr[49220] = -2147108043;
assign addr[49221] = -2147380486;
assign addr[49222] = -2147482655;
assign addr[49223] = -2147414542;
assign addr[49224] = -2147176152;
assign addr[49225] = -2146767505;
assign addr[49226] = -2146188631;
assign addr[49227] = -2145439578;
assign addr[49228] = -2144520405;
assign addr[49229] = -2143431184;
assign addr[49230] = -2142172003;
assign addr[49231] = -2140742960;
assign addr[49232] = -2139144169;
assign addr[49233] = -2137375758;
assign addr[49234] = -2135437865;
assign addr[49235] = -2133330646;
assign addr[49236] = -2131054266;
assign addr[49237] = -2128608907;
assign addr[49238] = -2125994762;
assign addr[49239] = -2123212038;
assign addr[49240] = -2120260957;
assign addr[49241] = -2117141752;
assign addr[49242] = -2113854671;
assign addr[49243] = -2110399974;
assign addr[49244] = -2106777935;
assign addr[49245] = -2102988841;
assign addr[49246] = -2099032994;
assign addr[49247] = -2094910706;
assign addr[49248] = -2090622304;
assign addr[49249] = -2086168128;
assign addr[49250] = -2081548533;
assign addr[49251] = -2076763883;
assign addr[49252] = -2071814558;
assign addr[49253] = -2066700952;
assign addr[49254] = -2061423468;
assign addr[49255] = -2055982526;
assign addr[49256] = -2050378558;
assign addr[49257] = -2044612007;
assign addr[49258] = -2038683330;
assign addr[49259] = -2032592999;
assign addr[49260] = -2026341495;
assign addr[49261] = -2019929315;
assign addr[49262] = -2013356967;
assign addr[49263] = -2006624971;
assign addr[49264] = -1999733863;
assign addr[49265] = -1992684188;
assign addr[49266] = -1985476506;
assign addr[49267] = -1978111387;
assign addr[49268] = -1970589416;
assign addr[49269] = -1962911189;
assign addr[49270] = -1955077316;
assign addr[49271] = -1947088417;
assign addr[49272] = -1938945125;
assign addr[49273] = -1930648088;
assign addr[49274] = -1922197961;
assign addr[49275] = -1913595416;
assign addr[49276] = -1904841135;
assign addr[49277] = -1895935811;
assign addr[49278] = -1886880151;
assign addr[49279] = -1877674873;
assign addr[49280] = -1868320707;
assign addr[49281] = -1858818395;
assign addr[49282] = -1849168689;
assign addr[49283] = -1839372356;
assign addr[49284] = -1829430172;
assign addr[49285] = -1819342925;
assign addr[49286] = -1809111415;
assign addr[49287] = -1798736454;
assign addr[49288] = -1788218865;
assign addr[49289] = -1777559480;
assign addr[49290] = -1766759146;
assign addr[49291] = -1755818718;
assign addr[49292] = -1744739065;
assign addr[49293] = -1733521064;
assign addr[49294] = -1722165606;
assign addr[49295] = -1710673591;
assign addr[49296] = -1699045930;
assign addr[49297] = -1687283545;
assign addr[49298] = -1675387369;
assign addr[49299] = -1663358344;
assign addr[49300] = -1651197426;
assign addr[49301] = -1638905577;
assign addr[49302] = -1626483774;
assign addr[49303] = -1613933000;
assign addr[49304] = -1601254251;
assign addr[49305] = -1588448533;
assign addr[49306] = -1575516860;
assign addr[49307] = -1562460258;
assign addr[49308] = -1549279763;
assign addr[49309] = -1535976419;
assign addr[49310] = -1522551282;
assign addr[49311] = -1509005416;
assign addr[49312] = -1495339895;
assign addr[49313] = -1481555802;
assign addr[49314] = -1467654232;
assign addr[49315] = -1453636285;
assign addr[49316] = -1439503074;
assign addr[49317] = -1425255719;
assign addr[49318] = -1410895350;
assign addr[49319] = -1396423105;
assign addr[49320] = -1381840133;
assign addr[49321] = -1367147589;
assign addr[49322] = -1352346639;
assign addr[49323] = -1337438456;
assign addr[49324] = -1322424222;
assign addr[49325] = -1307305128;
assign addr[49326] = -1292082373;
assign addr[49327] = -1276757164;
assign addr[49328] = -1261330715;
assign addr[49329] = -1245804251;
assign addr[49330] = -1230179002;
assign addr[49331] = -1214456207;
assign addr[49332] = -1198637114;
assign addr[49333] = -1182722976;
assign addr[49334] = -1166715055;
assign addr[49335] = -1150614620;
assign addr[49336] = -1134422949;
assign addr[49337] = -1118141326;
assign addr[49338] = -1101771040;
assign addr[49339] = -1085313391;
assign addr[49340] = -1068769683;
assign addr[49341] = -1052141228;
assign addr[49342] = -1035429345;
assign addr[49343] = -1018635358;
assign addr[49344] = -1001760600;
assign addr[49345] = -984806408;
assign addr[49346] = -967774128;
assign addr[49347] = -950665109;
assign addr[49348] = -933480707;
assign addr[49349] = -916222287;
assign addr[49350] = -898891215;
assign addr[49351] = -881488868;
assign addr[49352] = -864016623;
assign addr[49353] = -846475867;
assign addr[49354] = -828867991;
assign addr[49355] = -811194391;
assign addr[49356] = -793456467;
assign addr[49357] = -775655628;
assign addr[49358] = -757793284;
assign addr[49359] = -739870851;
assign addr[49360] = -721889752;
assign addr[49361] = -703851410;
assign addr[49362] = -685757258;
assign addr[49363] = -667608730;
assign addr[49364] = -649407264;
assign addr[49365] = -631154304;
assign addr[49366] = -612851297;
assign addr[49367] = -594499695;
assign addr[49368] = -576100953;
assign addr[49369] = -557656529;
assign addr[49370] = -539167887;
assign addr[49371] = -520636492;
assign addr[49372] = -502063814;
assign addr[49373] = -483451325;
assign addr[49374] = -464800501;
assign addr[49375] = -446112822;
assign addr[49376] = -427389768;
assign addr[49377] = -408632825;
assign addr[49378] = -389843480;
assign addr[49379] = -371023223;
assign addr[49380] = -352173546;
assign addr[49381] = -333295944;
assign addr[49382] = -314391913;
assign addr[49383] = -295462954;
assign addr[49384] = -276510565;
assign addr[49385] = -257536251;
assign addr[49386] = -238541516;
assign addr[49387] = -219527866;
assign addr[49388] = -200496809;
assign addr[49389] = -181449854;
assign addr[49390] = -162388511;
assign addr[49391] = -143314291;
assign addr[49392] = -124228708;
assign addr[49393] = -105133274;
assign addr[49394] = -86029503;
assign addr[49395] = -66918911;
assign addr[49396] = -47803013;
assign addr[49397] = -28683324;
assign addr[49398] = -9561361;
assign addr[49399] = 9561361;
assign addr[49400] = 28683324;
assign addr[49401] = 47803013;
assign addr[49402] = 66918911;
assign addr[49403] = 86029503;
assign addr[49404] = 105133274;
assign addr[49405] = 124228708;
assign addr[49406] = 143314291;
assign addr[49407] = 162388511;
assign addr[49408] = 181449854;
assign addr[49409] = 200496809;
assign addr[49410] = 219527866;
assign addr[49411] = 238541516;
assign addr[49412] = 257536251;
assign addr[49413] = 276510565;
assign addr[49414] = 295462953;
assign addr[49415] = 314391913;
assign addr[49416] = 333295944;
assign addr[49417] = 352173546;
assign addr[49418] = 371023223;
assign addr[49419] = 389843480;
assign addr[49420] = 408632825;
assign addr[49421] = 427389768;
assign addr[49422] = 446112822;
assign addr[49423] = 464800501;
assign addr[49424] = 483451325;
assign addr[49425] = 502063814;
assign addr[49426] = 520636492;
assign addr[49427] = 539167887;
assign addr[49428] = 557656529;
assign addr[49429] = 576100953;
assign addr[49430] = 594499695;
assign addr[49431] = 612851297;
assign addr[49432] = 631154304;
assign addr[49433] = 649407264;
assign addr[49434] = 667608730;
assign addr[49435] = 685757258;
assign addr[49436] = 703851410;
assign addr[49437] = 721889752;
assign addr[49438] = 739870851;
assign addr[49439] = 757793284;
assign addr[49440] = 775655628;
assign addr[49441] = 793456467;
assign addr[49442] = 811194391;
assign addr[49443] = 828867991;
assign addr[49444] = 846475867;
assign addr[49445] = 864016623;
assign addr[49446] = 881488868;
assign addr[49447] = 898891215;
assign addr[49448] = 916222287;
assign addr[49449] = 933480707;
assign addr[49450] = 950665109;
assign addr[49451] = 967774128;
assign addr[49452] = 984806408;
assign addr[49453] = 1001760600;
assign addr[49454] = 1018635358;
assign addr[49455] = 1035429345;
assign addr[49456] = 1052141228;
assign addr[49457] = 1068769683;
assign addr[49458] = 1085313391;
assign addr[49459] = 1101771040;
assign addr[49460] = 1118141326;
assign addr[49461] = 1134422949;
assign addr[49462] = 1150614620;
assign addr[49463] = 1166715055;
assign addr[49464] = 1182722976;
assign addr[49465] = 1198637114;
assign addr[49466] = 1214456207;
assign addr[49467] = 1230179002;
assign addr[49468] = 1245804251;
assign addr[49469] = 1261330715;
assign addr[49470] = 1276757164;
assign addr[49471] = 1292082373;
assign addr[49472] = 1307305128;
assign addr[49473] = 1322424222;
assign addr[49474] = 1337438456;
assign addr[49475] = 1352346639;
assign addr[49476] = 1367147589;
assign addr[49477] = 1381840133;
assign addr[49478] = 1396423105;
assign addr[49479] = 1410895350;
assign addr[49480] = 1425255719;
assign addr[49481] = 1439503074;
assign addr[49482] = 1453636285;
assign addr[49483] = 1467654232;
assign addr[49484] = 1481555802;
assign addr[49485] = 1495339895;
assign addr[49486] = 1509005416;
assign addr[49487] = 1522551282;
assign addr[49488] = 1535976419;
assign addr[49489] = 1549279763;
assign addr[49490] = 1562460258;
assign addr[49491] = 1575516860;
assign addr[49492] = 1588448533;
assign addr[49493] = 1601254251;
assign addr[49494] = 1613933000;
assign addr[49495] = 1626483774;
assign addr[49496] = 1638905577;
assign addr[49497] = 1651197426;
assign addr[49498] = 1663358344;
assign addr[49499] = 1675387369;
assign addr[49500] = 1687283545;
assign addr[49501] = 1699045930;
assign addr[49502] = 1710673591;
assign addr[49503] = 1722165606;
assign addr[49504] = 1733521064;
assign addr[49505] = 1744739065;
assign addr[49506] = 1755818718;
assign addr[49507] = 1766759146;
assign addr[49508] = 1777559480;
assign addr[49509] = 1788218865;
assign addr[49510] = 1798736454;
assign addr[49511] = 1809111415;
assign addr[49512] = 1819342925;
assign addr[49513] = 1829430172;
assign addr[49514] = 1839372356;
assign addr[49515] = 1849168689;
assign addr[49516] = 1858818395;
assign addr[49517] = 1868320707;
assign addr[49518] = 1877674873;
assign addr[49519] = 1886880151;
assign addr[49520] = 1895935811;
assign addr[49521] = 1904841135;
assign addr[49522] = 1913595416;
assign addr[49523] = 1922197961;
assign addr[49524] = 1930648088;
assign addr[49525] = 1938945125;
assign addr[49526] = 1947088417;
assign addr[49527] = 1955077316;
assign addr[49528] = 1962911189;
assign addr[49529] = 1970589416;
assign addr[49530] = 1978111387;
assign addr[49531] = 1985476506;
assign addr[49532] = 1992684188;
assign addr[49533] = 1999733863;
assign addr[49534] = 2006624971;
assign addr[49535] = 2013356967;
assign addr[49536] = 2019929315;
assign addr[49537] = 2026341495;
assign addr[49538] = 2032592999;
assign addr[49539] = 2038683330;
assign addr[49540] = 2044612007;
assign addr[49541] = 2050378558;
assign addr[49542] = 2055982526;
assign addr[49543] = 2061423468;
assign addr[49544] = 2066700952;
assign addr[49545] = 2071814558;
assign addr[49546] = 2076763883;
assign addr[49547] = 2081548533;
assign addr[49548] = 2086168128;
assign addr[49549] = 2090622304;
assign addr[49550] = 2094910706;
assign addr[49551] = 2099032994;
assign addr[49552] = 2102988841;
assign addr[49553] = 2106777935;
assign addr[49554] = 2110399974;
assign addr[49555] = 2113854671;
assign addr[49556] = 2117141752;
assign addr[49557] = 2120260957;
assign addr[49558] = 2123212038;
assign addr[49559] = 2125994762;
assign addr[49560] = 2128608907;
assign addr[49561] = 2131054266;
assign addr[49562] = 2133330646;
assign addr[49563] = 2135437865;
assign addr[49564] = 2137375758;
assign addr[49565] = 2139144169;
assign addr[49566] = 2140742960;
assign addr[49567] = 2142172003;
assign addr[49568] = 2143431184;
assign addr[49569] = 2144520405;
assign addr[49570] = 2145439578;
assign addr[49571] = 2146188631;
assign addr[49572] = 2146767505;
assign addr[49573] = 2147176152;
assign addr[49574] = 2147414542;
assign addr[49575] = 2147482655;
assign addr[49576] = 2147380486;
assign addr[49577] = 2147108043;
assign addr[49578] = 2146665347;
assign addr[49579] = 2146052433;
assign addr[49580] = 2145269351;
assign addr[49581] = 2144316162;
assign addr[49582] = 2143192942;
assign addr[49583] = 2141899780;
assign addr[49584] = 2140436778;
assign addr[49585] = 2138804053;
assign addr[49586] = 2137001733;
assign addr[49587] = 2135029962;
assign addr[49588] = 2132888897;
assign addr[49589] = 2130578706;
assign addr[49590] = 2128099574;
assign addr[49591] = 2125451696;
assign addr[49592] = 2122635283;
assign addr[49593] = 2119650558;
assign addr[49594] = 2116497758;
assign addr[49595] = 2113177132;
assign addr[49596] = 2109688944;
assign addr[49597] = 2106033471;
assign addr[49598] = 2102211002;
assign addr[49599] = 2098221841;
assign addr[49600] = 2094066304;
assign addr[49601] = 2089744719;
assign addr[49602] = 2085257431;
assign addr[49603] = 2080604795;
assign addr[49604] = 2075787180;
assign addr[49605] = 2070804967;
assign addr[49606] = 2065658552;
assign addr[49607] = 2060348343;
assign addr[49608] = 2054874761;
assign addr[49609] = 2049238240;
assign addr[49610] = 2043439226;
assign addr[49611] = 2037478181;
assign addr[49612] = 2031355576;
assign addr[49613] = 2025071897;
assign addr[49614] = 2018627642;
assign addr[49615] = 2012023322;
assign addr[49616] = 2005259462;
assign addr[49617] = 1998336596;
assign addr[49618] = 1991255274;
assign addr[49619] = 1984016058;
assign addr[49620] = 1976619522;
assign addr[49621] = 1969066252;
assign addr[49622] = 1961356847;
assign addr[49623] = 1953491918;
assign addr[49624] = 1945472089;
assign addr[49625] = 1937297997;
assign addr[49626] = 1928970288;
assign addr[49627] = 1920489624;
assign addr[49628] = 1911856677;
assign addr[49629] = 1903072131;
assign addr[49630] = 1894136683;
assign addr[49631] = 1885051042;
assign addr[49632] = 1875815927;
assign addr[49633] = 1866432072;
assign addr[49634] = 1856900221;
assign addr[49635] = 1847221128;
assign addr[49636] = 1837395562;
assign addr[49637] = 1827424302;
assign addr[49638] = 1817308138;
assign addr[49639] = 1807047873;
assign addr[49640] = 1796644320;
assign addr[49641] = 1786098304;
assign addr[49642] = 1775410662;
assign addr[49643] = 1764582240;
assign addr[49644] = 1753613897;
assign addr[49645] = 1742506504;
assign addr[49646] = 1731260941;
assign addr[49647] = 1719878099;
assign addr[49648] = 1708358881;
assign addr[49649] = 1696704201;
assign addr[49650] = 1684914983;
assign addr[49651] = 1672992161;
assign addr[49652] = 1660936681;
assign addr[49653] = 1648749499;
assign addr[49654] = 1636431582;
assign addr[49655] = 1623983905;
assign addr[49656] = 1611407456;
assign addr[49657] = 1598703233;
assign addr[49658] = 1585872242;
assign addr[49659] = 1572915501;
assign addr[49660] = 1559834037;
assign addr[49661] = 1546628888;
assign addr[49662] = 1533301101;
assign addr[49663] = 1519851733;
assign addr[49664] = 1506281850;
assign addr[49665] = 1492592527;
assign addr[49666] = 1478784851;
assign addr[49667] = 1464859917;
assign addr[49668] = 1450818828;
assign addr[49669] = 1436662698;
assign addr[49670] = 1422392650;
assign addr[49671] = 1408009814;
assign addr[49672] = 1393515332;
assign addr[49673] = 1378910353;
assign addr[49674] = 1364196034;
assign addr[49675] = 1349373543;
assign addr[49676] = 1334444055;
assign addr[49677] = 1319408754;
assign addr[49678] = 1304268832;
assign addr[49679] = 1289025489;
assign addr[49680] = 1273679934;
assign addr[49681] = 1258233384;
assign addr[49682] = 1242687064;
assign addr[49683] = 1227042207;
assign addr[49684] = 1211300053;
assign addr[49685] = 1195461849;
assign addr[49686] = 1179528853;
assign addr[49687] = 1163502328;
assign addr[49688] = 1147383544;
assign addr[49689] = 1131173780;
assign addr[49690] = 1114874320;
assign addr[49691] = 1098486458;
assign addr[49692] = 1082011492;
assign addr[49693] = 1065450729;
assign addr[49694] = 1048805483;
assign addr[49695] = 1032077073;
assign addr[49696] = 1015266825;
assign addr[49697] = 998376073;
assign addr[49698] = 981406156;
assign addr[49699] = 964358420;
assign addr[49700] = 947234215;
assign addr[49701] = 930034901;
assign addr[49702] = 912761841;
assign addr[49703] = 895416404;
assign addr[49704] = 877999966;
assign addr[49705] = 860513908;
assign addr[49706] = 842959617;
assign addr[49707] = 825338484;
assign addr[49708] = 807651907;
assign addr[49709] = 789901288;
assign addr[49710] = 772088034;
assign addr[49711] = 754213559;
assign addr[49712] = 736279279;
assign addr[49713] = 718286617;
assign addr[49714] = 700236999;
assign addr[49715] = 682131857;
assign addr[49716] = 663972625;
assign addr[49717] = 645760745;
assign addr[49718] = 627497660;
assign addr[49719] = 609184818;
assign addr[49720] = 590823671;
assign addr[49721] = 572415676;
assign addr[49722] = 553962291;
assign addr[49723] = 535464981;
assign addr[49724] = 516925212;
assign addr[49725] = 498344454;
assign addr[49726] = 479724180;
assign addr[49727] = 461065866;
assign addr[49728] = 442370993;
assign addr[49729] = 423641043;
assign addr[49730] = 404877501;
assign addr[49731] = 386081854;
assign addr[49732] = 367255594;
assign addr[49733] = 348400212;
assign addr[49734] = 329517204;
assign addr[49735] = 310608068;
assign addr[49736] = 291674302;
assign addr[49737] = 272717408;
assign addr[49738] = 253738890;
assign addr[49739] = 234740251;
assign addr[49740] = 215722999;
assign addr[49741] = 196688642;
assign addr[49742] = 177638688;
assign addr[49743] = 158574649;
assign addr[49744] = 139498035;
assign addr[49745] = 120410361;
assign addr[49746] = 101313138;
assign addr[49747] = 82207882;
assign addr[49748] = 63096108;
assign addr[49749] = 43979330;
assign addr[49750] = 24859065;
assign addr[49751] = 5736829;
assign addr[49752] = -13385863;
assign addr[49753] = -32507492;
assign addr[49754] = -51626544;
assign addr[49755] = -70741503;
assign addr[49756] = -89850852;
assign addr[49757] = -108953076;
assign addr[49758] = -128046661;
assign addr[49759] = -147130093;
assign addr[49760] = -166201858;
assign addr[49761] = -185260444;
assign addr[49762] = -204304341;
assign addr[49763] = -223332037;
assign addr[49764] = -242342025;
assign addr[49765] = -261332796;
assign addr[49766] = -280302845;
assign addr[49767] = -299250668;
assign addr[49768] = -318174762;
assign addr[49769] = -337073627;
assign addr[49770] = -355945764;
assign addr[49771] = -374789676;
assign addr[49772] = -393603870;
assign addr[49773] = -412386854;
assign addr[49774] = -431137138;
assign addr[49775] = -449853235;
assign addr[49776] = -468533662;
assign addr[49777] = -487176937;
assign addr[49778] = -505781581;
assign addr[49779] = -524346121;
assign addr[49780] = -542869083;
assign addr[49781] = -561348998;
assign addr[49782] = -579784402;
assign addr[49783] = -598173833;
assign addr[49784] = -616515832;
assign addr[49785] = -634808946;
assign addr[49786] = -653051723;
assign addr[49787] = -671242716;
assign addr[49788] = -689380485;
assign addr[49789] = -707463589;
assign addr[49790] = -725490597;
assign addr[49791] = -743460077;
assign addr[49792] = -761370605;
assign addr[49793] = -779220762;
assign addr[49794] = -797009130;
assign addr[49795] = -814734301;
assign addr[49796] = -832394869;
assign addr[49797] = -849989433;
assign addr[49798] = -867516597;
assign addr[49799] = -884974973;
assign addr[49800] = -902363176;
assign addr[49801] = -919679827;
assign addr[49802] = -936923553;
assign addr[49803] = -954092986;
assign addr[49804] = -971186766;
assign addr[49805] = -988203537;
assign addr[49806] = -1005141949;
assign addr[49807] = -1022000660;
assign addr[49808] = -1038778332;
assign addr[49809] = -1055473635;
assign addr[49810] = -1072085246;
assign addr[49811] = -1088611847;
assign addr[49812] = -1105052128;
assign addr[49813] = -1121404785;
assign addr[49814] = -1137668521;
assign addr[49815] = -1153842047;
assign addr[49816] = -1169924081;
assign addr[49817] = -1185913346;
assign addr[49818] = -1201808576;
assign addr[49819] = -1217608510;
assign addr[49820] = -1233311895;
assign addr[49821] = -1248917486;
assign addr[49822] = -1264424045;
assign addr[49823] = -1279830344;
assign addr[49824] = -1295135159;
assign addr[49825] = -1310337279;
assign addr[49826] = -1325435496;
assign addr[49827] = -1340428615;
assign addr[49828] = -1355315445;
assign addr[49829] = -1370094808;
assign addr[49830] = -1384765530;
assign addr[49831] = -1399326449;
assign addr[49832] = -1413776410;
assign addr[49833] = -1428114267;
assign addr[49834] = -1442338884;
assign addr[49835] = -1456449131;
assign addr[49836] = -1470443891;
assign addr[49837] = -1484322054;
assign addr[49838] = -1498082520;
assign addr[49839] = -1511724196;
assign addr[49840] = -1525246002;
assign addr[49841] = -1538646865;
assign addr[49842] = -1551925723;
assign addr[49843] = -1565081523;
assign addr[49844] = -1578113222;
assign addr[49845] = -1591019785;
assign addr[49846] = -1603800191;
assign addr[49847] = -1616453425;
assign addr[49848] = -1628978484;
assign addr[49849] = -1641374375;
assign addr[49850] = -1653640115;
assign addr[49851] = -1665774731;
assign addr[49852] = -1677777262;
assign addr[49853] = -1689646755;
assign addr[49854] = -1701382270;
assign addr[49855] = -1712982875;
assign addr[49856] = -1724447652;
assign addr[49857] = -1735775690;
assign addr[49858] = -1746966091;
assign addr[49859] = -1758017969;
assign addr[49860] = -1768930447;
assign addr[49861] = -1779702660;
assign addr[49862] = -1790333753;
assign addr[49863] = -1800822883;
assign addr[49864] = -1811169220;
assign addr[49865] = -1821371941;
assign addr[49866] = -1831430239;
assign addr[49867] = -1841343316;
assign addr[49868] = -1851110385;
assign addr[49869] = -1860730673;
assign addr[49870] = -1870203416;
assign addr[49871] = -1879527863;
assign addr[49872] = -1888703276;
assign addr[49873] = -1897728925;
assign addr[49874] = -1906604097;
assign addr[49875] = -1915328086;
assign addr[49876] = -1923900201;
assign addr[49877] = -1932319763;
assign addr[49878] = -1940586104;
assign addr[49879] = -1948698568;
assign addr[49880] = -1956656513;
assign addr[49881] = -1964459306;
assign addr[49882] = -1972106330;
assign addr[49883] = -1979596978;
assign addr[49884] = -1986930656;
assign addr[49885] = -1994106782;
assign addr[49886] = -2001124788;
assign addr[49887] = -2007984117;
assign addr[49888] = -2014684225;
assign addr[49889] = -2021224581;
assign addr[49890] = -2027604666;
assign addr[49891] = -2033823974;
assign addr[49892] = -2039882013;
assign addr[49893] = -2045778302;
assign addr[49894] = -2051512372;
assign addr[49895] = -2057083771;
assign addr[49896] = -2062492055;
assign addr[49897] = -2067736796;
assign addr[49898] = -2072817579;
assign addr[49899] = -2077733999;
assign addr[49900] = -2082485668;
assign addr[49901] = -2087072209;
assign addr[49902] = -2091493257;
assign addr[49903] = -2095748463;
assign addr[49904] = -2099837489;
assign addr[49905] = -2103760010;
assign addr[49906] = -2107515716;
assign addr[49907] = -2111104309;
assign addr[49908] = -2114525505;
assign addr[49909] = -2117779031;
assign addr[49910] = -2120864631;
assign addr[49911] = -2123782059;
assign addr[49912] = -2126531084;
assign addr[49913] = -2129111488;
assign addr[49914] = -2131523066;
assign addr[49915] = -2133765628;
assign addr[49916] = -2135838995;
assign addr[49917] = -2137743003;
assign addr[49918] = -2139477502;
assign addr[49919] = -2141042352;
assign addr[49920] = -2142437431;
assign addr[49921] = -2143662628;
assign addr[49922] = -2144717846;
assign addr[49923] = -2145603001;
assign addr[49924] = -2146318022;
assign addr[49925] = -2146862854;
assign addr[49926] = -2147237452;
assign addr[49927] = -2147441787;
assign addr[49928] = -2147475844;
assign addr[49929] = -2147339619;
assign addr[49930] = -2147033123;
assign addr[49931] = -2146556380;
assign addr[49932] = -2145909429;
assign addr[49933] = -2145092320;
assign addr[49934] = -2144105118;
assign addr[49935] = -2142947902;
assign addr[49936] = -2141620763;
assign addr[49937] = -2140123807;
assign addr[49938] = -2138457152;
assign addr[49939] = -2136620930;
assign addr[49940] = -2134615288;
assign addr[49941] = -2132440383;
assign addr[49942] = -2130096389;
assign addr[49943] = -2127583492;
assign addr[49944] = -2124901890;
assign addr[49945] = -2122051796;
assign addr[49946] = -2119033436;
assign addr[49947] = -2115847050;
assign addr[49948] = -2112492891;
assign addr[49949] = -2108971223;
assign addr[49950] = -2105282327;
assign addr[49951] = -2101426496;
assign addr[49952] = -2097404033;
assign addr[49953] = -2093215260;
assign addr[49954] = -2088860507;
assign addr[49955] = -2084340120;
assign addr[49956] = -2079654458;
assign addr[49957] = -2074803892;
assign addr[49958] = -2069788807;
assign addr[49959] = -2064609600;
assign addr[49960] = -2059266683;
assign addr[49961] = -2053760478;
assign addr[49962] = -2048091422;
assign addr[49963] = -2042259965;
assign addr[49964] = -2036266570;
assign addr[49965] = -2030111710;
assign addr[49966] = -2023795876;
assign addr[49967] = -2017319567;
assign addr[49968] = -2010683297;
assign addr[49969] = -2003887591;
assign addr[49970] = -1996932990;
assign addr[49971] = -1989820044;
assign addr[49972] = -1982549318;
assign addr[49973] = -1975121388;
assign addr[49974] = -1967536842;
assign addr[49975] = -1959796283;
assign addr[49976] = -1951900324;
assign addr[49977] = -1943849591;
assign addr[49978] = -1935644723;
assign addr[49979] = -1927286370;
assign addr[49980] = -1918775195;
assign addr[49981] = -1910111873;
assign addr[49982] = -1901297091;
assign addr[49983] = -1892331547;
assign addr[49984] = -1883215953;
assign addr[49985] = -1873951032;
assign addr[49986] = -1864537518;
assign addr[49987] = -1854976157;
assign addr[49988] = -1845267708;
assign addr[49989] = -1835412941;
assign addr[49990] = -1825412636;
assign addr[49991] = -1815267588;
assign addr[49992] = -1804978599;
assign addr[49993] = -1794546487;
assign addr[49994] = -1783972079;
assign addr[49995] = -1773256212;
assign addr[49996] = -1762399737;
assign addr[49997] = -1751403515;
assign addr[49998] = -1740268417;
assign addr[49999] = -1728995326;
assign addr[50000] = -1717585136;
assign addr[50001] = -1706038753;
assign addr[50002] = -1694357091;
assign addr[50003] = -1682541077;
assign addr[50004] = -1670591647;
assign addr[50005] = -1658509750;
assign addr[50006] = -1646296344;
assign addr[50007] = -1633952396;
assign addr[50008] = -1621478885;
assign addr[50009] = -1608876801;
assign addr[50010] = -1596147143;
assign addr[50011] = -1583290921;
assign addr[50012] = -1570309153;
assign addr[50013] = -1557202869;
assign addr[50014] = -1543973108;
assign addr[50015] = -1530620920;
assign addr[50016] = -1517147363;
assign addr[50017] = -1503553506;
assign addr[50018] = -1489840425;
assign addr[50019] = -1476009210;
assign addr[50020] = -1462060956;
assign addr[50021] = -1447996770;
assign addr[50022] = -1433817766;
assign addr[50023] = -1419525069;
assign addr[50024] = -1405119813;
assign addr[50025] = -1390603139;
assign addr[50026] = -1375976199;
assign addr[50027] = -1361240152;
assign addr[50028] = -1346396168;
assign addr[50029] = -1331445422;
assign addr[50030] = -1316389101;
assign addr[50031] = -1301228398;
assign addr[50032] = -1285964516;
assign addr[50033] = -1270598665;
assign addr[50034] = -1255132063;
assign addr[50035] = -1239565936;
assign addr[50036] = -1223901520;
assign addr[50037] = -1208140056;
assign addr[50038] = -1192282793;
assign addr[50039] = -1176330990;
assign addr[50040] = -1160285911;
assign addr[50041] = -1144148829;
assign addr[50042] = -1127921022;
assign addr[50043] = -1111603778;
assign addr[50044] = -1095198391;
assign addr[50045] = -1078706161;
assign addr[50046] = -1062128397;
assign addr[50047] = -1045466412;
assign addr[50048] = -1028721528;
assign addr[50049] = -1011895073;
assign addr[50050] = -994988380;
assign addr[50051] = -978002791;
assign addr[50052] = -960939653;
assign addr[50053] = -943800318;
assign addr[50054] = -926586145;
assign addr[50055] = -909298500;
assign addr[50056] = -891938752;
assign addr[50057] = -874508280;
assign addr[50058] = -857008464;
assign addr[50059] = -839440693;
assign addr[50060] = -821806359;
assign addr[50061] = -804106861;
assign addr[50062] = -786343603;
assign addr[50063] = -768517992;
assign addr[50064] = -750631442;
assign addr[50065] = -732685372;
assign addr[50066] = -714681204;
assign addr[50067] = -696620367;
assign addr[50068] = -678504291;
assign addr[50069] = -660334415;
assign addr[50070] = -642112178;
assign addr[50071] = -623839025;
assign addr[50072] = -605516406;
assign addr[50073] = -587145773;
assign addr[50074] = -568728583;
assign addr[50075] = -550266296;
assign addr[50076] = -531760377;
assign addr[50077] = -513212292;
assign addr[50078] = -494623513;
assign addr[50079] = -475995513;
assign addr[50080] = -457329769;
assign addr[50081] = -438627762;
assign addr[50082] = -419890975;
assign addr[50083] = -401120892;
assign addr[50084] = -382319004;
assign addr[50085] = -363486799;
assign addr[50086] = -344625773;
assign addr[50087] = -325737419;
assign addr[50088] = -306823237;
assign addr[50089] = -287884725;
assign addr[50090] = -268923386;
assign addr[50091] = -249940723;
assign addr[50092] = -230938242;
assign addr[50093] = -211917448;
assign addr[50094] = -192879850;
assign addr[50095] = -173826959;
assign addr[50096] = -154760284;
assign addr[50097] = -135681337;
assign addr[50098] = -116591632;
assign addr[50099] = -97492681;
assign addr[50100] = -78386000;
assign addr[50101] = -59273104;
assign addr[50102] = -40155507;
assign addr[50103] = -21034727;
assign addr[50104] = -1912278;
assign addr[50105] = 17210322;
assign addr[50106] = 36331557;
assign addr[50107] = 55449912;
assign addr[50108] = 74563870;
assign addr[50109] = 93671915;
assign addr[50110] = 112772533;
assign addr[50111] = 131864208;
assign addr[50112] = 150945428;
assign addr[50113] = 170014678;
assign addr[50114] = 189070447;
assign addr[50115] = 208111224;
assign addr[50116] = 227135500;
assign addr[50117] = 246141764;
assign addr[50118] = 265128512;
assign addr[50119] = 284094236;
assign addr[50120] = 303037433;
assign addr[50121] = 321956601;
assign addr[50122] = 340850240;
assign addr[50123] = 359716852;
assign addr[50124] = 378554940;
assign addr[50125] = 397363011;
assign addr[50126] = 416139574;
assign addr[50127] = 434883140;
assign addr[50128] = 453592221;
assign addr[50129] = 472265336;
assign addr[50130] = 490901003;
assign addr[50131] = 509497745;
assign addr[50132] = 528054086;
assign addr[50133] = 546568556;
assign addr[50134] = 565039687;
assign addr[50135] = 583466013;
assign addr[50136] = 601846074;
assign addr[50137] = 620178412;
assign addr[50138] = 638461574;
assign addr[50139] = 656694110;
assign addr[50140] = 674874574;
assign addr[50141] = 693001525;
assign addr[50142] = 711073524;
assign addr[50143] = 729089140;
assign addr[50144] = 747046944;
assign addr[50145] = 764945512;
assign addr[50146] = 782783424;
assign addr[50147] = 800559266;
assign addr[50148] = 818271628;
assign addr[50149] = 835919107;
assign addr[50150] = 853500302;
assign addr[50151] = 871013820;
assign addr[50152] = 888458272;
assign addr[50153] = 905832274;
assign addr[50154] = 923134450;
assign addr[50155] = 940363427;
assign addr[50156] = 957517838;
assign addr[50157] = 974596324;
assign addr[50158] = 991597531;
assign addr[50159] = 1008520110;
assign addr[50160] = 1025362720;
assign addr[50161] = 1042124025;
assign addr[50162] = 1058802695;
assign addr[50163] = 1075397409;
assign addr[50164] = 1091906851;
assign addr[50165] = 1108329711;
assign addr[50166] = 1124664687;
assign addr[50167] = 1140910484;
assign addr[50168] = 1157065814;
assign addr[50169] = 1173129396;
assign addr[50170] = 1189099956;
assign addr[50171] = 1204976227;
assign addr[50172] = 1220756951;
assign addr[50173] = 1236440877;
assign addr[50174] = 1252026760;
assign addr[50175] = 1267513365;
assign addr[50176] = 1282899464;
assign addr[50177] = 1298183838;
assign addr[50178] = 1313365273;
assign addr[50179] = 1328442566;
assign addr[50180] = 1343414522;
assign addr[50181] = 1358279953;
assign addr[50182] = 1373037681;
assign addr[50183] = 1387686535;
assign addr[50184] = 1402225355;
assign addr[50185] = 1416652986;
assign addr[50186] = 1430968286;
assign addr[50187] = 1445170118;
assign addr[50188] = 1459257358;
assign addr[50189] = 1473228887;
assign addr[50190] = 1487083598;
assign addr[50191] = 1500820393;
assign addr[50192] = 1514438181;
assign addr[50193] = 1527935884;
assign addr[50194] = 1541312431;
assign addr[50195] = 1554566762;
assign addr[50196] = 1567697824;
assign addr[50197] = 1580704578;
assign addr[50198] = 1593585992;
assign addr[50199] = 1606341043;
assign addr[50200] = 1618968722;
assign addr[50201] = 1631468027;
assign addr[50202] = 1643837966;
assign addr[50203] = 1656077559;
assign addr[50204] = 1668185835;
assign addr[50205] = 1680161834;
assign addr[50206] = 1692004606;
assign addr[50207] = 1703713213;
assign addr[50208] = 1715286726;
assign addr[50209] = 1726724227;
assign addr[50210] = 1738024810;
assign addr[50211] = 1749187577;
assign addr[50212] = 1760211645;
assign addr[50213] = 1771096139;
assign addr[50214] = 1781840195;
assign addr[50215] = 1792442963;
assign addr[50216] = 1802903601;
assign addr[50217] = 1813221279;
assign addr[50218] = 1823395180;
assign addr[50219] = 1833424497;
assign addr[50220] = 1843308435;
assign addr[50221] = 1853046210;
assign addr[50222] = 1862637049;
assign addr[50223] = 1872080193;
assign addr[50224] = 1881374892;
assign addr[50225] = 1890520410;
assign addr[50226] = 1899516021;
assign addr[50227] = 1908361011;
assign addr[50228] = 1917054681;
assign addr[50229] = 1925596340;
assign addr[50230] = 1933985310;
assign addr[50231] = 1942220928;
assign addr[50232] = 1950302539;
assign addr[50233] = 1958229503;
assign addr[50234] = 1966001192;
assign addr[50235] = 1973616989;
assign addr[50236] = 1981076290;
assign addr[50237] = 1988378503;
assign addr[50238] = 1995523051;
assign addr[50239] = 2002509365;
assign addr[50240] = 2009336893;
assign addr[50241] = 2016005093;
assign addr[50242] = 2022513436;
assign addr[50243] = 2028861406;
assign addr[50244] = 2035048499;
assign addr[50245] = 2041074226;
assign addr[50246] = 2046938108;
assign addr[50247] = 2052639680;
assign addr[50248] = 2058178491;
assign addr[50249] = 2063554100;
assign addr[50250] = 2068766083;
assign addr[50251] = 2073814024;
assign addr[50252] = 2078697525;
assign addr[50253] = 2083416198;
assign addr[50254] = 2087969669;
assign addr[50255] = 2092357577;
assign addr[50256] = 2096579573;
assign addr[50257] = 2100635323;
assign addr[50258] = 2104524506;
assign addr[50259] = 2108246813;
assign addr[50260] = 2111801949;
assign addr[50261] = 2115189632;
assign addr[50262] = 2118409593;
assign addr[50263] = 2121461578;
assign addr[50264] = 2124345343;
assign addr[50265] = 2127060661;
assign addr[50266] = 2129607316;
assign addr[50267] = 2131985106;
assign addr[50268] = 2134193842;
assign addr[50269] = 2136233350;
assign addr[50270] = 2138103468;
assign addr[50271] = 2139804048;
assign addr[50272] = 2141334954;
assign addr[50273] = 2142696065;
assign addr[50274] = 2143887273;
assign addr[50275] = 2144908484;
assign addr[50276] = 2145759618;
assign addr[50277] = 2146440605;
assign addr[50278] = 2146951393;
assign addr[50279] = 2147291941;
assign addr[50280] = 2147462221;
assign addr[50281] = 2147462221;
assign addr[50282] = 2147291941;
assign addr[50283] = 2146951393;
assign addr[50284] = 2146440605;
assign addr[50285] = 2145759618;
assign addr[50286] = 2144908484;
assign addr[50287] = 2143887273;
assign addr[50288] = 2142696065;
assign addr[50289] = 2141334954;
assign addr[50290] = 2139804048;
assign addr[50291] = 2138103468;
assign addr[50292] = 2136233350;
assign addr[50293] = 2134193842;
assign addr[50294] = 2131985106;
assign addr[50295] = 2129607316;
assign addr[50296] = 2127060661;
assign addr[50297] = 2124345343;
assign addr[50298] = 2121461578;
assign addr[50299] = 2118409593;
assign addr[50300] = 2115189632;
assign addr[50301] = 2111801949;
assign addr[50302] = 2108246813;
assign addr[50303] = 2104524506;
assign addr[50304] = 2100635323;
assign addr[50305] = 2096579573;
assign addr[50306] = 2092357577;
assign addr[50307] = 2087969669;
assign addr[50308] = 2083416198;
assign addr[50309] = 2078697525;
assign addr[50310] = 2073814024;
assign addr[50311] = 2068766083;
assign addr[50312] = 2063554100;
assign addr[50313] = 2058178491;
assign addr[50314] = 2052639680;
assign addr[50315] = 2046938108;
assign addr[50316] = 2041074226;
assign addr[50317] = 2035048499;
assign addr[50318] = 2028861406;
assign addr[50319] = 2022513436;
assign addr[50320] = 2016005093;
assign addr[50321] = 2009336893;
assign addr[50322] = 2002509365;
assign addr[50323] = 1995523051;
assign addr[50324] = 1988378503;
assign addr[50325] = 1981076290;
assign addr[50326] = 1973616989;
assign addr[50327] = 1966001192;
assign addr[50328] = 1958229503;
assign addr[50329] = 1950302539;
assign addr[50330] = 1942220928;
assign addr[50331] = 1933985310;
assign addr[50332] = 1925596340;
assign addr[50333] = 1917054681;
assign addr[50334] = 1908361011;
assign addr[50335] = 1899516021;
assign addr[50336] = 1890520410;
assign addr[50337] = 1881374892;
assign addr[50338] = 1872080193;
assign addr[50339] = 1862637049;
assign addr[50340] = 1853046210;
assign addr[50341] = 1843308435;
assign addr[50342] = 1833424497;
assign addr[50343] = 1823395180;
assign addr[50344] = 1813221279;
assign addr[50345] = 1802903601;
assign addr[50346] = 1792442963;
assign addr[50347] = 1781840195;
assign addr[50348] = 1771096139;
assign addr[50349] = 1760211645;
assign addr[50350] = 1749187577;
assign addr[50351] = 1738024810;
assign addr[50352] = 1726724227;
assign addr[50353] = 1715286726;
assign addr[50354] = 1703713213;
assign addr[50355] = 1692004606;
assign addr[50356] = 1680161834;
assign addr[50357] = 1668185835;
assign addr[50358] = 1656077559;
assign addr[50359] = 1643837966;
assign addr[50360] = 1631468027;
assign addr[50361] = 1618968722;
assign addr[50362] = 1606341043;
assign addr[50363] = 1593585992;
assign addr[50364] = 1580704578;
assign addr[50365] = 1567697824;
assign addr[50366] = 1554566762;
assign addr[50367] = 1541312431;
assign addr[50368] = 1527935884;
assign addr[50369] = 1514438181;
assign addr[50370] = 1500820393;
assign addr[50371] = 1487083598;
assign addr[50372] = 1473228887;
assign addr[50373] = 1459257358;
assign addr[50374] = 1445170118;
assign addr[50375] = 1430968286;
assign addr[50376] = 1416652986;
assign addr[50377] = 1402225355;
assign addr[50378] = 1387686535;
assign addr[50379] = 1373037681;
assign addr[50380] = 1358279953;
assign addr[50381] = 1343414522;
assign addr[50382] = 1328442566;
assign addr[50383] = 1313365273;
assign addr[50384] = 1298183838;
assign addr[50385] = 1282899464;
assign addr[50386] = 1267513365;
assign addr[50387] = 1252026760;
assign addr[50388] = 1236440877;
assign addr[50389] = 1220756951;
assign addr[50390] = 1204976227;
assign addr[50391] = 1189099956;
assign addr[50392] = 1173129396;
assign addr[50393] = 1157065814;
assign addr[50394] = 1140910484;
assign addr[50395] = 1124664687;
assign addr[50396] = 1108329711;
assign addr[50397] = 1091906851;
assign addr[50398] = 1075397409;
assign addr[50399] = 1058802695;
assign addr[50400] = 1042124025;
assign addr[50401] = 1025362720;
assign addr[50402] = 1008520110;
assign addr[50403] = 991597531;
assign addr[50404] = 974596324;
assign addr[50405] = 957517838;
assign addr[50406] = 940363427;
assign addr[50407] = 923134450;
assign addr[50408] = 905832274;
assign addr[50409] = 888458272;
assign addr[50410] = 871013820;
assign addr[50411] = 853500302;
assign addr[50412] = 835919107;
assign addr[50413] = 818271628;
assign addr[50414] = 800559266;
assign addr[50415] = 782783424;
assign addr[50416] = 764945512;
assign addr[50417] = 747046944;
assign addr[50418] = 729089140;
assign addr[50419] = 711073524;
assign addr[50420] = 693001525;
assign addr[50421] = 674874574;
assign addr[50422] = 656694110;
assign addr[50423] = 638461574;
assign addr[50424] = 620178412;
assign addr[50425] = 601846074;
assign addr[50426] = 583466013;
assign addr[50427] = 565039687;
assign addr[50428] = 546568556;
assign addr[50429] = 528054086;
assign addr[50430] = 509497745;
assign addr[50431] = 490901003;
assign addr[50432] = 472265336;
assign addr[50433] = 453592221;
assign addr[50434] = 434883140;
assign addr[50435] = 416139574;
assign addr[50436] = 397363011;
assign addr[50437] = 378554940;
assign addr[50438] = 359716852;
assign addr[50439] = 340850240;
assign addr[50440] = 321956601;
assign addr[50441] = 303037433;
assign addr[50442] = 284094236;
assign addr[50443] = 265128512;
assign addr[50444] = 246141764;
assign addr[50445] = 227135500;
assign addr[50446] = 208111224;
assign addr[50447] = 189070447;
assign addr[50448] = 170014678;
assign addr[50449] = 150945428;
assign addr[50450] = 131864208;
assign addr[50451] = 112772533;
assign addr[50452] = 93671915;
assign addr[50453] = 74563870;
assign addr[50454] = 55449912;
assign addr[50455] = 36331557;
assign addr[50456] = 17210322;
assign addr[50457] = -1912278;
assign addr[50458] = -21034727;
assign addr[50459] = -40155507;
assign addr[50460] = -59273104;
assign addr[50461] = -78386000;
assign addr[50462] = -97492681;
assign addr[50463] = -116591632;
assign addr[50464] = -135681337;
assign addr[50465] = -154760284;
assign addr[50466] = -173826959;
assign addr[50467] = -192879850;
assign addr[50468] = -211917448;
assign addr[50469] = -230938242;
assign addr[50470] = -249940723;
assign addr[50471] = -268923386;
assign addr[50472] = -287884725;
assign addr[50473] = -306823237;
assign addr[50474] = -325737419;
assign addr[50475] = -344625773;
assign addr[50476] = -363486799;
assign addr[50477] = -382319004;
assign addr[50478] = -401120892;
assign addr[50479] = -419890975;
assign addr[50480] = -438627762;
assign addr[50481] = -457329769;
assign addr[50482] = -475995513;
assign addr[50483] = -494623513;
assign addr[50484] = -513212292;
assign addr[50485] = -531760377;
assign addr[50486] = -550266296;
assign addr[50487] = -568728583;
assign addr[50488] = -587145773;
assign addr[50489] = -605516406;
assign addr[50490] = -623839025;
assign addr[50491] = -642112178;
assign addr[50492] = -660334415;
assign addr[50493] = -678504291;
assign addr[50494] = -696620367;
assign addr[50495] = -714681204;
assign addr[50496] = -732685372;
assign addr[50497] = -750631442;
assign addr[50498] = -768517992;
assign addr[50499] = -786343603;
assign addr[50500] = -804106861;
assign addr[50501] = -821806359;
assign addr[50502] = -839440693;
assign addr[50503] = -857008464;
assign addr[50504] = -874508280;
assign addr[50505] = -891938752;
assign addr[50506] = -909298500;
assign addr[50507] = -926586145;
assign addr[50508] = -943800318;
assign addr[50509] = -960939653;
assign addr[50510] = -978002791;
assign addr[50511] = -994988380;
assign addr[50512] = -1011895073;
assign addr[50513] = -1028721528;
assign addr[50514] = -1045466412;
assign addr[50515] = -1062128397;
assign addr[50516] = -1078706161;
assign addr[50517] = -1095198391;
assign addr[50518] = -1111603778;
assign addr[50519] = -1127921022;
assign addr[50520] = -1144148829;
assign addr[50521] = -1160285911;
assign addr[50522] = -1176330990;
assign addr[50523] = -1192282793;
assign addr[50524] = -1208140056;
assign addr[50525] = -1223901520;
assign addr[50526] = -1239565936;
assign addr[50527] = -1255132063;
assign addr[50528] = -1270598665;
assign addr[50529] = -1285964516;
assign addr[50530] = -1301228398;
assign addr[50531] = -1316389101;
assign addr[50532] = -1331445422;
assign addr[50533] = -1346396168;
assign addr[50534] = -1361240152;
assign addr[50535] = -1375976199;
assign addr[50536] = -1390603139;
assign addr[50537] = -1405119813;
assign addr[50538] = -1419525069;
assign addr[50539] = -1433817766;
assign addr[50540] = -1447996770;
assign addr[50541] = -1462060956;
assign addr[50542] = -1476009210;
assign addr[50543] = -1489840425;
assign addr[50544] = -1503553506;
assign addr[50545] = -1517147363;
assign addr[50546] = -1530620920;
assign addr[50547] = -1543973108;
assign addr[50548] = -1557202869;
assign addr[50549] = -1570309153;
assign addr[50550] = -1583290921;
assign addr[50551] = -1596147143;
assign addr[50552] = -1608876801;
assign addr[50553] = -1621478885;
assign addr[50554] = -1633952396;
assign addr[50555] = -1646296344;
assign addr[50556] = -1658509750;
assign addr[50557] = -1670591647;
assign addr[50558] = -1682541077;
assign addr[50559] = -1694357091;
assign addr[50560] = -1706038753;
assign addr[50561] = -1717585136;
assign addr[50562] = -1728995326;
assign addr[50563] = -1740268417;
assign addr[50564] = -1751403515;
assign addr[50565] = -1762399737;
assign addr[50566] = -1773256212;
assign addr[50567] = -1783972079;
assign addr[50568] = -1794546487;
assign addr[50569] = -1804978599;
assign addr[50570] = -1815267588;
assign addr[50571] = -1825412636;
assign addr[50572] = -1835412941;
assign addr[50573] = -1845267708;
assign addr[50574] = -1854976157;
assign addr[50575] = -1864537518;
assign addr[50576] = -1873951032;
assign addr[50577] = -1883215953;
assign addr[50578] = -1892331547;
assign addr[50579] = -1901297091;
assign addr[50580] = -1910111873;
assign addr[50581] = -1918775195;
assign addr[50582] = -1927286370;
assign addr[50583] = -1935644723;
assign addr[50584] = -1943849591;
assign addr[50585] = -1951900324;
assign addr[50586] = -1959796283;
assign addr[50587] = -1967536842;
assign addr[50588] = -1975121388;
assign addr[50589] = -1982549318;
assign addr[50590] = -1989820044;
assign addr[50591] = -1996932990;
assign addr[50592] = -2003887591;
assign addr[50593] = -2010683297;
assign addr[50594] = -2017319567;
assign addr[50595] = -2023795876;
assign addr[50596] = -2030111710;
assign addr[50597] = -2036266570;
assign addr[50598] = -2042259965;
assign addr[50599] = -2048091422;
assign addr[50600] = -2053760478;
assign addr[50601] = -2059266683;
assign addr[50602] = -2064609600;
assign addr[50603] = -2069788807;
assign addr[50604] = -2074803892;
assign addr[50605] = -2079654458;
assign addr[50606] = -2084340120;
assign addr[50607] = -2088860507;
assign addr[50608] = -2093215260;
assign addr[50609] = -2097404033;
assign addr[50610] = -2101426496;
assign addr[50611] = -2105282327;
assign addr[50612] = -2108971223;
assign addr[50613] = -2112492891;
assign addr[50614] = -2115847050;
assign addr[50615] = -2119033436;
assign addr[50616] = -2122051796;
assign addr[50617] = -2124901890;
assign addr[50618] = -2127583492;
assign addr[50619] = -2130096389;
assign addr[50620] = -2132440383;
assign addr[50621] = -2134615288;
assign addr[50622] = -2136620930;
assign addr[50623] = -2138457152;
assign addr[50624] = -2140123807;
assign addr[50625] = -2141620763;
assign addr[50626] = -2142947902;
assign addr[50627] = -2144105118;
assign addr[50628] = -2145092320;
assign addr[50629] = -2145909429;
assign addr[50630] = -2146556380;
assign addr[50631] = -2147033123;
assign addr[50632] = -2147339619;
assign addr[50633] = -2147475844;
assign addr[50634] = -2147441787;
assign addr[50635] = -2147237452;
assign addr[50636] = -2146862854;
assign addr[50637] = -2146318022;
assign addr[50638] = -2145603001;
assign addr[50639] = -2144717846;
assign addr[50640] = -2143662628;
assign addr[50641] = -2142437431;
assign addr[50642] = -2141042352;
assign addr[50643] = -2139477502;
assign addr[50644] = -2137743003;
assign addr[50645] = -2135838995;
assign addr[50646] = -2133765628;
assign addr[50647] = -2131523066;
assign addr[50648] = -2129111488;
assign addr[50649] = -2126531084;
assign addr[50650] = -2123782059;
assign addr[50651] = -2120864631;
assign addr[50652] = -2117779031;
assign addr[50653] = -2114525505;
assign addr[50654] = -2111104309;
assign addr[50655] = -2107515716;
assign addr[50656] = -2103760010;
assign addr[50657] = -2099837489;
assign addr[50658] = -2095748463;
assign addr[50659] = -2091493257;
assign addr[50660] = -2087072209;
assign addr[50661] = -2082485668;
assign addr[50662] = -2077733999;
assign addr[50663] = -2072817579;
assign addr[50664] = -2067736796;
assign addr[50665] = -2062492055;
assign addr[50666] = -2057083771;
assign addr[50667] = -2051512372;
assign addr[50668] = -2045778302;
assign addr[50669] = -2039882013;
assign addr[50670] = -2033823974;
assign addr[50671] = -2027604666;
assign addr[50672] = -2021224581;
assign addr[50673] = -2014684225;
assign addr[50674] = -2007984117;
assign addr[50675] = -2001124788;
assign addr[50676] = -1994106782;
assign addr[50677] = -1986930656;
assign addr[50678] = -1979596978;
assign addr[50679] = -1972106330;
assign addr[50680] = -1964459306;
assign addr[50681] = -1956656513;
assign addr[50682] = -1948698568;
assign addr[50683] = -1940586104;
assign addr[50684] = -1932319763;
assign addr[50685] = -1923900201;
assign addr[50686] = -1915328086;
assign addr[50687] = -1906604097;
assign addr[50688] = -1897728925;
assign addr[50689] = -1888703276;
assign addr[50690] = -1879527863;
assign addr[50691] = -1870203416;
assign addr[50692] = -1860730673;
assign addr[50693] = -1851110385;
assign addr[50694] = -1841343316;
assign addr[50695] = -1831430239;
assign addr[50696] = -1821371941;
assign addr[50697] = -1811169220;
assign addr[50698] = -1800822883;
assign addr[50699] = -1790333753;
assign addr[50700] = -1779702660;
assign addr[50701] = -1768930447;
assign addr[50702] = -1758017969;
assign addr[50703] = -1746966091;
assign addr[50704] = -1735775690;
assign addr[50705] = -1724447652;
assign addr[50706] = -1712982875;
assign addr[50707] = -1701382270;
assign addr[50708] = -1689646755;
assign addr[50709] = -1677777262;
assign addr[50710] = -1665774731;
assign addr[50711] = -1653640115;
assign addr[50712] = -1641374375;
assign addr[50713] = -1628978484;
assign addr[50714] = -1616453425;
assign addr[50715] = -1603800191;
assign addr[50716] = -1591019785;
assign addr[50717] = -1578113222;
assign addr[50718] = -1565081523;
assign addr[50719] = -1551925723;
assign addr[50720] = -1538646865;
assign addr[50721] = -1525246002;
assign addr[50722] = -1511724196;
assign addr[50723] = -1498082520;
assign addr[50724] = -1484322054;
assign addr[50725] = -1470443891;
assign addr[50726] = -1456449131;
assign addr[50727] = -1442338884;
assign addr[50728] = -1428114267;
assign addr[50729] = -1413776410;
assign addr[50730] = -1399326449;
assign addr[50731] = -1384765530;
assign addr[50732] = -1370094808;
assign addr[50733] = -1355315445;
assign addr[50734] = -1340428615;
assign addr[50735] = -1325435496;
assign addr[50736] = -1310337279;
assign addr[50737] = -1295135159;
assign addr[50738] = -1279830344;
assign addr[50739] = -1264424045;
assign addr[50740] = -1248917486;
assign addr[50741] = -1233311895;
assign addr[50742] = -1217608510;
assign addr[50743] = -1201808576;
assign addr[50744] = -1185913346;
assign addr[50745] = -1169924081;
assign addr[50746] = -1153842047;
assign addr[50747] = -1137668521;
assign addr[50748] = -1121404785;
assign addr[50749] = -1105052128;
assign addr[50750] = -1088611847;
assign addr[50751] = -1072085246;
assign addr[50752] = -1055473635;
assign addr[50753] = -1038778332;
assign addr[50754] = -1022000660;
assign addr[50755] = -1005141949;
assign addr[50756] = -988203537;
assign addr[50757] = -971186766;
assign addr[50758] = -954092986;
assign addr[50759] = -936923553;
assign addr[50760] = -919679827;
assign addr[50761] = -902363176;
assign addr[50762] = -884974973;
assign addr[50763] = -867516597;
assign addr[50764] = -849989433;
assign addr[50765] = -832394869;
assign addr[50766] = -814734301;
assign addr[50767] = -797009130;
assign addr[50768] = -779220762;
assign addr[50769] = -761370605;
assign addr[50770] = -743460077;
assign addr[50771] = -725490597;
assign addr[50772] = -707463589;
assign addr[50773] = -689380485;
assign addr[50774] = -671242716;
assign addr[50775] = -653051723;
assign addr[50776] = -634808946;
assign addr[50777] = -616515832;
assign addr[50778] = -598173833;
assign addr[50779] = -579784402;
assign addr[50780] = -561348998;
assign addr[50781] = -542869083;
assign addr[50782] = -524346121;
assign addr[50783] = -505781581;
assign addr[50784] = -487176937;
assign addr[50785] = -468533662;
assign addr[50786] = -449853235;
assign addr[50787] = -431137138;
assign addr[50788] = -412386854;
assign addr[50789] = -393603870;
assign addr[50790] = -374789676;
assign addr[50791] = -355945764;
assign addr[50792] = -337073627;
assign addr[50793] = -318174762;
assign addr[50794] = -299250668;
assign addr[50795] = -280302845;
assign addr[50796] = -261332796;
assign addr[50797] = -242342025;
assign addr[50798] = -223332037;
assign addr[50799] = -204304341;
assign addr[50800] = -185260444;
assign addr[50801] = -166201858;
assign addr[50802] = -147130093;
assign addr[50803] = -128046661;
assign addr[50804] = -108953076;
assign addr[50805] = -89850852;
assign addr[50806] = -70741503;
assign addr[50807] = -51626544;
assign addr[50808] = -32507492;
assign addr[50809] = -13385863;
assign addr[50810] = 5736829;
assign addr[50811] = 24859065;
assign addr[50812] = 43979330;
assign addr[50813] = 63096108;
assign addr[50814] = 82207882;
assign addr[50815] = 101313138;
assign addr[50816] = 120410361;
assign addr[50817] = 139498035;
assign addr[50818] = 158574649;
assign addr[50819] = 177638688;
assign addr[50820] = 196688642;
assign addr[50821] = 215722999;
assign addr[50822] = 234740251;
assign addr[50823] = 253738890;
assign addr[50824] = 272717408;
assign addr[50825] = 291674302;
assign addr[50826] = 310608068;
assign addr[50827] = 329517204;
assign addr[50828] = 348400212;
assign addr[50829] = 367255594;
assign addr[50830] = 386081854;
assign addr[50831] = 404877501;
assign addr[50832] = 423641043;
assign addr[50833] = 442370993;
assign addr[50834] = 461065866;
assign addr[50835] = 479724180;
assign addr[50836] = 498344454;
assign addr[50837] = 516925212;
assign addr[50838] = 535464981;
assign addr[50839] = 553962291;
assign addr[50840] = 572415676;
assign addr[50841] = 590823671;
assign addr[50842] = 609184818;
assign addr[50843] = 627497660;
assign addr[50844] = 645760745;
assign addr[50845] = 663972625;
assign addr[50846] = 682131857;
assign addr[50847] = 700236999;
assign addr[50848] = 718286617;
assign addr[50849] = 736279279;
assign addr[50850] = 754213559;
assign addr[50851] = 772088034;
assign addr[50852] = 789901288;
assign addr[50853] = 807651907;
assign addr[50854] = 825338484;
assign addr[50855] = 842959617;
assign addr[50856] = 860513908;
assign addr[50857] = 877999966;
assign addr[50858] = 895416404;
assign addr[50859] = 912761841;
assign addr[50860] = 930034901;
assign addr[50861] = 947234215;
assign addr[50862] = 964358420;
assign addr[50863] = 981406156;
assign addr[50864] = 998376073;
assign addr[50865] = 1015266825;
assign addr[50866] = 1032077073;
assign addr[50867] = 1048805483;
assign addr[50868] = 1065450729;
assign addr[50869] = 1082011492;
assign addr[50870] = 1098486458;
assign addr[50871] = 1114874320;
assign addr[50872] = 1131173780;
assign addr[50873] = 1147383544;
assign addr[50874] = 1163502328;
assign addr[50875] = 1179528853;
assign addr[50876] = 1195461849;
assign addr[50877] = 1211300053;
assign addr[50878] = 1227042207;
assign addr[50879] = 1242687064;
assign addr[50880] = 1258233384;
assign addr[50881] = 1273679934;
assign addr[50882] = 1289025489;
assign addr[50883] = 1304268832;
assign addr[50884] = 1319408754;
assign addr[50885] = 1334444055;
assign addr[50886] = 1349373543;
assign addr[50887] = 1364196034;
assign addr[50888] = 1378910353;
assign addr[50889] = 1393515332;
assign addr[50890] = 1408009814;
assign addr[50891] = 1422392650;
assign addr[50892] = 1436662698;
assign addr[50893] = 1450818828;
assign addr[50894] = 1464859917;
assign addr[50895] = 1478784851;
assign addr[50896] = 1492592527;
assign addr[50897] = 1506281850;
assign addr[50898] = 1519851733;
assign addr[50899] = 1533301101;
assign addr[50900] = 1546628888;
assign addr[50901] = 1559834037;
assign addr[50902] = 1572915501;
assign addr[50903] = 1585872242;
assign addr[50904] = 1598703233;
assign addr[50905] = 1611407456;
assign addr[50906] = 1623983905;
assign addr[50907] = 1636431582;
assign addr[50908] = 1648749499;
assign addr[50909] = 1660936681;
assign addr[50910] = 1672992161;
assign addr[50911] = 1684914983;
assign addr[50912] = 1696704201;
assign addr[50913] = 1708358881;
assign addr[50914] = 1719878099;
assign addr[50915] = 1731260941;
assign addr[50916] = 1742506504;
assign addr[50917] = 1753613897;
assign addr[50918] = 1764582240;
assign addr[50919] = 1775410662;
assign addr[50920] = 1786098304;
assign addr[50921] = 1796644320;
assign addr[50922] = 1807047873;
assign addr[50923] = 1817308138;
assign addr[50924] = 1827424302;
assign addr[50925] = 1837395562;
assign addr[50926] = 1847221128;
assign addr[50927] = 1856900221;
assign addr[50928] = 1866432072;
assign addr[50929] = 1875815927;
assign addr[50930] = 1885051042;
assign addr[50931] = 1894136683;
assign addr[50932] = 1903072131;
assign addr[50933] = 1911856677;
assign addr[50934] = 1920489624;
assign addr[50935] = 1928970288;
assign addr[50936] = 1937297997;
assign addr[50937] = 1945472089;
assign addr[50938] = 1953491918;
assign addr[50939] = 1961356847;
assign addr[50940] = 1969066252;
assign addr[50941] = 1976619522;
assign addr[50942] = 1984016058;
assign addr[50943] = 1991255274;
assign addr[50944] = 1998336596;
assign addr[50945] = 2005259462;
assign addr[50946] = 2012023322;
assign addr[50947] = 2018627642;
assign addr[50948] = 2025071897;
assign addr[50949] = 2031355576;
assign addr[50950] = 2037478181;
assign addr[50951] = 2043439226;
assign addr[50952] = 2049238240;
assign addr[50953] = 2054874761;
assign addr[50954] = 2060348343;
assign addr[50955] = 2065658552;
assign addr[50956] = 2070804967;
assign addr[50957] = 2075787180;
assign addr[50958] = 2080604795;
assign addr[50959] = 2085257431;
assign addr[50960] = 2089744719;
assign addr[50961] = 2094066304;
assign addr[50962] = 2098221841;
assign addr[50963] = 2102211002;
assign addr[50964] = 2106033471;
assign addr[50965] = 2109688944;
assign addr[50966] = 2113177132;
assign addr[50967] = 2116497758;
assign addr[50968] = 2119650558;
assign addr[50969] = 2122635283;
assign addr[50970] = 2125451696;
assign addr[50971] = 2128099574;
assign addr[50972] = 2130578706;
assign addr[50973] = 2132888897;
assign addr[50974] = 2135029962;
assign addr[50975] = 2137001733;
assign addr[50976] = 2138804053;
assign addr[50977] = 2140436778;
assign addr[50978] = 2141899780;
assign addr[50979] = 2143192942;
assign addr[50980] = 2144316162;
assign addr[50981] = 2145269351;
assign addr[50982] = 2146052433;
assign addr[50983] = 2146665347;
assign addr[50984] = 2147108043;
assign addr[50985] = 2147380486;
assign addr[50986] = 2147482655;
assign addr[50987] = 2147414542;
assign addr[50988] = 2147176152;
assign addr[50989] = 2146767505;
assign addr[50990] = 2146188631;
assign addr[50991] = 2145439578;
assign addr[50992] = 2144520405;
assign addr[50993] = 2143431184;
assign addr[50994] = 2142172003;
assign addr[50995] = 2140742960;
assign addr[50996] = 2139144169;
assign addr[50997] = 2137375758;
assign addr[50998] = 2135437865;
assign addr[50999] = 2133330646;
assign addr[51000] = 2131054266;
assign addr[51001] = 2128608907;
assign addr[51002] = 2125994762;
assign addr[51003] = 2123212038;
assign addr[51004] = 2120260957;
assign addr[51005] = 2117141752;
assign addr[51006] = 2113854671;
assign addr[51007] = 2110399974;
assign addr[51008] = 2106777935;
assign addr[51009] = 2102988841;
assign addr[51010] = 2099032994;
assign addr[51011] = 2094910706;
assign addr[51012] = 2090622304;
assign addr[51013] = 2086168128;
assign addr[51014] = 2081548533;
assign addr[51015] = 2076763883;
assign addr[51016] = 2071814558;
assign addr[51017] = 2066700952;
assign addr[51018] = 2061423468;
assign addr[51019] = 2055982526;
assign addr[51020] = 2050378558;
assign addr[51021] = 2044612007;
assign addr[51022] = 2038683330;
assign addr[51023] = 2032592999;
assign addr[51024] = 2026341495;
assign addr[51025] = 2019929315;
assign addr[51026] = 2013356967;
assign addr[51027] = 2006624971;
assign addr[51028] = 1999733863;
assign addr[51029] = 1992684188;
assign addr[51030] = 1985476506;
assign addr[51031] = 1978111387;
assign addr[51032] = 1970589416;
assign addr[51033] = 1962911189;
assign addr[51034] = 1955077316;
assign addr[51035] = 1947088417;
assign addr[51036] = 1938945125;
assign addr[51037] = 1930648088;
assign addr[51038] = 1922197961;
assign addr[51039] = 1913595416;
assign addr[51040] = 1904841135;
assign addr[51041] = 1895935811;
assign addr[51042] = 1886880151;
assign addr[51043] = 1877674873;
assign addr[51044] = 1868320707;
assign addr[51045] = 1858818395;
assign addr[51046] = 1849168689;
assign addr[51047] = 1839372356;
assign addr[51048] = 1829430172;
assign addr[51049] = 1819342925;
assign addr[51050] = 1809111415;
assign addr[51051] = 1798736454;
assign addr[51052] = 1788218865;
assign addr[51053] = 1777559480;
assign addr[51054] = 1766759146;
assign addr[51055] = 1755818718;
assign addr[51056] = 1744739065;
assign addr[51057] = 1733521064;
assign addr[51058] = 1722165606;
assign addr[51059] = 1710673591;
assign addr[51060] = 1699045930;
assign addr[51061] = 1687283545;
assign addr[51062] = 1675387369;
assign addr[51063] = 1663358344;
assign addr[51064] = 1651197426;
assign addr[51065] = 1638905577;
assign addr[51066] = 1626483774;
assign addr[51067] = 1613933000;
assign addr[51068] = 1601254251;
assign addr[51069] = 1588448533;
assign addr[51070] = 1575516860;
assign addr[51071] = 1562460258;
assign addr[51072] = 1549279763;
assign addr[51073] = 1535976419;
assign addr[51074] = 1522551282;
assign addr[51075] = 1509005416;
assign addr[51076] = 1495339895;
assign addr[51077] = 1481555802;
assign addr[51078] = 1467654232;
assign addr[51079] = 1453636285;
assign addr[51080] = 1439503074;
assign addr[51081] = 1425255719;
assign addr[51082] = 1410895350;
assign addr[51083] = 1396423105;
assign addr[51084] = 1381840133;
assign addr[51085] = 1367147589;
assign addr[51086] = 1352346639;
assign addr[51087] = 1337438456;
assign addr[51088] = 1322424222;
assign addr[51089] = 1307305128;
assign addr[51090] = 1292082373;
assign addr[51091] = 1276757164;
assign addr[51092] = 1261330715;
assign addr[51093] = 1245804251;
assign addr[51094] = 1230179002;
assign addr[51095] = 1214456207;
assign addr[51096] = 1198637114;
assign addr[51097] = 1182722976;
assign addr[51098] = 1166715055;
assign addr[51099] = 1150614620;
assign addr[51100] = 1134422949;
assign addr[51101] = 1118141326;
assign addr[51102] = 1101771040;
assign addr[51103] = 1085313391;
assign addr[51104] = 1068769683;
assign addr[51105] = 1052141228;
assign addr[51106] = 1035429345;
assign addr[51107] = 1018635358;
assign addr[51108] = 1001760600;
assign addr[51109] = 984806408;
assign addr[51110] = 967774128;
assign addr[51111] = 950665109;
assign addr[51112] = 933480707;
assign addr[51113] = 916222287;
assign addr[51114] = 898891215;
assign addr[51115] = 881488868;
assign addr[51116] = 864016623;
assign addr[51117] = 846475867;
assign addr[51118] = 828867991;
assign addr[51119] = 811194391;
assign addr[51120] = 793456467;
assign addr[51121] = 775655628;
assign addr[51122] = 757793284;
assign addr[51123] = 739870851;
assign addr[51124] = 721889752;
assign addr[51125] = 703851410;
assign addr[51126] = 685757258;
assign addr[51127] = 667608730;
assign addr[51128] = 649407264;
assign addr[51129] = 631154304;
assign addr[51130] = 612851297;
assign addr[51131] = 594499695;
assign addr[51132] = 576100953;
assign addr[51133] = 557656529;
assign addr[51134] = 539167887;
assign addr[51135] = 520636492;
assign addr[51136] = 502063814;
assign addr[51137] = 483451325;
assign addr[51138] = 464800501;
assign addr[51139] = 446112822;
assign addr[51140] = 427389768;
assign addr[51141] = 408632825;
assign addr[51142] = 389843480;
assign addr[51143] = 371023223;
assign addr[51144] = 352173546;
assign addr[51145] = 333295944;
assign addr[51146] = 314391913;
assign addr[51147] = 295462954;
assign addr[51148] = 276510565;
assign addr[51149] = 257536251;
assign addr[51150] = 238541516;
assign addr[51151] = 219527866;
assign addr[51152] = 200496809;
assign addr[51153] = 181449854;
assign addr[51154] = 162388511;
assign addr[51155] = 143314291;
assign addr[51156] = 124228708;
assign addr[51157] = 105133274;
assign addr[51158] = 86029503;
assign addr[51159] = 66918911;
assign addr[51160] = 47803013;
assign addr[51161] = 28683324;
assign addr[51162] = 9561361;
assign addr[51163] = -9561361;
assign addr[51164] = -28683324;
assign addr[51165] = -47803013;
assign addr[51166] = -66918911;
assign addr[51167] = -86029503;
assign addr[51168] = -105133274;
assign addr[51169] = -124228708;
assign addr[51170] = -143314291;
assign addr[51171] = -162388511;
assign addr[51172] = -181449854;
assign addr[51173] = -200496809;
assign addr[51174] = -219527866;
assign addr[51175] = -238541516;
assign addr[51176] = -257536251;
assign addr[51177] = -276510565;
assign addr[51178] = -295462953;
assign addr[51179] = -314391913;
assign addr[51180] = -333295944;
assign addr[51181] = -352173546;
assign addr[51182] = -371023223;
assign addr[51183] = -389843480;
assign addr[51184] = -408632825;
assign addr[51185] = -427389768;
assign addr[51186] = -446112822;
assign addr[51187] = -464800501;
assign addr[51188] = -483451325;
assign addr[51189] = -502063814;
assign addr[51190] = -520636492;
assign addr[51191] = -539167887;
assign addr[51192] = -557656529;
assign addr[51193] = -576100953;
assign addr[51194] = -594499695;
assign addr[51195] = -612851297;
assign addr[51196] = -631154304;
assign addr[51197] = -649407264;
assign addr[51198] = -667608730;
assign addr[51199] = -685757258;
assign addr[51200] = -703851410;
assign addr[51201] = -721889752;
assign addr[51202] = -739870851;
assign addr[51203] = -757793284;
assign addr[51204] = -775655628;
assign addr[51205] = -793456467;
assign addr[51206] = -811194391;
assign addr[51207] = -828867991;
assign addr[51208] = -846475867;
assign addr[51209] = -864016623;
assign addr[51210] = -881488868;
assign addr[51211] = -898891215;
assign addr[51212] = -916222287;
assign addr[51213] = -933480707;
assign addr[51214] = -950665109;
assign addr[51215] = -967774128;
assign addr[51216] = -984806408;
assign addr[51217] = -1001760600;
assign addr[51218] = -1018635358;
assign addr[51219] = -1035429345;
assign addr[51220] = -1052141228;
assign addr[51221] = -1068769683;
assign addr[51222] = -1085313391;
assign addr[51223] = -1101771040;
assign addr[51224] = -1118141326;
assign addr[51225] = -1134422949;
assign addr[51226] = -1150614620;
assign addr[51227] = -1166715055;
assign addr[51228] = -1182722976;
assign addr[51229] = -1198637114;
assign addr[51230] = -1214456207;
assign addr[51231] = -1230179002;
assign addr[51232] = -1245804251;
assign addr[51233] = -1261330715;
assign addr[51234] = -1276757164;
assign addr[51235] = -1292082373;
assign addr[51236] = -1307305128;
assign addr[51237] = -1322424222;
assign addr[51238] = -1337438456;
assign addr[51239] = -1352346639;
assign addr[51240] = -1367147589;
assign addr[51241] = -1381840133;
assign addr[51242] = -1396423105;
assign addr[51243] = -1410895350;
assign addr[51244] = -1425255719;
assign addr[51245] = -1439503074;
assign addr[51246] = -1453636285;
assign addr[51247] = -1467654232;
assign addr[51248] = -1481555802;
assign addr[51249] = -1495339895;
assign addr[51250] = -1509005416;
assign addr[51251] = -1522551282;
assign addr[51252] = -1535976419;
assign addr[51253] = -1549279763;
assign addr[51254] = -1562460258;
assign addr[51255] = -1575516860;
assign addr[51256] = -1588448533;
assign addr[51257] = -1601254251;
assign addr[51258] = -1613933000;
assign addr[51259] = -1626483774;
assign addr[51260] = -1638905577;
assign addr[51261] = -1651197426;
assign addr[51262] = -1663358344;
assign addr[51263] = -1675387369;
assign addr[51264] = -1687283545;
assign addr[51265] = -1699045930;
assign addr[51266] = -1710673591;
assign addr[51267] = -1722165606;
assign addr[51268] = -1733521064;
assign addr[51269] = -1744739065;
assign addr[51270] = -1755818718;
assign addr[51271] = -1766759146;
assign addr[51272] = -1777559480;
assign addr[51273] = -1788218865;
assign addr[51274] = -1798736454;
assign addr[51275] = -1809111415;
assign addr[51276] = -1819342925;
assign addr[51277] = -1829430172;
assign addr[51278] = -1839372356;
assign addr[51279] = -1849168689;
assign addr[51280] = -1858818395;
assign addr[51281] = -1868320707;
assign addr[51282] = -1877674873;
assign addr[51283] = -1886880151;
assign addr[51284] = -1895935811;
assign addr[51285] = -1904841135;
assign addr[51286] = -1913595416;
assign addr[51287] = -1922197961;
assign addr[51288] = -1930648088;
assign addr[51289] = -1938945125;
assign addr[51290] = -1947088417;
assign addr[51291] = -1955077316;
assign addr[51292] = -1962911189;
assign addr[51293] = -1970589416;
assign addr[51294] = -1978111387;
assign addr[51295] = -1985476506;
assign addr[51296] = -1992684188;
assign addr[51297] = -1999733863;
assign addr[51298] = -2006624971;
assign addr[51299] = -2013356967;
assign addr[51300] = -2019929315;
assign addr[51301] = -2026341495;
assign addr[51302] = -2032592999;
assign addr[51303] = -2038683330;
assign addr[51304] = -2044612007;
assign addr[51305] = -2050378558;
assign addr[51306] = -2055982526;
assign addr[51307] = -2061423468;
assign addr[51308] = -2066700952;
assign addr[51309] = -2071814558;
assign addr[51310] = -2076763883;
assign addr[51311] = -2081548533;
assign addr[51312] = -2086168128;
assign addr[51313] = -2090622304;
assign addr[51314] = -2094910706;
assign addr[51315] = -2099032994;
assign addr[51316] = -2102988841;
assign addr[51317] = -2106777935;
assign addr[51318] = -2110399974;
assign addr[51319] = -2113854671;
assign addr[51320] = -2117141752;
assign addr[51321] = -2120260957;
assign addr[51322] = -2123212038;
assign addr[51323] = -2125994762;
assign addr[51324] = -2128608907;
assign addr[51325] = -2131054266;
assign addr[51326] = -2133330646;
assign addr[51327] = -2135437865;
assign addr[51328] = -2137375758;
assign addr[51329] = -2139144169;
assign addr[51330] = -2140742960;
assign addr[51331] = -2142172003;
assign addr[51332] = -2143431184;
assign addr[51333] = -2144520405;
assign addr[51334] = -2145439578;
assign addr[51335] = -2146188631;
assign addr[51336] = -2146767505;
assign addr[51337] = -2147176152;
assign addr[51338] = -2147414542;
assign addr[51339] = -2147482655;
assign addr[51340] = -2147380486;
assign addr[51341] = -2147108043;
assign addr[51342] = -2146665347;
assign addr[51343] = -2146052433;
assign addr[51344] = -2145269351;
assign addr[51345] = -2144316162;
assign addr[51346] = -2143192942;
assign addr[51347] = -2141899780;
assign addr[51348] = -2140436778;
assign addr[51349] = -2138804053;
assign addr[51350] = -2137001733;
assign addr[51351] = -2135029962;
assign addr[51352] = -2132888897;
assign addr[51353] = -2130578706;
assign addr[51354] = -2128099574;
assign addr[51355] = -2125451696;
assign addr[51356] = -2122635283;
assign addr[51357] = -2119650558;
assign addr[51358] = -2116497758;
assign addr[51359] = -2113177132;
assign addr[51360] = -2109688944;
assign addr[51361] = -2106033471;
assign addr[51362] = -2102211002;
assign addr[51363] = -2098221841;
assign addr[51364] = -2094066304;
assign addr[51365] = -2089744719;
assign addr[51366] = -2085257431;
assign addr[51367] = -2080604795;
assign addr[51368] = -2075787180;
assign addr[51369] = -2070804967;
assign addr[51370] = -2065658552;
assign addr[51371] = -2060348343;
assign addr[51372] = -2054874761;
assign addr[51373] = -2049238240;
assign addr[51374] = -2043439226;
assign addr[51375] = -2037478181;
assign addr[51376] = -2031355576;
assign addr[51377] = -2025071897;
assign addr[51378] = -2018627642;
assign addr[51379] = -2012023322;
assign addr[51380] = -2005259462;
assign addr[51381] = -1998336596;
assign addr[51382] = -1991255274;
assign addr[51383] = -1984016058;
assign addr[51384] = -1976619522;
assign addr[51385] = -1969066252;
assign addr[51386] = -1961356847;
assign addr[51387] = -1953491918;
assign addr[51388] = -1945472089;
assign addr[51389] = -1937297997;
assign addr[51390] = -1928970288;
assign addr[51391] = -1920489624;
assign addr[51392] = -1911856677;
assign addr[51393] = -1903072131;
assign addr[51394] = -1894136683;
assign addr[51395] = -1885051042;
assign addr[51396] = -1875815927;
assign addr[51397] = -1866432072;
assign addr[51398] = -1856900221;
assign addr[51399] = -1847221128;
assign addr[51400] = -1837395562;
assign addr[51401] = -1827424302;
assign addr[51402] = -1817308138;
assign addr[51403] = -1807047873;
assign addr[51404] = -1796644320;
assign addr[51405] = -1786098304;
assign addr[51406] = -1775410662;
assign addr[51407] = -1764582240;
assign addr[51408] = -1753613897;
assign addr[51409] = -1742506504;
assign addr[51410] = -1731260941;
assign addr[51411] = -1719878099;
assign addr[51412] = -1708358881;
assign addr[51413] = -1696704201;
assign addr[51414] = -1684914983;
assign addr[51415] = -1672992161;
assign addr[51416] = -1660936681;
assign addr[51417] = -1648749499;
assign addr[51418] = -1636431582;
assign addr[51419] = -1623983905;
assign addr[51420] = -1611407456;
assign addr[51421] = -1598703233;
assign addr[51422] = -1585872242;
assign addr[51423] = -1572915501;
assign addr[51424] = -1559834037;
assign addr[51425] = -1546628888;
assign addr[51426] = -1533301101;
assign addr[51427] = -1519851733;
assign addr[51428] = -1506281850;
assign addr[51429] = -1492592527;
assign addr[51430] = -1478784851;
assign addr[51431] = -1464859917;
assign addr[51432] = -1450818828;
assign addr[51433] = -1436662698;
assign addr[51434] = -1422392650;
assign addr[51435] = -1408009814;
assign addr[51436] = -1393515332;
assign addr[51437] = -1378910353;
assign addr[51438] = -1364196034;
assign addr[51439] = -1349373543;
assign addr[51440] = -1334444055;
assign addr[51441] = -1319408754;
assign addr[51442] = -1304268832;
assign addr[51443] = -1289025489;
assign addr[51444] = -1273679934;
assign addr[51445] = -1258233384;
assign addr[51446] = -1242687064;
assign addr[51447] = -1227042207;
assign addr[51448] = -1211300053;
assign addr[51449] = -1195461849;
assign addr[51450] = -1179528853;
assign addr[51451] = -1163502328;
assign addr[51452] = -1147383544;
assign addr[51453] = -1131173780;
assign addr[51454] = -1114874320;
assign addr[51455] = -1098486458;
assign addr[51456] = -1082011492;
assign addr[51457] = -1065450729;
assign addr[51458] = -1048805483;
assign addr[51459] = -1032077073;
assign addr[51460] = -1015266825;
assign addr[51461] = -998376073;
assign addr[51462] = -981406156;
assign addr[51463] = -964358420;
assign addr[51464] = -947234215;
assign addr[51465] = -930034901;
assign addr[51466] = -912761841;
assign addr[51467] = -895416404;
assign addr[51468] = -877999966;
assign addr[51469] = -860513908;
assign addr[51470] = -842959617;
assign addr[51471] = -825338484;
assign addr[51472] = -807651907;
assign addr[51473] = -789901288;
assign addr[51474] = -772088034;
assign addr[51475] = -754213559;
assign addr[51476] = -736279279;
assign addr[51477] = -718286617;
assign addr[51478] = -700236999;
assign addr[51479] = -682131857;
assign addr[51480] = -663972625;
assign addr[51481] = -645760745;
assign addr[51482] = -627497660;
assign addr[51483] = -609184818;
assign addr[51484] = -590823671;
assign addr[51485] = -572415676;
assign addr[51486] = -553962291;
assign addr[51487] = -535464981;
assign addr[51488] = -516925212;
assign addr[51489] = -498344454;
assign addr[51490] = -479724180;
assign addr[51491] = -461065866;
assign addr[51492] = -442370993;
assign addr[51493] = -423641043;
assign addr[51494] = -404877501;
assign addr[51495] = -386081854;
assign addr[51496] = -367255594;
assign addr[51497] = -348400212;
assign addr[51498] = -329517204;
assign addr[51499] = -310608068;
assign addr[51500] = -291674302;
assign addr[51501] = -272717408;
assign addr[51502] = -253738890;
assign addr[51503] = -234740251;
assign addr[51504] = -215722999;
assign addr[51505] = -196688642;
assign addr[51506] = -177638688;
assign addr[51507] = -158574649;
assign addr[51508] = -139498035;
assign addr[51509] = -120410361;
assign addr[51510] = -101313138;
assign addr[51511] = -82207882;
assign addr[51512] = -63096108;
assign addr[51513] = -43979330;
assign addr[51514] = -24859065;
assign addr[51515] = -5736829;
assign addr[51516] = 13385863;
assign addr[51517] = 32507492;
assign addr[51518] = 51626544;
assign addr[51519] = 70741503;
assign addr[51520] = 89850852;
assign addr[51521] = 108953076;
assign addr[51522] = 128046661;
assign addr[51523] = 147130093;
assign addr[51524] = 166201858;
assign addr[51525] = 185260444;
assign addr[51526] = 204304341;
assign addr[51527] = 223332037;
assign addr[51528] = 242342025;
assign addr[51529] = 261332796;
assign addr[51530] = 280302845;
assign addr[51531] = 299250668;
assign addr[51532] = 318174762;
assign addr[51533] = 337073627;
assign addr[51534] = 355945764;
assign addr[51535] = 374789676;
assign addr[51536] = 393603870;
assign addr[51537] = 412386854;
assign addr[51538] = 431137138;
assign addr[51539] = 449853235;
assign addr[51540] = 468533662;
assign addr[51541] = 487176937;
assign addr[51542] = 505781581;
assign addr[51543] = 524346121;
assign addr[51544] = 542869083;
assign addr[51545] = 561348998;
assign addr[51546] = 579784402;
assign addr[51547] = 598173833;
assign addr[51548] = 616515832;
assign addr[51549] = 634808946;
assign addr[51550] = 653051723;
assign addr[51551] = 671242716;
assign addr[51552] = 689380485;
assign addr[51553] = 707463589;
assign addr[51554] = 725490597;
assign addr[51555] = 743460077;
assign addr[51556] = 761370605;
assign addr[51557] = 779220762;
assign addr[51558] = 797009130;
assign addr[51559] = 814734301;
assign addr[51560] = 832394869;
assign addr[51561] = 849989433;
assign addr[51562] = 867516597;
assign addr[51563] = 884974973;
assign addr[51564] = 902363176;
assign addr[51565] = 919679827;
assign addr[51566] = 936923553;
assign addr[51567] = 954092986;
assign addr[51568] = 971186766;
assign addr[51569] = 988203537;
assign addr[51570] = 1005141949;
assign addr[51571] = 1022000660;
assign addr[51572] = 1038778332;
assign addr[51573] = 1055473635;
assign addr[51574] = 1072085246;
assign addr[51575] = 1088611847;
assign addr[51576] = 1105052128;
assign addr[51577] = 1121404785;
assign addr[51578] = 1137668521;
assign addr[51579] = 1153842047;
assign addr[51580] = 1169924081;
assign addr[51581] = 1185913346;
assign addr[51582] = 1201808576;
assign addr[51583] = 1217608510;
assign addr[51584] = 1233311895;
assign addr[51585] = 1248917486;
assign addr[51586] = 1264424045;
assign addr[51587] = 1279830344;
assign addr[51588] = 1295135159;
assign addr[51589] = 1310337279;
assign addr[51590] = 1325435496;
assign addr[51591] = 1340428615;
assign addr[51592] = 1355315445;
assign addr[51593] = 1370094808;
assign addr[51594] = 1384765530;
assign addr[51595] = 1399326449;
assign addr[51596] = 1413776410;
assign addr[51597] = 1428114267;
assign addr[51598] = 1442338884;
assign addr[51599] = 1456449131;
assign addr[51600] = 1470443891;
assign addr[51601] = 1484322054;
assign addr[51602] = 1498082520;
assign addr[51603] = 1511724196;
assign addr[51604] = 1525246002;
assign addr[51605] = 1538646865;
assign addr[51606] = 1551925723;
assign addr[51607] = 1565081523;
assign addr[51608] = 1578113222;
assign addr[51609] = 1591019785;
assign addr[51610] = 1603800191;
assign addr[51611] = 1616453425;
assign addr[51612] = 1628978484;
assign addr[51613] = 1641374375;
assign addr[51614] = 1653640115;
assign addr[51615] = 1665774731;
assign addr[51616] = 1677777262;
assign addr[51617] = 1689646755;
assign addr[51618] = 1701382270;
assign addr[51619] = 1712982875;
assign addr[51620] = 1724447652;
assign addr[51621] = 1735775690;
assign addr[51622] = 1746966091;
assign addr[51623] = 1758017969;
assign addr[51624] = 1768930447;
assign addr[51625] = 1779702660;
assign addr[51626] = 1790333753;
assign addr[51627] = 1800822883;
assign addr[51628] = 1811169220;
assign addr[51629] = 1821371941;
assign addr[51630] = 1831430239;
assign addr[51631] = 1841343316;
assign addr[51632] = 1851110385;
assign addr[51633] = 1860730673;
assign addr[51634] = 1870203416;
assign addr[51635] = 1879527863;
assign addr[51636] = 1888703276;
assign addr[51637] = 1897728925;
assign addr[51638] = 1906604097;
assign addr[51639] = 1915328086;
assign addr[51640] = 1923900201;
assign addr[51641] = 1932319763;
assign addr[51642] = 1940586104;
assign addr[51643] = 1948698568;
assign addr[51644] = 1956656513;
assign addr[51645] = 1964459306;
assign addr[51646] = 1972106330;
assign addr[51647] = 1979596978;
assign addr[51648] = 1986930656;
assign addr[51649] = 1994106782;
assign addr[51650] = 2001124788;
assign addr[51651] = 2007984117;
assign addr[51652] = 2014684225;
assign addr[51653] = 2021224581;
assign addr[51654] = 2027604666;
assign addr[51655] = 2033823974;
assign addr[51656] = 2039882013;
assign addr[51657] = 2045778302;
assign addr[51658] = 2051512372;
assign addr[51659] = 2057083771;
assign addr[51660] = 2062492055;
assign addr[51661] = 2067736796;
assign addr[51662] = 2072817579;
assign addr[51663] = 2077733999;
assign addr[51664] = 2082485668;
assign addr[51665] = 2087072209;
assign addr[51666] = 2091493257;
assign addr[51667] = 2095748463;
assign addr[51668] = 2099837489;
assign addr[51669] = 2103760010;
assign addr[51670] = 2107515716;
assign addr[51671] = 2111104309;
assign addr[51672] = 2114525505;
assign addr[51673] = 2117779031;
assign addr[51674] = 2120864631;
assign addr[51675] = 2123782059;
assign addr[51676] = 2126531084;
assign addr[51677] = 2129111488;
assign addr[51678] = 2131523066;
assign addr[51679] = 2133765628;
assign addr[51680] = 2135838995;
assign addr[51681] = 2137743003;
assign addr[51682] = 2139477502;
assign addr[51683] = 2141042352;
assign addr[51684] = 2142437431;
assign addr[51685] = 2143662628;
assign addr[51686] = 2144717846;
assign addr[51687] = 2145603001;
assign addr[51688] = 2146318022;
assign addr[51689] = 2146862854;
assign addr[51690] = 2147237452;
assign addr[51691] = 2147441787;
assign addr[51692] = 2147475844;
assign addr[51693] = 2147339619;
assign addr[51694] = 2147033123;
assign addr[51695] = 2146556380;
assign addr[51696] = 2145909429;
assign addr[51697] = 2145092320;
assign addr[51698] = 2144105118;
assign addr[51699] = 2142947902;
assign addr[51700] = 2141620763;
assign addr[51701] = 2140123807;
assign addr[51702] = 2138457152;
assign addr[51703] = 2136620930;
assign addr[51704] = 2134615288;
assign addr[51705] = 2132440383;
assign addr[51706] = 2130096389;
assign addr[51707] = 2127583492;
assign addr[51708] = 2124901890;
assign addr[51709] = 2122051796;
assign addr[51710] = 2119033436;
assign addr[51711] = 2115847050;
assign addr[51712] = 2112492891;
assign addr[51713] = 2108971223;
assign addr[51714] = 2105282327;
assign addr[51715] = 2101426496;
assign addr[51716] = 2097404033;
assign addr[51717] = 2093215260;
assign addr[51718] = 2088860507;
assign addr[51719] = 2084340120;
assign addr[51720] = 2079654458;
assign addr[51721] = 2074803892;
assign addr[51722] = 2069788807;
assign addr[51723] = 2064609600;
assign addr[51724] = 2059266683;
assign addr[51725] = 2053760478;
assign addr[51726] = 2048091422;
assign addr[51727] = 2042259965;
assign addr[51728] = 2036266570;
assign addr[51729] = 2030111710;
assign addr[51730] = 2023795876;
assign addr[51731] = 2017319567;
assign addr[51732] = 2010683297;
assign addr[51733] = 2003887591;
assign addr[51734] = 1996932990;
assign addr[51735] = 1989820044;
assign addr[51736] = 1982549318;
assign addr[51737] = 1975121388;
assign addr[51738] = 1967536842;
assign addr[51739] = 1959796283;
assign addr[51740] = 1951900324;
assign addr[51741] = 1943849591;
assign addr[51742] = 1935644723;
assign addr[51743] = 1927286370;
assign addr[51744] = 1918775195;
assign addr[51745] = 1910111873;
assign addr[51746] = 1901297091;
assign addr[51747] = 1892331547;
assign addr[51748] = 1883215953;
assign addr[51749] = 1873951032;
assign addr[51750] = 1864537518;
assign addr[51751] = 1854976157;
assign addr[51752] = 1845267708;
assign addr[51753] = 1835412941;
assign addr[51754] = 1825412636;
assign addr[51755] = 1815267588;
assign addr[51756] = 1804978599;
assign addr[51757] = 1794546487;
assign addr[51758] = 1783972079;
assign addr[51759] = 1773256212;
assign addr[51760] = 1762399737;
assign addr[51761] = 1751403515;
assign addr[51762] = 1740268417;
assign addr[51763] = 1728995326;
assign addr[51764] = 1717585136;
assign addr[51765] = 1706038753;
assign addr[51766] = 1694357091;
assign addr[51767] = 1682541077;
assign addr[51768] = 1670591647;
assign addr[51769] = 1658509750;
assign addr[51770] = 1646296344;
assign addr[51771] = 1633952396;
assign addr[51772] = 1621478885;
assign addr[51773] = 1608876801;
assign addr[51774] = 1596147143;
assign addr[51775] = 1583290921;
assign addr[51776] = 1570309153;
assign addr[51777] = 1557202869;
assign addr[51778] = 1543973108;
assign addr[51779] = 1530620920;
assign addr[51780] = 1517147363;
assign addr[51781] = 1503553506;
assign addr[51782] = 1489840425;
assign addr[51783] = 1476009210;
assign addr[51784] = 1462060956;
assign addr[51785] = 1447996770;
assign addr[51786] = 1433817766;
assign addr[51787] = 1419525069;
assign addr[51788] = 1405119813;
assign addr[51789] = 1390603139;
assign addr[51790] = 1375976199;
assign addr[51791] = 1361240152;
assign addr[51792] = 1346396168;
assign addr[51793] = 1331445422;
assign addr[51794] = 1316389101;
assign addr[51795] = 1301228398;
assign addr[51796] = 1285964516;
assign addr[51797] = 1270598665;
assign addr[51798] = 1255132063;
assign addr[51799] = 1239565936;
assign addr[51800] = 1223901520;
assign addr[51801] = 1208140056;
assign addr[51802] = 1192282793;
assign addr[51803] = 1176330990;
assign addr[51804] = 1160285911;
assign addr[51805] = 1144148829;
assign addr[51806] = 1127921022;
assign addr[51807] = 1111603778;
assign addr[51808] = 1095198391;
assign addr[51809] = 1078706161;
assign addr[51810] = 1062128397;
assign addr[51811] = 1045466412;
assign addr[51812] = 1028721528;
assign addr[51813] = 1011895073;
assign addr[51814] = 994988380;
assign addr[51815] = 978002791;
assign addr[51816] = 960939653;
assign addr[51817] = 943800318;
assign addr[51818] = 926586145;
assign addr[51819] = 909298500;
assign addr[51820] = 891938752;
assign addr[51821] = 874508280;
assign addr[51822] = 857008464;
assign addr[51823] = 839440693;
assign addr[51824] = 821806359;
assign addr[51825] = 804106861;
assign addr[51826] = 786343603;
assign addr[51827] = 768517992;
assign addr[51828] = 750631442;
assign addr[51829] = 732685372;
assign addr[51830] = 714681204;
assign addr[51831] = 696620367;
assign addr[51832] = 678504291;
assign addr[51833] = 660334415;
assign addr[51834] = 642112178;
assign addr[51835] = 623839025;
assign addr[51836] = 605516406;
assign addr[51837] = 587145773;
assign addr[51838] = 568728583;
assign addr[51839] = 550266296;
assign addr[51840] = 531760377;
assign addr[51841] = 513212292;
assign addr[51842] = 494623513;
assign addr[51843] = 475995513;
assign addr[51844] = 457329769;
assign addr[51845] = 438627762;
assign addr[51846] = 419890975;
assign addr[51847] = 401120892;
assign addr[51848] = 382319004;
assign addr[51849] = 363486799;
assign addr[51850] = 344625773;
assign addr[51851] = 325737419;
assign addr[51852] = 306823237;
assign addr[51853] = 287884725;
assign addr[51854] = 268923386;
assign addr[51855] = 249940723;
assign addr[51856] = 230938242;
assign addr[51857] = 211917448;
assign addr[51858] = 192879850;
assign addr[51859] = 173826959;
assign addr[51860] = 154760284;
assign addr[51861] = 135681337;
assign addr[51862] = 116591632;
assign addr[51863] = 97492681;
assign addr[51864] = 78386000;
assign addr[51865] = 59273104;
assign addr[51866] = 40155507;
assign addr[51867] = 21034727;
assign addr[51868] = 1912278;
assign addr[51869] = -17210322;
assign addr[51870] = -36331557;
assign addr[51871] = -55449912;
assign addr[51872] = -74563870;
assign addr[51873] = -93671915;
assign addr[51874] = -112772533;
assign addr[51875] = -131864208;
assign addr[51876] = -150945428;
assign addr[51877] = -170014678;
assign addr[51878] = -189070447;
assign addr[51879] = -208111224;
assign addr[51880] = -227135500;
assign addr[51881] = -246141764;
assign addr[51882] = -265128512;
assign addr[51883] = -284094236;
assign addr[51884] = -303037433;
assign addr[51885] = -321956601;
assign addr[51886] = -340850240;
assign addr[51887] = -359716852;
assign addr[51888] = -378554940;
assign addr[51889] = -397363011;
assign addr[51890] = -416139574;
assign addr[51891] = -434883140;
assign addr[51892] = -453592221;
assign addr[51893] = -472265336;
assign addr[51894] = -490901003;
assign addr[51895] = -509497745;
assign addr[51896] = -528054086;
assign addr[51897] = -546568556;
assign addr[51898] = -565039687;
assign addr[51899] = -583466013;
assign addr[51900] = -601846074;
assign addr[51901] = -620178412;
assign addr[51902] = -638461574;
assign addr[51903] = -656694110;
assign addr[51904] = -674874574;
assign addr[51905] = -693001525;
assign addr[51906] = -711073524;
assign addr[51907] = -729089140;
assign addr[51908] = -747046944;
assign addr[51909] = -764945512;
assign addr[51910] = -782783424;
assign addr[51911] = -800559266;
assign addr[51912] = -818271628;
assign addr[51913] = -835919107;
assign addr[51914] = -853500302;
assign addr[51915] = -871013820;
assign addr[51916] = -888458272;
assign addr[51917] = -905832274;
assign addr[51918] = -923134450;
assign addr[51919] = -940363427;
assign addr[51920] = -957517838;
assign addr[51921] = -974596324;
assign addr[51922] = -991597531;
assign addr[51923] = -1008520110;
assign addr[51924] = -1025362720;
assign addr[51925] = -1042124025;
assign addr[51926] = -1058802695;
assign addr[51927] = -1075397409;
assign addr[51928] = -1091906851;
assign addr[51929] = -1108329711;
assign addr[51930] = -1124664687;
assign addr[51931] = -1140910484;
assign addr[51932] = -1157065814;
assign addr[51933] = -1173129396;
assign addr[51934] = -1189099956;
assign addr[51935] = -1204976227;
assign addr[51936] = -1220756951;
assign addr[51937] = -1236440877;
assign addr[51938] = -1252026760;
assign addr[51939] = -1267513365;
assign addr[51940] = -1282899464;
assign addr[51941] = -1298183838;
assign addr[51942] = -1313365273;
assign addr[51943] = -1328442566;
assign addr[51944] = -1343414522;
assign addr[51945] = -1358279953;
assign addr[51946] = -1373037681;
assign addr[51947] = -1387686535;
assign addr[51948] = -1402225355;
assign addr[51949] = -1416652986;
assign addr[51950] = -1430968286;
assign addr[51951] = -1445170118;
assign addr[51952] = -1459257358;
assign addr[51953] = -1473228887;
assign addr[51954] = -1487083598;
assign addr[51955] = -1500820393;
assign addr[51956] = -1514438181;
assign addr[51957] = -1527935884;
assign addr[51958] = -1541312431;
assign addr[51959] = -1554566762;
assign addr[51960] = -1567697824;
assign addr[51961] = -1580704578;
assign addr[51962] = -1593585992;
assign addr[51963] = -1606341043;
assign addr[51964] = -1618968722;
assign addr[51965] = -1631468027;
assign addr[51966] = -1643837966;
assign addr[51967] = -1656077559;
assign addr[51968] = -1668185835;
assign addr[51969] = -1680161834;
assign addr[51970] = -1692004606;
assign addr[51971] = -1703713213;
assign addr[51972] = -1715286726;
assign addr[51973] = -1726724227;
assign addr[51974] = -1738024810;
assign addr[51975] = -1749187577;
assign addr[51976] = -1760211645;
assign addr[51977] = -1771096139;
assign addr[51978] = -1781840195;
assign addr[51979] = -1792442963;
assign addr[51980] = -1802903601;
assign addr[51981] = -1813221279;
assign addr[51982] = -1823395180;
assign addr[51983] = -1833424497;
assign addr[51984] = -1843308435;
assign addr[51985] = -1853046210;
assign addr[51986] = -1862637049;
assign addr[51987] = -1872080193;
assign addr[51988] = -1881374892;
assign addr[51989] = -1890520410;
assign addr[51990] = -1899516021;
assign addr[51991] = -1908361011;
assign addr[51992] = -1917054681;
assign addr[51993] = -1925596340;
assign addr[51994] = -1933985310;
assign addr[51995] = -1942220928;
assign addr[51996] = -1950302539;
assign addr[51997] = -1958229503;
assign addr[51998] = -1966001192;
assign addr[51999] = -1973616989;
assign addr[52000] = -1981076290;
assign addr[52001] = -1988378503;
assign addr[52002] = -1995523051;
assign addr[52003] = -2002509365;
assign addr[52004] = -2009336893;
assign addr[52005] = -2016005093;
assign addr[52006] = -2022513436;
assign addr[52007] = -2028861406;
assign addr[52008] = -2035048499;
assign addr[52009] = -2041074226;
assign addr[52010] = -2046938108;
assign addr[52011] = -2052639680;
assign addr[52012] = -2058178491;
assign addr[52013] = -2063554100;
assign addr[52014] = -2068766083;
assign addr[52015] = -2073814024;
assign addr[52016] = -2078697525;
assign addr[52017] = -2083416198;
assign addr[52018] = -2087969669;
assign addr[52019] = -2092357577;
assign addr[52020] = -2096579573;
assign addr[52021] = -2100635323;
assign addr[52022] = -2104524506;
assign addr[52023] = -2108246813;
assign addr[52024] = -2111801949;
assign addr[52025] = -2115189632;
assign addr[52026] = -2118409593;
assign addr[52027] = -2121461578;
assign addr[52028] = -2124345343;
assign addr[52029] = -2127060661;
assign addr[52030] = -2129607316;
assign addr[52031] = -2131985106;
assign addr[52032] = -2134193842;
assign addr[52033] = -2136233350;
assign addr[52034] = -2138103468;
assign addr[52035] = -2139804048;
assign addr[52036] = -2141334954;
assign addr[52037] = -2142696065;
assign addr[52038] = -2143887273;
assign addr[52039] = -2144908484;
assign addr[52040] = -2145759618;
assign addr[52041] = -2146440605;
assign addr[52042] = -2146951393;
assign addr[52043] = -2147291941;
assign addr[52044] = -2147462221;
assign addr[52045] = -2147462221;
assign addr[52046] = -2147291941;
assign addr[52047] = -2146951393;
assign addr[52048] = -2146440605;
assign addr[52049] = -2145759618;
assign addr[52050] = -2144908484;
assign addr[52051] = -2143887273;
assign addr[52052] = -2142696065;
assign addr[52053] = -2141334954;
assign addr[52054] = -2139804048;
assign addr[52055] = -2138103468;
assign addr[52056] = -2136233350;
assign addr[52057] = -2134193842;
assign addr[52058] = -2131985106;
assign addr[52059] = -2129607316;
assign addr[52060] = -2127060661;
assign addr[52061] = -2124345343;
assign addr[52062] = -2121461578;
assign addr[52063] = -2118409593;
assign addr[52064] = -2115189632;
assign addr[52065] = -2111801949;
assign addr[52066] = -2108246813;
assign addr[52067] = -2104524506;
assign addr[52068] = -2100635323;
assign addr[52069] = -2096579573;
assign addr[52070] = -2092357577;
assign addr[52071] = -2087969669;
assign addr[52072] = -2083416198;
assign addr[52073] = -2078697525;
assign addr[52074] = -2073814024;
assign addr[52075] = -2068766083;
assign addr[52076] = -2063554100;
assign addr[52077] = -2058178491;
assign addr[52078] = -2052639680;
assign addr[52079] = -2046938108;
assign addr[52080] = -2041074226;
assign addr[52081] = -2035048499;
assign addr[52082] = -2028861406;
assign addr[52083] = -2022513436;
assign addr[52084] = -2016005093;
assign addr[52085] = -2009336893;
assign addr[52086] = -2002509365;
assign addr[52087] = -1995523051;
assign addr[52088] = -1988378503;
assign addr[52089] = -1981076290;
assign addr[52090] = -1973616989;
assign addr[52091] = -1966001192;
assign addr[52092] = -1958229503;
assign addr[52093] = -1950302539;
assign addr[52094] = -1942220928;
assign addr[52095] = -1933985310;
assign addr[52096] = -1925596340;
assign addr[52097] = -1917054681;
assign addr[52098] = -1908361011;
assign addr[52099] = -1899516021;
assign addr[52100] = -1890520410;
assign addr[52101] = -1881374892;
assign addr[52102] = -1872080193;
assign addr[52103] = -1862637049;
assign addr[52104] = -1853046210;
assign addr[52105] = -1843308435;
assign addr[52106] = -1833424497;
assign addr[52107] = -1823395180;
assign addr[52108] = -1813221279;
assign addr[52109] = -1802903601;
assign addr[52110] = -1792442963;
assign addr[52111] = -1781840195;
assign addr[52112] = -1771096139;
assign addr[52113] = -1760211645;
assign addr[52114] = -1749187577;
assign addr[52115] = -1738024810;
assign addr[52116] = -1726724227;
assign addr[52117] = -1715286726;
assign addr[52118] = -1703713213;
assign addr[52119] = -1692004606;
assign addr[52120] = -1680161834;
assign addr[52121] = -1668185835;
assign addr[52122] = -1656077559;
assign addr[52123] = -1643837966;
assign addr[52124] = -1631468027;
assign addr[52125] = -1618968722;
assign addr[52126] = -1606341043;
assign addr[52127] = -1593585992;
assign addr[52128] = -1580704578;
assign addr[52129] = -1567697824;
assign addr[52130] = -1554566762;
assign addr[52131] = -1541312431;
assign addr[52132] = -1527935884;
assign addr[52133] = -1514438181;
assign addr[52134] = -1500820393;
assign addr[52135] = -1487083598;
assign addr[52136] = -1473228887;
assign addr[52137] = -1459257358;
assign addr[52138] = -1445170118;
assign addr[52139] = -1430968286;
assign addr[52140] = -1416652986;
assign addr[52141] = -1402225355;
assign addr[52142] = -1387686535;
assign addr[52143] = -1373037681;
assign addr[52144] = -1358279953;
assign addr[52145] = -1343414522;
assign addr[52146] = -1328442566;
assign addr[52147] = -1313365273;
assign addr[52148] = -1298183838;
assign addr[52149] = -1282899464;
assign addr[52150] = -1267513365;
assign addr[52151] = -1252026760;
assign addr[52152] = -1236440877;
assign addr[52153] = -1220756951;
assign addr[52154] = -1204976227;
assign addr[52155] = -1189099956;
assign addr[52156] = -1173129396;
assign addr[52157] = -1157065814;
assign addr[52158] = -1140910484;
assign addr[52159] = -1124664687;
assign addr[52160] = -1108329711;
assign addr[52161] = -1091906851;
assign addr[52162] = -1075397409;
assign addr[52163] = -1058802695;
assign addr[52164] = -1042124025;
assign addr[52165] = -1025362720;
assign addr[52166] = -1008520110;
assign addr[52167] = -991597531;
assign addr[52168] = -974596324;
assign addr[52169] = -957517838;
assign addr[52170] = -940363427;
assign addr[52171] = -923134450;
assign addr[52172] = -905832274;
assign addr[52173] = -888458272;
assign addr[52174] = -871013820;
assign addr[52175] = -853500302;
assign addr[52176] = -835919107;
assign addr[52177] = -818271628;
assign addr[52178] = -800559266;
assign addr[52179] = -782783424;
assign addr[52180] = -764945512;
assign addr[52181] = -747046944;
assign addr[52182] = -729089140;
assign addr[52183] = -711073524;
assign addr[52184] = -693001525;
assign addr[52185] = -674874574;
assign addr[52186] = -656694110;
assign addr[52187] = -638461574;
assign addr[52188] = -620178412;
assign addr[52189] = -601846074;
assign addr[52190] = -583466013;
assign addr[52191] = -565039687;
assign addr[52192] = -546568556;
assign addr[52193] = -528054086;
assign addr[52194] = -509497745;
assign addr[52195] = -490901003;
assign addr[52196] = -472265336;
assign addr[52197] = -453592221;
assign addr[52198] = -434883140;
assign addr[52199] = -416139574;
assign addr[52200] = -397363011;
assign addr[52201] = -378554940;
assign addr[52202] = -359716852;
assign addr[52203] = -340850240;
assign addr[52204] = -321956601;
assign addr[52205] = -303037433;
assign addr[52206] = -284094236;
assign addr[52207] = -265128512;
assign addr[52208] = -246141764;
assign addr[52209] = -227135500;
assign addr[52210] = -208111224;
assign addr[52211] = -189070447;
assign addr[52212] = -170014678;
assign addr[52213] = -150945428;
assign addr[52214] = -131864208;
assign addr[52215] = -112772533;
assign addr[52216] = -93671915;
assign addr[52217] = -74563870;
assign addr[52218] = -55449912;
assign addr[52219] = -36331557;
assign addr[52220] = -17210322;
assign addr[52221] = 1912278;
assign addr[52222] = 21034727;
assign addr[52223] = 40155507;
assign addr[52224] = 59273104;
assign addr[52225] = 78386000;
assign addr[52226] = 97492681;
assign addr[52227] = 116591632;
assign addr[52228] = 135681337;
assign addr[52229] = 154760284;
assign addr[52230] = 173826959;
assign addr[52231] = 192879850;
assign addr[52232] = 211917448;
assign addr[52233] = 230938242;
assign addr[52234] = 249940723;
assign addr[52235] = 268923386;
assign addr[52236] = 287884725;
assign addr[52237] = 306823237;
assign addr[52238] = 325737419;
assign addr[52239] = 344625773;
assign addr[52240] = 363486799;
assign addr[52241] = 382319004;
assign addr[52242] = 401120892;
assign addr[52243] = 419890975;
assign addr[52244] = 438627762;
assign addr[52245] = 457329769;
assign addr[52246] = 475995513;
assign addr[52247] = 494623513;
assign addr[52248] = 513212292;
assign addr[52249] = 531760377;
assign addr[52250] = 550266296;
assign addr[52251] = 568728583;
assign addr[52252] = 587145773;
assign addr[52253] = 605516406;
assign addr[52254] = 623839025;
assign addr[52255] = 642112178;
assign addr[52256] = 660334415;
assign addr[52257] = 678504291;
assign addr[52258] = 696620367;
assign addr[52259] = 714681204;
assign addr[52260] = 732685372;
assign addr[52261] = 750631442;
assign addr[52262] = 768517992;
assign addr[52263] = 786343603;
assign addr[52264] = 804106861;
assign addr[52265] = 821806359;
assign addr[52266] = 839440693;
assign addr[52267] = 857008464;
assign addr[52268] = 874508280;
assign addr[52269] = 891938752;
assign addr[52270] = 909298500;
assign addr[52271] = 926586145;
assign addr[52272] = 943800318;
assign addr[52273] = 960939653;
assign addr[52274] = 978002791;
assign addr[52275] = 994988380;
assign addr[52276] = 1011895073;
assign addr[52277] = 1028721528;
assign addr[52278] = 1045466412;
assign addr[52279] = 1062128397;
assign addr[52280] = 1078706161;
assign addr[52281] = 1095198391;
assign addr[52282] = 1111603778;
assign addr[52283] = 1127921022;
assign addr[52284] = 1144148829;
assign addr[52285] = 1160285911;
assign addr[52286] = 1176330990;
assign addr[52287] = 1192282793;
assign addr[52288] = 1208140056;
assign addr[52289] = 1223901520;
assign addr[52290] = 1239565936;
assign addr[52291] = 1255132063;
assign addr[52292] = 1270598665;
assign addr[52293] = 1285964516;
assign addr[52294] = 1301228398;
assign addr[52295] = 1316389101;
assign addr[52296] = 1331445422;
assign addr[52297] = 1346396168;
assign addr[52298] = 1361240152;
assign addr[52299] = 1375976199;
assign addr[52300] = 1390603139;
assign addr[52301] = 1405119813;
assign addr[52302] = 1419525069;
assign addr[52303] = 1433817766;
assign addr[52304] = 1447996770;
assign addr[52305] = 1462060956;
assign addr[52306] = 1476009210;
assign addr[52307] = 1489840425;
assign addr[52308] = 1503553506;
assign addr[52309] = 1517147363;
assign addr[52310] = 1530620920;
assign addr[52311] = 1543973108;
assign addr[52312] = 1557202869;
assign addr[52313] = 1570309153;
assign addr[52314] = 1583290921;
assign addr[52315] = 1596147143;
assign addr[52316] = 1608876801;
assign addr[52317] = 1621478885;
assign addr[52318] = 1633952396;
assign addr[52319] = 1646296344;
assign addr[52320] = 1658509750;
assign addr[52321] = 1670591647;
assign addr[52322] = 1682541077;
assign addr[52323] = 1694357091;
assign addr[52324] = 1706038753;
assign addr[52325] = 1717585136;
assign addr[52326] = 1728995326;
assign addr[52327] = 1740268417;
assign addr[52328] = 1751403515;
assign addr[52329] = 1762399737;
assign addr[52330] = 1773256212;
assign addr[52331] = 1783972079;
assign addr[52332] = 1794546487;
assign addr[52333] = 1804978599;
assign addr[52334] = 1815267588;
assign addr[52335] = 1825412636;
assign addr[52336] = 1835412941;
assign addr[52337] = 1845267708;
assign addr[52338] = 1854976157;
assign addr[52339] = 1864537518;
assign addr[52340] = 1873951032;
assign addr[52341] = 1883215953;
assign addr[52342] = 1892331547;
assign addr[52343] = 1901297091;
assign addr[52344] = 1910111873;
assign addr[52345] = 1918775195;
assign addr[52346] = 1927286370;
assign addr[52347] = 1935644723;
assign addr[52348] = 1943849591;
assign addr[52349] = 1951900324;
assign addr[52350] = 1959796283;
assign addr[52351] = 1967536842;
assign addr[52352] = 1975121388;
assign addr[52353] = 1982549318;
assign addr[52354] = 1989820044;
assign addr[52355] = 1996932990;
assign addr[52356] = 2003887591;
assign addr[52357] = 2010683297;
assign addr[52358] = 2017319567;
assign addr[52359] = 2023795876;
assign addr[52360] = 2030111710;
assign addr[52361] = 2036266570;
assign addr[52362] = 2042259965;
assign addr[52363] = 2048091422;
assign addr[52364] = 2053760478;
assign addr[52365] = 2059266683;
assign addr[52366] = 2064609600;
assign addr[52367] = 2069788807;
assign addr[52368] = 2074803892;
assign addr[52369] = 2079654458;
assign addr[52370] = 2084340120;
assign addr[52371] = 2088860507;
assign addr[52372] = 2093215260;
assign addr[52373] = 2097404033;
assign addr[52374] = 2101426496;
assign addr[52375] = 2105282327;
assign addr[52376] = 2108971223;
assign addr[52377] = 2112492891;
assign addr[52378] = 2115847050;
assign addr[52379] = 2119033436;
assign addr[52380] = 2122051796;
assign addr[52381] = 2124901890;
assign addr[52382] = 2127583492;
assign addr[52383] = 2130096389;
assign addr[52384] = 2132440383;
assign addr[52385] = 2134615288;
assign addr[52386] = 2136620930;
assign addr[52387] = 2138457152;
assign addr[52388] = 2140123807;
assign addr[52389] = 2141620763;
assign addr[52390] = 2142947902;
assign addr[52391] = 2144105118;
assign addr[52392] = 2145092320;
assign addr[52393] = 2145909429;
assign addr[52394] = 2146556380;
assign addr[52395] = 2147033123;
assign addr[52396] = 2147339619;
assign addr[52397] = 2147475844;
assign addr[52398] = 2147441787;
assign addr[52399] = 2147237452;
assign addr[52400] = 2146862854;
assign addr[52401] = 2146318022;
assign addr[52402] = 2145603001;
assign addr[52403] = 2144717846;
assign addr[52404] = 2143662628;
assign addr[52405] = 2142437431;
assign addr[52406] = 2141042352;
assign addr[52407] = 2139477502;
assign addr[52408] = 2137743003;
assign addr[52409] = 2135838995;
assign addr[52410] = 2133765628;
assign addr[52411] = 2131523066;
assign addr[52412] = 2129111488;
assign addr[52413] = 2126531084;
assign addr[52414] = 2123782059;
assign addr[52415] = 2120864631;
assign addr[52416] = 2117779031;
assign addr[52417] = 2114525505;
assign addr[52418] = 2111104309;
assign addr[52419] = 2107515716;
assign addr[52420] = 2103760010;
assign addr[52421] = 2099837489;
assign addr[52422] = 2095748463;
assign addr[52423] = 2091493257;
assign addr[52424] = 2087072209;
assign addr[52425] = 2082485668;
assign addr[52426] = 2077733999;
assign addr[52427] = 2072817579;
assign addr[52428] = 2067736796;
assign addr[52429] = 2062492055;
assign addr[52430] = 2057083771;
assign addr[52431] = 2051512372;
assign addr[52432] = 2045778302;
assign addr[52433] = 2039882013;
assign addr[52434] = 2033823974;
assign addr[52435] = 2027604666;
assign addr[52436] = 2021224581;
assign addr[52437] = 2014684225;
assign addr[52438] = 2007984117;
assign addr[52439] = 2001124788;
assign addr[52440] = 1994106782;
assign addr[52441] = 1986930656;
assign addr[52442] = 1979596978;
assign addr[52443] = 1972106330;
assign addr[52444] = 1964459306;
assign addr[52445] = 1956656513;
assign addr[52446] = 1948698568;
assign addr[52447] = 1940586104;
assign addr[52448] = 1932319763;
assign addr[52449] = 1923900201;
assign addr[52450] = 1915328086;
assign addr[52451] = 1906604097;
assign addr[52452] = 1897728925;
assign addr[52453] = 1888703276;
assign addr[52454] = 1879527863;
assign addr[52455] = 1870203416;
assign addr[52456] = 1860730673;
assign addr[52457] = 1851110385;
assign addr[52458] = 1841343316;
assign addr[52459] = 1831430239;
assign addr[52460] = 1821371941;
assign addr[52461] = 1811169220;
assign addr[52462] = 1800822883;
assign addr[52463] = 1790333753;
assign addr[52464] = 1779702660;
assign addr[52465] = 1768930447;
assign addr[52466] = 1758017969;
assign addr[52467] = 1746966091;
assign addr[52468] = 1735775690;
assign addr[52469] = 1724447652;
assign addr[52470] = 1712982875;
assign addr[52471] = 1701382270;
assign addr[52472] = 1689646755;
assign addr[52473] = 1677777262;
assign addr[52474] = 1665774731;
assign addr[52475] = 1653640115;
assign addr[52476] = 1641374375;
assign addr[52477] = 1628978484;
assign addr[52478] = 1616453425;
assign addr[52479] = 1603800191;
assign addr[52480] = 1591019785;
assign addr[52481] = 1578113222;
assign addr[52482] = 1565081523;
assign addr[52483] = 1551925723;
assign addr[52484] = 1538646865;
assign addr[52485] = 1525246002;
assign addr[52486] = 1511724196;
assign addr[52487] = 1498082520;
assign addr[52488] = 1484322054;
assign addr[52489] = 1470443891;
assign addr[52490] = 1456449131;
assign addr[52491] = 1442338884;
assign addr[52492] = 1428114267;
assign addr[52493] = 1413776410;
assign addr[52494] = 1399326449;
assign addr[52495] = 1384765530;
assign addr[52496] = 1370094808;
assign addr[52497] = 1355315445;
assign addr[52498] = 1340428615;
assign addr[52499] = 1325435496;
assign addr[52500] = 1310337279;
assign addr[52501] = 1295135159;
assign addr[52502] = 1279830344;
assign addr[52503] = 1264424045;
assign addr[52504] = 1248917486;
assign addr[52505] = 1233311895;
assign addr[52506] = 1217608510;
assign addr[52507] = 1201808576;
assign addr[52508] = 1185913346;
assign addr[52509] = 1169924081;
assign addr[52510] = 1153842047;
assign addr[52511] = 1137668521;
assign addr[52512] = 1121404785;
assign addr[52513] = 1105052128;
assign addr[52514] = 1088611847;
assign addr[52515] = 1072085246;
assign addr[52516] = 1055473635;
assign addr[52517] = 1038778332;
assign addr[52518] = 1022000660;
assign addr[52519] = 1005141949;
assign addr[52520] = 988203537;
assign addr[52521] = 971186766;
assign addr[52522] = 954092986;
assign addr[52523] = 936923553;
assign addr[52524] = 919679827;
assign addr[52525] = 902363176;
assign addr[52526] = 884974973;
assign addr[52527] = 867516597;
assign addr[52528] = 849989433;
assign addr[52529] = 832394869;
assign addr[52530] = 814734301;
assign addr[52531] = 797009130;
assign addr[52532] = 779220762;
assign addr[52533] = 761370605;
assign addr[52534] = 743460077;
assign addr[52535] = 725490597;
assign addr[52536] = 707463589;
assign addr[52537] = 689380485;
assign addr[52538] = 671242716;
assign addr[52539] = 653051723;
assign addr[52540] = 634808946;
assign addr[52541] = 616515832;
assign addr[52542] = 598173833;
assign addr[52543] = 579784402;
assign addr[52544] = 561348998;
assign addr[52545] = 542869083;
assign addr[52546] = 524346121;
assign addr[52547] = 505781581;
assign addr[52548] = 487176937;
assign addr[52549] = 468533662;
assign addr[52550] = 449853235;
assign addr[52551] = 431137138;
assign addr[52552] = 412386854;
assign addr[52553] = 393603870;
assign addr[52554] = 374789676;
assign addr[52555] = 355945764;
assign addr[52556] = 337073627;
assign addr[52557] = 318174762;
assign addr[52558] = 299250668;
assign addr[52559] = 280302845;
assign addr[52560] = 261332796;
assign addr[52561] = 242342025;
assign addr[52562] = 223332037;
assign addr[52563] = 204304341;
assign addr[52564] = 185260444;
assign addr[52565] = 166201858;
assign addr[52566] = 147130093;
assign addr[52567] = 128046661;
assign addr[52568] = 108953076;
assign addr[52569] = 89850852;
assign addr[52570] = 70741503;
assign addr[52571] = 51626544;
assign addr[52572] = 32507492;
assign addr[52573] = 13385863;
assign addr[52574] = -5736829;
assign addr[52575] = -24859065;
assign addr[52576] = -43979330;
assign addr[52577] = -63096108;
assign addr[52578] = -82207882;
assign addr[52579] = -101313138;
assign addr[52580] = -120410361;
assign addr[52581] = -139498035;
assign addr[52582] = -158574649;
assign addr[52583] = -177638688;
assign addr[52584] = -196688642;
assign addr[52585] = -215722999;
assign addr[52586] = -234740251;
assign addr[52587] = -253738890;
assign addr[52588] = -272717408;
assign addr[52589] = -291674302;
assign addr[52590] = -310608068;
assign addr[52591] = -329517204;
assign addr[52592] = -348400212;
assign addr[52593] = -367255594;
assign addr[52594] = -386081854;
assign addr[52595] = -404877501;
assign addr[52596] = -423641043;
assign addr[52597] = -442370993;
assign addr[52598] = -461065866;
assign addr[52599] = -479724180;
assign addr[52600] = -498344454;
assign addr[52601] = -516925212;
assign addr[52602] = -535464981;
assign addr[52603] = -553962291;
assign addr[52604] = -572415676;
assign addr[52605] = -590823671;
assign addr[52606] = -609184818;
assign addr[52607] = -627497660;
assign addr[52608] = -645760745;
assign addr[52609] = -663972625;
assign addr[52610] = -682131857;
assign addr[52611] = -700236999;
assign addr[52612] = -718286617;
assign addr[52613] = -736279279;
assign addr[52614] = -754213559;
assign addr[52615] = -772088034;
assign addr[52616] = -789901288;
assign addr[52617] = -807651907;
assign addr[52618] = -825338484;
assign addr[52619] = -842959617;
assign addr[52620] = -860513908;
assign addr[52621] = -877999966;
assign addr[52622] = -895416404;
assign addr[52623] = -912761841;
assign addr[52624] = -930034901;
assign addr[52625] = -947234215;
assign addr[52626] = -964358420;
assign addr[52627] = -981406156;
assign addr[52628] = -998376073;
assign addr[52629] = -1015266825;
assign addr[52630] = -1032077073;
assign addr[52631] = -1048805483;
assign addr[52632] = -1065450729;
assign addr[52633] = -1082011492;
assign addr[52634] = -1098486458;
assign addr[52635] = -1114874320;
assign addr[52636] = -1131173780;
assign addr[52637] = -1147383544;
assign addr[52638] = -1163502328;
assign addr[52639] = -1179528853;
assign addr[52640] = -1195461849;
assign addr[52641] = -1211300053;
assign addr[52642] = -1227042207;
assign addr[52643] = -1242687064;
assign addr[52644] = -1258233384;
assign addr[52645] = -1273679934;
assign addr[52646] = -1289025489;
assign addr[52647] = -1304268832;
assign addr[52648] = -1319408754;
assign addr[52649] = -1334444055;
assign addr[52650] = -1349373543;
assign addr[52651] = -1364196034;
assign addr[52652] = -1378910353;
assign addr[52653] = -1393515332;
assign addr[52654] = -1408009814;
assign addr[52655] = -1422392650;
assign addr[52656] = -1436662698;
assign addr[52657] = -1450818828;
assign addr[52658] = -1464859917;
assign addr[52659] = -1478784851;
assign addr[52660] = -1492592527;
assign addr[52661] = -1506281850;
assign addr[52662] = -1519851733;
assign addr[52663] = -1533301101;
assign addr[52664] = -1546628888;
assign addr[52665] = -1559834037;
assign addr[52666] = -1572915501;
assign addr[52667] = -1585872242;
assign addr[52668] = -1598703233;
assign addr[52669] = -1611407456;
assign addr[52670] = -1623983905;
assign addr[52671] = -1636431582;
assign addr[52672] = -1648749499;
assign addr[52673] = -1660936681;
assign addr[52674] = -1672992161;
assign addr[52675] = -1684914983;
assign addr[52676] = -1696704201;
assign addr[52677] = -1708358881;
assign addr[52678] = -1719878099;
assign addr[52679] = -1731260941;
assign addr[52680] = -1742506504;
assign addr[52681] = -1753613897;
assign addr[52682] = -1764582240;
assign addr[52683] = -1775410662;
assign addr[52684] = -1786098304;
assign addr[52685] = -1796644320;
assign addr[52686] = -1807047873;
assign addr[52687] = -1817308138;
assign addr[52688] = -1827424302;
assign addr[52689] = -1837395562;
assign addr[52690] = -1847221128;
assign addr[52691] = -1856900221;
assign addr[52692] = -1866432072;
assign addr[52693] = -1875815927;
assign addr[52694] = -1885051042;
assign addr[52695] = -1894136683;
assign addr[52696] = -1903072131;
assign addr[52697] = -1911856677;
assign addr[52698] = -1920489624;
assign addr[52699] = -1928970288;
assign addr[52700] = -1937297997;
assign addr[52701] = -1945472089;
assign addr[52702] = -1953491918;
assign addr[52703] = -1961356847;
assign addr[52704] = -1969066252;
assign addr[52705] = -1976619522;
assign addr[52706] = -1984016058;
assign addr[52707] = -1991255274;
assign addr[52708] = -1998336596;
assign addr[52709] = -2005259462;
assign addr[52710] = -2012023322;
assign addr[52711] = -2018627642;
assign addr[52712] = -2025071897;
assign addr[52713] = -2031355576;
assign addr[52714] = -2037478181;
assign addr[52715] = -2043439226;
assign addr[52716] = -2049238240;
assign addr[52717] = -2054874761;
assign addr[52718] = -2060348343;
assign addr[52719] = -2065658552;
assign addr[52720] = -2070804967;
assign addr[52721] = -2075787180;
assign addr[52722] = -2080604795;
assign addr[52723] = -2085257431;
assign addr[52724] = -2089744719;
assign addr[52725] = -2094066304;
assign addr[52726] = -2098221841;
assign addr[52727] = -2102211002;
assign addr[52728] = -2106033471;
assign addr[52729] = -2109688944;
assign addr[52730] = -2113177132;
assign addr[52731] = -2116497758;
assign addr[52732] = -2119650558;
assign addr[52733] = -2122635283;
assign addr[52734] = -2125451696;
assign addr[52735] = -2128099574;
assign addr[52736] = -2130578706;
assign addr[52737] = -2132888897;
assign addr[52738] = -2135029962;
assign addr[52739] = -2137001733;
assign addr[52740] = -2138804053;
assign addr[52741] = -2140436778;
assign addr[52742] = -2141899780;
assign addr[52743] = -2143192942;
assign addr[52744] = -2144316162;
assign addr[52745] = -2145269351;
assign addr[52746] = -2146052433;
assign addr[52747] = -2146665347;
assign addr[52748] = -2147108043;
assign addr[52749] = -2147380486;
assign addr[52750] = -2147482655;
assign addr[52751] = -2147414542;
assign addr[52752] = -2147176152;
assign addr[52753] = -2146767505;
assign addr[52754] = -2146188631;
assign addr[52755] = -2145439578;
assign addr[52756] = -2144520405;
assign addr[52757] = -2143431184;
assign addr[52758] = -2142172003;
assign addr[52759] = -2140742960;
assign addr[52760] = -2139144169;
assign addr[52761] = -2137375758;
assign addr[52762] = -2135437865;
assign addr[52763] = -2133330646;
assign addr[52764] = -2131054266;
assign addr[52765] = -2128608907;
assign addr[52766] = -2125994762;
assign addr[52767] = -2123212038;
assign addr[52768] = -2120260957;
assign addr[52769] = -2117141752;
assign addr[52770] = -2113854671;
assign addr[52771] = -2110399974;
assign addr[52772] = -2106777935;
assign addr[52773] = -2102988841;
assign addr[52774] = -2099032994;
assign addr[52775] = -2094910706;
assign addr[52776] = -2090622304;
assign addr[52777] = -2086168128;
assign addr[52778] = -2081548533;
assign addr[52779] = -2076763883;
assign addr[52780] = -2071814558;
assign addr[52781] = -2066700952;
assign addr[52782] = -2061423468;
assign addr[52783] = -2055982526;
assign addr[52784] = -2050378558;
assign addr[52785] = -2044612007;
assign addr[52786] = -2038683330;
assign addr[52787] = -2032592999;
assign addr[52788] = -2026341495;
assign addr[52789] = -2019929315;
assign addr[52790] = -2013356967;
assign addr[52791] = -2006624971;
assign addr[52792] = -1999733863;
assign addr[52793] = -1992684188;
assign addr[52794] = -1985476506;
assign addr[52795] = -1978111387;
assign addr[52796] = -1970589416;
assign addr[52797] = -1962911189;
assign addr[52798] = -1955077316;
assign addr[52799] = -1947088417;
assign addr[52800] = -1938945125;
assign addr[52801] = -1930648088;
assign addr[52802] = -1922197961;
assign addr[52803] = -1913595416;
assign addr[52804] = -1904841135;
assign addr[52805] = -1895935811;
assign addr[52806] = -1886880151;
assign addr[52807] = -1877674873;
assign addr[52808] = -1868320707;
assign addr[52809] = -1858818395;
assign addr[52810] = -1849168689;
assign addr[52811] = -1839372356;
assign addr[52812] = -1829430172;
assign addr[52813] = -1819342925;
assign addr[52814] = -1809111415;
assign addr[52815] = -1798736454;
assign addr[52816] = -1788218865;
assign addr[52817] = -1777559480;
assign addr[52818] = -1766759146;
assign addr[52819] = -1755818718;
assign addr[52820] = -1744739065;
assign addr[52821] = -1733521064;
assign addr[52822] = -1722165606;
assign addr[52823] = -1710673591;
assign addr[52824] = -1699045930;
assign addr[52825] = -1687283545;
assign addr[52826] = -1675387369;
assign addr[52827] = -1663358344;
assign addr[52828] = -1651197426;
assign addr[52829] = -1638905577;
assign addr[52830] = -1626483774;
assign addr[52831] = -1613933000;
assign addr[52832] = -1601254251;
assign addr[52833] = -1588448533;
assign addr[52834] = -1575516860;
assign addr[52835] = -1562460258;
assign addr[52836] = -1549279763;
assign addr[52837] = -1535976419;
assign addr[52838] = -1522551282;
assign addr[52839] = -1509005416;
assign addr[52840] = -1495339895;
assign addr[52841] = -1481555802;
assign addr[52842] = -1467654232;
assign addr[52843] = -1453636285;
assign addr[52844] = -1439503074;
assign addr[52845] = -1425255719;
assign addr[52846] = -1410895350;
assign addr[52847] = -1396423105;
assign addr[52848] = -1381840133;
assign addr[52849] = -1367147589;
assign addr[52850] = -1352346639;
assign addr[52851] = -1337438456;
assign addr[52852] = -1322424222;
assign addr[52853] = -1307305128;
assign addr[52854] = -1292082373;
assign addr[52855] = -1276757164;
assign addr[52856] = -1261330715;
assign addr[52857] = -1245804251;
assign addr[52858] = -1230179002;
assign addr[52859] = -1214456207;
assign addr[52860] = -1198637114;
assign addr[52861] = -1182722976;
assign addr[52862] = -1166715055;
assign addr[52863] = -1150614620;
assign addr[52864] = -1134422949;
assign addr[52865] = -1118141326;
assign addr[52866] = -1101771040;
assign addr[52867] = -1085313391;
assign addr[52868] = -1068769683;
assign addr[52869] = -1052141228;
assign addr[52870] = -1035429345;
assign addr[52871] = -1018635358;
assign addr[52872] = -1001760600;
assign addr[52873] = -984806408;
assign addr[52874] = -967774128;
assign addr[52875] = -950665109;
assign addr[52876] = -933480707;
assign addr[52877] = -916222287;
assign addr[52878] = -898891215;
assign addr[52879] = -881488868;
assign addr[52880] = -864016623;
assign addr[52881] = -846475867;
assign addr[52882] = -828867991;
assign addr[52883] = -811194391;
assign addr[52884] = -793456467;
assign addr[52885] = -775655628;
assign addr[52886] = -757793284;
assign addr[52887] = -739870851;
assign addr[52888] = -721889752;
assign addr[52889] = -703851410;
assign addr[52890] = -685757258;
assign addr[52891] = -667608730;
assign addr[52892] = -649407264;
assign addr[52893] = -631154304;
assign addr[52894] = -612851297;
assign addr[52895] = -594499695;
assign addr[52896] = -576100953;
assign addr[52897] = -557656529;
assign addr[52898] = -539167887;
assign addr[52899] = -520636492;
assign addr[52900] = -502063814;
assign addr[52901] = -483451325;
assign addr[52902] = -464800501;
assign addr[52903] = -446112822;
assign addr[52904] = -427389768;
assign addr[52905] = -408632825;
assign addr[52906] = -389843480;
assign addr[52907] = -371023223;
assign addr[52908] = -352173546;
assign addr[52909] = -333295944;
assign addr[52910] = -314391913;
assign addr[52911] = -295462954;
assign addr[52912] = -276510565;
assign addr[52913] = -257536251;
assign addr[52914] = -238541516;
assign addr[52915] = -219527866;
assign addr[52916] = -200496809;
assign addr[52917] = -181449854;
assign addr[52918] = -162388511;
assign addr[52919] = -143314291;
assign addr[52920] = -124228708;
assign addr[52921] = -105133274;
assign addr[52922] = -86029503;
assign addr[52923] = -66918911;
assign addr[52924] = -47803013;
assign addr[52925] = -28683324;
assign addr[52926] = -9561361;
assign addr[52927] = 9561361;
assign addr[52928] = 28683324;
assign addr[52929] = 47803013;
assign addr[52930] = 66918911;
assign addr[52931] = 86029503;
assign addr[52932] = 105133274;
assign addr[52933] = 124228708;
assign addr[52934] = 143314291;
assign addr[52935] = 162388511;
assign addr[52936] = 181449854;
assign addr[52937] = 200496809;
assign addr[52938] = 219527866;
assign addr[52939] = 238541516;
assign addr[52940] = 257536251;
assign addr[52941] = 276510565;
assign addr[52942] = 295462953;
assign addr[52943] = 314391913;
assign addr[52944] = 333295944;
assign addr[52945] = 352173546;
assign addr[52946] = 371023223;
assign addr[52947] = 389843480;
assign addr[52948] = 408632825;
assign addr[52949] = 427389768;
assign addr[52950] = 446112822;
assign addr[52951] = 464800501;
assign addr[52952] = 483451325;
assign addr[52953] = 502063814;
assign addr[52954] = 520636492;
assign addr[52955] = 539167887;
assign addr[52956] = 557656529;
assign addr[52957] = 576100953;
assign addr[52958] = 594499695;
assign addr[52959] = 612851297;
assign addr[52960] = 631154304;
assign addr[52961] = 649407264;
assign addr[52962] = 667608730;
assign addr[52963] = 685757258;
assign addr[52964] = 703851410;
assign addr[52965] = 721889752;
assign addr[52966] = 739870851;
assign addr[52967] = 757793284;
assign addr[52968] = 775655628;
assign addr[52969] = 793456467;
assign addr[52970] = 811194391;
assign addr[52971] = 828867991;
assign addr[52972] = 846475867;
assign addr[52973] = 864016623;
assign addr[52974] = 881488868;
assign addr[52975] = 898891215;
assign addr[52976] = 916222287;
assign addr[52977] = 933480707;
assign addr[52978] = 950665109;
assign addr[52979] = 967774128;
assign addr[52980] = 984806408;
assign addr[52981] = 1001760600;
assign addr[52982] = 1018635358;
assign addr[52983] = 1035429345;
assign addr[52984] = 1052141228;
assign addr[52985] = 1068769683;
assign addr[52986] = 1085313391;
assign addr[52987] = 1101771040;
assign addr[52988] = 1118141326;
assign addr[52989] = 1134422949;
assign addr[52990] = 1150614620;
assign addr[52991] = 1166715055;
assign addr[52992] = 1182722976;
assign addr[52993] = 1198637114;
assign addr[52994] = 1214456207;
assign addr[52995] = 1230179002;
assign addr[52996] = 1245804251;
assign addr[52997] = 1261330715;
assign addr[52998] = 1276757164;
assign addr[52999] = 1292082373;
assign addr[53000] = 1307305128;
assign addr[53001] = 1322424222;
assign addr[53002] = 1337438456;
assign addr[53003] = 1352346639;
assign addr[53004] = 1367147589;
assign addr[53005] = 1381840133;
assign addr[53006] = 1396423105;
assign addr[53007] = 1410895350;
assign addr[53008] = 1425255719;
assign addr[53009] = 1439503074;
assign addr[53010] = 1453636285;
assign addr[53011] = 1467654232;
assign addr[53012] = 1481555802;
assign addr[53013] = 1495339895;
assign addr[53014] = 1509005416;
assign addr[53015] = 1522551282;
assign addr[53016] = 1535976419;
assign addr[53017] = 1549279763;
assign addr[53018] = 1562460258;
assign addr[53019] = 1575516860;
assign addr[53020] = 1588448533;
assign addr[53021] = 1601254251;
assign addr[53022] = 1613933000;
assign addr[53023] = 1626483774;
assign addr[53024] = 1638905577;
assign addr[53025] = 1651197426;
assign addr[53026] = 1663358344;
assign addr[53027] = 1675387369;
assign addr[53028] = 1687283545;
assign addr[53029] = 1699045930;
assign addr[53030] = 1710673591;
assign addr[53031] = 1722165606;
assign addr[53032] = 1733521064;
assign addr[53033] = 1744739065;
assign addr[53034] = 1755818718;
assign addr[53035] = 1766759146;
assign addr[53036] = 1777559480;
assign addr[53037] = 1788218865;
assign addr[53038] = 1798736454;
assign addr[53039] = 1809111415;
assign addr[53040] = 1819342925;
assign addr[53041] = 1829430172;
assign addr[53042] = 1839372356;
assign addr[53043] = 1849168689;
assign addr[53044] = 1858818395;
assign addr[53045] = 1868320707;
assign addr[53046] = 1877674873;
assign addr[53047] = 1886880151;
assign addr[53048] = 1895935811;
assign addr[53049] = 1904841135;
assign addr[53050] = 1913595416;
assign addr[53051] = 1922197961;
assign addr[53052] = 1930648088;
assign addr[53053] = 1938945125;
assign addr[53054] = 1947088417;
assign addr[53055] = 1955077316;
assign addr[53056] = 1962911189;
assign addr[53057] = 1970589416;
assign addr[53058] = 1978111387;
assign addr[53059] = 1985476506;
assign addr[53060] = 1992684188;
assign addr[53061] = 1999733863;
assign addr[53062] = 2006624971;
assign addr[53063] = 2013356967;
assign addr[53064] = 2019929315;
assign addr[53065] = 2026341495;
assign addr[53066] = 2032592999;
assign addr[53067] = 2038683330;
assign addr[53068] = 2044612007;
assign addr[53069] = 2050378558;
assign addr[53070] = 2055982526;
assign addr[53071] = 2061423468;
assign addr[53072] = 2066700952;
assign addr[53073] = 2071814558;
assign addr[53074] = 2076763883;
assign addr[53075] = 2081548533;
assign addr[53076] = 2086168128;
assign addr[53077] = 2090622304;
assign addr[53078] = 2094910706;
assign addr[53079] = 2099032994;
assign addr[53080] = 2102988841;
assign addr[53081] = 2106777935;
assign addr[53082] = 2110399974;
assign addr[53083] = 2113854671;
assign addr[53084] = 2117141752;
assign addr[53085] = 2120260957;
assign addr[53086] = 2123212038;
assign addr[53087] = 2125994762;
assign addr[53088] = 2128608907;
assign addr[53089] = 2131054266;
assign addr[53090] = 2133330646;
assign addr[53091] = 2135437865;
assign addr[53092] = 2137375758;
assign addr[53093] = 2139144169;
assign addr[53094] = 2140742960;
assign addr[53095] = 2142172003;
assign addr[53096] = 2143431184;
assign addr[53097] = 2144520405;
assign addr[53098] = 2145439578;
assign addr[53099] = 2146188631;
assign addr[53100] = 2146767505;
assign addr[53101] = 2147176152;
assign addr[53102] = 2147414542;
assign addr[53103] = 2147482655;
assign addr[53104] = 2147380486;
assign addr[53105] = 2147108043;
assign addr[53106] = 2146665347;
assign addr[53107] = 2146052433;
assign addr[53108] = 2145269351;
assign addr[53109] = 2144316162;
assign addr[53110] = 2143192942;
assign addr[53111] = 2141899780;
assign addr[53112] = 2140436778;
assign addr[53113] = 2138804053;
assign addr[53114] = 2137001733;
assign addr[53115] = 2135029962;
assign addr[53116] = 2132888897;
assign addr[53117] = 2130578706;
assign addr[53118] = 2128099574;
assign addr[53119] = 2125451696;
assign addr[53120] = 2122635283;
assign addr[53121] = 2119650558;
assign addr[53122] = 2116497758;
assign addr[53123] = 2113177132;
assign addr[53124] = 2109688944;
assign addr[53125] = 2106033471;
assign addr[53126] = 2102211002;
assign addr[53127] = 2098221841;
assign addr[53128] = 2094066304;
assign addr[53129] = 2089744719;
assign addr[53130] = 2085257431;
assign addr[53131] = 2080604795;
assign addr[53132] = 2075787180;
assign addr[53133] = 2070804967;
assign addr[53134] = 2065658552;
assign addr[53135] = 2060348343;
assign addr[53136] = 2054874761;
assign addr[53137] = 2049238240;
assign addr[53138] = 2043439226;
assign addr[53139] = 2037478181;
assign addr[53140] = 2031355576;
assign addr[53141] = 2025071897;
assign addr[53142] = 2018627642;
assign addr[53143] = 2012023322;
assign addr[53144] = 2005259462;
assign addr[53145] = 1998336596;
assign addr[53146] = 1991255274;
assign addr[53147] = 1984016058;
assign addr[53148] = 1976619522;
assign addr[53149] = 1969066252;
assign addr[53150] = 1961356847;
assign addr[53151] = 1953491918;
assign addr[53152] = 1945472089;
assign addr[53153] = 1937297997;
assign addr[53154] = 1928970288;
assign addr[53155] = 1920489624;
assign addr[53156] = 1911856677;
assign addr[53157] = 1903072131;
assign addr[53158] = 1894136683;
assign addr[53159] = 1885051042;
assign addr[53160] = 1875815927;
assign addr[53161] = 1866432072;
assign addr[53162] = 1856900221;
assign addr[53163] = 1847221128;
assign addr[53164] = 1837395562;
assign addr[53165] = 1827424302;
assign addr[53166] = 1817308138;
assign addr[53167] = 1807047873;
assign addr[53168] = 1796644320;
assign addr[53169] = 1786098304;
assign addr[53170] = 1775410662;
assign addr[53171] = 1764582240;
assign addr[53172] = 1753613897;
assign addr[53173] = 1742506504;
assign addr[53174] = 1731260941;
assign addr[53175] = 1719878099;
assign addr[53176] = 1708358881;
assign addr[53177] = 1696704201;
assign addr[53178] = 1684914983;
assign addr[53179] = 1672992161;
assign addr[53180] = 1660936681;
assign addr[53181] = 1648749499;
assign addr[53182] = 1636431582;
assign addr[53183] = 1623983905;
assign addr[53184] = 1611407456;
assign addr[53185] = 1598703233;
assign addr[53186] = 1585872242;
assign addr[53187] = 1572915501;
assign addr[53188] = 1559834037;
assign addr[53189] = 1546628888;
assign addr[53190] = 1533301101;
assign addr[53191] = 1519851733;
assign addr[53192] = 1506281850;
assign addr[53193] = 1492592527;
assign addr[53194] = 1478784851;
assign addr[53195] = 1464859917;
assign addr[53196] = 1450818828;
assign addr[53197] = 1436662698;
assign addr[53198] = 1422392650;
assign addr[53199] = 1408009814;
assign addr[53200] = 1393515332;
assign addr[53201] = 1378910353;
assign addr[53202] = 1364196034;
assign addr[53203] = 1349373543;
assign addr[53204] = 1334444055;
assign addr[53205] = 1319408754;
assign addr[53206] = 1304268832;
assign addr[53207] = 1289025489;
assign addr[53208] = 1273679934;
assign addr[53209] = 1258233384;
assign addr[53210] = 1242687064;
assign addr[53211] = 1227042207;
assign addr[53212] = 1211300053;
assign addr[53213] = 1195461849;
assign addr[53214] = 1179528853;
assign addr[53215] = 1163502328;
assign addr[53216] = 1147383544;
assign addr[53217] = 1131173780;
assign addr[53218] = 1114874320;
assign addr[53219] = 1098486458;
assign addr[53220] = 1082011492;
assign addr[53221] = 1065450729;
assign addr[53222] = 1048805483;
assign addr[53223] = 1032077073;
assign addr[53224] = 1015266825;
assign addr[53225] = 998376073;
assign addr[53226] = 981406156;
assign addr[53227] = 964358420;
assign addr[53228] = 947234215;
assign addr[53229] = 930034901;
assign addr[53230] = 912761841;
assign addr[53231] = 895416404;
assign addr[53232] = 877999966;
assign addr[53233] = 860513908;
assign addr[53234] = 842959617;
assign addr[53235] = 825338484;
assign addr[53236] = 807651907;
assign addr[53237] = 789901288;
assign addr[53238] = 772088034;
assign addr[53239] = 754213559;
assign addr[53240] = 736279279;
assign addr[53241] = 718286617;
assign addr[53242] = 700236999;
assign addr[53243] = 682131857;
assign addr[53244] = 663972625;
assign addr[53245] = 645760745;
assign addr[53246] = 627497660;
assign addr[53247] = 609184818;
assign addr[53248] = 590823671;
assign addr[53249] = 572415676;
assign addr[53250] = 553962291;
assign addr[53251] = 535464981;
assign addr[53252] = 516925212;
assign addr[53253] = 498344454;
assign addr[53254] = 479724180;
assign addr[53255] = 461065866;
assign addr[53256] = 442370993;
assign addr[53257] = 423641043;
assign addr[53258] = 404877501;
assign addr[53259] = 386081854;
assign addr[53260] = 367255594;
assign addr[53261] = 348400212;
assign addr[53262] = 329517204;
assign addr[53263] = 310608068;
assign addr[53264] = 291674302;
assign addr[53265] = 272717408;
assign addr[53266] = 253738890;
assign addr[53267] = 234740251;
assign addr[53268] = 215722999;
assign addr[53269] = 196688642;
assign addr[53270] = 177638688;
assign addr[53271] = 158574649;
assign addr[53272] = 139498035;
assign addr[53273] = 120410361;
assign addr[53274] = 101313138;
assign addr[53275] = 82207882;
assign addr[53276] = 63096108;
assign addr[53277] = 43979330;
assign addr[53278] = 24859065;
assign addr[53279] = 5736829;
assign addr[53280] = -13385863;
assign addr[53281] = -32507492;
assign addr[53282] = -51626544;
assign addr[53283] = -70741503;
assign addr[53284] = -89850852;
assign addr[53285] = -108953076;
assign addr[53286] = -128046661;
assign addr[53287] = -147130093;
assign addr[53288] = -166201858;
assign addr[53289] = -185260444;
assign addr[53290] = -204304341;
assign addr[53291] = -223332037;
assign addr[53292] = -242342025;
assign addr[53293] = -261332796;
assign addr[53294] = -280302845;
assign addr[53295] = -299250668;
assign addr[53296] = -318174762;
assign addr[53297] = -337073627;
assign addr[53298] = -355945764;
assign addr[53299] = -374789676;
assign addr[53300] = -393603870;
assign addr[53301] = -412386854;
assign addr[53302] = -431137138;
assign addr[53303] = -449853235;
assign addr[53304] = -468533662;
assign addr[53305] = -487176937;
assign addr[53306] = -505781581;
assign addr[53307] = -524346121;
assign addr[53308] = -542869083;
assign addr[53309] = -561348998;
assign addr[53310] = -579784402;
assign addr[53311] = -598173833;
assign addr[53312] = -616515832;
assign addr[53313] = -634808946;
assign addr[53314] = -653051723;
assign addr[53315] = -671242716;
assign addr[53316] = -689380485;
assign addr[53317] = -707463589;
assign addr[53318] = -725490597;
assign addr[53319] = -743460077;
assign addr[53320] = -761370605;
assign addr[53321] = -779220762;
assign addr[53322] = -797009130;
assign addr[53323] = -814734301;
assign addr[53324] = -832394869;
assign addr[53325] = -849989433;
assign addr[53326] = -867516597;
assign addr[53327] = -884974973;
assign addr[53328] = -902363176;
assign addr[53329] = -919679827;
assign addr[53330] = -936923553;
assign addr[53331] = -954092986;
assign addr[53332] = -971186766;
assign addr[53333] = -988203537;
assign addr[53334] = -1005141949;
assign addr[53335] = -1022000660;
assign addr[53336] = -1038778332;
assign addr[53337] = -1055473635;
assign addr[53338] = -1072085246;
assign addr[53339] = -1088611847;
assign addr[53340] = -1105052128;
assign addr[53341] = -1121404785;
assign addr[53342] = -1137668521;
assign addr[53343] = -1153842047;
assign addr[53344] = -1169924081;
assign addr[53345] = -1185913346;
assign addr[53346] = -1201808576;
assign addr[53347] = -1217608510;
assign addr[53348] = -1233311895;
assign addr[53349] = -1248917486;
assign addr[53350] = -1264424045;
assign addr[53351] = -1279830344;
assign addr[53352] = -1295135159;
assign addr[53353] = -1310337279;
assign addr[53354] = -1325435496;
assign addr[53355] = -1340428615;
assign addr[53356] = -1355315445;
assign addr[53357] = -1370094808;
assign addr[53358] = -1384765530;
assign addr[53359] = -1399326449;
assign addr[53360] = -1413776410;
assign addr[53361] = -1428114267;
assign addr[53362] = -1442338884;
assign addr[53363] = -1456449131;
assign addr[53364] = -1470443891;
assign addr[53365] = -1484322054;
assign addr[53366] = -1498082520;
assign addr[53367] = -1511724196;
assign addr[53368] = -1525246002;
assign addr[53369] = -1538646865;
assign addr[53370] = -1551925723;
assign addr[53371] = -1565081523;
assign addr[53372] = -1578113222;
assign addr[53373] = -1591019785;
assign addr[53374] = -1603800191;
assign addr[53375] = -1616453425;
assign addr[53376] = -1628978484;
assign addr[53377] = -1641374375;
assign addr[53378] = -1653640115;
assign addr[53379] = -1665774731;
assign addr[53380] = -1677777262;
assign addr[53381] = -1689646755;
assign addr[53382] = -1701382270;
assign addr[53383] = -1712982875;
assign addr[53384] = -1724447652;
assign addr[53385] = -1735775690;
assign addr[53386] = -1746966091;
assign addr[53387] = -1758017969;
assign addr[53388] = -1768930447;
assign addr[53389] = -1779702660;
assign addr[53390] = -1790333753;
assign addr[53391] = -1800822883;
assign addr[53392] = -1811169220;
assign addr[53393] = -1821371941;
assign addr[53394] = -1831430239;
assign addr[53395] = -1841343316;
assign addr[53396] = -1851110385;
assign addr[53397] = -1860730673;
assign addr[53398] = -1870203416;
assign addr[53399] = -1879527863;
assign addr[53400] = -1888703276;
assign addr[53401] = -1897728925;
assign addr[53402] = -1906604097;
assign addr[53403] = -1915328086;
assign addr[53404] = -1923900201;
assign addr[53405] = -1932319763;
assign addr[53406] = -1940586104;
assign addr[53407] = -1948698568;
assign addr[53408] = -1956656513;
assign addr[53409] = -1964459306;
assign addr[53410] = -1972106330;
assign addr[53411] = -1979596978;
assign addr[53412] = -1986930656;
assign addr[53413] = -1994106782;
assign addr[53414] = -2001124788;
assign addr[53415] = -2007984117;
assign addr[53416] = -2014684225;
assign addr[53417] = -2021224581;
assign addr[53418] = -2027604666;
assign addr[53419] = -2033823974;
assign addr[53420] = -2039882013;
assign addr[53421] = -2045778302;
assign addr[53422] = -2051512372;
assign addr[53423] = -2057083771;
assign addr[53424] = -2062492055;
assign addr[53425] = -2067736796;
assign addr[53426] = -2072817579;
assign addr[53427] = -2077733999;
assign addr[53428] = -2082485668;
assign addr[53429] = -2087072209;
assign addr[53430] = -2091493257;
assign addr[53431] = -2095748463;
assign addr[53432] = -2099837489;
assign addr[53433] = -2103760010;
assign addr[53434] = -2107515716;
assign addr[53435] = -2111104309;
assign addr[53436] = -2114525505;
assign addr[53437] = -2117779031;
assign addr[53438] = -2120864631;
assign addr[53439] = -2123782059;
assign addr[53440] = -2126531084;
assign addr[53441] = -2129111488;
assign addr[53442] = -2131523066;
assign addr[53443] = -2133765628;
assign addr[53444] = -2135838995;
assign addr[53445] = -2137743003;
assign addr[53446] = -2139477502;
assign addr[53447] = -2141042352;
assign addr[53448] = -2142437431;
assign addr[53449] = -2143662628;
assign addr[53450] = -2144717846;
assign addr[53451] = -2145603001;
assign addr[53452] = -2146318022;
assign addr[53453] = -2146862854;
assign addr[53454] = -2147237452;
assign addr[53455] = -2147441787;
assign addr[53456] = -2147475844;
assign addr[53457] = -2147339619;
assign addr[53458] = -2147033123;
assign addr[53459] = -2146556380;
assign addr[53460] = -2145909429;
assign addr[53461] = -2145092320;
assign addr[53462] = -2144105118;
assign addr[53463] = -2142947902;
assign addr[53464] = -2141620763;
assign addr[53465] = -2140123807;
assign addr[53466] = -2138457152;
assign addr[53467] = -2136620930;
assign addr[53468] = -2134615288;
assign addr[53469] = -2132440383;
assign addr[53470] = -2130096389;
assign addr[53471] = -2127583492;
assign addr[53472] = -2124901890;
assign addr[53473] = -2122051796;
assign addr[53474] = -2119033436;
assign addr[53475] = -2115847050;
assign addr[53476] = -2112492891;
assign addr[53477] = -2108971223;
assign addr[53478] = -2105282327;
assign addr[53479] = -2101426496;
assign addr[53480] = -2097404033;
assign addr[53481] = -2093215260;
assign addr[53482] = -2088860507;
assign addr[53483] = -2084340120;
assign addr[53484] = -2079654458;
assign addr[53485] = -2074803892;
assign addr[53486] = -2069788807;
assign addr[53487] = -2064609600;
assign addr[53488] = -2059266683;
assign addr[53489] = -2053760478;
assign addr[53490] = -2048091422;
assign addr[53491] = -2042259965;
assign addr[53492] = -2036266570;
assign addr[53493] = -2030111710;
assign addr[53494] = -2023795876;
assign addr[53495] = -2017319567;
assign addr[53496] = -2010683297;
assign addr[53497] = -2003887591;
assign addr[53498] = -1996932990;
assign addr[53499] = -1989820044;
assign addr[53500] = -1982549318;
assign addr[53501] = -1975121388;
assign addr[53502] = -1967536842;
assign addr[53503] = -1959796283;
assign addr[53504] = -1951900324;
assign addr[53505] = -1943849591;
assign addr[53506] = -1935644723;
assign addr[53507] = -1927286370;
assign addr[53508] = -1918775195;
assign addr[53509] = -1910111873;
assign addr[53510] = -1901297091;
assign addr[53511] = -1892331547;
assign addr[53512] = -1883215953;
assign addr[53513] = -1873951032;
assign addr[53514] = -1864537518;
assign addr[53515] = -1854976157;
assign addr[53516] = -1845267708;
assign addr[53517] = -1835412941;
assign addr[53518] = -1825412636;
assign addr[53519] = -1815267588;
assign addr[53520] = -1804978599;
assign addr[53521] = -1794546487;
assign addr[53522] = -1783972079;
assign addr[53523] = -1773256212;
assign addr[53524] = -1762399737;
assign addr[53525] = -1751403515;
assign addr[53526] = -1740268417;
assign addr[53527] = -1728995326;
assign addr[53528] = -1717585136;
assign addr[53529] = -1706038753;
assign addr[53530] = -1694357091;
assign addr[53531] = -1682541077;
assign addr[53532] = -1670591647;
assign addr[53533] = -1658509750;
assign addr[53534] = -1646296344;
assign addr[53535] = -1633952396;
assign addr[53536] = -1621478885;
assign addr[53537] = -1608876801;
assign addr[53538] = -1596147143;
assign addr[53539] = -1583290921;
assign addr[53540] = -1570309153;
assign addr[53541] = -1557202869;
assign addr[53542] = -1543973108;
assign addr[53543] = -1530620920;
assign addr[53544] = -1517147363;
assign addr[53545] = -1503553506;
assign addr[53546] = -1489840425;
assign addr[53547] = -1476009210;
assign addr[53548] = -1462060956;
assign addr[53549] = -1447996770;
assign addr[53550] = -1433817766;
assign addr[53551] = -1419525069;
assign addr[53552] = -1405119813;
assign addr[53553] = -1390603139;
assign addr[53554] = -1375976199;
assign addr[53555] = -1361240152;
assign addr[53556] = -1346396168;
assign addr[53557] = -1331445422;
assign addr[53558] = -1316389101;
assign addr[53559] = -1301228398;
assign addr[53560] = -1285964516;
assign addr[53561] = -1270598665;
assign addr[53562] = -1255132063;
assign addr[53563] = -1239565936;
assign addr[53564] = -1223901520;
assign addr[53565] = -1208140056;
assign addr[53566] = -1192282793;
assign addr[53567] = -1176330990;
assign addr[53568] = -1160285911;
assign addr[53569] = -1144148829;
assign addr[53570] = -1127921022;
assign addr[53571] = -1111603778;
assign addr[53572] = -1095198391;
assign addr[53573] = -1078706161;
assign addr[53574] = -1062128397;
assign addr[53575] = -1045466412;
assign addr[53576] = -1028721528;
assign addr[53577] = -1011895073;
assign addr[53578] = -994988380;
assign addr[53579] = -978002791;
assign addr[53580] = -960939653;
assign addr[53581] = -943800318;
assign addr[53582] = -926586145;
assign addr[53583] = -909298500;
assign addr[53584] = -891938752;
assign addr[53585] = -874508280;
assign addr[53586] = -857008464;
assign addr[53587] = -839440693;
assign addr[53588] = -821806359;
assign addr[53589] = -804106861;
assign addr[53590] = -786343603;
assign addr[53591] = -768517992;
assign addr[53592] = -750631442;
assign addr[53593] = -732685372;
assign addr[53594] = -714681204;
assign addr[53595] = -696620367;
assign addr[53596] = -678504291;
assign addr[53597] = -660334415;
assign addr[53598] = -642112178;
assign addr[53599] = -623839025;
assign addr[53600] = -605516406;
assign addr[53601] = -587145773;
assign addr[53602] = -568728583;
assign addr[53603] = -550266296;
assign addr[53604] = -531760377;
assign addr[53605] = -513212292;
assign addr[53606] = -494623513;
assign addr[53607] = -475995513;
assign addr[53608] = -457329769;
assign addr[53609] = -438627762;
assign addr[53610] = -419890975;
assign addr[53611] = -401120892;
assign addr[53612] = -382319004;
assign addr[53613] = -363486799;
assign addr[53614] = -344625773;
assign addr[53615] = -325737419;
assign addr[53616] = -306823237;
assign addr[53617] = -287884725;
assign addr[53618] = -268923386;
assign addr[53619] = -249940723;
assign addr[53620] = -230938242;
assign addr[53621] = -211917448;
assign addr[53622] = -192879850;
assign addr[53623] = -173826959;
assign addr[53624] = -154760284;
assign addr[53625] = -135681337;
assign addr[53626] = -116591632;
assign addr[53627] = -97492681;
assign addr[53628] = -78386000;
assign addr[53629] = -59273104;
assign addr[53630] = -40155507;
assign addr[53631] = -21034727;
assign addr[53632] = -1912278;
assign addr[53633] = 17210322;
assign addr[53634] = 36331557;
assign addr[53635] = 55449912;
assign addr[53636] = 74563870;
assign addr[53637] = 93671915;
assign addr[53638] = 112772533;
assign addr[53639] = 131864208;
assign addr[53640] = 150945428;
assign addr[53641] = 170014678;
assign addr[53642] = 189070447;
assign addr[53643] = 208111224;
assign addr[53644] = 227135500;
assign addr[53645] = 246141764;
assign addr[53646] = 265128512;
assign addr[53647] = 284094236;
assign addr[53648] = 303037433;
assign addr[53649] = 321956601;
assign addr[53650] = 340850240;
assign addr[53651] = 359716852;
assign addr[53652] = 378554940;
assign addr[53653] = 397363011;
assign addr[53654] = 416139574;
assign addr[53655] = 434883140;
assign addr[53656] = 453592221;
assign addr[53657] = 472265336;
assign addr[53658] = 490901003;
assign addr[53659] = 509497745;
assign addr[53660] = 528054086;
assign addr[53661] = 546568556;
assign addr[53662] = 565039687;
assign addr[53663] = 583466013;
assign addr[53664] = 601846074;
assign addr[53665] = 620178412;
assign addr[53666] = 638461574;
assign addr[53667] = 656694110;
assign addr[53668] = 674874574;
assign addr[53669] = 693001525;
assign addr[53670] = 711073524;
assign addr[53671] = 729089140;
assign addr[53672] = 747046944;
assign addr[53673] = 764945512;
assign addr[53674] = 782783424;
assign addr[53675] = 800559266;
assign addr[53676] = 818271628;
assign addr[53677] = 835919107;
assign addr[53678] = 853500302;
assign addr[53679] = 871013820;
assign addr[53680] = 888458272;
assign addr[53681] = 905832274;
assign addr[53682] = 923134450;
assign addr[53683] = 940363427;
assign addr[53684] = 957517838;
assign addr[53685] = 974596324;
assign addr[53686] = 991597531;
assign addr[53687] = 1008520110;
assign addr[53688] = 1025362720;
assign addr[53689] = 1042124025;
assign addr[53690] = 1058802695;
assign addr[53691] = 1075397409;
assign addr[53692] = 1091906851;
assign addr[53693] = 1108329711;
assign addr[53694] = 1124664687;
assign addr[53695] = 1140910484;
assign addr[53696] = 1157065814;
assign addr[53697] = 1173129396;
assign addr[53698] = 1189099956;
assign addr[53699] = 1204976227;
assign addr[53700] = 1220756951;
assign addr[53701] = 1236440877;
assign addr[53702] = 1252026760;
assign addr[53703] = 1267513365;
assign addr[53704] = 1282899464;
assign addr[53705] = 1298183838;
assign addr[53706] = 1313365273;
assign addr[53707] = 1328442566;
assign addr[53708] = 1343414522;
assign addr[53709] = 1358279953;
assign addr[53710] = 1373037681;
assign addr[53711] = 1387686535;
assign addr[53712] = 1402225355;
assign addr[53713] = 1416652986;
assign addr[53714] = 1430968286;
assign addr[53715] = 1445170118;
assign addr[53716] = 1459257358;
assign addr[53717] = 1473228887;
assign addr[53718] = 1487083598;
assign addr[53719] = 1500820393;
assign addr[53720] = 1514438181;
assign addr[53721] = 1527935884;
assign addr[53722] = 1541312431;
assign addr[53723] = 1554566762;
assign addr[53724] = 1567697824;
assign addr[53725] = 1580704578;
assign addr[53726] = 1593585992;
assign addr[53727] = 1606341043;
assign addr[53728] = 1618968722;
assign addr[53729] = 1631468027;
assign addr[53730] = 1643837966;
assign addr[53731] = 1656077559;
assign addr[53732] = 1668185835;
assign addr[53733] = 1680161834;
assign addr[53734] = 1692004606;
assign addr[53735] = 1703713213;
assign addr[53736] = 1715286726;
assign addr[53737] = 1726724227;
assign addr[53738] = 1738024810;
assign addr[53739] = 1749187577;
assign addr[53740] = 1760211645;
assign addr[53741] = 1771096139;
assign addr[53742] = 1781840195;
assign addr[53743] = 1792442963;
assign addr[53744] = 1802903601;
assign addr[53745] = 1813221279;
assign addr[53746] = 1823395180;
assign addr[53747] = 1833424497;
assign addr[53748] = 1843308435;
assign addr[53749] = 1853046210;
assign addr[53750] = 1862637049;
assign addr[53751] = 1872080193;
assign addr[53752] = 1881374892;
assign addr[53753] = 1890520410;
assign addr[53754] = 1899516021;
assign addr[53755] = 1908361011;
assign addr[53756] = 1917054681;
assign addr[53757] = 1925596340;
assign addr[53758] = 1933985310;
assign addr[53759] = 1942220928;
assign addr[53760] = 1950302539;
assign addr[53761] = 1958229503;
assign addr[53762] = 1966001192;
assign addr[53763] = 1973616989;
assign addr[53764] = 1981076290;
assign addr[53765] = 1988378503;
assign addr[53766] = 1995523051;
assign addr[53767] = 2002509365;
assign addr[53768] = 2009336893;
assign addr[53769] = 2016005093;
assign addr[53770] = 2022513436;
assign addr[53771] = 2028861406;
assign addr[53772] = 2035048499;
assign addr[53773] = 2041074226;
assign addr[53774] = 2046938108;
assign addr[53775] = 2052639680;
assign addr[53776] = 2058178491;
assign addr[53777] = 2063554100;
assign addr[53778] = 2068766083;
assign addr[53779] = 2073814024;
assign addr[53780] = 2078697525;
assign addr[53781] = 2083416198;
assign addr[53782] = 2087969669;
assign addr[53783] = 2092357577;
assign addr[53784] = 2096579573;
assign addr[53785] = 2100635323;
assign addr[53786] = 2104524506;
assign addr[53787] = 2108246813;
assign addr[53788] = 2111801949;
assign addr[53789] = 2115189632;
assign addr[53790] = 2118409593;
assign addr[53791] = 2121461578;
assign addr[53792] = 2124345343;
assign addr[53793] = 2127060661;
assign addr[53794] = 2129607316;
assign addr[53795] = 2131985106;
assign addr[53796] = 2134193842;
assign addr[53797] = 2136233350;
assign addr[53798] = 2138103468;
assign addr[53799] = 2139804048;
assign addr[53800] = 2141334954;
assign addr[53801] = 2142696065;
assign addr[53802] = 2143887273;
assign addr[53803] = 2144908484;
assign addr[53804] = 2145759618;
assign addr[53805] = 2146440605;
assign addr[53806] = 2146951393;
assign addr[53807] = 2147291941;
assign addr[53808] = 2147462221;
assign addr[53809] = 2147462221;
assign addr[53810] = 2147291941;
assign addr[53811] = 2146951393;
assign addr[53812] = 2146440605;
assign addr[53813] = 2145759618;
assign addr[53814] = 2144908484;
assign addr[53815] = 2143887273;
assign addr[53816] = 2142696065;
assign addr[53817] = 2141334954;
assign addr[53818] = 2139804048;
assign addr[53819] = 2138103468;
assign addr[53820] = 2136233350;
assign addr[53821] = 2134193842;
assign addr[53822] = 2131985106;
assign addr[53823] = 2129607316;
assign addr[53824] = 2127060661;
assign addr[53825] = 2124345343;
assign addr[53826] = 2121461578;
assign addr[53827] = 2118409593;
assign addr[53828] = 2115189632;
assign addr[53829] = 2111801949;
assign addr[53830] = 2108246813;
assign addr[53831] = 2104524506;
assign addr[53832] = 2100635323;
assign addr[53833] = 2096579573;
assign addr[53834] = 2092357577;
assign addr[53835] = 2087969669;
assign addr[53836] = 2083416198;
assign addr[53837] = 2078697525;
assign addr[53838] = 2073814024;
assign addr[53839] = 2068766083;
assign addr[53840] = 2063554100;
assign addr[53841] = 2058178491;
assign addr[53842] = 2052639680;
assign addr[53843] = 2046938108;
assign addr[53844] = 2041074226;
assign addr[53845] = 2035048499;
assign addr[53846] = 2028861406;
assign addr[53847] = 2022513436;
assign addr[53848] = 2016005093;
assign addr[53849] = 2009336893;
assign addr[53850] = 2002509365;
assign addr[53851] = 1995523051;
assign addr[53852] = 1988378503;
assign addr[53853] = 1981076290;
assign addr[53854] = 1973616989;
assign addr[53855] = 1966001192;
assign addr[53856] = 1958229503;
assign addr[53857] = 1950302539;
assign addr[53858] = 1942220928;
assign addr[53859] = 1933985310;
assign addr[53860] = 1925596340;
assign addr[53861] = 1917054681;
assign addr[53862] = 1908361011;
assign addr[53863] = 1899516021;
assign addr[53864] = 1890520410;
assign addr[53865] = 1881374892;
assign addr[53866] = 1872080193;
assign addr[53867] = 1862637049;
assign addr[53868] = 1853046210;
assign addr[53869] = 1843308435;
assign addr[53870] = 1833424497;
assign addr[53871] = 1823395180;
assign addr[53872] = 1813221279;
assign addr[53873] = 1802903601;
assign addr[53874] = 1792442963;
assign addr[53875] = 1781840195;
assign addr[53876] = 1771096139;
assign addr[53877] = 1760211645;
assign addr[53878] = 1749187577;
assign addr[53879] = 1738024810;
assign addr[53880] = 1726724227;
assign addr[53881] = 1715286726;
assign addr[53882] = 1703713213;
assign addr[53883] = 1692004606;
assign addr[53884] = 1680161834;
assign addr[53885] = 1668185835;
assign addr[53886] = 1656077559;
assign addr[53887] = 1643837966;
assign addr[53888] = 1631468027;
assign addr[53889] = 1618968722;
assign addr[53890] = 1606341043;
assign addr[53891] = 1593585992;
assign addr[53892] = 1580704578;
assign addr[53893] = 1567697824;
assign addr[53894] = 1554566762;
assign addr[53895] = 1541312431;
assign addr[53896] = 1527935884;
assign addr[53897] = 1514438181;
assign addr[53898] = 1500820393;
assign addr[53899] = 1487083598;
assign addr[53900] = 1473228887;
assign addr[53901] = 1459257358;
assign addr[53902] = 1445170118;
assign addr[53903] = 1430968286;
assign addr[53904] = 1416652986;
assign addr[53905] = 1402225355;
assign addr[53906] = 1387686535;
assign addr[53907] = 1373037681;
assign addr[53908] = 1358279953;
assign addr[53909] = 1343414522;
assign addr[53910] = 1328442566;
assign addr[53911] = 1313365273;
assign addr[53912] = 1298183838;
assign addr[53913] = 1282899464;
assign addr[53914] = 1267513365;
assign addr[53915] = 1252026760;
assign addr[53916] = 1236440877;
assign addr[53917] = 1220756951;
assign addr[53918] = 1204976227;
assign addr[53919] = 1189099956;
assign addr[53920] = 1173129396;
assign addr[53921] = 1157065814;
assign addr[53922] = 1140910484;
assign addr[53923] = 1124664687;
assign addr[53924] = 1108329711;
assign addr[53925] = 1091906851;
assign addr[53926] = 1075397409;
assign addr[53927] = 1058802695;
assign addr[53928] = 1042124025;
assign addr[53929] = 1025362720;
assign addr[53930] = 1008520110;
assign addr[53931] = 991597531;
assign addr[53932] = 974596324;
assign addr[53933] = 957517838;
assign addr[53934] = 940363427;
assign addr[53935] = 923134450;
assign addr[53936] = 905832274;
assign addr[53937] = 888458272;
assign addr[53938] = 871013820;
assign addr[53939] = 853500302;
assign addr[53940] = 835919107;
assign addr[53941] = 818271628;
assign addr[53942] = 800559266;
assign addr[53943] = 782783424;
assign addr[53944] = 764945512;
assign addr[53945] = 747046944;
assign addr[53946] = 729089140;
assign addr[53947] = 711073524;
assign addr[53948] = 693001525;
assign addr[53949] = 674874574;
assign addr[53950] = 656694110;
assign addr[53951] = 638461574;
assign addr[53952] = 620178412;
assign addr[53953] = 601846074;
assign addr[53954] = 583466013;
assign addr[53955] = 565039687;
assign addr[53956] = 546568556;
assign addr[53957] = 528054086;
assign addr[53958] = 509497745;
assign addr[53959] = 490901003;
assign addr[53960] = 472265336;
assign addr[53961] = 453592221;
assign addr[53962] = 434883140;
assign addr[53963] = 416139574;
assign addr[53964] = 397363011;
assign addr[53965] = 378554940;
assign addr[53966] = 359716852;
assign addr[53967] = 340850240;
assign addr[53968] = 321956601;
assign addr[53969] = 303037433;
assign addr[53970] = 284094236;
assign addr[53971] = 265128512;
assign addr[53972] = 246141764;
assign addr[53973] = 227135500;
assign addr[53974] = 208111224;
assign addr[53975] = 189070447;
assign addr[53976] = 170014678;
assign addr[53977] = 150945428;
assign addr[53978] = 131864208;
assign addr[53979] = 112772533;
assign addr[53980] = 93671915;
assign addr[53981] = 74563870;
assign addr[53982] = 55449912;
assign addr[53983] = 36331557;
assign addr[53984] = 17210322;
assign addr[53985] = -1912278;
assign addr[53986] = -21034727;
assign addr[53987] = -40155507;
assign addr[53988] = -59273104;
assign addr[53989] = -78386000;
assign addr[53990] = -97492681;
assign addr[53991] = -116591632;
assign addr[53992] = -135681337;
assign addr[53993] = -154760284;
assign addr[53994] = -173826959;
assign addr[53995] = -192879850;
assign addr[53996] = -211917448;
assign addr[53997] = -230938242;
assign addr[53998] = -249940723;
assign addr[53999] = -268923386;
assign addr[54000] = -287884725;
assign addr[54001] = -306823237;
assign addr[54002] = -325737419;
assign addr[54003] = -344625773;
assign addr[54004] = -363486799;
assign addr[54005] = -382319004;
assign addr[54006] = -401120892;
assign addr[54007] = -419890975;
assign addr[54008] = -438627762;
assign addr[54009] = -457329769;
assign addr[54010] = -475995513;
assign addr[54011] = -494623513;
assign addr[54012] = -513212292;
assign addr[54013] = -531760377;
assign addr[54014] = -550266296;
assign addr[54015] = -568728583;
assign addr[54016] = -587145773;
assign addr[54017] = -605516406;
assign addr[54018] = -623839025;
assign addr[54019] = -642112178;
assign addr[54020] = -660334415;
assign addr[54021] = -678504291;
assign addr[54022] = -696620367;
assign addr[54023] = -714681204;
assign addr[54024] = -732685372;
assign addr[54025] = -750631442;
assign addr[54026] = -768517992;
assign addr[54027] = -786343603;
assign addr[54028] = -804106861;
assign addr[54029] = -821806359;
assign addr[54030] = -839440693;
assign addr[54031] = -857008464;
assign addr[54032] = -874508280;
assign addr[54033] = -891938752;
assign addr[54034] = -909298500;
assign addr[54035] = -926586145;
assign addr[54036] = -943800318;
assign addr[54037] = -960939653;
assign addr[54038] = -978002791;
assign addr[54039] = -994988380;
assign addr[54040] = -1011895073;
assign addr[54041] = -1028721528;
assign addr[54042] = -1045466412;
assign addr[54043] = -1062128397;
assign addr[54044] = -1078706161;
assign addr[54045] = -1095198391;
assign addr[54046] = -1111603778;
assign addr[54047] = -1127921022;
assign addr[54048] = -1144148829;
assign addr[54049] = -1160285911;
assign addr[54050] = -1176330990;
assign addr[54051] = -1192282793;
assign addr[54052] = -1208140056;
assign addr[54053] = -1223901520;
assign addr[54054] = -1239565936;
assign addr[54055] = -1255132063;
assign addr[54056] = -1270598665;
assign addr[54057] = -1285964516;
assign addr[54058] = -1301228398;
assign addr[54059] = -1316389101;
assign addr[54060] = -1331445422;
assign addr[54061] = -1346396168;
assign addr[54062] = -1361240152;
assign addr[54063] = -1375976199;
assign addr[54064] = -1390603139;
assign addr[54065] = -1405119813;
assign addr[54066] = -1419525069;
assign addr[54067] = -1433817766;
assign addr[54068] = -1447996770;
assign addr[54069] = -1462060956;
assign addr[54070] = -1476009210;
assign addr[54071] = -1489840425;
assign addr[54072] = -1503553506;
assign addr[54073] = -1517147363;
assign addr[54074] = -1530620920;
assign addr[54075] = -1543973108;
assign addr[54076] = -1557202869;
assign addr[54077] = -1570309153;
assign addr[54078] = -1583290921;
assign addr[54079] = -1596147143;
assign addr[54080] = -1608876801;
assign addr[54081] = -1621478885;
assign addr[54082] = -1633952396;
assign addr[54083] = -1646296344;
assign addr[54084] = -1658509750;
assign addr[54085] = -1670591647;
assign addr[54086] = -1682541077;
assign addr[54087] = -1694357091;
assign addr[54088] = -1706038753;
assign addr[54089] = -1717585136;
assign addr[54090] = -1728995326;
assign addr[54091] = -1740268417;
assign addr[54092] = -1751403515;
assign addr[54093] = -1762399737;
assign addr[54094] = -1773256212;
assign addr[54095] = -1783972079;
assign addr[54096] = -1794546487;
assign addr[54097] = -1804978599;
assign addr[54098] = -1815267588;
assign addr[54099] = -1825412636;
assign addr[54100] = -1835412941;
assign addr[54101] = -1845267708;
assign addr[54102] = -1854976157;
assign addr[54103] = -1864537518;
assign addr[54104] = -1873951032;
assign addr[54105] = -1883215953;
assign addr[54106] = -1892331547;
assign addr[54107] = -1901297091;
assign addr[54108] = -1910111873;
assign addr[54109] = -1918775195;
assign addr[54110] = -1927286370;
assign addr[54111] = -1935644723;
assign addr[54112] = -1943849591;
assign addr[54113] = -1951900324;
assign addr[54114] = -1959796283;
assign addr[54115] = -1967536842;
assign addr[54116] = -1975121388;
assign addr[54117] = -1982549318;
assign addr[54118] = -1989820044;
assign addr[54119] = -1996932990;
assign addr[54120] = -2003887591;
assign addr[54121] = -2010683297;
assign addr[54122] = -2017319567;
assign addr[54123] = -2023795876;
assign addr[54124] = -2030111710;
assign addr[54125] = -2036266570;
assign addr[54126] = -2042259965;
assign addr[54127] = -2048091422;
assign addr[54128] = -2053760478;
assign addr[54129] = -2059266683;
assign addr[54130] = -2064609600;
assign addr[54131] = -2069788807;
assign addr[54132] = -2074803892;
assign addr[54133] = -2079654458;
assign addr[54134] = -2084340120;
assign addr[54135] = -2088860507;
assign addr[54136] = -2093215260;
assign addr[54137] = -2097404033;
assign addr[54138] = -2101426496;
assign addr[54139] = -2105282327;
assign addr[54140] = -2108971223;
assign addr[54141] = -2112492891;
assign addr[54142] = -2115847050;
assign addr[54143] = -2119033436;
assign addr[54144] = -2122051796;
assign addr[54145] = -2124901890;
assign addr[54146] = -2127583492;
assign addr[54147] = -2130096389;
assign addr[54148] = -2132440383;
assign addr[54149] = -2134615288;
assign addr[54150] = -2136620930;
assign addr[54151] = -2138457152;
assign addr[54152] = -2140123807;
assign addr[54153] = -2141620763;
assign addr[54154] = -2142947902;
assign addr[54155] = -2144105118;
assign addr[54156] = -2145092320;
assign addr[54157] = -2145909429;
assign addr[54158] = -2146556380;
assign addr[54159] = -2147033123;
assign addr[54160] = -2147339619;
assign addr[54161] = -2147475844;
assign addr[54162] = -2147441787;
assign addr[54163] = -2147237452;
assign addr[54164] = -2146862854;
assign addr[54165] = -2146318022;
assign addr[54166] = -2145603001;
assign addr[54167] = -2144717846;
assign addr[54168] = -2143662628;
assign addr[54169] = -2142437431;
assign addr[54170] = -2141042352;
assign addr[54171] = -2139477502;
assign addr[54172] = -2137743003;
assign addr[54173] = -2135838995;
assign addr[54174] = -2133765628;
assign addr[54175] = -2131523066;
assign addr[54176] = -2129111488;
assign addr[54177] = -2126531084;
assign addr[54178] = -2123782059;
assign addr[54179] = -2120864631;
assign addr[54180] = -2117779031;
assign addr[54181] = -2114525505;
assign addr[54182] = -2111104309;
assign addr[54183] = -2107515716;
assign addr[54184] = -2103760010;
assign addr[54185] = -2099837489;
assign addr[54186] = -2095748463;
assign addr[54187] = -2091493257;
assign addr[54188] = -2087072209;
assign addr[54189] = -2082485668;
assign addr[54190] = -2077733999;
assign addr[54191] = -2072817579;
assign addr[54192] = -2067736796;
assign addr[54193] = -2062492055;
assign addr[54194] = -2057083771;
assign addr[54195] = -2051512372;
assign addr[54196] = -2045778302;
assign addr[54197] = -2039882013;
assign addr[54198] = -2033823974;
assign addr[54199] = -2027604666;
assign addr[54200] = -2021224581;
assign addr[54201] = -2014684225;
assign addr[54202] = -2007984117;
assign addr[54203] = -2001124788;
assign addr[54204] = -1994106782;
assign addr[54205] = -1986930656;
assign addr[54206] = -1979596978;
assign addr[54207] = -1972106330;
assign addr[54208] = -1964459306;
assign addr[54209] = -1956656513;
assign addr[54210] = -1948698568;
assign addr[54211] = -1940586104;
assign addr[54212] = -1932319763;
assign addr[54213] = -1923900201;
assign addr[54214] = -1915328086;
assign addr[54215] = -1906604097;
assign addr[54216] = -1897728925;
assign addr[54217] = -1888703276;
assign addr[54218] = -1879527863;
assign addr[54219] = -1870203416;
assign addr[54220] = -1860730673;
assign addr[54221] = -1851110385;
assign addr[54222] = -1841343316;
assign addr[54223] = -1831430239;
assign addr[54224] = -1821371941;
assign addr[54225] = -1811169220;
assign addr[54226] = -1800822883;
assign addr[54227] = -1790333753;
assign addr[54228] = -1779702660;
assign addr[54229] = -1768930447;
assign addr[54230] = -1758017969;
assign addr[54231] = -1746966091;
assign addr[54232] = -1735775690;
assign addr[54233] = -1724447652;
assign addr[54234] = -1712982875;
assign addr[54235] = -1701382270;
assign addr[54236] = -1689646755;
assign addr[54237] = -1677777262;
assign addr[54238] = -1665774731;
assign addr[54239] = -1653640115;
assign addr[54240] = -1641374375;
assign addr[54241] = -1628978484;
assign addr[54242] = -1616453425;
assign addr[54243] = -1603800191;
assign addr[54244] = -1591019785;
assign addr[54245] = -1578113222;
assign addr[54246] = -1565081523;
assign addr[54247] = -1551925723;
assign addr[54248] = -1538646865;
assign addr[54249] = -1525246002;
assign addr[54250] = -1511724196;
assign addr[54251] = -1498082520;
assign addr[54252] = -1484322054;
assign addr[54253] = -1470443891;
assign addr[54254] = -1456449131;
assign addr[54255] = -1442338884;
assign addr[54256] = -1428114267;
assign addr[54257] = -1413776410;
assign addr[54258] = -1399326449;
assign addr[54259] = -1384765530;
assign addr[54260] = -1370094808;
assign addr[54261] = -1355315445;
assign addr[54262] = -1340428615;
assign addr[54263] = -1325435496;
assign addr[54264] = -1310337279;
assign addr[54265] = -1295135159;
assign addr[54266] = -1279830344;
assign addr[54267] = -1264424045;
assign addr[54268] = -1248917486;
assign addr[54269] = -1233311895;
assign addr[54270] = -1217608510;
assign addr[54271] = -1201808576;
assign addr[54272] = -1185913346;
assign addr[54273] = -1169924081;
assign addr[54274] = -1153842047;
assign addr[54275] = -1137668521;
assign addr[54276] = -1121404785;
assign addr[54277] = -1105052128;
assign addr[54278] = -1088611847;
assign addr[54279] = -1072085246;
assign addr[54280] = -1055473635;
assign addr[54281] = -1038778332;
assign addr[54282] = -1022000660;
assign addr[54283] = -1005141949;
assign addr[54284] = -988203537;
assign addr[54285] = -971186766;
assign addr[54286] = -954092986;
assign addr[54287] = -936923553;
assign addr[54288] = -919679827;
assign addr[54289] = -902363176;
assign addr[54290] = -884974973;
assign addr[54291] = -867516597;
assign addr[54292] = -849989433;
assign addr[54293] = -832394869;
assign addr[54294] = -814734301;
assign addr[54295] = -797009130;
assign addr[54296] = -779220762;
assign addr[54297] = -761370605;
assign addr[54298] = -743460077;
assign addr[54299] = -725490597;
assign addr[54300] = -707463589;
assign addr[54301] = -689380485;
assign addr[54302] = -671242716;
assign addr[54303] = -653051723;
assign addr[54304] = -634808946;
assign addr[54305] = -616515832;
assign addr[54306] = -598173833;
assign addr[54307] = -579784402;
assign addr[54308] = -561348998;
assign addr[54309] = -542869083;
assign addr[54310] = -524346121;
assign addr[54311] = -505781581;
assign addr[54312] = -487176937;
assign addr[54313] = -468533662;
assign addr[54314] = -449853235;
assign addr[54315] = -431137138;
assign addr[54316] = -412386854;
assign addr[54317] = -393603870;
assign addr[54318] = -374789676;
assign addr[54319] = -355945764;
assign addr[54320] = -337073627;
assign addr[54321] = -318174762;
assign addr[54322] = -299250668;
assign addr[54323] = -280302845;
assign addr[54324] = -261332796;
assign addr[54325] = -242342025;
assign addr[54326] = -223332037;
assign addr[54327] = -204304341;
assign addr[54328] = -185260444;
assign addr[54329] = -166201858;
assign addr[54330] = -147130093;
assign addr[54331] = -128046661;
assign addr[54332] = -108953076;
assign addr[54333] = -89850852;
assign addr[54334] = -70741503;
assign addr[54335] = -51626544;
assign addr[54336] = -32507492;
assign addr[54337] = -13385863;
assign addr[54338] = 5736829;
assign addr[54339] = 24859065;
assign addr[54340] = 43979330;
assign addr[54341] = 63096108;
assign addr[54342] = 82207882;
assign addr[54343] = 101313138;
assign addr[54344] = 120410361;
assign addr[54345] = 139498035;
assign addr[54346] = 158574649;
assign addr[54347] = 177638688;
assign addr[54348] = 196688642;
assign addr[54349] = 215722999;
assign addr[54350] = 234740251;
assign addr[54351] = 253738890;
assign addr[54352] = 272717408;
assign addr[54353] = 291674302;
assign addr[54354] = 310608068;
assign addr[54355] = 329517204;
assign addr[54356] = 348400212;
assign addr[54357] = 367255594;
assign addr[54358] = 386081854;
assign addr[54359] = 404877501;
assign addr[54360] = 423641043;
assign addr[54361] = 442370993;
assign addr[54362] = 461065866;
assign addr[54363] = 479724180;
assign addr[54364] = 498344454;
assign addr[54365] = 516925212;
assign addr[54366] = 535464981;
assign addr[54367] = 553962291;
assign addr[54368] = 572415676;
assign addr[54369] = 590823671;
assign addr[54370] = 609184818;
assign addr[54371] = 627497660;
assign addr[54372] = 645760745;
assign addr[54373] = 663972625;
assign addr[54374] = 682131857;
assign addr[54375] = 700236999;
assign addr[54376] = 718286617;
assign addr[54377] = 736279279;
assign addr[54378] = 754213559;
assign addr[54379] = 772088034;
assign addr[54380] = 789901288;
assign addr[54381] = 807651907;
assign addr[54382] = 825338484;
assign addr[54383] = 842959617;
assign addr[54384] = 860513908;
assign addr[54385] = 877999966;
assign addr[54386] = 895416404;
assign addr[54387] = 912761841;
assign addr[54388] = 930034901;
assign addr[54389] = 947234215;
assign addr[54390] = 964358420;
assign addr[54391] = 981406156;
assign addr[54392] = 998376073;
assign addr[54393] = 1015266825;
assign addr[54394] = 1032077073;
assign addr[54395] = 1048805483;
assign addr[54396] = 1065450729;
assign addr[54397] = 1082011492;
assign addr[54398] = 1098486458;
assign addr[54399] = 1114874320;
assign addr[54400] = 1131173780;
assign addr[54401] = 1147383544;
assign addr[54402] = 1163502328;
assign addr[54403] = 1179528853;
assign addr[54404] = 1195461849;
assign addr[54405] = 1211300053;
assign addr[54406] = 1227042207;
assign addr[54407] = 1242687064;
assign addr[54408] = 1258233384;
assign addr[54409] = 1273679934;
assign addr[54410] = 1289025489;
assign addr[54411] = 1304268832;
assign addr[54412] = 1319408754;
assign addr[54413] = 1334444055;
assign addr[54414] = 1349373543;
assign addr[54415] = 1364196034;
assign addr[54416] = 1378910353;
assign addr[54417] = 1393515332;
assign addr[54418] = 1408009814;
assign addr[54419] = 1422392650;
assign addr[54420] = 1436662698;
assign addr[54421] = 1450818828;
assign addr[54422] = 1464859917;
assign addr[54423] = 1478784851;
assign addr[54424] = 1492592527;
assign addr[54425] = 1506281850;
assign addr[54426] = 1519851733;
assign addr[54427] = 1533301101;
assign addr[54428] = 1546628888;
assign addr[54429] = 1559834037;
assign addr[54430] = 1572915501;
assign addr[54431] = 1585872242;
assign addr[54432] = 1598703233;
assign addr[54433] = 1611407456;
assign addr[54434] = 1623983905;
assign addr[54435] = 1636431582;
assign addr[54436] = 1648749499;
assign addr[54437] = 1660936681;
assign addr[54438] = 1672992161;
assign addr[54439] = 1684914983;
assign addr[54440] = 1696704201;
assign addr[54441] = 1708358881;
assign addr[54442] = 1719878099;
assign addr[54443] = 1731260941;
assign addr[54444] = 1742506504;
assign addr[54445] = 1753613897;
assign addr[54446] = 1764582240;
assign addr[54447] = 1775410662;
assign addr[54448] = 1786098304;
assign addr[54449] = 1796644320;
assign addr[54450] = 1807047873;
assign addr[54451] = 1817308138;
assign addr[54452] = 1827424302;
assign addr[54453] = 1837395562;
assign addr[54454] = 1847221128;
assign addr[54455] = 1856900221;
assign addr[54456] = 1866432072;
assign addr[54457] = 1875815927;
assign addr[54458] = 1885051042;
assign addr[54459] = 1894136683;
assign addr[54460] = 1903072131;
assign addr[54461] = 1911856677;
assign addr[54462] = 1920489624;
assign addr[54463] = 1928970288;
assign addr[54464] = 1937297997;
assign addr[54465] = 1945472089;
assign addr[54466] = 1953491918;
assign addr[54467] = 1961356847;
assign addr[54468] = 1969066252;
assign addr[54469] = 1976619522;
assign addr[54470] = 1984016058;
assign addr[54471] = 1991255274;
assign addr[54472] = 1998336596;
assign addr[54473] = 2005259462;
assign addr[54474] = 2012023322;
assign addr[54475] = 2018627642;
assign addr[54476] = 2025071897;
assign addr[54477] = 2031355576;
assign addr[54478] = 2037478181;
assign addr[54479] = 2043439226;
assign addr[54480] = 2049238240;
assign addr[54481] = 2054874761;
assign addr[54482] = 2060348343;
assign addr[54483] = 2065658552;
assign addr[54484] = 2070804967;
assign addr[54485] = 2075787180;
assign addr[54486] = 2080604795;
assign addr[54487] = 2085257431;
assign addr[54488] = 2089744719;
assign addr[54489] = 2094066304;
assign addr[54490] = 2098221841;
assign addr[54491] = 2102211002;
assign addr[54492] = 2106033471;
assign addr[54493] = 2109688944;
assign addr[54494] = 2113177132;
assign addr[54495] = 2116497758;
assign addr[54496] = 2119650558;
assign addr[54497] = 2122635283;
assign addr[54498] = 2125451696;
assign addr[54499] = 2128099574;
assign addr[54500] = 2130578706;
assign addr[54501] = 2132888897;
assign addr[54502] = 2135029962;
assign addr[54503] = 2137001733;
assign addr[54504] = 2138804053;
assign addr[54505] = 2140436778;
assign addr[54506] = 2141899780;
assign addr[54507] = 2143192942;
assign addr[54508] = 2144316162;
assign addr[54509] = 2145269351;
assign addr[54510] = 2146052433;
assign addr[54511] = 2146665347;
assign addr[54512] = 2147108043;
assign addr[54513] = 2147380486;
assign addr[54514] = 2147482655;
assign addr[54515] = 2147414542;
assign addr[54516] = 2147176152;
assign addr[54517] = 2146767505;
assign addr[54518] = 2146188631;
assign addr[54519] = 2145439578;
assign addr[54520] = 2144520405;
assign addr[54521] = 2143431184;
assign addr[54522] = 2142172003;
assign addr[54523] = 2140742960;
assign addr[54524] = 2139144169;
assign addr[54525] = 2137375758;
assign addr[54526] = 2135437865;
assign addr[54527] = 2133330646;
assign addr[54528] = 2131054266;
assign addr[54529] = 2128608907;
assign addr[54530] = 2125994762;
assign addr[54531] = 2123212038;
assign addr[54532] = 2120260957;
assign addr[54533] = 2117141752;
assign addr[54534] = 2113854671;
assign addr[54535] = 2110399974;
assign addr[54536] = 2106777935;
assign addr[54537] = 2102988841;
assign addr[54538] = 2099032994;
assign addr[54539] = 2094910706;
assign addr[54540] = 2090622304;
assign addr[54541] = 2086168128;
assign addr[54542] = 2081548533;
assign addr[54543] = 2076763883;
assign addr[54544] = 2071814558;
assign addr[54545] = 2066700952;
assign addr[54546] = 2061423468;
assign addr[54547] = 2055982526;
assign addr[54548] = 2050378558;
assign addr[54549] = 2044612007;
assign addr[54550] = 2038683330;
assign addr[54551] = 2032592999;
assign addr[54552] = 2026341495;
assign addr[54553] = 2019929315;
assign addr[54554] = 2013356967;
assign addr[54555] = 2006624971;
assign addr[54556] = 1999733863;
assign addr[54557] = 1992684188;
assign addr[54558] = 1985476506;
assign addr[54559] = 1978111387;
assign addr[54560] = 1970589416;
assign addr[54561] = 1962911189;
assign addr[54562] = 1955077316;
assign addr[54563] = 1947088417;
assign addr[54564] = 1938945125;
assign addr[54565] = 1930648088;
assign addr[54566] = 1922197961;
assign addr[54567] = 1913595416;
assign addr[54568] = 1904841135;
assign addr[54569] = 1895935811;
assign addr[54570] = 1886880151;
assign addr[54571] = 1877674873;
assign addr[54572] = 1868320707;
assign addr[54573] = 1858818395;
assign addr[54574] = 1849168689;
assign addr[54575] = 1839372356;
assign addr[54576] = 1829430172;
assign addr[54577] = 1819342925;
assign addr[54578] = 1809111415;
assign addr[54579] = 1798736454;
assign addr[54580] = 1788218865;
assign addr[54581] = 1777559480;
assign addr[54582] = 1766759146;
assign addr[54583] = 1755818718;
assign addr[54584] = 1744739065;
assign addr[54585] = 1733521064;
assign addr[54586] = 1722165606;
assign addr[54587] = 1710673591;
assign addr[54588] = 1699045930;
assign addr[54589] = 1687283545;
assign addr[54590] = 1675387369;
assign addr[54591] = 1663358344;
assign addr[54592] = 1651197426;
assign addr[54593] = 1638905577;
assign addr[54594] = 1626483774;
assign addr[54595] = 1613933000;
assign addr[54596] = 1601254251;
assign addr[54597] = 1588448533;
assign addr[54598] = 1575516860;
assign addr[54599] = 1562460258;
assign addr[54600] = 1549279763;
assign addr[54601] = 1535976419;
assign addr[54602] = 1522551282;
assign addr[54603] = 1509005416;
assign addr[54604] = 1495339895;
assign addr[54605] = 1481555802;
assign addr[54606] = 1467654232;
assign addr[54607] = 1453636285;
assign addr[54608] = 1439503074;
assign addr[54609] = 1425255719;
assign addr[54610] = 1410895350;
assign addr[54611] = 1396423105;
assign addr[54612] = 1381840133;
assign addr[54613] = 1367147589;
assign addr[54614] = 1352346639;
assign addr[54615] = 1337438456;
assign addr[54616] = 1322424222;
assign addr[54617] = 1307305128;
assign addr[54618] = 1292082373;
assign addr[54619] = 1276757164;
assign addr[54620] = 1261330715;
assign addr[54621] = 1245804251;
assign addr[54622] = 1230179002;
assign addr[54623] = 1214456207;
assign addr[54624] = 1198637114;
assign addr[54625] = 1182722976;
assign addr[54626] = 1166715055;
assign addr[54627] = 1150614620;
assign addr[54628] = 1134422949;
assign addr[54629] = 1118141326;
assign addr[54630] = 1101771040;
assign addr[54631] = 1085313391;
assign addr[54632] = 1068769683;
assign addr[54633] = 1052141228;
assign addr[54634] = 1035429345;
assign addr[54635] = 1018635358;
assign addr[54636] = 1001760600;
assign addr[54637] = 984806408;
assign addr[54638] = 967774128;
assign addr[54639] = 950665109;
assign addr[54640] = 933480707;
assign addr[54641] = 916222287;
assign addr[54642] = 898891215;
assign addr[54643] = 881488868;
assign addr[54644] = 864016623;
assign addr[54645] = 846475867;
assign addr[54646] = 828867991;
assign addr[54647] = 811194391;
assign addr[54648] = 793456467;
assign addr[54649] = 775655628;
assign addr[54650] = 757793284;
assign addr[54651] = 739870851;
assign addr[54652] = 721889752;
assign addr[54653] = 703851410;
assign addr[54654] = 685757258;
assign addr[54655] = 667608730;
assign addr[54656] = 649407264;
assign addr[54657] = 631154304;
assign addr[54658] = 612851297;
assign addr[54659] = 594499695;
assign addr[54660] = 576100953;
assign addr[54661] = 557656529;
assign addr[54662] = 539167887;
assign addr[54663] = 520636492;
assign addr[54664] = 502063814;
assign addr[54665] = 483451325;
assign addr[54666] = 464800501;
assign addr[54667] = 446112822;
assign addr[54668] = 427389768;
assign addr[54669] = 408632825;
assign addr[54670] = 389843480;
assign addr[54671] = 371023223;
assign addr[54672] = 352173546;
assign addr[54673] = 333295944;
assign addr[54674] = 314391913;
assign addr[54675] = 295462954;
assign addr[54676] = 276510565;
assign addr[54677] = 257536251;
assign addr[54678] = 238541516;
assign addr[54679] = 219527866;
assign addr[54680] = 200496809;
assign addr[54681] = 181449854;
assign addr[54682] = 162388511;
assign addr[54683] = 143314291;
assign addr[54684] = 124228708;
assign addr[54685] = 105133274;
assign addr[54686] = 86029503;
assign addr[54687] = 66918911;
assign addr[54688] = 47803013;
assign addr[54689] = 28683324;
assign addr[54690] = 9561361;
assign addr[54691] = -9561361;
assign addr[54692] = -28683324;
assign addr[54693] = -47803013;
assign addr[54694] = -66918911;
assign addr[54695] = -86029503;
assign addr[54696] = -105133274;
assign addr[54697] = -124228708;
assign addr[54698] = -143314291;
assign addr[54699] = -162388511;
assign addr[54700] = -181449854;
assign addr[54701] = -200496809;
assign addr[54702] = -219527866;
assign addr[54703] = -238541516;
assign addr[54704] = -257536251;
assign addr[54705] = -276510565;
assign addr[54706] = -295462953;
assign addr[54707] = -314391913;
assign addr[54708] = -333295944;
assign addr[54709] = -352173546;
assign addr[54710] = -371023223;
assign addr[54711] = -389843480;
assign addr[54712] = -408632825;
assign addr[54713] = -427389768;
assign addr[54714] = -446112822;
assign addr[54715] = -464800501;
assign addr[54716] = -483451325;
assign addr[54717] = -502063814;
assign addr[54718] = -520636492;
assign addr[54719] = -539167887;
assign addr[54720] = -557656529;
assign addr[54721] = -576100953;
assign addr[54722] = -594499695;
assign addr[54723] = -612851297;
assign addr[54724] = -631154304;
assign addr[54725] = -649407264;
assign addr[54726] = -667608730;
assign addr[54727] = -685757258;
assign addr[54728] = -703851410;
assign addr[54729] = -721889752;
assign addr[54730] = -739870851;
assign addr[54731] = -757793284;
assign addr[54732] = -775655628;
assign addr[54733] = -793456467;
assign addr[54734] = -811194391;
assign addr[54735] = -828867991;
assign addr[54736] = -846475867;
assign addr[54737] = -864016623;
assign addr[54738] = -881488868;
assign addr[54739] = -898891215;
assign addr[54740] = -916222287;
assign addr[54741] = -933480707;
assign addr[54742] = -950665109;
assign addr[54743] = -967774128;
assign addr[54744] = -984806408;
assign addr[54745] = -1001760600;
assign addr[54746] = -1018635358;
assign addr[54747] = -1035429345;
assign addr[54748] = -1052141228;
assign addr[54749] = -1068769683;
assign addr[54750] = -1085313391;
assign addr[54751] = -1101771040;
assign addr[54752] = -1118141326;
assign addr[54753] = -1134422949;
assign addr[54754] = -1150614620;
assign addr[54755] = -1166715055;
assign addr[54756] = -1182722976;
assign addr[54757] = -1198637114;
assign addr[54758] = -1214456207;
assign addr[54759] = -1230179002;
assign addr[54760] = -1245804251;
assign addr[54761] = -1261330715;
assign addr[54762] = -1276757164;
assign addr[54763] = -1292082373;
assign addr[54764] = -1307305128;
assign addr[54765] = -1322424222;
assign addr[54766] = -1337438456;
assign addr[54767] = -1352346639;
assign addr[54768] = -1367147589;
assign addr[54769] = -1381840133;
assign addr[54770] = -1396423105;
assign addr[54771] = -1410895350;
assign addr[54772] = -1425255719;
assign addr[54773] = -1439503074;
assign addr[54774] = -1453636285;
assign addr[54775] = -1467654232;
assign addr[54776] = -1481555802;
assign addr[54777] = -1495339895;
assign addr[54778] = -1509005416;
assign addr[54779] = -1522551282;
assign addr[54780] = -1535976419;
assign addr[54781] = -1549279763;
assign addr[54782] = -1562460258;
assign addr[54783] = -1575516860;
assign addr[54784] = -1588448533;
assign addr[54785] = -1601254251;
assign addr[54786] = -1613933000;
assign addr[54787] = -1626483774;
assign addr[54788] = -1638905577;
assign addr[54789] = -1651197426;
assign addr[54790] = -1663358344;
assign addr[54791] = -1675387369;
assign addr[54792] = -1687283545;
assign addr[54793] = -1699045930;
assign addr[54794] = -1710673591;
assign addr[54795] = -1722165606;
assign addr[54796] = -1733521064;
assign addr[54797] = -1744739065;
assign addr[54798] = -1755818718;
assign addr[54799] = -1766759146;
assign addr[54800] = -1777559480;
assign addr[54801] = -1788218865;
assign addr[54802] = -1798736454;
assign addr[54803] = -1809111415;
assign addr[54804] = -1819342925;
assign addr[54805] = -1829430172;
assign addr[54806] = -1839372356;
assign addr[54807] = -1849168689;
assign addr[54808] = -1858818395;
assign addr[54809] = -1868320707;
assign addr[54810] = -1877674873;
assign addr[54811] = -1886880151;
assign addr[54812] = -1895935811;
assign addr[54813] = -1904841135;
assign addr[54814] = -1913595416;
assign addr[54815] = -1922197961;
assign addr[54816] = -1930648088;
assign addr[54817] = -1938945125;
assign addr[54818] = -1947088417;
assign addr[54819] = -1955077316;
assign addr[54820] = -1962911189;
assign addr[54821] = -1970589416;
assign addr[54822] = -1978111387;
assign addr[54823] = -1985476506;
assign addr[54824] = -1992684188;
assign addr[54825] = -1999733863;
assign addr[54826] = -2006624971;
assign addr[54827] = -2013356967;
assign addr[54828] = -2019929315;
assign addr[54829] = -2026341495;
assign addr[54830] = -2032592999;
assign addr[54831] = -2038683330;
assign addr[54832] = -2044612007;
assign addr[54833] = -2050378558;
assign addr[54834] = -2055982526;
assign addr[54835] = -2061423468;
assign addr[54836] = -2066700952;
assign addr[54837] = -2071814558;
assign addr[54838] = -2076763883;
assign addr[54839] = -2081548533;
assign addr[54840] = -2086168128;
assign addr[54841] = -2090622304;
assign addr[54842] = -2094910706;
assign addr[54843] = -2099032994;
assign addr[54844] = -2102988841;
assign addr[54845] = -2106777935;
assign addr[54846] = -2110399974;
assign addr[54847] = -2113854671;
assign addr[54848] = -2117141752;
assign addr[54849] = -2120260957;
assign addr[54850] = -2123212038;
assign addr[54851] = -2125994762;
assign addr[54852] = -2128608907;
assign addr[54853] = -2131054266;
assign addr[54854] = -2133330646;
assign addr[54855] = -2135437865;
assign addr[54856] = -2137375758;
assign addr[54857] = -2139144169;
assign addr[54858] = -2140742960;
assign addr[54859] = -2142172003;
assign addr[54860] = -2143431184;
assign addr[54861] = -2144520405;
assign addr[54862] = -2145439578;
assign addr[54863] = -2146188631;
assign addr[54864] = -2146767505;
assign addr[54865] = -2147176152;
assign addr[54866] = -2147414542;
assign addr[54867] = -2147482655;
assign addr[54868] = -2147380486;
assign addr[54869] = -2147108043;
assign addr[54870] = -2146665347;
assign addr[54871] = -2146052433;
assign addr[54872] = -2145269351;
assign addr[54873] = -2144316162;
assign addr[54874] = -2143192942;
assign addr[54875] = -2141899780;
assign addr[54876] = -2140436778;
assign addr[54877] = -2138804053;
assign addr[54878] = -2137001733;
assign addr[54879] = -2135029962;
assign addr[54880] = -2132888897;
assign addr[54881] = -2130578706;
assign addr[54882] = -2128099574;
assign addr[54883] = -2125451696;
assign addr[54884] = -2122635283;
assign addr[54885] = -2119650558;
assign addr[54886] = -2116497758;
assign addr[54887] = -2113177132;
assign addr[54888] = -2109688944;
assign addr[54889] = -2106033471;
assign addr[54890] = -2102211002;
assign addr[54891] = -2098221841;
assign addr[54892] = -2094066304;
assign addr[54893] = -2089744719;
assign addr[54894] = -2085257431;
assign addr[54895] = -2080604795;
assign addr[54896] = -2075787180;
assign addr[54897] = -2070804967;
assign addr[54898] = -2065658552;
assign addr[54899] = -2060348343;
assign addr[54900] = -2054874761;
assign addr[54901] = -2049238240;
assign addr[54902] = -2043439226;
assign addr[54903] = -2037478181;
assign addr[54904] = -2031355576;
assign addr[54905] = -2025071897;
assign addr[54906] = -2018627642;
assign addr[54907] = -2012023322;
assign addr[54908] = -2005259462;
assign addr[54909] = -1998336596;
assign addr[54910] = -1991255274;
assign addr[54911] = -1984016058;
assign addr[54912] = -1976619522;
assign addr[54913] = -1969066252;
assign addr[54914] = -1961356847;
assign addr[54915] = -1953491918;
assign addr[54916] = -1945472089;
assign addr[54917] = -1937297997;
assign addr[54918] = -1928970288;
assign addr[54919] = -1920489624;
assign addr[54920] = -1911856677;
assign addr[54921] = -1903072131;
assign addr[54922] = -1894136683;
assign addr[54923] = -1885051042;
assign addr[54924] = -1875815927;
assign addr[54925] = -1866432072;
assign addr[54926] = -1856900221;
assign addr[54927] = -1847221128;
assign addr[54928] = -1837395562;
assign addr[54929] = -1827424302;
assign addr[54930] = -1817308138;
assign addr[54931] = -1807047873;
assign addr[54932] = -1796644320;
assign addr[54933] = -1786098304;
assign addr[54934] = -1775410662;
assign addr[54935] = -1764582240;
assign addr[54936] = -1753613897;
assign addr[54937] = -1742506504;
assign addr[54938] = -1731260941;
assign addr[54939] = -1719878099;
assign addr[54940] = -1708358881;
assign addr[54941] = -1696704201;
assign addr[54942] = -1684914983;
assign addr[54943] = -1672992161;
assign addr[54944] = -1660936681;
assign addr[54945] = -1648749499;
assign addr[54946] = -1636431582;
assign addr[54947] = -1623983905;
assign addr[54948] = -1611407456;
assign addr[54949] = -1598703233;
assign addr[54950] = -1585872242;
assign addr[54951] = -1572915501;
assign addr[54952] = -1559834037;
assign addr[54953] = -1546628888;
assign addr[54954] = -1533301101;
assign addr[54955] = -1519851733;
assign addr[54956] = -1506281850;
assign addr[54957] = -1492592527;
assign addr[54958] = -1478784851;
assign addr[54959] = -1464859917;
assign addr[54960] = -1450818828;
assign addr[54961] = -1436662698;
assign addr[54962] = -1422392650;
assign addr[54963] = -1408009814;
assign addr[54964] = -1393515332;
assign addr[54965] = -1378910353;
assign addr[54966] = -1364196034;
assign addr[54967] = -1349373543;
assign addr[54968] = -1334444055;
assign addr[54969] = -1319408754;
assign addr[54970] = -1304268832;
assign addr[54971] = -1289025489;
assign addr[54972] = -1273679934;
assign addr[54973] = -1258233384;
assign addr[54974] = -1242687064;
assign addr[54975] = -1227042207;
assign addr[54976] = -1211300053;
assign addr[54977] = -1195461849;
assign addr[54978] = -1179528853;
assign addr[54979] = -1163502328;
assign addr[54980] = -1147383544;
assign addr[54981] = -1131173780;
assign addr[54982] = -1114874320;
assign addr[54983] = -1098486458;
assign addr[54984] = -1082011492;
assign addr[54985] = -1065450729;
assign addr[54986] = -1048805483;
assign addr[54987] = -1032077073;
assign addr[54988] = -1015266825;
assign addr[54989] = -998376073;
assign addr[54990] = -981406156;
assign addr[54991] = -964358420;
assign addr[54992] = -947234215;
assign addr[54993] = -930034901;
assign addr[54994] = -912761841;
assign addr[54995] = -895416404;
assign addr[54996] = -877999966;
assign addr[54997] = -860513908;
assign addr[54998] = -842959617;
assign addr[54999] = -825338484;
assign addr[55000] = -807651907;
assign addr[55001] = -789901288;
assign addr[55002] = -772088034;
assign addr[55003] = -754213559;
assign addr[55004] = -736279279;
assign addr[55005] = -718286617;
assign addr[55006] = -700236999;
assign addr[55007] = -682131857;
assign addr[55008] = -663972625;
assign addr[55009] = -645760745;
assign addr[55010] = -627497660;
assign addr[55011] = -609184818;
assign addr[55012] = -590823671;
assign addr[55013] = -572415676;
assign addr[55014] = -553962291;
assign addr[55015] = -535464981;
assign addr[55016] = -516925212;
assign addr[55017] = -498344454;
assign addr[55018] = -479724180;
assign addr[55019] = -461065866;
assign addr[55020] = -442370993;
assign addr[55021] = -423641043;
assign addr[55022] = -404877501;
assign addr[55023] = -386081854;
assign addr[55024] = -367255594;
assign addr[55025] = -348400212;
assign addr[55026] = -329517204;
assign addr[55027] = -310608068;
assign addr[55028] = -291674302;
assign addr[55029] = -272717408;
assign addr[55030] = -253738890;
assign addr[55031] = -234740251;
assign addr[55032] = -215722999;
assign addr[55033] = -196688642;
assign addr[55034] = -177638688;
assign addr[55035] = -158574649;
assign addr[55036] = -139498035;
assign addr[55037] = -120410361;
assign addr[55038] = -101313138;
assign addr[55039] = -82207882;
assign addr[55040] = -63096108;
assign addr[55041] = -43979330;
assign addr[55042] = -24859065;
assign addr[55043] = -5736829;
assign addr[55044] = 13385863;
assign addr[55045] = 32507492;
assign addr[55046] = 51626544;
assign addr[55047] = 70741503;
assign addr[55048] = 89850852;
assign addr[55049] = 108953076;
assign addr[55050] = 128046661;
assign addr[55051] = 147130093;
assign addr[55052] = 166201858;
assign addr[55053] = 185260444;
assign addr[55054] = 204304341;
assign addr[55055] = 223332037;
assign addr[55056] = 242342025;
assign addr[55057] = 261332796;
assign addr[55058] = 280302845;
assign addr[55059] = 299250668;
assign addr[55060] = 318174762;
assign addr[55061] = 337073627;
assign addr[55062] = 355945764;
assign addr[55063] = 374789676;
assign addr[55064] = 393603870;
assign addr[55065] = 412386854;
assign addr[55066] = 431137138;
assign addr[55067] = 449853235;
assign addr[55068] = 468533662;
assign addr[55069] = 487176937;
assign addr[55070] = 505781581;
assign addr[55071] = 524346121;
assign addr[55072] = 542869083;
assign addr[55073] = 561348998;
assign addr[55074] = 579784402;
assign addr[55075] = 598173833;
assign addr[55076] = 616515832;
assign addr[55077] = 634808946;
assign addr[55078] = 653051723;
assign addr[55079] = 671242716;
assign addr[55080] = 689380485;
assign addr[55081] = 707463589;
assign addr[55082] = 725490597;
assign addr[55083] = 743460077;
assign addr[55084] = 761370605;
assign addr[55085] = 779220762;
assign addr[55086] = 797009130;
assign addr[55087] = 814734301;
assign addr[55088] = 832394869;
assign addr[55089] = 849989433;
assign addr[55090] = 867516597;
assign addr[55091] = 884974973;
assign addr[55092] = 902363176;
assign addr[55093] = 919679827;
assign addr[55094] = 936923553;
assign addr[55095] = 954092986;
assign addr[55096] = 971186766;
assign addr[55097] = 988203537;
assign addr[55098] = 1005141949;
assign addr[55099] = 1022000660;
assign addr[55100] = 1038778332;
assign addr[55101] = 1055473635;
assign addr[55102] = 1072085246;
assign addr[55103] = 1088611847;
assign addr[55104] = 1105052128;
assign addr[55105] = 1121404785;
assign addr[55106] = 1137668521;
assign addr[55107] = 1153842047;
assign addr[55108] = 1169924081;
assign addr[55109] = 1185913346;
assign addr[55110] = 1201808576;
assign addr[55111] = 1217608510;
assign addr[55112] = 1233311895;
assign addr[55113] = 1248917486;
assign addr[55114] = 1264424045;
assign addr[55115] = 1279830344;
assign addr[55116] = 1295135159;
assign addr[55117] = 1310337279;
assign addr[55118] = 1325435496;
assign addr[55119] = 1340428615;
assign addr[55120] = 1355315445;
assign addr[55121] = 1370094808;
assign addr[55122] = 1384765530;
assign addr[55123] = 1399326449;
assign addr[55124] = 1413776410;
assign addr[55125] = 1428114267;
assign addr[55126] = 1442338884;
assign addr[55127] = 1456449131;
assign addr[55128] = 1470443891;
assign addr[55129] = 1484322054;
assign addr[55130] = 1498082520;
assign addr[55131] = 1511724196;
assign addr[55132] = 1525246002;
assign addr[55133] = 1538646865;
assign addr[55134] = 1551925723;
assign addr[55135] = 1565081523;
assign addr[55136] = 1578113222;
assign addr[55137] = 1591019785;
assign addr[55138] = 1603800191;
assign addr[55139] = 1616453425;
assign addr[55140] = 1628978484;
assign addr[55141] = 1641374375;
assign addr[55142] = 1653640115;
assign addr[55143] = 1665774731;
assign addr[55144] = 1677777262;
assign addr[55145] = 1689646755;
assign addr[55146] = 1701382270;
assign addr[55147] = 1712982875;
assign addr[55148] = 1724447652;
assign addr[55149] = 1735775690;
assign addr[55150] = 1746966091;
assign addr[55151] = 1758017969;
assign addr[55152] = 1768930447;
assign addr[55153] = 1779702660;
assign addr[55154] = 1790333753;
assign addr[55155] = 1800822883;
assign addr[55156] = 1811169220;
assign addr[55157] = 1821371941;
assign addr[55158] = 1831430239;
assign addr[55159] = 1841343316;
assign addr[55160] = 1851110385;
assign addr[55161] = 1860730673;
assign addr[55162] = 1870203416;
assign addr[55163] = 1879527863;
assign addr[55164] = 1888703276;
assign addr[55165] = 1897728925;
assign addr[55166] = 1906604097;
assign addr[55167] = 1915328086;
assign addr[55168] = 1923900201;
assign addr[55169] = 1932319763;
assign addr[55170] = 1940586104;
assign addr[55171] = 1948698568;
assign addr[55172] = 1956656513;
assign addr[55173] = 1964459306;
assign addr[55174] = 1972106330;
assign addr[55175] = 1979596978;
assign addr[55176] = 1986930656;
assign addr[55177] = 1994106782;
assign addr[55178] = 2001124788;
assign addr[55179] = 2007984117;
assign addr[55180] = 2014684225;
assign addr[55181] = 2021224581;
assign addr[55182] = 2027604666;
assign addr[55183] = 2033823974;
assign addr[55184] = 2039882013;
assign addr[55185] = 2045778302;
assign addr[55186] = 2051512372;
assign addr[55187] = 2057083771;
assign addr[55188] = 2062492055;
assign addr[55189] = 2067736796;
assign addr[55190] = 2072817579;
assign addr[55191] = 2077733999;
assign addr[55192] = 2082485668;
assign addr[55193] = 2087072209;
assign addr[55194] = 2091493257;
assign addr[55195] = 2095748463;
assign addr[55196] = 2099837489;
assign addr[55197] = 2103760010;
assign addr[55198] = 2107515716;
assign addr[55199] = 2111104309;
assign addr[55200] = 2114525505;
assign addr[55201] = 2117779031;
assign addr[55202] = 2120864631;
assign addr[55203] = 2123782059;
assign addr[55204] = 2126531084;
assign addr[55205] = 2129111488;
assign addr[55206] = 2131523066;
assign addr[55207] = 2133765628;
assign addr[55208] = 2135838995;
assign addr[55209] = 2137743003;
assign addr[55210] = 2139477502;
assign addr[55211] = 2141042352;
assign addr[55212] = 2142437431;
assign addr[55213] = 2143662628;
assign addr[55214] = 2144717846;
assign addr[55215] = 2145603001;
assign addr[55216] = 2146318022;
assign addr[55217] = 2146862854;
assign addr[55218] = 2147237452;
assign addr[55219] = 2147441787;
assign addr[55220] = 2147475844;
assign addr[55221] = 2147339619;
assign addr[55222] = 2147033123;
assign addr[55223] = 2146556380;
assign addr[55224] = 2145909429;
assign addr[55225] = 2145092320;
assign addr[55226] = 2144105118;
assign addr[55227] = 2142947902;
assign addr[55228] = 2141620763;
assign addr[55229] = 2140123807;
assign addr[55230] = 2138457152;
assign addr[55231] = 2136620930;
assign addr[55232] = 2134615288;
assign addr[55233] = 2132440383;
assign addr[55234] = 2130096389;
assign addr[55235] = 2127583492;
assign addr[55236] = 2124901890;
assign addr[55237] = 2122051796;
assign addr[55238] = 2119033436;
assign addr[55239] = 2115847050;
assign addr[55240] = 2112492891;
assign addr[55241] = 2108971223;
assign addr[55242] = 2105282327;
assign addr[55243] = 2101426496;
assign addr[55244] = 2097404033;
assign addr[55245] = 2093215260;
assign addr[55246] = 2088860507;
assign addr[55247] = 2084340120;
assign addr[55248] = 2079654458;
assign addr[55249] = 2074803892;
assign addr[55250] = 2069788807;
assign addr[55251] = 2064609600;
assign addr[55252] = 2059266683;
assign addr[55253] = 2053760478;
assign addr[55254] = 2048091422;
assign addr[55255] = 2042259965;
assign addr[55256] = 2036266570;
assign addr[55257] = 2030111710;
assign addr[55258] = 2023795876;
assign addr[55259] = 2017319567;
assign addr[55260] = 2010683297;
assign addr[55261] = 2003887591;
assign addr[55262] = 1996932990;
assign addr[55263] = 1989820044;
assign addr[55264] = 1982549318;
assign addr[55265] = 1975121388;
assign addr[55266] = 1967536842;
assign addr[55267] = 1959796283;
assign addr[55268] = 1951900324;
assign addr[55269] = 1943849591;
assign addr[55270] = 1935644723;
assign addr[55271] = 1927286370;
assign addr[55272] = 1918775195;
assign addr[55273] = 1910111873;
assign addr[55274] = 1901297091;
assign addr[55275] = 1892331547;
assign addr[55276] = 1883215953;
assign addr[55277] = 1873951032;
assign addr[55278] = 1864537518;
assign addr[55279] = 1854976157;
assign addr[55280] = 1845267708;
assign addr[55281] = 1835412941;
assign addr[55282] = 1825412636;
assign addr[55283] = 1815267588;
assign addr[55284] = 1804978599;
assign addr[55285] = 1794546487;
assign addr[55286] = 1783972079;
assign addr[55287] = 1773256212;
assign addr[55288] = 1762399737;
assign addr[55289] = 1751403515;
assign addr[55290] = 1740268417;
assign addr[55291] = 1728995326;
assign addr[55292] = 1717585136;
assign addr[55293] = 1706038753;
assign addr[55294] = 1694357091;
assign addr[55295] = 1682541077;
assign addr[55296] = 1670591647;
assign addr[55297] = 1658509750;
assign addr[55298] = 1646296344;
assign addr[55299] = 1633952396;
assign addr[55300] = 1621478885;
assign addr[55301] = 1608876801;
assign addr[55302] = 1596147143;
assign addr[55303] = 1583290921;
assign addr[55304] = 1570309153;
assign addr[55305] = 1557202869;
assign addr[55306] = 1543973108;
assign addr[55307] = 1530620920;
assign addr[55308] = 1517147363;
assign addr[55309] = 1503553506;
assign addr[55310] = 1489840425;
assign addr[55311] = 1476009210;
assign addr[55312] = 1462060956;
assign addr[55313] = 1447996770;
assign addr[55314] = 1433817766;
assign addr[55315] = 1419525069;
assign addr[55316] = 1405119813;
assign addr[55317] = 1390603139;
assign addr[55318] = 1375976199;
assign addr[55319] = 1361240152;
assign addr[55320] = 1346396168;
assign addr[55321] = 1331445422;
assign addr[55322] = 1316389101;
assign addr[55323] = 1301228398;
assign addr[55324] = 1285964516;
assign addr[55325] = 1270598665;
assign addr[55326] = 1255132063;
assign addr[55327] = 1239565936;
assign addr[55328] = 1223901520;
assign addr[55329] = 1208140056;
assign addr[55330] = 1192282793;
assign addr[55331] = 1176330990;
assign addr[55332] = 1160285911;
assign addr[55333] = 1144148829;
assign addr[55334] = 1127921022;
assign addr[55335] = 1111603778;
assign addr[55336] = 1095198391;
assign addr[55337] = 1078706161;
assign addr[55338] = 1062128397;
assign addr[55339] = 1045466412;
assign addr[55340] = 1028721528;
assign addr[55341] = 1011895073;
assign addr[55342] = 994988380;
assign addr[55343] = 978002791;
assign addr[55344] = 960939653;
assign addr[55345] = 943800318;
assign addr[55346] = 926586145;
assign addr[55347] = 909298500;
assign addr[55348] = 891938752;
assign addr[55349] = 874508280;
assign addr[55350] = 857008464;
assign addr[55351] = 839440693;
assign addr[55352] = 821806359;
assign addr[55353] = 804106861;
assign addr[55354] = 786343603;
assign addr[55355] = 768517992;
assign addr[55356] = 750631442;
assign addr[55357] = 732685372;
assign addr[55358] = 714681204;
assign addr[55359] = 696620367;
assign addr[55360] = 678504291;
assign addr[55361] = 660334415;
assign addr[55362] = 642112178;
assign addr[55363] = 623839025;
assign addr[55364] = 605516406;
assign addr[55365] = 587145773;
assign addr[55366] = 568728583;
assign addr[55367] = 550266296;
assign addr[55368] = 531760377;
assign addr[55369] = 513212292;
assign addr[55370] = 494623513;
assign addr[55371] = 475995513;
assign addr[55372] = 457329769;
assign addr[55373] = 438627762;
assign addr[55374] = 419890975;
assign addr[55375] = 401120892;
assign addr[55376] = 382319004;
assign addr[55377] = 363486799;
assign addr[55378] = 344625773;
assign addr[55379] = 325737419;
assign addr[55380] = 306823237;
assign addr[55381] = 287884725;
assign addr[55382] = 268923386;
assign addr[55383] = 249940723;
assign addr[55384] = 230938242;
assign addr[55385] = 211917448;
assign addr[55386] = 192879850;
assign addr[55387] = 173826959;
assign addr[55388] = 154760284;
assign addr[55389] = 135681337;
assign addr[55390] = 116591632;
assign addr[55391] = 97492681;
assign addr[55392] = 78386000;
assign addr[55393] = 59273104;
assign addr[55394] = 40155507;
assign addr[55395] = 21034727;
assign addr[55396] = 1912278;
assign addr[55397] = -17210322;
assign addr[55398] = -36331557;
assign addr[55399] = -55449912;
assign addr[55400] = -74563870;
assign addr[55401] = -93671915;
assign addr[55402] = -112772533;
assign addr[55403] = -131864208;
assign addr[55404] = -150945428;
assign addr[55405] = -170014678;
assign addr[55406] = -189070447;
assign addr[55407] = -208111224;
assign addr[55408] = -227135500;
assign addr[55409] = -246141764;
assign addr[55410] = -265128512;
assign addr[55411] = -284094236;
assign addr[55412] = -303037433;
assign addr[55413] = -321956601;
assign addr[55414] = -340850240;
assign addr[55415] = -359716852;
assign addr[55416] = -378554940;
assign addr[55417] = -397363011;
assign addr[55418] = -416139574;
assign addr[55419] = -434883140;
assign addr[55420] = -453592221;
assign addr[55421] = -472265336;
assign addr[55422] = -490901003;
assign addr[55423] = -509497745;
assign addr[55424] = -528054086;
assign addr[55425] = -546568556;
assign addr[55426] = -565039687;
assign addr[55427] = -583466013;
assign addr[55428] = -601846074;
assign addr[55429] = -620178412;
assign addr[55430] = -638461574;
assign addr[55431] = -656694110;
assign addr[55432] = -674874574;
assign addr[55433] = -693001525;
assign addr[55434] = -711073524;
assign addr[55435] = -729089140;
assign addr[55436] = -747046944;
assign addr[55437] = -764945512;
assign addr[55438] = -782783424;
assign addr[55439] = -800559266;
assign addr[55440] = -818271628;
assign addr[55441] = -835919107;
assign addr[55442] = -853500302;
assign addr[55443] = -871013820;
assign addr[55444] = -888458272;
assign addr[55445] = -905832274;
assign addr[55446] = -923134450;
assign addr[55447] = -940363427;
assign addr[55448] = -957517838;
assign addr[55449] = -974596324;
assign addr[55450] = -991597531;
assign addr[55451] = -1008520110;
assign addr[55452] = -1025362720;
assign addr[55453] = -1042124025;
assign addr[55454] = -1058802695;
assign addr[55455] = -1075397409;
assign addr[55456] = -1091906851;
assign addr[55457] = -1108329711;
assign addr[55458] = -1124664687;
assign addr[55459] = -1140910484;
assign addr[55460] = -1157065814;
assign addr[55461] = -1173129396;
assign addr[55462] = -1189099956;
assign addr[55463] = -1204976227;
assign addr[55464] = -1220756951;
assign addr[55465] = -1236440877;
assign addr[55466] = -1252026760;
assign addr[55467] = -1267513365;
assign addr[55468] = -1282899464;
assign addr[55469] = -1298183838;
assign addr[55470] = -1313365273;
assign addr[55471] = -1328442566;
assign addr[55472] = -1343414522;
assign addr[55473] = -1358279953;
assign addr[55474] = -1373037681;
assign addr[55475] = -1387686535;
assign addr[55476] = -1402225355;
assign addr[55477] = -1416652986;
assign addr[55478] = -1430968286;
assign addr[55479] = -1445170118;
assign addr[55480] = -1459257358;
assign addr[55481] = -1473228887;
assign addr[55482] = -1487083598;
assign addr[55483] = -1500820393;
assign addr[55484] = -1514438181;
assign addr[55485] = -1527935884;
assign addr[55486] = -1541312431;
assign addr[55487] = -1554566762;
assign addr[55488] = -1567697824;
assign addr[55489] = -1580704578;
assign addr[55490] = -1593585992;
assign addr[55491] = -1606341043;
assign addr[55492] = -1618968722;
assign addr[55493] = -1631468027;
assign addr[55494] = -1643837966;
assign addr[55495] = -1656077559;
assign addr[55496] = -1668185835;
assign addr[55497] = -1680161834;
assign addr[55498] = -1692004606;
assign addr[55499] = -1703713213;
assign addr[55500] = -1715286726;
assign addr[55501] = -1726724227;
assign addr[55502] = -1738024810;
assign addr[55503] = -1749187577;
assign addr[55504] = -1760211645;
assign addr[55505] = -1771096139;
assign addr[55506] = -1781840195;
assign addr[55507] = -1792442963;
assign addr[55508] = -1802903601;
assign addr[55509] = -1813221279;
assign addr[55510] = -1823395180;
assign addr[55511] = -1833424497;
assign addr[55512] = -1843308435;
assign addr[55513] = -1853046210;
assign addr[55514] = -1862637049;
assign addr[55515] = -1872080193;
assign addr[55516] = -1881374892;
assign addr[55517] = -1890520410;
assign addr[55518] = -1899516021;
assign addr[55519] = -1908361011;
assign addr[55520] = -1917054681;
assign addr[55521] = -1925596340;
assign addr[55522] = -1933985310;
assign addr[55523] = -1942220928;
assign addr[55524] = -1950302539;
assign addr[55525] = -1958229503;
assign addr[55526] = -1966001192;
assign addr[55527] = -1973616989;
assign addr[55528] = -1981076290;
assign addr[55529] = -1988378503;
assign addr[55530] = -1995523051;
assign addr[55531] = -2002509365;
assign addr[55532] = -2009336893;
assign addr[55533] = -2016005093;
assign addr[55534] = -2022513436;
assign addr[55535] = -2028861406;
assign addr[55536] = -2035048499;
assign addr[55537] = -2041074226;
assign addr[55538] = -2046938108;
assign addr[55539] = -2052639680;
assign addr[55540] = -2058178491;
assign addr[55541] = -2063554100;
assign addr[55542] = -2068766083;
assign addr[55543] = -2073814024;
assign addr[55544] = -2078697525;
assign addr[55545] = -2083416198;
assign addr[55546] = -2087969669;
assign addr[55547] = -2092357577;
assign addr[55548] = -2096579573;
assign addr[55549] = -2100635323;
assign addr[55550] = -2104524506;
assign addr[55551] = -2108246813;
assign addr[55552] = -2111801949;
assign addr[55553] = -2115189632;
assign addr[55554] = -2118409593;
assign addr[55555] = -2121461578;
assign addr[55556] = -2124345343;
assign addr[55557] = -2127060661;
assign addr[55558] = -2129607316;
assign addr[55559] = -2131985106;
assign addr[55560] = -2134193842;
assign addr[55561] = -2136233350;
assign addr[55562] = -2138103468;
assign addr[55563] = -2139804048;
assign addr[55564] = -2141334954;
assign addr[55565] = -2142696065;
assign addr[55566] = -2143887273;
assign addr[55567] = -2144908484;
assign addr[55568] = -2145759618;
assign addr[55569] = -2146440605;
assign addr[55570] = -2146951393;
assign addr[55571] = -2147291941;
assign addr[55572] = -2147462221;
assign addr[55573] = -2147462221;
assign addr[55574] = -2147291941;
assign addr[55575] = -2146951393;
assign addr[55576] = -2146440605;
assign addr[55577] = -2145759618;
assign addr[55578] = -2144908484;
assign addr[55579] = -2143887273;
assign addr[55580] = -2142696065;
assign addr[55581] = -2141334954;
assign addr[55582] = -2139804048;
assign addr[55583] = -2138103468;
assign addr[55584] = -2136233350;
assign addr[55585] = -2134193842;
assign addr[55586] = -2131985106;
assign addr[55587] = -2129607316;
assign addr[55588] = -2127060661;
assign addr[55589] = -2124345343;
assign addr[55590] = -2121461578;
assign addr[55591] = -2118409593;
assign addr[55592] = -2115189632;
assign addr[55593] = -2111801949;
assign addr[55594] = -2108246813;
assign addr[55595] = -2104524506;
assign addr[55596] = -2100635323;
assign addr[55597] = -2096579573;
assign addr[55598] = -2092357577;
assign addr[55599] = -2087969669;
assign addr[55600] = -2083416198;
assign addr[55601] = -2078697525;
assign addr[55602] = -2073814024;
assign addr[55603] = -2068766083;
assign addr[55604] = -2063554100;
assign addr[55605] = -2058178491;
assign addr[55606] = -2052639680;
assign addr[55607] = -2046938108;
assign addr[55608] = -2041074226;
assign addr[55609] = -2035048499;
assign addr[55610] = -2028861406;
assign addr[55611] = -2022513436;
assign addr[55612] = -2016005093;
assign addr[55613] = -2009336893;
assign addr[55614] = -2002509365;
assign addr[55615] = -1995523051;
assign addr[55616] = -1988378503;
assign addr[55617] = -1981076290;
assign addr[55618] = -1973616989;
assign addr[55619] = -1966001192;
assign addr[55620] = -1958229503;
assign addr[55621] = -1950302539;
assign addr[55622] = -1942220928;
assign addr[55623] = -1933985310;
assign addr[55624] = -1925596340;
assign addr[55625] = -1917054681;
assign addr[55626] = -1908361011;
assign addr[55627] = -1899516021;
assign addr[55628] = -1890520410;
assign addr[55629] = -1881374892;
assign addr[55630] = -1872080193;
assign addr[55631] = -1862637049;
assign addr[55632] = -1853046210;
assign addr[55633] = -1843308435;
assign addr[55634] = -1833424497;
assign addr[55635] = -1823395180;
assign addr[55636] = -1813221279;
assign addr[55637] = -1802903601;
assign addr[55638] = -1792442963;
assign addr[55639] = -1781840195;
assign addr[55640] = -1771096139;
assign addr[55641] = -1760211645;
assign addr[55642] = -1749187577;
assign addr[55643] = -1738024810;
assign addr[55644] = -1726724227;
assign addr[55645] = -1715286726;
assign addr[55646] = -1703713213;
assign addr[55647] = -1692004606;
assign addr[55648] = -1680161834;
assign addr[55649] = -1668185835;
assign addr[55650] = -1656077559;
assign addr[55651] = -1643837966;
assign addr[55652] = -1631468027;
assign addr[55653] = -1618968722;
assign addr[55654] = -1606341043;
assign addr[55655] = -1593585992;
assign addr[55656] = -1580704578;
assign addr[55657] = -1567697824;
assign addr[55658] = -1554566762;
assign addr[55659] = -1541312431;
assign addr[55660] = -1527935884;
assign addr[55661] = -1514438181;
assign addr[55662] = -1500820393;
assign addr[55663] = -1487083598;
assign addr[55664] = -1473228887;
assign addr[55665] = -1459257358;
assign addr[55666] = -1445170118;
assign addr[55667] = -1430968286;
assign addr[55668] = -1416652986;
assign addr[55669] = -1402225355;
assign addr[55670] = -1387686535;
assign addr[55671] = -1373037681;
assign addr[55672] = -1358279953;
assign addr[55673] = -1343414522;
assign addr[55674] = -1328442566;
assign addr[55675] = -1313365273;
assign addr[55676] = -1298183838;
assign addr[55677] = -1282899464;
assign addr[55678] = -1267513365;
assign addr[55679] = -1252026760;
assign addr[55680] = -1236440877;
assign addr[55681] = -1220756951;
assign addr[55682] = -1204976227;
assign addr[55683] = -1189099956;
assign addr[55684] = -1173129396;
assign addr[55685] = -1157065814;
assign addr[55686] = -1140910484;
assign addr[55687] = -1124664687;
assign addr[55688] = -1108329711;
assign addr[55689] = -1091906851;
assign addr[55690] = -1075397409;
assign addr[55691] = -1058802695;
assign addr[55692] = -1042124025;
assign addr[55693] = -1025362720;
assign addr[55694] = -1008520110;
assign addr[55695] = -991597531;
assign addr[55696] = -974596324;
assign addr[55697] = -957517838;
assign addr[55698] = -940363427;
assign addr[55699] = -923134450;
assign addr[55700] = -905832274;
assign addr[55701] = -888458272;
assign addr[55702] = -871013820;
assign addr[55703] = -853500302;
assign addr[55704] = -835919107;
assign addr[55705] = -818271628;
assign addr[55706] = -800559266;
assign addr[55707] = -782783424;
assign addr[55708] = -764945512;
assign addr[55709] = -747046944;
assign addr[55710] = -729089140;
assign addr[55711] = -711073525;
assign addr[55712] = -693001525;
assign addr[55713] = -674874574;
assign addr[55714] = -656694110;
assign addr[55715] = -638461574;
assign addr[55716] = -620178412;
assign addr[55717] = -601846074;
assign addr[55718] = -583466013;
assign addr[55719] = -565039687;
assign addr[55720] = -546568556;
assign addr[55721] = -528054086;
assign addr[55722] = -509497745;
assign addr[55723] = -490901003;
assign addr[55724] = -472265336;
assign addr[55725] = -453592221;
assign addr[55726] = -434883140;
assign addr[55727] = -416139574;
assign addr[55728] = -397363011;
assign addr[55729] = -378554940;
assign addr[55730] = -359716852;
assign addr[55731] = -340850240;
assign addr[55732] = -321956601;
assign addr[55733] = -303037433;
assign addr[55734] = -284094236;
assign addr[55735] = -265128512;
assign addr[55736] = -246141764;
assign addr[55737] = -227135500;
assign addr[55738] = -208111224;
assign addr[55739] = -189070447;
assign addr[55740] = -170014678;
assign addr[55741] = -150945428;
assign addr[55742] = -131864208;
assign addr[55743] = -112772533;
assign addr[55744] = -93671915;
assign addr[55745] = -74563870;
assign addr[55746] = -55449912;
assign addr[55747] = -36331557;
assign addr[55748] = -17210322;
assign addr[55749] = 1912278;
assign addr[55750] = 21034727;
assign addr[55751] = 40155507;
assign addr[55752] = 59273104;
assign addr[55753] = 78386000;
assign addr[55754] = 97492681;
assign addr[55755] = 116591632;
assign addr[55756] = 135681337;
assign addr[55757] = 154760284;
assign addr[55758] = 173826959;
assign addr[55759] = 192879850;
assign addr[55760] = 211917448;
assign addr[55761] = 230938242;
assign addr[55762] = 249940723;
assign addr[55763] = 268923386;
assign addr[55764] = 287884725;
assign addr[55765] = 306823237;
assign addr[55766] = 325737419;
assign addr[55767] = 344625773;
assign addr[55768] = 363486799;
assign addr[55769] = 382319004;
assign addr[55770] = 401120892;
assign addr[55771] = 419890975;
assign addr[55772] = 438627762;
assign addr[55773] = 457329769;
assign addr[55774] = 475995513;
assign addr[55775] = 494623513;
assign addr[55776] = 513212292;
assign addr[55777] = 531760377;
assign addr[55778] = 550266296;
assign addr[55779] = 568728583;
assign addr[55780] = 587145773;
assign addr[55781] = 605516406;
assign addr[55782] = 623839025;
assign addr[55783] = 642112178;
assign addr[55784] = 660334415;
assign addr[55785] = 678504291;
assign addr[55786] = 696620367;
assign addr[55787] = 714681204;
assign addr[55788] = 732685372;
assign addr[55789] = 750631442;
assign addr[55790] = 768517992;
assign addr[55791] = 786343603;
assign addr[55792] = 804106861;
assign addr[55793] = 821806359;
assign addr[55794] = 839440693;
assign addr[55795] = 857008464;
assign addr[55796] = 874508280;
assign addr[55797] = 891938752;
assign addr[55798] = 909298500;
assign addr[55799] = 926586145;
assign addr[55800] = 943800318;
assign addr[55801] = 960939653;
assign addr[55802] = 978002791;
assign addr[55803] = 994988380;
assign addr[55804] = 1011895073;
assign addr[55805] = 1028721528;
assign addr[55806] = 1045466412;
assign addr[55807] = 1062128397;
assign addr[55808] = 1078706161;
assign addr[55809] = 1095198391;
assign addr[55810] = 1111603778;
assign addr[55811] = 1127921022;
assign addr[55812] = 1144148829;
assign addr[55813] = 1160285911;
assign addr[55814] = 1176330990;
assign addr[55815] = 1192282793;
assign addr[55816] = 1208140056;
assign addr[55817] = 1223901520;
assign addr[55818] = 1239565936;
assign addr[55819] = 1255132063;
assign addr[55820] = 1270598665;
assign addr[55821] = 1285964516;
assign addr[55822] = 1301228398;
assign addr[55823] = 1316389101;
assign addr[55824] = 1331445422;
assign addr[55825] = 1346396168;
assign addr[55826] = 1361240152;
assign addr[55827] = 1375976199;
assign addr[55828] = 1390603139;
assign addr[55829] = 1405119813;
assign addr[55830] = 1419525069;
assign addr[55831] = 1433817766;
assign addr[55832] = 1447996770;
assign addr[55833] = 1462060956;
assign addr[55834] = 1476009210;
assign addr[55835] = 1489840425;
assign addr[55836] = 1503553506;
assign addr[55837] = 1517147363;
assign addr[55838] = 1530620920;
assign addr[55839] = 1543973108;
assign addr[55840] = 1557202869;
assign addr[55841] = 1570309153;
assign addr[55842] = 1583290921;
assign addr[55843] = 1596147143;
assign addr[55844] = 1608876801;
assign addr[55845] = 1621478885;
assign addr[55846] = 1633952396;
assign addr[55847] = 1646296344;
assign addr[55848] = 1658509750;
assign addr[55849] = 1670591647;
assign addr[55850] = 1682541077;
assign addr[55851] = 1694357091;
assign addr[55852] = 1706038753;
assign addr[55853] = 1717585136;
assign addr[55854] = 1728995326;
assign addr[55855] = 1740268417;
assign addr[55856] = 1751403515;
assign addr[55857] = 1762399737;
assign addr[55858] = 1773256212;
assign addr[55859] = 1783972079;
assign addr[55860] = 1794546487;
assign addr[55861] = 1804978599;
assign addr[55862] = 1815267588;
assign addr[55863] = 1825412636;
assign addr[55864] = 1835412941;
assign addr[55865] = 1845267708;
assign addr[55866] = 1854976157;
assign addr[55867] = 1864537518;
assign addr[55868] = 1873951032;
assign addr[55869] = 1883215953;
assign addr[55870] = 1892331547;
assign addr[55871] = 1901297091;
assign addr[55872] = 1910111873;
assign addr[55873] = 1918775195;
assign addr[55874] = 1927286370;
assign addr[55875] = 1935644723;
assign addr[55876] = 1943849591;
assign addr[55877] = 1951900324;
assign addr[55878] = 1959796283;
assign addr[55879] = 1967536842;
assign addr[55880] = 1975121388;
assign addr[55881] = 1982549318;
assign addr[55882] = 1989820044;
assign addr[55883] = 1996932990;
assign addr[55884] = 2003887591;
assign addr[55885] = 2010683297;
assign addr[55886] = 2017319567;
assign addr[55887] = 2023795876;
assign addr[55888] = 2030111710;
assign addr[55889] = 2036266570;
assign addr[55890] = 2042259965;
assign addr[55891] = 2048091422;
assign addr[55892] = 2053760478;
assign addr[55893] = 2059266683;
assign addr[55894] = 2064609600;
assign addr[55895] = 2069788807;
assign addr[55896] = 2074803892;
assign addr[55897] = 2079654458;
assign addr[55898] = 2084340120;
assign addr[55899] = 2088860507;
assign addr[55900] = 2093215260;
assign addr[55901] = 2097404033;
assign addr[55902] = 2101426496;
assign addr[55903] = 2105282327;
assign addr[55904] = 2108971223;
assign addr[55905] = 2112492891;
assign addr[55906] = 2115847050;
assign addr[55907] = 2119033436;
assign addr[55908] = 2122051796;
assign addr[55909] = 2124901890;
assign addr[55910] = 2127583492;
assign addr[55911] = 2130096389;
assign addr[55912] = 2132440383;
assign addr[55913] = 2134615288;
assign addr[55914] = 2136620930;
assign addr[55915] = 2138457152;
assign addr[55916] = 2140123807;
assign addr[55917] = 2141620763;
assign addr[55918] = 2142947902;
assign addr[55919] = 2144105118;
assign addr[55920] = 2145092320;
assign addr[55921] = 2145909429;
assign addr[55922] = 2146556380;
assign addr[55923] = 2147033123;
assign addr[55924] = 2147339619;
assign addr[55925] = 2147475844;
assign addr[55926] = 2147441787;
assign addr[55927] = 2147237452;
assign addr[55928] = 2146862854;
assign addr[55929] = 2146318022;
assign addr[55930] = 2145603001;
assign addr[55931] = 2144717846;
assign addr[55932] = 2143662628;
assign addr[55933] = 2142437431;
assign addr[55934] = 2141042352;
assign addr[55935] = 2139477502;
assign addr[55936] = 2137743003;
assign addr[55937] = 2135838995;
assign addr[55938] = 2133765628;
assign addr[55939] = 2131523066;
assign addr[55940] = 2129111488;
assign addr[55941] = 2126531084;
assign addr[55942] = 2123782059;
assign addr[55943] = 2120864631;
assign addr[55944] = 2117779031;
assign addr[55945] = 2114525505;
assign addr[55946] = 2111104309;
assign addr[55947] = 2107515716;
assign addr[55948] = 2103760010;
assign addr[55949] = 2099837489;
assign addr[55950] = 2095748463;
assign addr[55951] = 2091493257;
assign addr[55952] = 2087072209;
assign addr[55953] = 2082485668;
assign addr[55954] = 2077733999;
assign addr[55955] = 2072817579;
assign addr[55956] = 2067736796;
assign addr[55957] = 2062492055;
assign addr[55958] = 2057083771;
assign addr[55959] = 2051512372;
assign addr[55960] = 2045778302;
assign addr[55961] = 2039882013;
assign addr[55962] = 2033823974;
assign addr[55963] = 2027604666;
assign addr[55964] = 2021224581;
assign addr[55965] = 2014684225;
assign addr[55966] = 2007984117;
assign addr[55967] = 2001124788;
assign addr[55968] = 1994106782;
assign addr[55969] = 1986930656;
assign addr[55970] = 1979596978;
assign addr[55971] = 1972106330;
assign addr[55972] = 1964459306;
assign addr[55973] = 1956656513;
assign addr[55974] = 1948698568;
assign addr[55975] = 1940586104;
assign addr[55976] = 1932319763;
assign addr[55977] = 1923900201;
assign addr[55978] = 1915328086;
assign addr[55979] = 1906604097;
assign addr[55980] = 1897728925;
assign addr[55981] = 1888703276;
assign addr[55982] = 1879527863;
assign addr[55983] = 1870203416;
assign addr[55984] = 1860730673;
assign addr[55985] = 1851110385;
assign addr[55986] = 1841343316;
assign addr[55987] = 1831430239;
assign addr[55988] = 1821371941;
assign addr[55989] = 1811169220;
assign addr[55990] = 1800822883;
assign addr[55991] = 1790333753;
assign addr[55992] = 1779702660;
assign addr[55993] = 1768930447;
assign addr[55994] = 1758017969;
assign addr[55995] = 1746966091;
assign addr[55996] = 1735775690;
assign addr[55997] = 1724447652;
assign addr[55998] = 1712982875;
assign addr[55999] = 1701382270;
assign addr[56000] = 1689646755;
assign addr[56001] = 1677777262;
assign addr[56002] = 1665774731;
assign addr[56003] = 1653640115;
assign addr[56004] = 1641374375;
assign addr[56005] = 1628978484;
assign addr[56006] = 1616453425;
assign addr[56007] = 1603800191;
assign addr[56008] = 1591019785;
assign addr[56009] = 1578113222;
assign addr[56010] = 1565081523;
assign addr[56011] = 1551925723;
assign addr[56012] = 1538646865;
assign addr[56013] = 1525246002;
assign addr[56014] = 1511724196;
assign addr[56015] = 1498082520;
assign addr[56016] = 1484322054;
assign addr[56017] = 1470443891;
assign addr[56018] = 1456449131;
assign addr[56019] = 1442338884;
assign addr[56020] = 1428114267;
assign addr[56021] = 1413776410;
assign addr[56022] = 1399326449;
assign addr[56023] = 1384765530;
assign addr[56024] = 1370094808;
assign addr[56025] = 1355315445;
assign addr[56026] = 1340428615;
assign addr[56027] = 1325435496;
assign addr[56028] = 1310337279;
assign addr[56029] = 1295135159;
assign addr[56030] = 1279830344;
assign addr[56031] = 1264424045;
assign addr[56032] = 1248917486;
assign addr[56033] = 1233311895;
assign addr[56034] = 1217608510;
assign addr[56035] = 1201808576;
assign addr[56036] = 1185913346;
assign addr[56037] = 1169924081;
assign addr[56038] = 1153842047;
assign addr[56039] = 1137668521;
assign addr[56040] = 1121404785;
assign addr[56041] = 1105052128;
assign addr[56042] = 1088611847;
assign addr[56043] = 1072085246;
assign addr[56044] = 1055473635;
assign addr[56045] = 1038778332;
assign addr[56046] = 1022000660;
assign addr[56047] = 1005141949;
assign addr[56048] = 988203537;
assign addr[56049] = 971186766;
assign addr[56050] = 954092986;
assign addr[56051] = 936923553;
assign addr[56052] = 919679827;
assign addr[56053] = 902363176;
assign addr[56054] = 884974973;
assign addr[56055] = 867516597;
assign addr[56056] = 849989433;
assign addr[56057] = 832394869;
assign addr[56058] = 814734301;
assign addr[56059] = 797009130;
assign addr[56060] = 779220762;
assign addr[56061] = 761370605;
assign addr[56062] = 743460077;
assign addr[56063] = 725490597;
assign addr[56064] = 707463589;
assign addr[56065] = 689380485;
assign addr[56066] = 671242716;
assign addr[56067] = 653051723;
assign addr[56068] = 634808946;
assign addr[56069] = 616515832;
assign addr[56070] = 598173833;
assign addr[56071] = 579784402;
assign addr[56072] = 561348998;
assign addr[56073] = 542869083;
assign addr[56074] = 524346121;
assign addr[56075] = 505781581;
assign addr[56076] = 487176937;
assign addr[56077] = 468533662;
assign addr[56078] = 449853235;
assign addr[56079] = 431137138;
assign addr[56080] = 412386854;
assign addr[56081] = 393603870;
assign addr[56082] = 374789676;
assign addr[56083] = 355945764;
assign addr[56084] = 337073627;
assign addr[56085] = 318174762;
assign addr[56086] = 299250668;
assign addr[56087] = 280302845;
assign addr[56088] = 261332796;
assign addr[56089] = 242342025;
assign addr[56090] = 223332037;
assign addr[56091] = 204304341;
assign addr[56092] = 185260444;
assign addr[56093] = 166201858;
assign addr[56094] = 147130093;
assign addr[56095] = 128046661;
assign addr[56096] = 108953076;
assign addr[56097] = 89850852;
assign addr[56098] = 70741503;
assign addr[56099] = 51626544;
assign addr[56100] = 32507492;
assign addr[56101] = 13385863;
assign addr[56102] = -5736829;
assign addr[56103] = -24859065;
assign addr[56104] = -43979330;
assign addr[56105] = -63096108;
assign addr[56106] = -82207882;
assign addr[56107] = -101313138;
assign addr[56108] = -120410361;
assign addr[56109] = -139498035;
assign addr[56110] = -158574649;
assign addr[56111] = -177638688;
assign addr[56112] = -196688642;
assign addr[56113] = -215722999;
assign addr[56114] = -234740251;
assign addr[56115] = -253738890;
assign addr[56116] = -272717408;
assign addr[56117] = -291674302;
assign addr[56118] = -310608068;
assign addr[56119] = -329517204;
assign addr[56120] = -348400212;
assign addr[56121] = -367255594;
assign addr[56122] = -386081854;
assign addr[56123] = -404877501;
assign addr[56124] = -423641043;
assign addr[56125] = -442370993;
assign addr[56126] = -461065866;
assign addr[56127] = -479724180;
assign addr[56128] = -498344454;
assign addr[56129] = -516925212;
assign addr[56130] = -535464981;
assign addr[56131] = -553962291;
assign addr[56132] = -572415676;
assign addr[56133] = -590823671;
assign addr[56134] = -609184818;
assign addr[56135] = -627497660;
assign addr[56136] = -645760745;
assign addr[56137] = -663972625;
assign addr[56138] = -682131857;
assign addr[56139] = -700236999;
assign addr[56140] = -718286617;
assign addr[56141] = -736279279;
assign addr[56142] = -754213559;
assign addr[56143] = -772088034;
assign addr[56144] = -789901288;
assign addr[56145] = -807651907;
assign addr[56146] = -825338484;
assign addr[56147] = -842959617;
assign addr[56148] = -860513908;
assign addr[56149] = -877999966;
assign addr[56150] = -895416404;
assign addr[56151] = -912761841;
assign addr[56152] = -930034901;
assign addr[56153] = -947234215;
assign addr[56154] = -964358420;
assign addr[56155] = -981406156;
assign addr[56156] = -998376073;
assign addr[56157] = -1015266825;
assign addr[56158] = -1032077073;
assign addr[56159] = -1048805483;
assign addr[56160] = -1065450729;
assign addr[56161] = -1082011492;
assign addr[56162] = -1098486458;
assign addr[56163] = -1114874320;
assign addr[56164] = -1131173780;
assign addr[56165] = -1147383544;
assign addr[56166] = -1163502328;
assign addr[56167] = -1179528853;
assign addr[56168] = -1195461849;
assign addr[56169] = -1211300053;
assign addr[56170] = -1227042207;
assign addr[56171] = -1242687064;
assign addr[56172] = -1258233384;
assign addr[56173] = -1273679934;
assign addr[56174] = -1289025489;
assign addr[56175] = -1304268832;
assign addr[56176] = -1319408754;
assign addr[56177] = -1334444055;
assign addr[56178] = -1349373543;
assign addr[56179] = -1364196034;
assign addr[56180] = -1378910353;
assign addr[56181] = -1393515332;
assign addr[56182] = -1408009814;
assign addr[56183] = -1422392650;
assign addr[56184] = -1436662698;
assign addr[56185] = -1450818828;
assign addr[56186] = -1464859917;
assign addr[56187] = -1478784851;
assign addr[56188] = -1492592527;
assign addr[56189] = -1506281850;
assign addr[56190] = -1519851733;
assign addr[56191] = -1533301101;
assign addr[56192] = -1546628888;
assign addr[56193] = -1559834037;
assign addr[56194] = -1572915501;
assign addr[56195] = -1585872242;
assign addr[56196] = -1598703233;
assign addr[56197] = -1611407456;
assign addr[56198] = -1623983905;
assign addr[56199] = -1636431582;
assign addr[56200] = -1648749499;
assign addr[56201] = -1660936681;
assign addr[56202] = -1672992161;
assign addr[56203] = -1684914983;
assign addr[56204] = -1696704201;
assign addr[56205] = -1708358881;
assign addr[56206] = -1719878099;
assign addr[56207] = -1731260941;
assign addr[56208] = -1742506504;
assign addr[56209] = -1753613897;
assign addr[56210] = -1764582240;
assign addr[56211] = -1775410662;
assign addr[56212] = -1786098304;
assign addr[56213] = -1796644320;
assign addr[56214] = -1807047873;
assign addr[56215] = -1817308138;
assign addr[56216] = -1827424302;
assign addr[56217] = -1837395562;
assign addr[56218] = -1847221128;
assign addr[56219] = -1856900221;
assign addr[56220] = -1866432072;
assign addr[56221] = -1875815927;
assign addr[56222] = -1885051042;
assign addr[56223] = -1894136683;
assign addr[56224] = -1903072131;
assign addr[56225] = -1911856677;
assign addr[56226] = -1920489624;
assign addr[56227] = -1928970288;
assign addr[56228] = -1937297997;
assign addr[56229] = -1945472089;
assign addr[56230] = -1953491918;
assign addr[56231] = -1961356847;
assign addr[56232] = -1969066252;
assign addr[56233] = -1976619522;
assign addr[56234] = -1984016058;
assign addr[56235] = -1991255274;
assign addr[56236] = -1998336596;
assign addr[56237] = -2005259462;
assign addr[56238] = -2012023322;
assign addr[56239] = -2018627642;
assign addr[56240] = -2025071897;
assign addr[56241] = -2031355576;
assign addr[56242] = -2037478181;
assign addr[56243] = -2043439226;
assign addr[56244] = -2049238240;
assign addr[56245] = -2054874761;
assign addr[56246] = -2060348343;
assign addr[56247] = -2065658552;
assign addr[56248] = -2070804967;
assign addr[56249] = -2075787180;
assign addr[56250] = -2080604795;
assign addr[56251] = -2085257431;
assign addr[56252] = -2089744719;
assign addr[56253] = -2094066304;
assign addr[56254] = -2098221841;
assign addr[56255] = -2102211002;
assign addr[56256] = -2106033471;
assign addr[56257] = -2109688944;
assign addr[56258] = -2113177132;
assign addr[56259] = -2116497758;
assign addr[56260] = -2119650558;
assign addr[56261] = -2122635283;
assign addr[56262] = -2125451696;
assign addr[56263] = -2128099574;
assign addr[56264] = -2130578706;
assign addr[56265] = -2132888897;
assign addr[56266] = -2135029962;
assign addr[56267] = -2137001733;
assign addr[56268] = -2138804053;
assign addr[56269] = -2140436778;
assign addr[56270] = -2141899780;
assign addr[56271] = -2143192942;
assign addr[56272] = -2144316162;
assign addr[56273] = -2145269351;
assign addr[56274] = -2146052433;
assign addr[56275] = -2146665347;
assign addr[56276] = -2147108043;
assign addr[56277] = -2147380486;
assign addr[56278] = -2147482655;
assign addr[56279] = -2147414542;
assign addr[56280] = -2147176152;
assign addr[56281] = -2146767505;
assign addr[56282] = -2146188631;
assign addr[56283] = -2145439578;
assign addr[56284] = -2144520405;
assign addr[56285] = -2143431184;
assign addr[56286] = -2142172003;
assign addr[56287] = -2140742960;
assign addr[56288] = -2139144169;
assign addr[56289] = -2137375758;
assign addr[56290] = -2135437865;
assign addr[56291] = -2133330646;
assign addr[56292] = -2131054266;
assign addr[56293] = -2128608907;
assign addr[56294] = -2125994762;
assign addr[56295] = -2123212038;
assign addr[56296] = -2120260957;
assign addr[56297] = -2117141752;
assign addr[56298] = -2113854671;
assign addr[56299] = -2110399974;
assign addr[56300] = -2106777935;
assign addr[56301] = -2102988841;
assign addr[56302] = -2099032994;
assign addr[56303] = -2094910706;
assign addr[56304] = -2090622304;
assign addr[56305] = -2086168128;
assign addr[56306] = -2081548533;
assign addr[56307] = -2076763883;
assign addr[56308] = -2071814558;
assign addr[56309] = -2066700952;
assign addr[56310] = -2061423468;
assign addr[56311] = -2055982526;
assign addr[56312] = -2050378558;
assign addr[56313] = -2044612007;
assign addr[56314] = -2038683330;
assign addr[56315] = -2032592999;
assign addr[56316] = -2026341495;
assign addr[56317] = -2019929315;
assign addr[56318] = -2013356967;
assign addr[56319] = -2006624971;
assign addr[56320] = -1999733863;
assign addr[56321] = -1992684188;
assign addr[56322] = -1985476506;
assign addr[56323] = -1978111387;
assign addr[56324] = -1970589416;
assign addr[56325] = -1962911189;
assign addr[56326] = -1955077316;
assign addr[56327] = -1947088417;
assign addr[56328] = -1938945125;
assign addr[56329] = -1930648088;
assign addr[56330] = -1922197961;
assign addr[56331] = -1913595416;
assign addr[56332] = -1904841135;
assign addr[56333] = -1895935811;
assign addr[56334] = -1886880151;
assign addr[56335] = -1877674873;
assign addr[56336] = -1868320707;
assign addr[56337] = -1858818395;
assign addr[56338] = -1849168689;
assign addr[56339] = -1839372356;
assign addr[56340] = -1829430172;
assign addr[56341] = -1819342925;
assign addr[56342] = -1809111415;
assign addr[56343] = -1798736454;
assign addr[56344] = -1788218865;
assign addr[56345] = -1777559480;
assign addr[56346] = -1766759146;
assign addr[56347] = -1755818718;
assign addr[56348] = -1744739065;
assign addr[56349] = -1733521064;
assign addr[56350] = -1722165606;
assign addr[56351] = -1710673591;
assign addr[56352] = -1699045930;
assign addr[56353] = -1687283545;
assign addr[56354] = -1675387369;
assign addr[56355] = -1663358344;
assign addr[56356] = -1651197426;
assign addr[56357] = -1638905577;
assign addr[56358] = -1626483774;
assign addr[56359] = -1613933000;
assign addr[56360] = -1601254251;
assign addr[56361] = -1588448533;
assign addr[56362] = -1575516860;
assign addr[56363] = -1562460258;
assign addr[56364] = -1549279763;
assign addr[56365] = -1535976419;
assign addr[56366] = -1522551282;
assign addr[56367] = -1509005416;
assign addr[56368] = -1495339895;
assign addr[56369] = -1481555802;
assign addr[56370] = -1467654232;
assign addr[56371] = -1453636285;
assign addr[56372] = -1439503074;
assign addr[56373] = -1425255719;
assign addr[56374] = -1410895350;
assign addr[56375] = -1396423105;
assign addr[56376] = -1381840133;
assign addr[56377] = -1367147589;
assign addr[56378] = -1352346639;
assign addr[56379] = -1337438456;
assign addr[56380] = -1322424222;
assign addr[56381] = -1307305128;
assign addr[56382] = -1292082373;
assign addr[56383] = -1276757164;
assign addr[56384] = -1261330715;
assign addr[56385] = -1245804251;
assign addr[56386] = -1230179002;
assign addr[56387] = -1214456207;
assign addr[56388] = -1198637114;
assign addr[56389] = -1182722976;
assign addr[56390] = -1166715055;
assign addr[56391] = -1150614620;
assign addr[56392] = -1134422949;
assign addr[56393] = -1118141326;
assign addr[56394] = -1101771040;
assign addr[56395] = -1085313391;
assign addr[56396] = -1068769683;
assign addr[56397] = -1052141228;
assign addr[56398] = -1035429345;
assign addr[56399] = -1018635358;
assign addr[56400] = -1001760600;
assign addr[56401] = -984806408;
assign addr[56402] = -967774128;
assign addr[56403] = -950665109;
assign addr[56404] = -933480707;
assign addr[56405] = -916222287;
assign addr[56406] = -898891215;
assign addr[56407] = -881488868;
assign addr[56408] = -864016623;
assign addr[56409] = -846475867;
assign addr[56410] = -828867991;
assign addr[56411] = -811194391;
assign addr[56412] = -793456467;
assign addr[56413] = -775655628;
assign addr[56414] = -757793284;
assign addr[56415] = -739870851;
assign addr[56416] = -721889752;
assign addr[56417] = -703851410;
assign addr[56418] = -685757258;
assign addr[56419] = -667608730;
assign addr[56420] = -649407264;
assign addr[56421] = -631154304;
assign addr[56422] = -612851297;
assign addr[56423] = -594499695;
assign addr[56424] = -576100953;
assign addr[56425] = -557656529;
assign addr[56426] = -539167887;
assign addr[56427] = -520636492;
assign addr[56428] = -502063814;
assign addr[56429] = -483451325;
assign addr[56430] = -464800501;
assign addr[56431] = -446112822;
assign addr[56432] = -427389768;
assign addr[56433] = -408632825;
assign addr[56434] = -389843480;
assign addr[56435] = -371023223;
assign addr[56436] = -352173546;
assign addr[56437] = -333295944;
assign addr[56438] = -314391913;
assign addr[56439] = -295462954;
assign addr[56440] = -276510565;
assign addr[56441] = -257536251;
assign addr[56442] = -238541516;
assign addr[56443] = -219527866;
assign addr[56444] = -200496809;
assign addr[56445] = -181449854;
assign addr[56446] = -162388511;
assign addr[56447] = -143314291;
assign addr[56448] = -124228708;
assign addr[56449] = -105133274;
assign addr[56450] = -86029503;
assign addr[56451] = -66918911;
assign addr[56452] = -47803013;
assign addr[56453] = -28683324;
assign addr[56454] = -9561361;
assign addr[56455] = 9561361;
assign addr[56456] = 28683324;
assign addr[56457] = 47803013;
assign addr[56458] = 66918911;
assign addr[56459] = 86029503;
assign addr[56460] = 105133274;
assign addr[56461] = 124228708;
assign addr[56462] = 143314291;
assign addr[56463] = 162388511;
assign addr[56464] = 181449854;
assign addr[56465] = 200496809;
assign addr[56466] = 219527866;
assign addr[56467] = 238541516;
assign addr[56468] = 257536251;
assign addr[56469] = 276510565;
assign addr[56470] = 295462953;
assign addr[56471] = 314391913;
assign addr[56472] = 333295944;
assign addr[56473] = 352173546;
assign addr[56474] = 371023223;
assign addr[56475] = 389843480;
assign addr[56476] = 408632825;
assign addr[56477] = 427389768;
assign addr[56478] = 446112822;
assign addr[56479] = 464800501;
assign addr[56480] = 483451325;
assign addr[56481] = 502063814;
assign addr[56482] = 520636492;
assign addr[56483] = 539167887;
assign addr[56484] = 557656529;
assign addr[56485] = 576100953;
assign addr[56486] = 594499695;
assign addr[56487] = 612851297;
assign addr[56488] = 631154304;
assign addr[56489] = 649407264;
assign addr[56490] = 667608730;
assign addr[56491] = 685757258;
assign addr[56492] = 703851410;
assign addr[56493] = 721889752;
assign addr[56494] = 739870851;
assign addr[56495] = 757793284;
assign addr[56496] = 775655628;
assign addr[56497] = 793456467;
assign addr[56498] = 811194391;
assign addr[56499] = 828867991;
assign addr[56500] = 846475867;
assign addr[56501] = 864016623;
assign addr[56502] = 881488868;
assign addr[56503] = 898891215;
assign addr[56504] = 916222287;
assign addr[56505] = 933480707;
assign addr[56506] = 950665109;
assign addr[56507] = 967774128;
assign addr[56508] = 984806408;
assign addr[56509] = 1001760600;
assign addr[56510] = 1018635358;
assign addr[56511] = 1035429345;
assign addr[56512] = 1052141228;
assign addr[56513] = 1068769683;
assign addr[56514] = 1085313391;
assign addr[56515] = 1101771040;
assign addr[56516] = 1118141326;
assign addr[56517] = 1134422949;
assign addr[56518] = 1150614620;
assign addr[56519] = 1166715055;
assign addr[56520] = 1182722976;
assign addr[56521] = 1198637114;
assign addr[56522] = 1214456207;
assign addr[56523] = 1230179002;
assign addr[56524] = 1245804251;
assign addr[56525] = 1261330715;
assign addr[56526] = 1276757164;
assign addr[56527] = 1292082373;
assign addr[56528] = 1307305128;
assign addr[56529] = 1322424222;
assign addr[56530] = 1337438456;
assign addr[56531] = 1352346639;
assign addr[56532] = 1367147589;
assign addr[56533] = 1381840133;
assign addr[56534] = 1396423105;
assign addr[56535] = 1410895350;
assign addr[56536] = 1425255719;
assign addr[56537] = 1439503074;
assign addr[56538] = 1453636285;
assign addr[56539] = 1467654232;
assign addr[56540] = 1481555802;
assign addr[56541] = 1495339895;
assign addr[56542] = 1509005416;
assign addr[56543] = 1522551282;
assign addr[56544] = 1535976419;
assign addr[56545] = 1549279763;
assign addr[56546] = 1562460258;
assign addr[56547] = 1575516860;
assign addr[56548] = 1588448533;
assign addr[56549] = 1601254251;
assign addr[56550] = 1613933000;
assign addr[56551] = 1626483774;
assign addr[56552] = 1638905577;
assign addr[56553] = 1651197426;
assign addr[56554] = 1663358344;
assign addr[56555] = 1675387369;
assign addr[56556] = 1687283545;
assign addr[56557] = 1699045930;
assign addr[56558] = 1710673591;
assign addr[56559] = 1722165606;
assign addr[56560] = 1733521064;
assign addr[56561] = 1744739065;
assign addr[56562] = 1755818718;
assign addr[56563] = 1766759146;
assign addr[56564] = 1777559480;
assign addr[56565] = 1788218865;
assign addr[56566] = 1798736454;
assign addr[56567] = 1809111415;
assign addr[56568] = 1819342925;
assign addr[56569] = 1829430172;
assign addr[56570] = 1839372356;
assign addr[56571] = 1849168689;
assign addr[56572] = 1858818395;
assign addr[56573] = 1868320707;
assign addr[56574] = 1877674873;
assign addr[56575] = 1886880151;
assign addr[56576] = 1895935811;
assign addr[56577] = 1904841135;
assign addr[56578] = 1913595416;
assign addr[56579] = 1922197961;
assign addr[56580] = 1930648088;
assign addr[56581] = 1938945125;
assign addr[56582] = 1947088417;
assign addr[56583] = 1955077316;
assign addr[56584] = 1962911189;
assign addr[56585] = 1970589416;
assign addr[56586] = 1978111387;
assign addr[56587] = 1985476506;
assign addr[56588] = 1992684188;
assign addr[56589] = 1999733863;
assign addr[56590] = 2006624971;
assign addr[56591] = 2013356967;
assign addr[56592] = 2019929315;
assign addr[56593] = 2026341495;
assign addr[56594] = 2032592999;
assign addr[56595] = 2038683330;
assign addr[56596] = 2044612007;
assign addr[56597] = 2050378558;
assign addr[56598] = 2055982526;
assign addr[56599] = 2061423468;
assign addr[56600] = 2066700952;
assign addr[56601] = 2071814558;
assign addr[56602] = 2076763883;
assign addr[56603] = 2081548533;
assign addr[56604] = 2086168128;
assign addr[56605] = 2090622304;
assign addr[56606] = 2094910706;
assign addr[56607] = 2099032994;
assign addr[56608] = 2102988841;
assign addr[56609] = 2106777935;
assign addr[56610] = 2110399974;
assign addr[56611] = 2113854671;
assign addr[56612] = 2117141752;
assign addr[56613] = 2120260957;
assign addr[56614] = 2123212038;
assign addr[56615] = 2125994762;
assign addr[56616] = 2128608907;
assign addr[56617] = 2131054266;
assign addr[56618] = 2133330646;
assign addr[56619] = 2135437865;
assign addr[56620] = 2137375758;
assign addr[56621] = 2139144169;
assign addr[56622] = 2140742960;
assign addr[56623] = 2142172003;
assign addr[56624] = 2143431184;
assign addr[56625] = 2144520405;
assign addr[56626] = 2145439578;
assign addr[56627] = 2146188631;
assign addr[56628] = 2146767505;
assign addr[56629] = 2147176152;
assign addr[56630] = 2147414542;
assign addr[56631] = 2147482655;
assign addr[56632] = 2147380486;
assign addr[56633] = 2147108043;
assign addr[56634] = 2146665347;
assign addr[56635] = 2146052433;
assign addr[56636] = 2145269351;
assign addr[56637] = 2144316162;
assign addr[56638] = 2143192942;
assign addr[56639] = 2141899780;
assign addr[56640] = 2140436778;
assign addr[56641] = 2138804053;
assign addr[56642] = 2137001733;
assign addr[56643] = 2135029962;
assign addr[56644] = 2132888897;
assign addr[56645] = 2130578706;
assign addr[56646] = 2128099574;
assign addr[56647] = 2125451696;
assign addr[56648] = 2122635283;
assign addr[56649] = 2119650558;
assign addr[56650] = 2116497758;
assign addr[56651] = 2113177132;
assign addr[56652] = 2109688944;
assign addr[56653] = 2106033471;
assign addr[56654] = 2102211002;
assign addr[56655] = 2098221841;
assign addr[56656] = 2094066304;
assign addr[56657] = 2089744719;
assign addr[56658] = 2085257431;
assign addr[56659] = 2080604795;
assign addr[56660] = 2075787180;
assign addr[56661] = 2070804967;
assign addr[56662] = 2065658552;
assign addr[56663] = 2060348343;
assign addr[56664] = 2054874761;
assign addr[56665] = 2049238240;
assign addr[56666] = 2043439226;
assign addr[56667] = 2037478181;
assign addr[56668] = 2031355576;
assign addr[56669] = 2025071897;
assign addr[56670] = 2018627642;
assign addr[56671] = 2012023322;
assign addr[56672] = 2005259462;
assign addr[56673] = 1998336596;
assign addr[56674] = 1991255274;
assign addr[56675] = 1984016058;
assign addr[56676] = 1976619522;
assign addr[56677] = 1969066252;
assign addr[56678] = 1961356847;
assign addr[56679] = 1953491918;
assign addr[56680] = 1945472089;
assign addr[56681] = 1937297997;
assign addr[56682] = 1928970288;
assign addr[56683] = 1920489624;
assign addr[56684] = 1911856677;
assign addr[56685] = 1903072131;
assign addr[56686] = 1894136683;
assign addr[56687] = 1885051042;
assign addr[56688] = 1875815927;
assign addr[56689] = 1866432072;
assign addr[56690] = 1856900221;
assign addr[56691] = 1847221128;
assign addr[56692] = 1837395562;
assign addr[56693] = 1827424302;
assign addr[56694] = 1817308138;
assign addr[56695] = 1807047873;
assign addr[56696] = 1796644320;
assign addr[56697] = 1786098304;
assign addr[56698] = 1775410662;
assign addr[56699] = 1764582240;
assign addr[56700] = 1753613897;
assign addr[56701] = 1742506504;
assign addr[56702] = 1731260941;
assign addr[56703] = 1719878099;
assign addr[56704] = 1708358881;
assign addr[56705] = 1696704201;
assign addr[56706] = 1684914983;
assign addr[56707] = 1672992161;
assign addr[56708] = 1660936681;
assign addr[56709] = 1648749499;
assign addr[56710] = 1636431582;
assign addr[56711] = 1623983905;
assign addr[56712] = 1611407456;
assign addr[56713] = 1598703233;
assign addr[56714] = 1585872242;
assign addr[56715] = 1572915501;
assign addr[56716] = 1559834037;
assign addr[56717] = 1546628888;
assign addr[56718] = 1533301101;
assign addr[56719] = 1519851733;
assign addr[56720] = 1506281850;
assign addr[56721] = 1492592527;
assign addr[56722] = 1478784851;
assign addr[56723] = 1464859917;
assign addr[56724] = 1450818828;
assign addr[56725] = 1436662698;
assign addr[56726] = 1422392650;
assign addr[56727] = 1408009814;
assign addr[56728] = 1393515332;
assign addr[56729] = 1378910353;
assign addr[56730] = 1364196034;
assign addr[56731] = 1349373543;
assign addr[56732] = 1334444055;
assign addr[56733] = 1319408754;
assign addr[56734] = 1304268832;
assign addr[56735] = 1289025489;
assign addr[56736] = 1273679934;
assign addr[56737] = 1258233384;
assign addr[56738] = 1242687064;
assign addr[56739] = 1227042207;
assign addr[56740] = 1211300053;
assign addr[56741] = 1195461849;
assign addr[56742] = 1179528853;
assign addr[56743] = 1163502328;
assign addr[56744] = 1147383544;
assign addr[56745] = 1131173780;
assign addr[56746] = 1114874320;
assign addr[56747] = 1098486458;
assign addr[56748] = 1082011492;
assign addr[56749] = 1065450729;
assign addr[56750] = 1048805483;
assign addr[56751] = 1032077073;
assign addr[56752] = 1015266825;
assign addr[56753] = 998376073;
assign addr[56754] = 981406156;
assign addr[56755] = 964358420;
assign addr[56756] = 947234215;
assign addr[56757] = 930034901;
assign addr[56758] = 912761841;
assign addr[56759] = 895416404;
assign addr[56760] = 877999966;
assign addr[56761] = 860513908;
assign addr[56762] = 842959617;
assign addr[56763] = 825338484;
assign addr[56764] = 807651907;
assign addr[56765] = 789901288;
assign addr[56766] = 772088034;
assign addr[56767] = 754213559;
assign addr[56768] = 736279279;
assign addr[56769] = 718286617;
assign addr[56770] = 700236999;
assign addr[56771] = 682131857;
assign addr[56772] = 663972625;
assign addr[56773] = 645760745;
assign addr[56774] = 627497660;
assign addr[56775] = 609184818;
assign addr[56776] = 590823671;
assign addr[56777] = 572415676;
assign addr[56778] = 553962291;
assign addr[56779] = 535464981;
assign addr[56780] = 516925212;
assign addr[56781] = 498344454;
assign addr[56782] = 479724180;
assign addr[56783] = 461065866;
assign addr[56784] = 442370993;
assign addr[56785] = 423641043;
assign addr[56786] = 404877501;
assign addr[56787] = 386081854;
assign addr[56788] = 367255594;
assign addr[56789] = 348400212;
assign addr[56790] = 329517204;
assign addr[56791] = 310608068;
assign addr[56792] = 291674302;
assign addr[56793] = 272717408;
assign addr[56794] = 253738890;
assign addr[56795] = 234740251;
assign addr[56796] = 215722999;
assign addr[56797] = 196688642;
assign addr[56798] = 177638688;
assign addr[56799] = 158574649;
assign addr[56800] = 139498035;
assign addr[56801] = 120410361;
assign addr[56802] = 101313138;
assign addr[56803] = 82207882;
assign addr[56804] = 63096108;
assign addr[56805] = 43979330;
assign addr[56806] = 24859065;
assign addr[56807] = 5736829;
assign addr[56808] = -13385863;
assign addr[56809] = -32507492;
assign addr[56810] = -51626544;
assign addr[56811] = -70741503;
assign addr[56812] = -89850852;
assign addr[56813] = -108953076;
assign addr[56814] = -128046661;
assign addr[56815] = -147130093;
assign addr[56816] = -166201858;
assign addr[56817] = -185260444;
assign addr[56818] = -204304341;
assign addr[56819] = -223332037;
assign addr[56820] = -242342025;
assign addr[56821] = -261332796;
assign addr[56822] = -280302845;
assign addr[56823] = -299250668;
assign addr[56824] = -318174762;
assign addr[56825] = -337073627;
assign addr[56826] = -355945764;
assign addr[56827] = -374789676;
assign addr[56828] = -393603870;
assign addr[56829] = -412386854;
assign addr[56830] = -431137138;
assign addr[56831] = -449853235;
assign addr[56832] = -468533662;
assign addr[56833] = -487176937;
assign addr[56834] = -505781581;
assign addr[56835] = -524346121;
assign addr[56836] = -542869083;
assign addr[56837] = -561348998;
assign addr[56838] = -579784402;
assign addr[56839] = -598173833;
assign addr[56840] = -616515832;
assign addr[56841] = -634808946;
assign addr[56842] = -653051723;
assign addr[56843] = -671242716;
assign addr[56844] = -689380485;
assign addr[56845] = -707463589;
assign addr[56846] = -725490597;
assign addr[56847] = -743460077;
assign addr[56848] = -761370605;
assign addr[56849] = -779220762;
assign addr[56850] = -797009130;
assign addr[56851] = -814734301;
assign addr[56852] = -832394869;
assign addr[56853] = -849989433;
assign addr[56854] = -867516597;
assign addr[56855] = -884974973;
assign addr[56856] = -902363176;
assign addr[56857] = -919679827;
assign addr[56858] = -936923553;
assign addr[56859] = -954092986;
assign addr[56860] = -971186766;
assign addr[56861] = -988203537;
assign addr[56862] = -1005141949;
assign addr[56863] = -1022000660;
assign addr[56864] = -1038778332;
assign addr[56865] = -1055473635;
assign addr[56866] = -1072085246;
assign addr[56867] = -1088611847;
assign addr[56868] = -1105052128;
assign addr[56869] = -1121404785;
assign addr[56870] = -1137668521;
assign addr[56871] = -1153842047;
assign addr[56872] = -1169924081;
assign addr[56873] = -1185913346;
assign addr[56874] = -1201808576;
assign addr[56875] = -1217608510;
assign addr[56876] = -1233311895;
assign addr[56877] = -1248917486;
assign addr[56878] = -1264424045;
assign addr[56879] = -1279830344;
assign addr[56880] = -1295135159;
assign addr[56881] = -1310337279;
assign addr[56882] = -1325435496;
assign addr[56883] = -1340428615;
assign addr[56884] = -1355315445;
assign addr[56885] = -1370094808;
assign addr[56886] = -1384765530;
assign addr[56887] = -1399326449;
assign addr[56888] = -1413776410;
assign addr[56889] = -1428114267;
assign addr[56890] = -1442338884;
assign addr[56891] = -1456449131;
assign addr[56892] = -1470443891;
assign addr[56893] = -1484322054;
assign addr[56894] = -1498082520;
assign addr[56895] = -1511724196;
assign addr[56896] = -1525246002;
assign addr[56897] = -1538646865;
assign addr[56898] = -1551925723;
assign addr[56899] = -1565081523;
assign addr[56900] = -1578113222;
assign addr[56901] = -1591019785;
assign addr[56902] = -1603800191;
assign addr[56903] = -1616453425;
assign addr[56904] = -1628978484;
assign addr[56905] = -1641374375;
assign addr[56906] = -1653640115;
assign addr[56907] = -1665774731;
assign addr[56908] = -1677777262;
assign addr[56909] = -1689646755;
assign addr[56910] = -1701382270;
assign addr[56911] = -1712982875;
assign addr[56912] = -1724447652;
assign addr[56913] = -1735775690;
assign addr[56914] = -1746966091;
assign addr[56915] = -1758017969;
assign addr[56916] = -1768930447;
assign addr[56917] = -1779702660;
assign addr[56918] = -1790333753;
assign addr[56919] = -1800822883;
assign addr[56920] = -1811169220;
assign addr[56921] = -1821371941;
assign addr[56922] = -1831430239;
assign addr[56923] = -1841343316;
assign addr[56924] = -1851110385;
assign addr[56925] = -1860730673;
assign addr[56926] = -1870203416;
assign addr[56927] = -1879527863;
assign addr[56928] = -1888703276;
assign addr[56929] = -1897728925;
assign addr[56930] = -1906604097;
assign addr[56931] = -1915328086;
assign addr[56932] = -1923900201;
assign addr[56933] = -1932319763;
assign addr[56934] = -1940586104;
assign addr[56935] = -1948698568;
assign addr[56936] = -1956656513;
assign addr[56937] = -1964459306;
assign addr[56938] = -1972106330;
assign addr[56939] = -1979596978;
assign addr[56940] = -1986930656;
assign addr[56941] = -1994106782;
assign addr[56942] = -2001124788;
assign addr[56943] = -2007984117;
assign addr[56944] = -2014684225;
assign addr[56945] = -2021224581;
assign addr[56946] = -2027604666;
assign addr[56947] = -2033823974;
assign addr[56948] = -2039882013;
assign addr[56949] = -2045778302;
assign addr[56950] = -2051512372;
assign addr[56951] = -2057083771;
assign addr[56952] = -2062492055;
assign addr[56953] = -2067736796;
assign addr[56954] = -2072817579;
assign addr[56955] = -2077733999;
assign addr[56956] = -2082485668;
assign addr[56957] = -2087072209;
assign addr[56958] = -2091493257;
assign addr[56959] = -2095748463;
assign addr[56960] = -2099837489;
assign addr[56961] = -2103760010;
assign addr[56962] = -2107515716;
assign addr[56963] = -2111104309;
assign addr[56964] = -2114525505;
assign addr[56965] = -2117779031;
assign addr[56966] = -2120864631;
assign addr[56967] = -2123782059;
assign addr[56968] = -2126531084;
assign addr[56969] = -2129111488;
assign addr[56970] = -2131523066;
assign addr[56971] = -2133765628;
assign addr[56972] = -2135838995;
assign addr[56973] = -2137743003;
assign addr[56974] = -2139477502;
assign addr[56975] = -2141042352;
assign addr[56976] = -2142437431;
assign addr[56977] = -2143662628;
assign addr[56978] = -2144717846;
assign addr[56979] = -2145603001;
assign addr[56980] = -2146318022;
assign addr[56981] = -2146862854;
assign addr[56982] = -2147237452;
assign addr[56983] = -2147441787;
assign addr[56984] = -2147475844;
assign addr[56985] = -2147339619;
assign addr[56986] = -2147033123;
assign addr[56987] = -2146556380;
assign addr[56988] = -2145909429;
assign addr[56989] = -2145092320;
assign addr[56990] = -2144105118;
assign addr[56991] = -2142947902;
assign addr[56992] = -2141620763;
assign addr[56993] = -2140123807;
assign addr[56994] = -2138457152;
assign addr[56995] = -2136620930;
assign addr[56996] = -2134615288;
assign addr[56997] = -2132440383;
assign addr[56998] = -2130096389;
assign addr[56999] = -2127583492;
assign addr[57000] = -2124901890;
assign addr[57001] = -2122051796;
assign addr[57002] = -2119033436;
assign addr[57003] = -2115847050;
assign addr[57004] = -2112492891;
assign addr[57005] = -2108971223;
assign addr[57006] = -2105282327;
assign addr[57007] = -2101426496;
assign addr[57008] = -2097404033;
assign addr[57009] = -2093215260;
assign addr[57010] = -2088860507;
assign addr[57011] = -2084340120;
assign addr[57012] = -2079654458;
assign addr[57013] = -2074803892;
assign addr[57014] = -2069788807;
assign addr[57015] = -2064609600;
assign addr[57016] = -2059266683;
assign addr[57017] = -2053760478;
assign addr[57018] = -2048091422;
assign addr[57019] = -2042259965;
assign addr[57020] = -2036266570;
assign addr[57021] = -2030111710;
assign addr[57022] = -2023795876;
assign addr[57023] = -2017319567;
assign addr[57024] = -2010683297;
assign addr[57025] = -2003887591;
assign addr[57026] = -1996932990;
assign addr[57027] = -1989820044;
assign addr[57028] = -1982549318;
assign addr[57029] = -1975121388;
assign addr[57030] = -1967536842;
assign addr[57031] = -1959796283;
assign addr[57032] = -1951900324;
assign addr[57033] = -1943849591;
assign addr[57034] = -1935644723;
assign addr[57035] = -1927286370;
assign addr[57036] = -1918775195;
assign addr[57037] = -1910111873;
assign addr[57038] = -1901297091;
assign addr[57039] = -1892331547;
assign addr[57040] = -1883215953;
assign addr[57041] = -1873951032;
assign addr[57042] = -1864537518;
assign addr[57043] = -1854976157;
assign addr[57044] = -1845267708;
assign addr[57045] = -1835412941;
assign addr[57046] = -1825412636;
assign addr[57047] = -1815267588;
assign addr[57048] = -1804978599;
assign addr[57049] = -1794546487;
assign addr[57050] = -1783972079;
assign addr[57051] = -1773256212;
assign addr[57052] = -1762399737;
assign addr[57053] = -1751403515;
assign addr[57054] = -1740268417;
assign addr[57055] = -1728995326;
assign addr[57056] = -1717585136;
assign addr[57057] = -1706038753;
assign addr[57058] = -1694357091;
assign addr[57059] = -1682541077;
assign addr[57060] = -1670591647;
assign addr[57061] = -1658509750;
assign addr[57062] = -1646296344;
assign addr[57063] = -1633952396;
assign addr[57064] = -1621478885;
assign addr[57065] = -1608876801;
assign addr[57066] = -1596147143;
assign addr[57067] = -1583290921;
assign addr[57068] = -1570309153;
assign addr[57069] = -1557202869;
assign addr[57070] = -1543973108;
assign addr[57071] = -1530620920;
assign addr[57072] = -1517147363;
assign addr[57073] = -1503553506;
assign addr[57074] = -1489840425;
assign addr[57075] = -1476009210;
assign addr[57076] = -1462060956;
assign addr[57077] = -1447996770;
assign addr[57078] = -1433817766;
assign addr[57079] = -1419525069;
assign addr[57080] = -1405119813;
assign addr[57081] = -1390603139;
assign addr[57082] = -1375976199;
assign addr[57083] = -1361240152;
assign addr[57084] = -1346396168;
assign addr[57085] = -1331445422;
assign addr[57086] = -1316389101;
assign addr[57087] = -1301228398;
assign addr[57088] = -1285964516;
assign addr[57089] = -1270598665;
assign addr[57090] = -1255132063;
assign addr[57091] = -1239565936;
assign addr[57092] = -1223901520;
assign addr[57093] = -1208140056;
assign addr[57094] = -1192282793;
assign addr[57095] = -1176330990;
assign addr[57096] = -1160285911;
assign addr[57097] = -1144148829;
assign addr[57098] = -1127921022;
assign addr[57099] = -1111603778;
assign addr[57100] = -1095198391;
assign addr[57101] = -1078706161;
assign addr[57102] = -1062128397;
assign addr[57103] = -1045466412;
assign addr[57104] = -1028721528;
assign addr[57105] = -1011895073;
assign addr[57106] = -994988380;
assign addr[57107] = -978002791;
assign addr[57108] = -960939653;
assign addr[57109] = -943800318;
assign addr[57110] = -926586145;
assign addr[57111] = -909298500;
assign addr[57112] = -891938752;
assign addr[57113] = -874508280;
assign addr[57114] = -857008464;
assign addr[57115] = -839440693;
assign addr[57116] = -821806359;
assign addr[57117] = -804106861;
assign addr[57118] = -786343603;
assign addr[57119] = -768517992;
assign addr[57120] = -750631442;
assign addr[57121] = -732685372;
assign addr[57122] = -714681204;
assign addr[57123] = -696620367;
assign addr[57124] = -678504291;
assign addr[57125] = -660334415;
assign addr[57126] = -642112178;
assign addr[57127] = -623839025;
assign addr[57128] = -605516406;
assign addr[57129] = -587145773;
assign addr[57130] = -568728583;
assign addr[57131] = -550266296;
assign addr[57132] = -531760377;
assign addr[57133] = -513212292;
assign addr[57134] = -494623513;
assign addr[57135] = -475995513;
assign addr[57136] = -457329769;
assign addr[57137] = -438627762;
assign addr[57138] = -419890975;
assign addr[57139] = -401120892;
assign addr[57140] = -382319004;
assign addr[57141] = -363486799;
assign addr[57142] = -344625773;
assign addr[57143] = -325737419;
assign addr[57144] = -306823237;
assign addr[57145] = -287884725;
assign addr[57146] = -268923386;
assign addr[57147] = -249940723;
assign addr[57148] = -230938242;
assign addr[57149] = -211917448;
assign addr[57150] = -192879850;
assign addr[57151] = -173826959;
assign addr[57152] = -154760284;
assign addr[57153] = -135681337;
assign addr[57154] = -116591632;
assign addr[57155] = -97492681;
assign addr[57156] = -78386000;
assign addr[57157] = -59273104;
assign addr[57158] = -40155507;
assign addr[57159] = -21034727;
assign addr[57160] = -1912278;
assign addr[57161] = 17210322;
assign addr[57162] = 36331557;
assign addr[57163] = 55449912;
assign addr[57164] = 74563870;
assign addr[57165] = 93671915;
assign addr[57166] = 112772533;
assign addr[57167] = 131864208;
assign addr[57168] = 150945428;
assign addr[57169] = 170014678;
assign addr[57170] = 189070447;
assign addr[57171] = 208111224;
assign addr[57172] = 227135500;
assign addr[57173] = 246141764;
assign addr[57174] = 265128512;
assign addr[57175] = 284094236;
assign addr[57176] = 303037433;
assign addr[57177] = 321956601;
assign addr[57178] = 340850240;
assign addr[57179] = 359716852;
assign addr[57180] = 378554940;
assign addr[57181] = 397363011;
assign addr[57182] = 416139574;
assign addr[57183] = 434883140;
assign addr[57184] = 453592221;
assign addr[57185] = 472265336;
assign addr[57186] = 490901003;
assign addr[57187] = 509497745;
assign addr[57188] = 528054086;
assign addr[57189] = 546568556;
assign addr[57190] = 565039687;
assign addr[57191] = 583466013;
assign addr[57192] = 601846074;
assign addr[57193] = 620178412;
assign addr[57194] = 638461574;
assign addr[57195] = 656694110;
assign addr[57196] = 674874574;
assign addr[57197] = 693001525;
assign addr[57198] = 711073524;
assign addr[57199] = 729089140;
assign addr[57200] = 747046944;
assign addr[57201] = 764945512;
assign addr[57202] = 782783424;
assign addr[57203] = 800559266;
assign addr[57204] = 818271628;
assign addr[57205] = 835919107;
assign addr[57206] = 853500302;
assign addr[57207] = 871013820;
assign addr[57208] = 888458272;
assign addr[57209] = 905832274;
assign addr[57210] = 923134450;
assign addr[57211] = 940363427;
assign addr[57212] = 957517838;
assign addr[57213] = 974596324;
assign addr[57214] = 991597531;
assign addr[57215] = 1008520110;
assign addr[57216] = 1025362720;
assign addr[57217] = 1042124025;
assign addr[57218] = 1058802695;
assign addr[57219] = 1075397409;
assign addr[57220] = 1091906851;
assign addr[57221] = 1108329711;
assign addr[57222] = 1124664687;
assign addr[57223] = 1140910484;
assign addr[57224] = 1157065814;
assign addr[57225] = 1173129396;
assign addr[57226] = 1189099956;
assign addr[57227] = 1204976227;
assign addr[57228] = 1220756951;
assign addr[57229] = 1236440877;
assign addr[57230] = 1252026760;
assign addr[57231] = 1267513365;
assign addr[57232] = 1282899464;
assign addr[57233] = 1298183838;
assign addr[57234] = 1313365273;
assign addr[57235] = 1328442566;
assign addr[57236] = 1343414522;
assign addr[57237] = 1358279953;
assign addr[57238] = 1373037681;
assign addr[57239] = 1387686535;
assign addr[57240] = 1402225355;
assign addr[57241] = 1416652986;
assign addr[57242] = 1430968286;
assign addr[57243] = 1445170118;
assign addr[57244] = 1459257358;
assign addr[57245] = 1473228887;
assign addr[57246] = 1487083598;
assign addr[57247] = 1500820393;
assign addr[57248] = 1514438181;
assign addr[57249] = 1527935884;
assign addr[57250] = 1541312431;
assign addr[57251] = 1554566762;
assign addr[57252] = 1567697824;
assign addr[57253] = 1580704578;
assign addr[57254] = 1593585992;
assign addr[57255] = 1606341043;
assign addr[57256] = 1618968722;
assign addr[57257] = 1631468027;
assign addr[57258] = 1643837966;
assign addr[57259] = 1656077559;
assign addr[57260] = 1668185835;
assign addr[57261] = 1680161834;
assign addr[57262] = 1692004606;
assign addr[57263] = 1703713213;
assign addr[57264] = 1715286726;
assign addr[57265] = 1726724227;
assign addr[57266] = 1738024810;
assign addr[57267] = 1749187577;
assign addr[57268] = 1760211645;
assign addr[57269] = 1771096139;
assign addr[57270] = 1781840195;
assign addr[57271] = 1792442963;
assign addr[57272] = 1802903601;
assign addr[57273] = 1813221279;
assign addr[57274] = 1823395180;
assign addr[57275] = 1833424497;
assign addr[57276] = 1843308435;
assign addr[57277] = 1853046210;
assign addr[57278] = 1862637049;
assign addr[57279] = 1872080193;
assign addr[57280] = 1881374892;
assign addr[57281] = 1890520410;
assign addr[57282] = 1899516021;
assign addr[57283] = 1908361011;
assign addr[57284] = 1917054681;
assign addr[57285] = 1925596340;
assign addr[57286] = 1933985310;
assign addr[57287] = 1942220928;
assign addr[57288] = 1950302539;
assign addr[57289] = 1958229503;
assign addr[57290] = 1966001192;
assign addr[57291] = 1973616989;
assign addr[57292] = 1981076290;
assign addr[57293] = 1988378503;
assign addr[57294] = 1995523051;
assign addr[57295] = 2002509365;
assign addr[57296] = 2009336893;
assign addr[57297] = 2016005093;
assign addr[57298] = 2022513436;
assign addr[57299] = 2028861406;
assign addr[57300] = 2035048499;
assign addr[57301] = 2041074226;
assign addr[57302] = 2046938108;
assign addr[57303] = 2052639680;
assign addr[57304] = 2058178491;
assign addr[57305] = 2063554100;
assign addr[57306] = 2068766083;
assign addr[57307] = 2073814024;
assign addr[57308] = 2078697525;
assign addr[57309] = 2083416198;
assign addr[57310] = 2087969669;
assign addr[57311] = 2092357577;
assign addr[57312] = 2096579573;
assign addr[57313] = 2100635323;
assign addr[57314] = 2104524506;
assign addr[57315] = 2108246813;
assign addr[57316] = 2111801949;
assign addr[57317] = 2115189632;
assign addr[57318] = 2118409593;
assign addr[57319] = 2121461578;
assign addr[57320] = 2124345343;
assign addr[57321] = 2127060661;
assign addr[57322] = 2129607316;
assign addr[57323] = 2131985106;
assign addr[57324] = 2134193842;
assign addr[57325] = 2136233350;
assign addr[57326] = 2138103468;
assign addr[57327] = 2139804048;
assign addr[57328] = 2141334954;
assign addr[57329] = 2142696065;
assign addr[57330] = 2143887273;
assign addr[57331] = 2144908484;
assign addr[57332] = 2145759618;
assign addr[57333] = 2146440605;
assign addr[57334] = 2146951393;
assign addr[57335] = 2147291941;
assign addr[57336] = 2147462221;
assign addr[57337] = 2147462221;
assign addr[57338] = 2147291941;
assign addr[57339] = 2146951393;
assign addr[57340] = 2146440605;
assign addr[57341] = 2145759618;
assign addr[57342] = 2144908484;
assign addr[57343] = 2143887273;
assign addr[57344] = 2142696065;
assign addr[57345] = 2141334954;
assign addr[57346] = 2139804048;
assign addr[57347] = 2138103468;
assign addr[57348] = 2136233350;
assign addr[57349] = 2134193842;
assign addr[57350] = 2131985106;
assign addr[57351] = 2129607316;
assign addr[57352] = 2127060661;
assign addr[57353] = 2124345343;
assign addr[57354] = 2121461578;
assign addr[57355] = 2118409593;
assign addr[57356] = 2115189632;
assign addr[57357] = 2111801949;
assign addr[57358] = 2108246813;
assign addr[57359] = 2104524506;
assign addr[57360] = 2100635323;
assign addr[57361] = 2096579573;
assign addr[57362] = 2092357577;
assign addr[57363] = 2087969669;
assign addr[57364] = 2083416198;
assign addr[57365] = 2078697525;
assign addr[57366] = 2073814024;
assign addr[57367] = 2068766083;
assign addr[57368] = 2063554100;
assign addr[57369] = 2058178491;
assign addr[57370] = 2052639680;
assign addr[57371] = 2046938108;
assign addr[57372] = 2041074226;
assign addr[57373] = 2035048499;
assign addr[57374] = 2028861406;
assign addr[57375] = 2022513436;
assign addr[57376] = 2016005093;
assign addr[57377] = 2009336893;
assign addr[57378] = 2002509365;
assign addr[57379] = 1995523051;
assign addr[57380] = 1988378503;
assign addr[57381] = 1981076290;
assign addr[57382] = 1973616989;
assign addr[57383] = 1966001192;
assign addr[57384] = 1958229503;
assign addr[57385] = 1950302539;
assign addr[57386] = 1942220928;
assign addr[57387] = 1933985310;
assign addr[57388] = 1925596340;
assign addr[57389] = 1917054681;
assign addr[57390] = 1908361011;
assign addr[57391] = 1899516021;
assign addr[57392] = 1890520410;
assign addr[57393] = 1881374892;
assign addr[57394] = 1872080193;
assign addr[57395] = 1862637049;
assign addr[57396] = 1853046210;
assign addr[57397] = 1843308435;
assign addr[57398] = 1833424497;
assign addr[57399] = 1823395180;
assign addr[57400] = 1813221279;
assign addr[57401] = 1802903601;
assign addr[57402] = 1792442963;
assign addr[57403] = 1781840195;
assign addr[57404] = 1771096139;
assign addr[57405] = 1760211645;
assign addr[57406] = 1749187577;
assign addr[57407] = 1738024810;
assign addr[57408] = 1726724227;
assign addr[57409] = 1715286726;
assign addr[57410] = 1703713213;
assign addr[57411] = 1692004606;
assign addr[57412] = 1680161834;
assign addr[57413] = 1668185835;
assign addr[57414] = 1656077559;
assign addr[57415] = 1643837966;
assign addr[57416] = 1631468027;
assign addr[57417] = 1618968722;
assign addr[57418] = 1606341043;
assign addr[57419] = 1593585992;
assign addr[57420] = 1580704578;
assign addr[57421] = 1567697824;
assign addr[57422] = 1554566762;
assign addr[57423] = 1541312431;
assign addr[57424] = 1527935884;
assign addr[57425] = 1514438181;
assign addr[57426] = 1500820393;
assign addr[57427] = 1487083598;
assign addr[57428] = 1473228887;
assign addr[57429] = 1459257358;
assign addr[57430] = 1445170118;
assign addr[57431] = 1430968286;
assign addr[57432] = 1416652986;
assign addr[57433] = 1402225355;
assign addr[57434] = 1387686535;
assign addr[57435] = 1373037681;
assign addr[57436] = 1358279953;
assign addr[57437] = 1343414522;
assign addr[57438] = 1328442566;
assign addr[57439] = 1313365273;
assign addr[57440] = 1298183838;
assign addr[57441] = 1282899464;
assign addr[57442] = 1267513365;
assign addr[57443] = 1252026760;
assign addr[57444] = 1236440877;
assign addr[57445] = 1220756951;
assign addr[57446] = 1204976227;
assign addr[57447] = 1189099956;
assign addr[57448] = 1173129396;
assign addr[57449] = 1157065814;
assign addr[57450] = 1140910484;
assign addr[57451] = 1124664687;
assign addr[57452] = 1108329711;
assign addr[57453] = 1091906851;
assign addr[57454] = 1075397409;
assign addr[57455] = 1058802695;
assign addr[57456] = 1042124025;
assign addr[57457] = 1025362720;
assign addr[57458] = 1008520110;
assign addr[57459] = 991597531;
assign addr[57460] = 974596324;
assign addr[57461] = 957517838;
assign addr[57462] = 940363427;
assign addr[57463] = 923134450;
assign addr[57464] = 905832274;
assign addr[57465] = 888458272;
assign addr[57466] = 871013820;
assign addr[57467] = 853500302;
assign addr[57468] = 835919107;
assign addr[57469] = 818271628;
assign addr[57470] = 800559266;
assign addr[57471] = 782783424;
assign addr[57472] = 764945512;
assign addr[57473] = 747046944;
assign addr[57474] = 729089140;
assign addr[57475] = 711073525;
assign addr[57476] = 693001525;
assign addr[57477] = 674874574;
assign addr[57478] = 656694110;
assign addr[57479] = 638461574;
assign addr[57480] = 620178412;
assign addr[57481] = 601846074;
assign addr[57482] = 583466013;
assign addr[57483] = 565039687;
assign addr[57484] = 546568556;
assign addr[57485] = 528054086;
assign addr[57486] = 509497745;
assign addr[57487] = 490901003;
assign addr[57488] = 472265336;
assign addr[57489] = 453592221;
assign addr[57490] = 434883140;
assign addr[57491] = 416139574;
assign addr[57492] = 397363011;
assign addr[57493] = 378554940;
assign addr[57494] = 359716852;
assign addr[57495] = 340850240;
assign addr[57496] = 321956601;
assign addr[57497] = 303037433;
assign addr[57498] = 284094236;
assign addr[57499] = 265128512;
assign addr[57500] = 246141764;
assign addr[57501] = 227135500;
assign addr[57502] = 208111224;
assign addr[57503] = 189070447;
assign addr[57504] = 170014678;
assign addr[57505] = 150945428;
assign addr[57506] = 131864208;
assign addr[57507] = 112772533;
assign addr[57508] = 93671915;
assign addr[57509] = 74563870;
assign addr[57510] = 55449912;
assign addr[57511] = 36331557;
assign addr[57512] = 17210322;
assign addr[57513] = -1912278;
assign addr[57514] = -21034727;
assign addr[57515] = -40155507;
assign addr[57516] = -59273104;
assign addr[57517] = -78386000;
assign addr[57518] = -97492681;
assign addr[57519] = -116591632;
assign addr[57520] = -135681337;
assign addr[57521] = -154760284;
assign addr[57522] = -173826959;
assign addr[57523] = -192879850;
assign addr[57524] = -211917448;
assign addr[57525] = -230938242;
assign addr[57526] = -249940723;
assign addr[57527] = -268923386;
assign addr[57528] = -287884725;
assign addr[57529] = -306823237;
assign addr[57530] = -325737419;
assign addr[57531] = -344625773;
assign addr[57532] = -363486799;
assign addr[57533] = -382319004;
assign addr[57534] = -401120892;
assign addr[57535] = -419890975;
assign addr[57536] = -438627762;
assign addr[57537] = -457329769;
assign addr[57538] = -475995513;
assign addr[57539] = -494623513;
assign addr[57540] = -513212292;
assign addr[57541] = -531760377;
assign addr[57542] = -550266296;
assign addr[57543] = -568728583;
assign addr[57544] = -587145773;
assign addr[57545] = -605516406;
assign addr[57546] = -623839025;
assign addr[57547] = -642112178;
assign addr[57548] = -660334415;
assign addr[57549] = -678504291;
assign addr[57550] = -696620367;
assign addr[57551] = -714681204;
assign addr[57552] = -732685372;
assign addr[57553] = -750631442;
assign addr[57554] = -768517992;
assign addr[57555] = -786343603;
assign addr[57556] = -804106861;
assign addr[57557] = -821806359;
assign addr[57558] = -839440693;
assign addr[57559] = -857008464;
assign addr[57560] = -874508280;
assign addr[57561] = -891938752;
assign addr[57562] = -909298500;
assign addr[57563] = -926586145;
assign addr[57564] = -943800318;
assign addr[57565] = -960939653;
assign addr[57566] = -978002791;
assign addr[57567] = -994988380;
assign addr[57568] = -1011895073;
assign addr[57569] = -1028721528;
assign addr[57570] = -1045466412;
assign addr[57571] = -1062128397;
assign addr[57572] = -1078706161;
assign addr[57573] = -1095198391;
assign addr[57574] = -1111603778;
assign addr[57575] = -1127921022;
assign addr[57576] = -1144148829;
assign addr[57577] = -1160285911;
assign addr[57578] = -1176330990;
assign addr[57579] = -1192282793;
assign addr[57580] = -1208140056;
assign addr[57581] = -1223901520;
assign addr[57582] = -1239565936;
assign addr[57583] = -1255132063;
assign addr[57584] = -1270598665;
assign addr[57585] = -1285964516;
assign addr[57586] = -1301228398;
assign addr[57587] = -1316389101;
assign addr[57588] = -1331445422;
assign addr[57589] = -1346396168;
assign addr[57590] = -1361240152;
assign addr[57591] = -1375976199;
assign addr[57592] = -1390603139;
assign addr[57593] = -1405119813;
assign addr[57594] = -1419525069;
assign addr[57595] = -1433817766;
assign addr[57596] = -1447996770;
assign addr[57597] = -1462060956;
assign addr[57598] = -1476009210;
assign addr[57599] = -1489840425;
assign addr[57600] = -1503553506;
assign addr[57601] = -1517147363;
assign addr[57602] = -1530620920;
assign addr[57603] = -1543973108;
assign addr[57604] = -1557202869;
assign addr[57605] = -1570309153;
assign addr[57606] = -1583290921;
assign addr[57607] = -1596147143;
assign addr[57608] = -1608876801;
assign addr[57609] = -1621478885;
assign addr[57610] = -1633952396;
assign addr[57611] = -1646296344;
assign addr[57612] = -1658509750;
assign addr[57613] = -1670591647;
assign addr[57614] = -1682541077;
assign addr[57615] = -1694357091;
assign addr[57616] = -1706038753;
assign addr[57617] = -1717585136;
assign addr[57618] = -1728995326;
assign addr[57619] = -1740268417;
assign addr[57620] = -1751403515;
assign addr[57621] = -1762399737;
assign addr[57622] = -1773256212;
assign addr[57623] = -1783972079;
assign addr[57624] = -1794546487;
assign addr[57625] = -1804978599;
assign addr[57626] = -1815267588;
assign addr[57627] = -1825412636;
assign addr[57628] = -1835412941;
assign addr[57629] = -1845267708;
assign addr[57630] = -1854976157;
assign addr[57631] = -1864537518;
assign addr[57632] = -1873951032;
assign addr[57633] = -1883215953;
assign addr[57634] = -1892331547;
assign addr[57635] = -1901297091;
assign addr[57636] = -1910111873;
assign addr[57637] = -1918775195;
assign addr[57638] = -1927286370;
assign addr[57639] = -1935644723;
assign addr[57640] = -1943849591;
assign addr[57641] = -1951900324;
assign addr[57642] = -1959796283;
assign addr[57643] = -1967536842;
assign addr[57644] = -1975121388;
assign addr[57645] = -1982549318;
assign addr[57646] = -1989820044;
assign addr[57647] = -1996932990;
assign addr[57648] = -2003887591;
assign addr[57649] = -2010683297;
assign addr[57650] = -2017319567;
assign addr[57651] = -2023795876;
assign addr[57652] = -2030111710;
assign addr[57653] = -2036266570;
assign addr[57654] = -2042259965;
assign addr[57655] = -2048091422;
assign addr[57656] = -2053760478;
assign addr[57657] = -2059266683;
assign addr[57658] = -2064609600;
assign addr[57659] = -2069788807;
assign addr[57660] = -2074803892;
assign addr[57661] = -2079654458;
assign addr[57662] = -2084340120;
assign addr[57663] = -2088860507;
assign addr[57664] = -2093215260;
assign addr[57665] = -2097404033;
assign addr[57666] = -2101426496;
assign addr[57667] = -2105282327;
assign addr[57668] = -2108971223;
assign addr[57669] = -2112492891;
assign addr[57670] = -2115847050;
assign addr[57671] = -2119033436;
assign addr[57672] = -2122051796;
assign addr[57673] = -2124901890;
assign addr[57674] = -2127583492;
assign addr[57675] = -2130096389;
assign addr[57676] = -2132440383;
assign addr[57677] = -2134615288;
assign addr[57678] = -2136620930;
assign addr[57679] = -2138457152;
assign addr[57680] = -2140123807;
assign addr[57681] = -2141620763;
assign addr[57682] = -2142947902;
assign addr[57683] = -2144105118;
assign addr[57684] = -2145092320;
assign addr[57685] = -2145909429;
assign addr[57686] = -2146556380;
assign addr[57687] = -2147033123;
assign addr[57688] = -2147339619;
assign addr[57689] = -2147475844;
assign addr[57690] = -2147441787;
assign addr[57691] = -2147237452;
assign addr[57692] = -2146862854;
assign addr[57693] = -2146318022;
assign addr[57694] = -2145603001;
assign addr[57695] = -2144717846;
assign addr[57696] = -2143662628;
assign addr[57697] = -2142437431;
assign addr[57698] = -2141042352;
assign addr[57699] = -2139477502;
assign addr[57700] = -2137743003;
assign addr[57701] = -2135838995;
assign addr[57702] = -2133765628;
assign addr[57703] = -2131523066;
assign addr[57704] = -2129111488;
assign addr[57705] = -2126531084;
assign addr[57706] = -2123782059;
assign addr[57707] = -2120864631;
assign addr[57708] = -2117779031;
assign addr[57709] = -2114525505;
assign addr[57710] = -2111104309;
assign addr[57711] = -2107515716;
assign addr[57712] = -2103760010;
assign addr[57713] = -2099837489;
assign addr[57714] = -2095748463;
assign addr[57715] = -2091493257;
assign addr[57716] = -2087072209;
assign addr[57717] = -2082485668;
assign addr[57718] = -2077733999;
assign addr[57719] = -2072817579;
assign addr[57720] = -2067736796;
assign addr[57721] = -2062492055;
assign addr[57722] = -2057083771;
assign addr[57723] = -2051512372;
assign addr[57724] = -2045778302;
assign addr[57725] = -2039882013;
assign addr[57726] = -2033823974;
assign addr[57727] = -2027604666;
assign addr[57728] = -2021224581;
assign addr[57729] = -2014684225;
assign addr[57730] = -2007984117;
assign addr[57731] = -2001124788;
assign addr[57732] = -1994106782;
assign addr[57733] = -1986930656;
assign addr[57734] = -1979596978;
assign addr[57735] = -1972106330;
assign addr[57736] = -1964459306;
assign addr[57737] = -1956656513;
assign addr[57738] = -1948698568;
assign addr[57739] = -1940586104;
assign addr[57740] = -1932319763;
assign addr[57741] = -1923900201;
assign addr[57742] = -1915328086;
assign addr[57743] = -1906604097;
assign addr[57744] = -1897728925;
assign addr[57745] = -1888703276;
assign addr[57746] = -1879527863;
assign addr[57747] = -1870203416;
assign addr[57748] = -1860730673;
assign addr[57749] = -1851110385;
assign addr[57750] = -1841343316;
assign addr[57751] = -1831430239;
assign addr[57752] = -1821371941;
assign addr[57753] = -1811169220;
assign addr[57754] = -1800822883;
assign addr[57755] = -1790333753;
assign addr[57756] = -1779702660;
assign addr[57757] = -1768930447;
assign addr[57758] = -1758017969;
assign addr[57759] = -1746966091;
assign addr[57760] = -1735775690;
assign addr[57761] = -1724447652;
assign addr[57762] = -1712982875;
assign addr[57763] = -1701382270;
assign addr[57764] = -1689646755;
assign addr[57765] = -1677777262;
assign addr[57766] = -1665774731;
assign addr[57767] = -1653640115;
assign addr[57768] = -1641374375;
assign addr[57769] = -1628978484;
assign addr[57770] = -1616453425;
assign addr[57771] = -1603800191;
assign addr[57772] = -1591019785;
assign addr[57773] = -1578113222;
assign addr[57774] = -1565081523;
assign addr[57775] = -1551925723;
assign addr[57776] = -1538646865;
assign addr[57777] = -1525246002;
assign addr[57778] = -1511724196;
assign addr[57779] = -1498082520;
assign addr[57780] = -1484322054;
assign addr[57781] = -1470443891;
assign addr[57782] = -1456449131;
assign addr[57783] = -1442338884;
assign addr[57784] = -1428114267;
assign addr[57785] = -1413776410;
assign addr[57786] = -1399326449;
assign addr[57787] = -1384765530;
assign addr[57788] = -1370094808;
assign addr[57789] = -1355315445;
assign addr[57790] = -1340428615;
assign addr[57791] = -1325435496;
assign addr[57792] = -1310337279;
assign addr[57793] = -1295135159;
assign addr[57794] = -1279830344;
assign addr[57795] = -1264424045;
assign addr[57796] = -1248917486;
assign addr[57797] = -1233311895;
assign addr[57798] = -1217608510;
assign addr[57799] = -1201808576;
assign addr[57800] = -1185913346;
assign addr[57801] = -1169924081;
assign addr[57802] = -1153842047;
assign addr[57803] = -1137668521;
assign addr[57804] = -1121404785;
assign addr[57805] = -1105052128;
assign addr[57806] = -1088611847;
assign addr[57807] = -1072085246;
assign addr[57808] = -1055473635;
assign addr[57809] = -1038778332;
assign addr[57810] = -1022000660;
assign addr[57811] = -1005141949;
assign addr[57812] = -988203537;
assign addr[57813] = -971186766;
assign addr[57814] = -954092986;
assign addr[57815] = -936923553;
assign addr[57816] = -919679827;
assign addr[57817] = -902363176;
assign addr[57818] = -884974973;
assign addr[57819] = -867516597;
assign addr[57820] = -849989433;
assign addr[57821] = -832394869;
assign addr[57822] = -814734301;
assign addr[57823] = -797009130;
assign addr[57824] = -779220762;
assign addr[57825] = -761370605;
assign addr[57826] = -743460077;
assign addr[57827] = -725490597;
assign addr[57828] = -707463589;
assign addr[57829] = -689380485;
assign addr[57830] = -671242716;
assign addr[57831] = -653051723;
assign addr[57832] = -634808946;
assign addr[57833] = -616515832;
assign addr[57834] = -598173833;
assign addr[57835] = -579784402;
assign addr[57836] = -561348998;
assign addr[57837] = -542869083;
assign addr[57838] = -524346121;
assign addr[57839] = -505781581;
assign addr[57840] = -487176937;
assign addr[57841] = -468533662;
assign addr[57842] = -449853235;
assign addr[57843] = -431137138;
assign addr[57844] = -412386854;
assign addr[57845] = -393603870;
assign addr[57846] = -374789676;
assign addr[57847] = -355945764;
assign addr[57848] = -337073627;
assign addr[57849] = -318174762;
assign addr[57850] = -299250668;
assign addr[57851] = -280302845;
assign addr[57852] = -261332796;
assign addr[57853] = -242342025;
assign addr[57854] = -223332037;
assign addr[57855] = -204304341;
assign addr[57856] = -185260444;
assign addr[57857] = -166201858;
assign addr[57858] = -147130093;
assign addr[57859] = -128046661;
assign addr[57860] = -108953076;
assign addr[57861] = -89850852;
assign addr[57862] = -70741503;
assign addr[57863] = -51626544;
assign addr[57864] = -32507492;
assign addr[57865] = -13385863;
assign addr[57866] = 5736829;
assign addr[57867] = 24859065;
assign addr[57868] = 43979330;
assign addr[57869] = 63096108;
assign addr[57870] = 82207882;
assign addr[57871] = 101313138;
assign addr[57872] = 120410361;
assign addr[57873] = 139498035;
assign addr[57874] = 158574649;
assign addr[57875] = 177638688;
assign addr[57876] = 196688642;
assign addr[57877] = 215722999;
assign addr[57878] = 234740251;
assign addr[57879] = 253738890;
assign addr[57880] = 272717408;
assign addr[57881] = 291674302;
assign addr[57882] = 310608068;
assign addr[57883] = 329517204;
assign addr[57884] = 348400212;
assign addr[57885] = 367255594;
assign addr[57886] = 386081854;
assign addr[57887] = 404877501;
assign addr[57888] = 423641043;
assign addr[57889] = 442370993;
assign addr[57890] = 461065866;
assign addr[57891] = 479724180;
assign addr[57892] = 498344454;
assign addr[57893] = 516925212;
assign addr[57894] = 535464981;
assign addr[57895] = 553962291;
assign addr[57896] = 572415676;
assign addr[57897] = 590823671;
assign addr[57898] = 609184818;
assign addr[57899] = 627497660;
assign addr[57900] = 645760745;
assign addr[57901] = 663972625;
assign addr[57902] = 682131857;
assign addr[57903] = 700236999;
assign addr[57904] = 718286617;
assign addr[57905] = 736279279;
assign addr[57906] = 754213559;
assign addr[57907] = 772088034;
assign addr[57908] = 789901288;
assign addr[57909] = 807651907;
assign addr[57910] = 825338484;
assign addr[57911] = 842959617;
assign addr[57912] = 860513908;
assign addr[57913] = 877999966;
assign addr[57914] = 895416404;
assign addr[57915] = 912761841;
assign addr[57916] = 930034901;
assign addr[57917] = 947234215;
assign addr[57918] = 964358420;
assign addr[57919] = 981406156;
assign addr[57920] = 998376073;
assign addr[57921] = 1015266825;
assign addr[57922] = 1032077073;
assign addr[57923] = 1048805483;
assign addr[57924] = 1065450729;
assign addr[57925] = 1082011492;
assign addr[57926] = 1098486458;
assign addr[57927] = 1114874320;
assign addr[57928] = 1131173780;
assign addr[57929] = 1147383544;
assign addr[57930] = 1163502328;
assign addr[57931] = 1179528853;
assign addr[57932] = 1195461849;
assign addr[57933] = 1211300053;
assign addr[57934] = 1227042207;
assign addr[57935] = 1242687064;
assign addr[57936] = 1258233384;
assign addr[57937] = 1273679934;
assign addr[57938] = 1289025489;
assign addr[57939] = 1304268832;
assign addr[57940] = 1319408754;
assign addr[57941] = 1334444055;
assign addr[57942] = 1349373543;
assign addr[57943] = 1364196034;
assign addr[57944] = 1378910353;
assign addr[57945] = 1393515332;
assign addr[57946] = 1408009814;
assign addr[57947] = 1422392650;
assign addr[57948] = 1436662698;
assign addr[57949] = 1450818828;
assign addr[57950] = 1464859917;
assign addr[57951] = 1478784851;
assign addr[57952] = 1492592527;
assign addr[57953] = 1506281850;
assign addr[57954] = 1519851733;
assign addr[57955] = 1533301101;
assign addr[57956] = 1546628888;
assign addr[57957] = 1559834037;
assign addr[57958] = 1572915501;
assign addr[57959] = 1585872242;
assign addr[57960] = 1598703233;
assign addr[57961] = 1611407456;
assign addr[57962] = 1623983905;
assign addr[57963] = 1636431582;
assign addr[57964] = 1648749499;
assign addr[57965] = 1660936681;
assign addr[57966] = 1672992161;
assign addr[57967] = 1684914983;
assign addr[57968] = 1696704201;
assign addr[57969] = 1708358881;
assign addr[57970] = 1719878099;
assign addr[57971] = 1731260941;
assign addr[57972] = 1742506504;
assign addr[57973] = 1753613897;
assign addr[57974] = 1764582240;
assign addr[57975] = 1775410662;
assign addr[57976] = 1786098304;
assign addr[57977] = 1796644320;
assign addr[57978] = 1807047873;
assign addr[57979] = 1817308138;
assign addr[57980] = 1827424302;
assign addr[57981] = 1837395562;
assign addr[57982] = 1847221128;
assign addr[57983] = 1856900221;
assign addr[57984] = 1866432072;
assign addr[57985] = 1875815927;
assign addr[57986] = 1885051042;
assign addr[57987] = 1894136683;
assign addr[57988] = 1903072131;
assign addr[57989] = 1911856677;
assign addr[57990] = 1920489624;
assign addr[57991] = 1928970288;
assign addr[57992] = 1937297997;
assign addr[57993] = 1945472089;
assign addr[57994] = 1953491918;
assign addr[57995] = 1961356847;
assign addr[57996] = 1969066252;
assign addr[57997] = 1976619522;
assign addr[57998] = 1984016058;
assign addr[57999] = 1991255274;
assign addr[58000] = 1998336596;
assign addr[58001] = 2005259462;
assign addr[58002] = 2012023322;
assign addr[58003] = 2018627642;
assign addr[58004] = 2025071897;
assign addr[58005] = 2031355576;
assign addr[58006] = 2037478181;
assign addr[58007] = 2043439226;
assign addr[58008] = 2049238240;
assign addr[58009] = 2054874761;
assign addr[58010] = 2060348343;
assign addr[58011] = 2065658552;
assign addr[58012] = 2070804967;
assign addr[58013] = 2075787180;
assign addr[58014] = 2080604795;
assign addr[58015] = 2085257431;
assign addr[58016] = 2089744719;
assign addr[58017] = 2094066304;
assign addr[58018] = 2098221841;
assign addr[58019] = 2102211002;
assign addr[58020] = 2106033471;
assign addr[58021] = 2109688944;
assign addr[58022] = 2113177132;
assign addr[58023] = 2116497758;
assign addr[58024] = 2119650558;
assign addr[58025] = 2122635283;
assign addr[58026] = 2125451696;
assign addr[58027] = 2128099574;
assign addr[58028] = 2130578706;
assign addr[58029] = 2132888897;
assign addr[58030] = 2135029962;
assign addr[58031] = 2137001733;
assign addr[58032] = 2138804053;
assign addr[58033] = 2140436778;
assign addr[58034] = 2141899780;
assign addr[58035] = 2143192942;
assign addr[58036] = 2144316162;
assign addr[58037] = 2145269351;
assign addr[58038] = 2146052433;
assign addr[58039] = 2146665347;
assign addr[58040] = 2147108043;
assign addr[58041] = 2147380486;
assign addr[58042] = 2147482655;
assign addr[58043] = 2147414542;
assign addr[58044] = 2147176152;
assign addr[58045] = 2146767505;
assign addr[58046] = 2146188631;
assign addr[58047] = 2145439578;
assign addr[58048] = 2144520405;
assign addr[58049] = 2143431184;
assign addr[58050] = 2142172003;
assign addr[58051] = 2140742960;
assign addr[58052] = 2139144169;
assign addr[58053] = 2137375758;
assign addr[58054] = 2135437865;
assign addr[58055] = 2133330646;
assign addr[58056] = 2131054266;
assign addr[58057] = 2128608907;
assign addr[58058] = 2125994762;
assign addr[58059] = 2123212038;
assign addr[58060] = 2120260957;
assign addr[58061] = 2117141752;
assign addr[58062] = 2113854671;
assign addr[58063] = 2110399974;
assign addr[58064] = 2106777935;
assign addr[58065] = 2102988841;
assign addr[58066] = 2099032994;
assign addr[58067] = 2094910706;
assign addr[58068] = 2090622304;
assign addr[58069] = 2086168128;
assign addr[58070] = 2081548533;
assign addr[58071] = 2076763883;
assign addr[58072] = 2071814558;
assign addr[58073] = 2066700952;
assign addr[58074] = 2061423468;
assign addr[58075] = 2055982526;
assign addr[58076] = 2050378558;
assign addr[58077] = 2044612007;
assign addr[58078] = 2038683330;
assign addr[58079] = 2032592999;
assign addr[58080] = 2026341495;
assign addr[58081] = 2019929315;
assign addr[58082] = 2013356967;
assign addr[58083] = 2006624971;
assign addr[58084] = 1999733863;
assign addr[58085] = 1992684188;
assign addr[58086] = 1985476506;
assign addr[58087] = 1978111387;
assign addr[58088] = 1970589416;
assign addr[58089] = 1962911189;
assign addr[58090] = 1955077316;
assign addr[58091] = 1947088417;
assign addr[58092] = 1938945125;
assign addr[58093] = 1930648088;
assign addr[58094] = 1922197961;
assign addr[58095] = 1913595416;
assign addr[58096] = 1904841135;
assign addr[58097] = 1895935811;
assign addr[58098] = 1886880151;
assign addr[58099] = 1877674873;
assign addr[58100] = 1868320707;
assign addr[58101] = 1858818395;
assign addr[58102] = 1849168689;
assign addr[58103] = 1839372356;
assign addr[58104] = 1829430172;
assign addr[58105] = 1819342925;
assign addr[58106] = 1809111415;
assign addr[58107] = 1798736454;
assign addr[58108] = 1788218865;
assign addr[58109] = 1777559480;
assign addr[58110] = 1766759146;
assign addr[58111] = 1755818718;
assign addr[58112] = 1744739065;
assign addr[58113] = 1733521064;
assign addr[58114] = 1722165606;
assign addr[58115] = 1710673591;
assign addr[58116] = 1699045930;
assign addr[58117] = 1687283545;
assign addr[58118] = 1675387369;
assign addr[58119] = 1663358344;
assign addr[58120] = 1651197426;
assign addr[58121] = 1638905577;
assign addr[58122] = 1626483774;
assign addr[58123] = 1613933000;
assign addr[58124] = 1601254251;
assign addr[58125] = 1588448533;
assign addr[58126] = 1575516860;
assign addr[58127] = 1562460258;
assign addr[58128] = 1549279763;
assign addr[58129] = 1535976419;
assign addr[58130] = 1522551282;
assign addr[58131] = 1509005416;
assign addr[58132] = 1495339895;
assign addr[58133] = 1481555802;
assign addr[58134] = 1467654232;
assign addr[58135] = 1453636285;
assign addr[58136] = 1439503074;
assign addr[58137] = 1425255719;
assign addr[58138] = 1410895350;
assign addr[58139] = 1396423105;
assign addr[58140] = 1381840133;
assign addr[58141] = 1367147589;
assign addr[58142] = 1352346639;
assign addr[58143] = 1337438456;
assign addr[58144] = 1322424222;
assign addr[58145] = 1307305128;
assign addr[58146] = 1292082373;
assign addr[58147] = 1276757164;
assign addr[58148] = 1261330715;
assign addr[58149] = 1245804251;
assign addr[58150] = 1230179002;
assign addr[58151] = 1214456207;
assign addr[58152] = 1198637114;
assign addr[58153] = 1182722976;
assign addr[58154] = 1166715055;
assign addr[58155] = 1150614620;
assign addr[58156] = 1134422949;
assign addr[58157] = 1118141326;
assign addr[58158] = 1101771040;
assign addr[58159] = 1085313391;
assign addr[58160] = 1068769683;
assign addr[58161] = 1052141228;
assign addr[58162] = 1035429345;
assign addr[58163] = 1018635358;
assign addr[58164] = 1001760600;
assign addr[58165] = 984806408;
assign addr[58166] = 967774128;
assign addr[58167] = 950665109;
assign addr[58168] = 933480707;
assign addr[58169] = 916222287;
assign addr[58170] = 898891215;
assign addr[58171] = 881488868;
assign addr[58172] = 864016623;
assign addr[58173] = 846475867;
assign addr[58174] = 828867991;
assign addr[58175] = 811194391;
assign addr[58176] = 793456467;
assign addr[58177] = 775655628;
assign addr[58178] = 757793284;
assign addr[58179] = 739870851;
assign addr[58180] = 721889752;
assign addr[58181] = 703851410;
assign addr[58182] = 685757258;
assign addr[58183] = 667608730;
assign addr[58184] = 649407264;
assign addr[58185] = 631154304;
assign addr[58186] = 612851297;
assign addr[58187] = 594499695;
assign addr[58188] = 576100953;
assign addr[58189] = 557656529;
assign addr[58190] = 539167887;
assign addr[58191] = 520636492;
assign addr[58192] = 502063814;
assign addr[58193] = 483451325;
assign addr[58194] = 464800501;
assign addr[58195] = 446112822;
assign addr[58196] = 427389768;
assign addr[58197] = 408632825;
assign addr[58198] = 389843480;
assign addr[58199] = 371023223;
assign addr[58200] = 352173546;
assign addr[58201] = 333295944;
assign addr[58202] = 314391913;
assign addr[58203] = 295462954;
assign addr[58204] = 276510565;
assign addr[58205] = 257536251;
assign addr[58206] = 238541516;
assign addr[58207] = 219527866;
assign addr[58208] = 200496809;
assign addr[58209] = 181449854;
assign addr[58210] = 162388511;
assign addr[58211] = 143314291;
assign addr[58212] = 124228708;
assign addr[58213] = 105133274;
assign addr[58214] = 86029503;
assign addr[58215] = 66918911;
assign addr[58216] = 47803013;
assign addr[58217] = 28683324;
assign addr[58218] = 9561361;
assign addr[58219] = -9561361;
assign addr[58220] = -28683324;
assign addr[58221] = -47803013;
assign addr[58222] = -66918911;
assign addr[58223] = -86029503;
assign addr[58224] = -105133274;
assign addr[58225] = -124228708;
assign addr[58226] = -143314291;
assign addr[58227] = -162388511;
assign addr[58228] = -181449854;
assign addr[58229] = -200496809;
assign addr[58230] = -219527866;
assign addr[58231] = -238541516;
assign addr[58232] = -257536251;
assign addr[58233] = -276510565;
assign addr[58234] = -295462953;
assign addr[58235] = -314391913;
assign addr[58236] = -333295944;
assign addr[58237] = -352173546;
assign addr[58238] = -371023223;
assign addr[58239] = -389843480;
assign addr[58240] = -408632825;
assign addr[58241] = -427389768;
assign addr[58242] = -446112822;
assign addr[58243] = -464800501;
assign addr[58244] = -483451325;
assign addr[58245] = -502063814;
assign addr[58246] = -520636492;
assign addr[58247] = -539167887;
assign addr[58248] = -557656529;
assign addr[58249] = -576100953;
assign addr[58250] = -594499695;
assign addr[58251] = -612851297;
assign addr[58252] = -631154304;
assign addr[58253] = -649407264;
assign addr[58254] = -667608730;
assign addr[58255] = -685757258;
assign addr[58256] = -703851410;
assign addr[58257] = -721889752;
assign addr[58258] = -739870851;
assign addr[58259] = -757793284;
assign addr[58260] = -775655628;
assign addr[58261] = -793456467;
assign addr[58262] = -811194391;
assign addr[58263] = -828867991;
assign addr[58264] = -846475867;
assign addr[58265] = -864016623;
assign addr[58266] = -881488868;
assign addr[58267] = -898891215;
assign addr[58268] = -916222287;
assign addr[58269] = -933480707;
assign addr[58270] = -950665109;
assign addr[58271] = -967774128;
assign addr[58272] = -984806408;
assign addr[58273] = -1001760600;
assign addr[58274] = -1018635358;
assign addr[58275] = -1035429345;
assign addr[58276] = -1052141228;
assign addr[58277] = -1068769683;
assign addr[58278] = -1085313391;
assign addr[58279] = -1101771040;
assign addr[58280] = -1118141326;
assign addr[58281] = -1134422949;
assign addr[58282] = -1150614620;
assign addr[58283] = -1166715055;
assign addr[58284] = -1182722976;
assign addr[58285] = -1198637114;
assign addr[58286] = -1214456207;
assign addr[58287] = -1230179002;
assign addr[58288] = -1245804251;
assign addr[58289] = -1261330715;
assign addr[58290] = -1276757164;
assign addr[58291] = -1292082373;
assign addr[58292] = -1307305128;
assign addr[58293] = -1322424222;
assign addr[58294] = -1337438456;
assign addr[58295] = -1352346639;
assign addr[58296] = -1367147589;
assign addr[58297] = -1381840133;
assign addr[58298] = -1396423105;
assign addr[58299] = -1410895350;
assign addr[58300] = -1425255719;
assign addr[58301] = -1439503074;
assign addr[58302] = -1453636285;
assign addr[58303] = -1467654232;
assign addr[58304] = -1481555802;
assign addr[58305] = -1495339895;
assign addr[58306] = -1509005416;
assign addr[58307] = -1522551282;
assign addr[58308] = -1535976419;
assign addr[58309] = -1549279763;
assign addr[58310] = -1562460258;
assign addr[58311] = -1575516860;
assign addr[58312] = -1588448533;
assign addr[58313] = -1601254251;
assign addr[58314] = -1613933000;
assign addr[58315] = -1626483774;
assign addr[58316] = -1638905577;
assign addr[58317] = -1651197426;
assign addr[58318] = -1663358344;
assign addr[58319] = -1675387369;
assign addr[58320] = -1687283545;
assign addr[58321] = -1699045930;
assign addr[58322] = -1710673591;
assign addr[58323] = -1722165606;
assign addr[58324] = -1733521064;
assign addr[58325] = -1744739065;
assign addr[58326] = -1755818718;
assign addr[58327] = -1766759146;
assign addr[58328] = -1777559480;
assign addr[58329] = -1788218865;
assign addr[58330] = -1798736454;
assign addr[58331] = -1809111415;
assign addr[58332] = -1819342925;
assign addr[58333] = -1829430172;
assign addr[58334] = -1839372356;
assign addr[58335] = -1849168689;
assign addr[58336] = -1858818395;
assign addr[58337] = -1868320707;
assign addr[58338] = -1877674873;
assign addr[58339] = -1886880151;
assign addr[58340] = -1895935811;
assign addr[58341] = -1904841135;
assign addr[58342] = -1913595416;
assign addr[58343] = -1922197961;
assign addr[58344] = -1930648088;
assign addr[58345] = -1938945125;
assign addr[58346] = -1947088417;
assign addr[58347] = -1955077316;
assign addr[58348] = -1962911189;
assign addr[58349] = -1970589416;
assign addr[58350] = -1978111387;
assign addr[58351] = -1985476506;
assign addr[58352] = -1992684188;
assign addr[58353] = -1999733863;
assign addr[58354] = -2006624971;
assign addr[58355] = -2013356967;
assign addr[58356] = -2019929315;
assign addr[58357] = -2026341495;
assign addr[58358] = -2032592999;
assign addr[58359] = -2038683330;
assign addr[58360] = -2044612007;
assign addr[58361] = -2050378558;
assign addr[58362] = -2055982526;
assign addr[58363] = -2061423468;
assign addr[58364] = -2066700952;
assign addr[58365] = -2071814558;
assign addr[58366] = -2076763883;
assign addr[58367] = -2081548533;
assign addr[58368] = -2086168128;
assign addr[58369] = -2090622304;
assign addr[58370] = -2094910706;
assign addr[58371] = -2099032994;
assign addr[58372] = -2102988841;
assign addr[58373] = -2106777935;
assign addr[58374] = -2110399974;
assign addr[58375] = -2113854671;
assign addr[58376] = -2117141752;
assign addr[58377] = -2120260957;
assign addr[58378] = -2123212038;
assign addr[58379] = -2125994762;
assign addr[58380] = -2128608907;
assign addr[58381] = -2131054266;
assign addr[58382] = -2133330646;
assign addr[58383] = -2135437865;
assign addr[58384] = -2137375758;
assign addr[58385] = -2139144169;
assign addr[58386] = -2140742960;
assign addr[58387] = -2142172003;
assign addr[58388] = -2143431184;
assign addr[58389] = -2144520405;
assign addr[58390] = -2145439578;
assign addr[58391] = -2146188631;
assign addr[58392] = -2146767505;
assign addr[58393] = -2147176152;
assign addr[58394] = -2147414542;
assign addr[58395] = -2147482655;
assign addr[58396] = -2147380486;
assign addr[58397] = -2147108043;
assign addr[58398] = -2146665347;
assign addr[58399] = -2146052433;
assign addr[58400] = -2145269351;
assign addr[58401] = -2144316162;
assign addr[58402] = -2143192942;
assign addr[58403] = -2141899780;
assign addr[58404] = -2140436778;
assign addr[58405] = -2138804053;
assign addr[58406] = -2137001733;
assign addr[58407] = -2135029962;
assign addr[58408] = -2132888897;
assign addr[58409] = -2130578706;
assign addr[58410] = -2128099574;
assign addr[58411] = -2125451696;
assign addr[58412] = -2122635283;
assign addr[58413] = -2119650558;
assign addr[58414] = -2116497758;
assign addr[58415] = -2113177132;
assign addr[58416] = -2109688944;
assign addr[58417] = -2106033471;
assign addr[58418] = -2102211002;
assign addr[58419] = -2098221841;
assign addr[58420] = -2094066304;
assign addr[58421] = -2089744719;
assign addr[58422] = -2085257431;
assign addr[58423] = -2080604795;
assign addr[58424] = -2075787180;
assign addr[58425] = -2070804967;
assign addr[58426] = -2065658552;
assign addr[58427] = -2060348343;
assign addr[58428] = -2054874761;
assign addr[58429] = -2049238240;
assign addr[58430] = -2043439226;
assign addr[58431] = -2037478181;
assign addr[58432] = -2031355576;
assign addr[58433] = -2025071897;
assign addr[58434] = -2018627642;
assign addr[58435] = -2012023322;
assign addr[58436] = -2005259462;
assign addr[58437] = -1998336596;
assign addr[58438] = -1991255274;
assign addr[58439] = -1984016058;
assign addr[58440] = -1976619522;
assign addr[58441] = -1969066252;
assign addr[58442] = -1961356847;
assign addr[58443] = -1953491918;
assign addr[58444] = -1945472089;
assign addr[58445] = -1937297997;
assign addr[58446] = -1928970288;
assign addr[58447] = -1920489624;
assign addr[58448] = -1911856677;
assign addr[58449] = -1903072131;
assign addr[58450] = -1894136683;
assign addr[58451] = -1885051042;
assign addr[58452] = -1875815927;
assign addr[58453] = -1866432072;
assign addr[58454] = -1856900221;
assign addr[58455] = -1847221128;
assign addr[58456] = -1837395562;
assign addr[58457] = -1827424302;
assign addr[58458] = -1817308138;
assign addr[58459] = -1807047873;
assign addr[58460] = -1796644320;
assign addr[58461] = -1786098304;
assign addr[58462] = -1775410662;
assign addr[58463] = -1764582240;
assign addr[58464] = -1753613897;
assign addr[58465] = -1742506504;
assign addr[58466] = -1731260941;
assign addr[58467] = -1719878099;
assign addr[58468] = -1708358881;
assign addr[58469] = -1696704201;
assign addr[58470] = -1684914983;
assign addr[58471] = -1672992161;
assign addr[58472] = -1660936681;
assign addr[58473] = -1648749499;
assign addr[58474] = -1636431582;
assign addr[58475] = -1623983905;
assign addr[58476] = -1611407456;
assign addr[58477] = -1598703233;
assign addr[58478] = -1585872242;
assign addr[58479] = -1572915501;
assign addr[58480] = -1559834037;
assign addr[58481] = -1546628888;
assign addr[58482] = -1533301101;
assign addr[58483] = -1519851733;
assign addr[58484] = -1506281850;
assign addr[58485] = -1492592527;
assign addr[58486] = -1478784851;
assign addr[58487] = -1464859917;
assign addr[58488] = -1450818828;
assign addr[58489] = -1436662698;
assign addr[58490] = -1422392650;
assign addr[58491] = -1408009814;
assign addr[58492] = -1393515332;
assign addr[58493] = -1378910353;
assign addr[58494] = -1364196034;
assign addr[58495] = -1349373543;
assign addr[58496] = -1334444055;
assign addr[58497] = -1319408754;
assign addr[58498] = -1304268832;
assign addr[58499] = -1289025489;
assign addr[58500] = -1273679934;
assign addr[58501] = -1258233384;
assign addr[58502] = -1242687064;
assign addr[58503] = -1227042207;
assign addr[58504] = -1211300053;
assign addr[58505] = -1195461849;
assign addr[58506] = -1179528853;
assign addr[58507] = -1163502328;
assign addr[58508] = -1147383544;
assign addr[58509] = -1131173780;
assign addr[58510] = -1114874320;
assign addr[58511] = -1098486458;
assign addr[58512] = -1082011492;
assign addr[58513] = -1065450729;
assign addr[58514] = -1048805483;
assign addr[58515] = -1032077073;
assign addr[58516] = -1015266825;
assign addr[58517] = -998376073;
assign addr[58518] = -981406156;
assign addr[58519] = -964358420;
assign addr[58520] = -947234215;
assign addr[58521] = -930034901;
assign addr[58522] = -912761841;
assign addr[58523] = -895416404;
assign addr[58524] = -877999966;
assign addr[58525] = -860513908;
assign addr[58526] = -842959617;
assign addr[58527] = -825338484;
assign addr[58528] = -807651907;
assign addr[58529] = -789901288;
assign addr[58530] = -772088034;
assign addr[58531] = -754213559;
assign addr[58532] = -736279279;
assign addr[58533] = -718286617;
assign addr[58534] = -700236999;
assign addr[58535] = -682131857;
assign addr[58536] = -663972625;
assign addr[58537] = -645760745;
assign addr[58538] = -627497660;
assign addr[58539] = -609184818;
assign addr[58540] = -590823671;
assign addr[58541] = -572415676;
assign addr[58542] = -553962291;
assign addr[58543] = -535464981;
assign addr[58544] = -516925212;
assign addr[58545] = -498344454;
assign addr[58546] = -479724180;
assign addr[58547] = -461065866;
assign addr[58548] = -442370993;
assign addr[58549] = -423641043;
assign addr[58550] = -404877501;
assign addr[58551] = -386081854;
assign addr[58552] = -367255594;
assign addr[58553] = -348400212;
assign addr[58554] = -329517204;
assign addr[58555] = -310608068;
assign addr[58556] = -291674302;
assign addr[58557] = -272717408;
assign addr[58558] = -253738890;
assign addr[58559] = -234740251;
assign addr[58560] = -215722999;
assign addr[58561] = -196688642;
assign addr[58562] = -177638688;
assign addr[58563] = -158574649;
assign addr[58564] = -139498035;
assign addr[58565] = -120410361;
assign addr[58566] = -101313138;
assign addr[58567] = -82207882;
assign addr[58568] = -63096108;
assign addr[58569] = -43979330;
assign addr[58570] = -24859065;
assign addr[58571] = -5736829;
assign addr[58572] = 13385863;
assign addr[58573] = 32507492;
assign addr[58574] = 51626544;
assign addr[58575] = 70741503;
assign addr[58576] = 89850852;
assign addr[58577] = 108953076;
assign addr[58578] = 128046661;
assign addr[58579] = 147130093;
assign addr[58580] = 166201858;
assign addr[58581] = 185260444;
assign addr[58582] = 204304341;
assign addr[58583] = 223332037;
assign addr[58584] = 242342025;
assign addr[58585] = 261332796;
assign addr[58586] = 280302845;
assign addr[58587] = 299250668;
assign addr[58588] = 318174762;
assign addr[58589] = 337073627;
assign addr[58590] = 355945764;
assign addr[58591] = 374789676;
assign addr[58592] = 393603870;
assign addr[58593] = 412386854;
assign addr[58594] = 431137138;
assign addr[58595] = 449853235;
assign addr[58596] = 468533662;
assign addr[58597] = 487176937;
assign addr[58598] = 505781581;
assign addr[58599] = 524346121;
assign addr[58600] = 542869083;
assign addr[58601] = 561348998;
assign addr[58602] = 579784402;
assign addr[58603] = 598173833;
assign addr[58604] = 616515832;
assign addr[58605] = 634808946;
assign addr[58606] = 653051723;
assign addr[58607] = 671242716;
assign addr[58608] = 689380485;
assign addr[58609] = 707463589;
assign addr[58610] = 725490597;
assign addr[58611] = 743460077;
assign addr[58612] = 761370605;
assign addr[58613] = 779220762;
assign addr[58614] = 797009130;
assign addr[58615] = 814734301;
assign addr[58616] = 832394869;
assign addr[58617] = 849989433;
assign addr[58618] = 867516597;
assign addr[58619] = 884974973;
assign addr[58620] = 902363176;
assign addr[58621] = 919679827;
assign addr[58622] = 936923553;
assign addr[58623] = 954092986;
assign addr[58624] = 971186766;
assign addr[58625] = 988203537;
assign addr[58626] = 1005141949;
assign addr[58627] = 1022000660;
assign addr[58628] = 1038778332;
assign addr[58629] = 1055473635;
assign addr[58630] = 1072085246;
assign addr[58631] = 1088611847;
assign addr[58632] = 1105052128;
assign addr[58633] = 1121404785;
assign addr[58634] = 1137668521;
assign addr[58635] = 1153842047;
assign addr[58636] = 1169924081;
assign addr[58637] = 1185913346;
assign addr[58638] = 1201808576;
assign addr[58639] = 1217608510;
assign addr[58640] = 1233311895;
assign addr[58641] = 1248917486;
assign addr[58642] = 1264424045;
assign addr[58643] = 1279830344;
assign addr[58644] = 1295135159;
assign addr[58645] = 1310337279;
assign addr[58646] = 1325435496;
assign addr[58647] = 1340428615;
assign addr[58648] = 1355315445;
assign addr[58649] = 1370094808;
assign addr[58650] = 1384765530;
assign addr[58651] = 1399326449;
assign addr[58652] = 1413776410;
assign addr[58653] = 1428114267;
assign addr[58654] = 1442338884;
assign addr[58655] = 1456449131;
assign addr[58656] = 1470443891;
assign addr[58657] = 1484322054;
assign addr[58658] = 1498082520;
assign addr[58659] = 1511724196;
assign addr[58660] = 1525246002;
assign addr[58661] = 1538646865;
assign addr[58662] = 1551925723;
assign addr[58663] = 1565081523;
assign addr[58664] = 1578113222;
assign addr[58665] = 1591019785;
assign addr[58666] = 1603800191;
assign addr[58667] = 1616453425;
assign addr[58668] = 1628978484;
assign addr[58669] = 1641374375;
assign addr[58670] = 1653640115;
assign addr[58671] = 1665774731;
assign addr[58672] = 1677777262;
assign addr[58673] = 1689646755;
assign addr[58674] = 1701382270;
assign addr[58675] = 1712982875;
assign addr[58676] = 1724447652;
assign addr[58677] = 1735775690;
assign addr[58678] = 1746966091;
assign addr[58679] = 1758017969;
assign addr[58680] = 1768930447;
assign addr[58681] = 1779702660;
assign addr[58682] = 1790333753;
assign addr[58683] = 1800822883;
assign addr[58684] = 1811169220;
assign addr[58685] = 1821371941;
assign addr[58686] = 1831430239;
assign addr[58687] = 1841343316;
assign addr[58688] = 1851110385;
assign addr[58689] = 1860730673;
assign addr[58690] = 1870203416;
assign addr[58691] = 1879527863;
assign addr[58692] = 1888703276;
assign addr[58693] = 1897728925;
assign addr[58694] = 1906604097;
assign addr[58695] = 1915328086;
assign addr[58696] = 1923900201;
assign addr[58697] = 1932319763;
assign addr[58698] = 1940586104;
assign addr[58699] = 1948698568;
assign addr[58700] = 1956656513;
assign addr[58701] = 1964459306;
assign addr[58702] = 1972106330;
assign addr[58703] = 1979596978;
assign addr[58704] = 1986930656;
assign addr[58705] = 1994106782;
assign addr[58706] = 2001124788;
assign addr[58707] = 2007984117;
assign addr[58708] = 2014684225;
assign addr[58709] = 2021224581;
assign addr[58710] = 2027604666;
assign addr[58711] = 2033823974;
assign addr[58712] = 2039882013;
assign addr[58713] = 2045778302;
assign addr[58714] = 2051512372;
assign addr[58715] = 2057083771;
assign addr[58716] = 2062492055;
assign addr[58717] = 2067736796;
assign addr[58718] = 2072817579;
assign addr[58719] = 2077733999;
assign addr[58720] = 2082485668;
assign addr[58721] = 2087072209;
assign addr[58722] = 2091493257;
assign addr[58723] = 2095748463;
assign addr[58724] = 2099837489;
assign addr[58725] = 2103760010;
assign addr[58726] = 2107515716;
assign addr[58727] = 2111104309;
assign addr[58728] = 2114525505;
assign addr[58729] = 2117779031;
assign addr[58730] = 2120864631;
assign addr[58731] = 2123782059;
assign addr[58732] = 2126531084;
assign addr[58733] = 2129111488;
assign addr[58734] = 2131523066;
assign addr[58735] = 2133765628;
assign addr[58736] = 2135838995;
assign addr[58737] = 2137743003;
assign addr[58738] = 2139477502;
assign addr[58739] = 2141042352;
assign addr[58740] = 2142437431;
assign addr[58741] = 2143662628;
assign addr[58742] = 2144717846;
assign addr[58743] = 2145603001;
assign addr[58744] = 2146318022;
assign addr[58745] = 2146862854;
assign addr[58746] = 2147237452;
assign addr[58747] = 2147441787;
assign addr[58748] = 2147475844;
assign addr[58749] = 2147339619;
assign addr[58750] = 2147033123;
assign addr[58751] = 2146556380;
assign addr[58752] = 2145909429;
assign addr[58753] = 2145092320;
assign addr[58754] = 2144105118;
assign addr[58755] = 2142947902;
assign addr[58756] = 2141620763;
assign addr[58757] = 2140123807;
assign addr[58758] = 2138457152;
assign addr[58759] = 2136620930;
assign addr[58760] = 2134615288;
assign addr[58761] = 2132440383;
assign addr[58762] = 2130096389;
assign addr[58763] = 2127583492;
assign addr[58764] = 2124901890;
assign addr[58765] = 2122051796;
assign addr[58766] = 2119033436;
assign addr[58767] = 2115847050;
assign addr[58768] = 2112492891;
assign addr[58769] = 2108971223;
assign addr[58770] = 2105282327;
assign addr[58771] = 2101426496;
assign addr[58772] = 2097404033;
assign addr[58773] = 2093215260;
assign addr[58774] = 2088860507;
assign addr[58775] = 2084340120;
assign addr[58776] = 2079654458;
assign addr[58777] = 2074803892;
assign addr[58778] = 2069788807;
assign addr[58779] = 2064609600;
assign addr[58780] = 2059266683;
assign addr[58781] = 2053760478;
assign addr[58782] = 2048091422;
assign addr[58783] = 2042259965;
assign addr[58784] = 2036266570;
assign addr[58785] = 2030111710;
assign addr[58786] = 2023795876;
assign addr[58787] = 2017319567;
assign addr[58788] = 2010683297;
assign addr[58789] = 2003887591;
assign addr[58790] = 1996932990;
assign addr[58791] = 1989820044;
assign addr[58792] = 1982549318;
assign addr[58793] = 1975121388;
assign addr[58794] = 1967536842;
assign addr[58795] = 1959796283;
assign addr[58796] = 1951900324;
assign addr[58797] = 1943849591;
assign addr[58798] = 1935644723;
assign addr[58799] = 1927286370;
assign addr[58800] = 1918775195;
assign addr[58801] = 1910111873;
assign addr[58802] = 1901297091;
assign addr[58803] = 1892331547;
assign addr[58804] = 1883215953;
assign addr[58805] = 1873951032;
assign addr[58806] = 1864537518;
assign addr[58807] = 1854976157;
assign addr[58808] = 1845267708;
assign addr[58809] = 1835412941;
assign addr[58810] = 1825412636;
assign addr[58811] = 1815267588;
assign addr[58812] = 1804978599;
assign addr[58813] = 1794546487;
assign addr[58814] = 1783972079;
assign addr[58815] = 1773256212;
assign addr[58816] = 1762399737;
assign addr[58817] = 1751403515;
assign addr[58818] = 1740268417;
assign addr[58819] = 1728995326;
assign addr[58820] = 1717585136;
assign addr[58821] = 1706038753;
assign addr[58822] = 1694357091;
assign addr[58823] = 1682541077;
assign addr[58824] = 1670591647;
assign addr[58825] = 1658509750;
assign addr[58826] = 1646296344;
assign addr[58827] = 1633952396;
assign addr[58828] = 1621478885;
assign addr[58829] = 1608876801;
assign addr[58830] = 1596147143;
assign addr[58831] = 1583290921;
assign addr[58832] = 1570309153;
assign addr[58833] = 1557202869;
assign addr[58834] = 1543973108;
assign addr[58835] = 1530620920;
assign addr[58836] = 1517147363;
assign addr[58837] = 1503553506;
assign addr[58838] = 1489840425;
assign addr[58839] = 1476009210;
assign addr[58840] = 1462060956;
assign addr[58841] = 1447996770;
assign addr[58842] = 1433817766;
assign addr[58843] = 1419525069;
assign addr[58844] = 1405119813;
assign addr[58845] = 1390603139;
assign addr[58846] = 1375976199;
assign addr[58847] = 1361240152;
assign addr[58848] = 1346396168;
assign addr[58849] = 1331445422;
assign addr[58850] = 1316389101;
assign addr[58851] = 1301228398;
assign addr[58852] = 1285964516;
assign addr[58853] = 1270598665;
assign addr[58854] = 1255132063;
assign addr[58855] = 1239565936;
assign addr[58856] = 1223901520;
assign addr[58857] = 1208140056;
assign addr[58858] = 1192282793;
assign addr[58859] = 1176330990;
assign addr[58860] = 1160285911;
assign addr[58861] = 1144148829;
assign addr[58862] = 1127921022;
assign addr[58863] = 1111603778;
assign addr[58864] = 1095198391;
assign addr[58865] = 1078706161;
assign addr[58866] = 1062128397;
assign addr[58867] = 1045466412;
assign addr[58868] = 1028721528;
assign addr[58869] = 1011895073;
assign addr[58870] = 994988380;
assign addr[58871] = 978002791;
assign addr[58872] = 960939653;
assign addr[58873] = 943800318;
assign addr[58874] = 926586145;
assign addr[58875] = 909298500;
assign addr[58876] = 891938752;
assign addr[58877] = 874508280;
assign addr[58878] = 857008464;
assign addr[58879] = 839440693;
assign addr[58880] = 821806359;
assign addr[58881] = 804106861;
assign addr[58882] = 786343603;
assign addr[58883] = 768517992;
assign addr[58884] = 750631442;
assign addr[58885] = 732685372;
assign addr[58886] = 714681204;
assign addr[58887] = 696620367;
assign addr[58888] = 678504291;
assign addr[58889] = 660334415;
assign addr[58890] = 642112178;
assign addr[58891] = 623839025;
assign addr[58892] = 605516406;
assign addr[58893] = 587145773;
assign addr[58894] = 568728583;
assign addr[58895] = 550266296;
assign addr[58896] = 531760377;
assign addr[58897] = 513212292;
assign addr[58898] = 494623513;
assign addr[58899] = 475995513;
assign addr[58900] = 457329769;
assign addr[58901] = 438627762;
assign addr[58902] = 419890975;
assign addr[58903] = 401120892;
assign addr[58904] = 382319004;
assign addr[58905] = 363486799;
assign addr[58906] = 344625773;
assign addr[58907] = 325737419;
assign addr[58908] = 306823237;
assign addr[58909] = 287884725;
assign addr[58910] = 268923386;
assign addr[58911] = 249940723;
assign addr[58912] = 230938242;
assign addr[58913] = 211917448;
assign addr[58914] = 192879850;
assign addr[58915] = 173826959;
assign addr[58916] = 154760284;
assign addr[58917] = 135681337;
assign addr[58918] = 116591632;
assign addr[58919] = 97492681;
assign addr[58920] = 78386000;
assign addr[58921] = 59273104;
assign addr[58922] = 40155507;
assign addr[58923] = 21034727;
assign addr[58924] = 1912278;
assign addr[58925] = -17210322;
assign addr[58926] = -36331557;
assign addr[58927] = -55449912;
assign addr[58928] = -74563870;
assign addr[58929] = -93671915;
assign addr[58930] = -112772533;
assign addr[58931] = -131864208;
assign addr[58932] = -150945428;
assign addr[58933] = -170014678;
assign addr[58934] = -189070447;
assign addr[58935] = -208111224;
assign addr[58936] = -227135500;
assign addr[58937] = -246141764;
assign addr[58938] = -265128512;
assign addr[58939] = -284094236;
assign addr[58940] = -303037433;
assign addr[58941] = -321956601;
assign addr[58942] = -340850240;
assign addr[58943] = -359716852;
assign addr[58944] = -378554940;
assign addr[58945] = -397363011;
assign addr[58946] = -416139574;
assign addr[58947] = -434883140;
assign addr[58948] = -453592221;
assign addr[58949] = -472265336;
assign addr[58950] = -490901003;
assign addr[58951] = -509497745;
assign addr[58952] = -528054086;
assign addr[58953] = -546568556;
assign addr[58954] = -565039687;
assign addr[58955] = -583466013;
assign addr[58956] = -601846074;
assign addr[58957] = -620178412;
assign addr[58958] = -638461574;
assign addr[58959] = -656694110;
assign addr[58960] = -674874574;
assign addr[58961] = -693001525;
assign addr[58962] = -711073524;
assign addr[58963] = -729089140;
assign addr[58964] = -747046944;
assign addr[58965] = -764945512;
assign addr[58966] = -782783424;
assign addr[58967] = -800559266;
assign addr[58968] = -818271628;
assign addr[58969] = -835919107;
assign addr[58970] = -853500302;
assign addr[58971] = -871013820;
assign addr[58972] = -888458272;
assign addr[58973] = -905832274;
assign addr[58974] = -923134450;
assign addr[58975] = -940363427;
assign addr[58976] = -957517838;
assign addr[58977] = -974596324;
assign addr[58978] = -991597531;
assign addr[58979] = -1008520110;
assign addr[58980] = -1025362720;
assign addr[58981] = -1042124025;
assign addr[58982] = -1058802695;
assign addr[58983] = -1075397409;
assign addr[58984] = -1091906851;
assign addr[58985] = -1108329711;
assign addr[58986] = -1124664687;
assign addr[58987] = -1140910484;
assign addr[58988] = -1157065814;
assign addr[58989] = -1173129396;
assign addr[58990] = -1189099956;
assign addr[58991] = -1204976227;
assign addr[58992] = -1220756951;
assign addr[58993] = -1236440877;
assign addr[58994] = -1252026760;
assign addr[58995] = -1267513365;
assign addr[58996] = -1282899464;
assign addr[58997] = -1298183838;
assign addr[58998] = -1313365273;
assign addr[58999] = -1328442566;
assign addr[59000] = -1343414522;
assign addr[59001] = -1358279953;
assign addr[59002] = -1373037681;
assign addr[59003] = -1387686535;
assign addr[59004] = -1402225355;
assign addr[59005] = -1416652986;
assign addr[59006] = -1430968286;
assign addr[59007] = -1445170118;
assign addr[59008] = -1459257358;
assign addr[59009] = -1473228887;
assign addr[59010] = -1487083598;
assign addr[59011] = -1500820393;
assign addr[59012] = -1514438181;
assign addr[59013] = -1527935884;
assign addr[59014] = -1541312431;
assign addr[59015] = -1554566762;
assign addr[59016] = -1567697824;
assign addr[59017] = -1580704578;
assign addr[59018] = -1593585992;
assign addr[59019] = -1606341043;
assign addr[59020] = -1618968722;
assign addr[59021] = -1631468027;
assign addr[59022] = -1643837966;
assign addr[59023] = -1656077559;
assign addr[59024] = -1668185835;
assign addr[59025] = -1680161834;
assign addr[59026] = -1692004606;
assign addr[59027] = -1703713213;
assign addr[59028] = -1715286726;
assign addr[59029] = -1726724227;
assign addr[59030] = -1738024810;
assign addr[59031] = -1749187577;
assign addr[59032] = -1760211645;
assign addr[59033] = -1771096139;
assign addr[59034] = -1781840195;
assign addr[59035] = -1792442963;
assign addr[59036] = -1802903601;
assign addr[59037] = -1813221279;
assign addr[59038] = -1823395180;
assign addr[59039] = -1833424497;
assign addr[59040] = -1843308435;
assign addr[59041] = -1853046210;
assign addr[59042] = -1862637049;
assign addr[59043] = -1872080193;
assign addr[59044] = -1881374892;
assign addr[59045] = -1890520410;
assign addr[59046] = -1899516021;
assign addr[59047] = -1908361011;
assign addr[59048] = -1917054681;
assign addr[59049] = -1925596340;
assign addr[59050] = -1933985310;
assign addr[59051] = -1942220928;
assign addr[59052] = -1950302539;
assign addr[59053] = -1958229503;
assign addr[59054] = -1966001192;
assign addr[59055] = -1973616989;
assign addr[59056] = -1981076290;
assign addr[59057] = -1988378503;
assign addr[59058] = -1995523051;
assign addr[59059] = -2002509365;
assign addr[59060] = -2009336893;
assign addr[59061] = -2016005093;
assign addr[59062] = -2022513436;
assign addr[59063] = -2028861406;
assign addr[59064] = -2035048499;
assign addr[59065] = -2041074226;
assign addr[59066] = -2046938108;
assign addr[59067] = -2052639680;
assign addr[59068] = -2058178491;
assign addr[59069] = -2063554100;
assign addr[59070] = -2068766083;
assign addr[59071] = -2073814024;
assign addr[59072] = -2078697525;
assign addr[59073] = -2083416198;
assign addr[59074] = -2087969669;
assign addr[59075] = -2092357577;
assign addr[59076] = -2096579573;
assign addr[59077] = -2100635323;
assign addr[59078] = -2104524506;
assign addr[59079] = -2108246813;
assign addr[59080] = -2111801949;
assign addr[59081] = -2115189632;
assign addr[59082] = -2118409593;
assign addr[59083] = -2121461578;
assign addr[59084] = -2124345343;
assign addr[59085] = -2127060661;
assign addr[59086] = -2129607316;
assign addr[59087] = -2131985106;
assign addr[59088] = -2134193842;
assign addr[59089] = -2136233350;
assign addr[59090] = -2138103468;
assign addr[59091] = -2139804048;
assign addr[59092] = -2141334954;
assign addr[59093] = -2142696065;
assign addr[59094] = -2143887273;
assign addr[59095] = -2144908484;
assign addr[59096] = -2145759618;
assign addr[59097] = -2146440605;
assign addr[59098] = -2146951393;
assign addr[59099] = -2147291941;
assign addr[59100] = -2147462221;
assign addr[59101] = -2147462221;
assign addr[59102] = -2147291941;
assign addr[59103] = -2146951393;
assign addr[59104] = -2146440605;
assign addr[59105] = -2145759618;
assign addr[59106] = -2144908484;
assign addr[59107] = -2143887273;
assign addr[59108] = -2142696065;
assign addr[59109] = -2141334954;
assign addr[59110] = -2139804048;
assign addr[59111] = -2138103468;
assign addr[59112] = -2136233350;
assign addr[59113] = -2134193842;
assign addr[59114] = -2131985106;
assign addr[59115] = -2129607316;
assign addr[59116] = -2127060661;
assign addr[59117] = -2124345343;
assign addr[59118] = -2121461578;
assign addr[59119] = -2118409593;
assign addr[59120] = -2115189632;
assign addr[59121] = -2111801949;
assign addr[59122] = -2108246813;
assign addr[59123] = -2104524506;
assign addr[59124] = -2100635323;
assign addr[59125] = -2096579573;
assign addr[59126] = -2092357577;
assign addr[59127] = -2087969669;
assign addr[59128] = -2083416198;
assign addr[59129] = -2078697525;
assign addr[59130] = -2073814024;
assign addr[59131] = -2068766083;
assign addr[59132] = -2063554100;
assign addr[59133] = -2058178491;
assign addr[59134] = -2052639680;
assign addr[59135] = -2046938108;
assign addr[59136] = -2041074226;
assign addr[59137] = -2035048499;
assign addr[59138] = -2028861406;
assign addr[59139] = -2022513436;
assign addr[59140] = -2016005093;
assign addr[59141] = -2009336893;
assign addr[59142] = -2002509365;
assign addr[59143] = -1995523051;
assign addr[59144] = -1988378503;
assign addr[59145] = -1981076290;
assign addr[59146] = -1973616989;
assign addr[59147] = -1966001192;
assign addr[59148] = -1958229503;
assign addr[59149] = -1950302539;
assign addr[59150] = -1942220928;
assign addr[59151] = -1933985310;
assign addr[59152] = -1925596340;
assign addr[59153] = -1917054681;
assign addr[59154] = -1908361011;
assign addr[59155] = -1899516021;
assign addr[59156] = -1890520410;
assign addr[59157] = -1881374892;
assign addr[59158] = -1872080193;
assign addr[59159] = -1862637049;
assign addr[59160] = -1853046210;
assign addr[59161] = -1843308435;
assign addr[59162] = -1833424497;
assign addr[59163] = -1823395180;
assign addr[59164] = -1813221279;
assign addr[59165] = -1802903601;
assign addr[59166] = -1792442963;
assign addr[59167] = -1781840195;
assign addr[59168] = -1771096139;
assign addr[59169] = -1760211645;
assign addr[59170] = -1749187577;
assign addr[59171] = -1738024810;
assign addr[59172] = -1726724227;
assign addr[59173] = -1715286726;
assign addr[59174] = -1703713213;
assign addr[59175] = -1692004606;
assign addr[59176] = -1680161834;
assign addr[59177] = -1668185835;
assign addr[59178] = -1656077559;
assign addr[59179] = -1643837966;
assign addr[59180] = -1631468027;
assign addr[59181] = -1618968722;
assign addr[59182] = -1606341043;
assign addr[59183] = -1593585992;
assign addr[59184] = -1580704578;
assign addr[59185] = -1567697824;
assign addr[59186] = -1554566762;
assign addr[59187] = -1541312431;
assign addr[59188] = -1527935884;
assign addr[59189] = -1514438181;
assign addr[59190] = -1500820393;
assign addr[59191] = -1487083598;
assign addr[59192] = -1473228887;
assign addr[59193] = -1459257358;
assign addr[59194] = -1445170118;
assign addr[59195] = -1430968286;
assign addr[59196] = -1416652986;
assign addr[59197] = -1402225355;
assign addr[59198] = -1387686535;
assign addr[59199] = -1373037681;
assign addr[59200] = -1358279953;
assign addr[59201] = -1343414522;
assign addr[59202] = -1328442566;
assign addr[59203] = -1313365273;
assign addr[59204] = -1298183838;
assign addr[59205] = -1282899464;
assign addr[59206] = -1267513365;
assign addr[59207] = -1252026760;
assign addr[59208] = -1236440877;
assign addr[59209] = -1220756951;
assign addr[59210] = -1204976227;
assign addr[59211] = -1189099956;
assign addr[59212] = -1173129396;
assign addr[59213] = -1157065814;
assign addr[59214] = -1140910484;
assign addr[59215] = -1124664687;
assign addr[59216] = -1108329711;
assign addr[59217] = -1091906851;
assign addr[59218] = -1075397409;
assign addr[59219] = -1058802695;
assign addr[59220] = -1042124025;
assign addr[59221] = -1025362720;
assign addr[59222] = -1008520110;
assign addr[59223] = -991597531;
assign addr[59224] = -974596324;
assign addr[59225] = -957517838;
assign addr[59226] = -940363427;
assign addr[59227] = -923134450;
assign addr[59228] = -905832274;
assign addr[59229] = -888458272;
assign addr[59230] = -871013820;
assign addr[59231] = -853500302;
assign addr[59232] = -835919107;
assign addr[59233] = -818271628;
assign addr[59234] = -800559266;
assign addr[59235] = -782783424;
assign addr[59236] = -764945512;
assign addr[59237] = -747046944;
assign addr[59238] = -729089140;
assign addr[59239] = -711073524;
assign addr[59240] = -693001525;
assign addr[59241] = -674874574;
assign addr[59242] = -656694110;
assign addr[59243] = -638461574;
assign addr[59244] = -620178412;
assign addr[59245] = -601846074;
assign addr[59246] = -583466013;
assign addr[59247] = -565039687;
assign addr[59248] = -546568556;
assign addr[59249] = -528054086;
assign addr[59250] = -509497745;
assign addr[59251] = -490901003;
assign addr[59252] = -472265336;
assign addr[59253] = -453592221;
assign addr[59254] = -434883140;
assign addr[59255] = -416139574;
assign addr[59256] = -397363011;
assign addr[59257] = -378554940;
assign addr[59258] = -359716852;
assign addr[59259] = -340850240;
assign addr[59260] = -321956601;
assign addr[59261] = -303037433;
assign addr[59262] = -284094236;
assign addr[59263] = -265128512;
assign addr[59264] = -246141764;
assign addr[59265] = -227135500;
assign addr[59266] = -208111224;
assign addr[59267] = -189070447;
assign addr[59268] = -170014678;
assign addr[59269] = -150945428;
assign addr[59270] = -131864208;
assign addr[59271] = -112772533;
assign addr[59272] = -93671915;
assign addr[59273] = -74563870;
assign addr[59274] = -55449912;
assign addr[59275] = -36331557;
assign addr[59276] = -17210322;
assign addr[59277] = 1912278;
assign addr[59278] = 21034727;
assign addr[59279] = 40155507;
assign addr[59280] = 59273104;
assign addr[59281] = 78386000;
assign addr[59282] = 97492681;
assign addr[59283] = 116591632;
assign addr[59284] = 135681337;
assign addr[59285] = 154760284;
assign addr[59286] = 173826959;
assign addr[59287] = 192879850;
assign addr[59288] = 211917448;
assign addr[59289] = 230938242;
assign addr[59290] = 249940723;
assign addr[59291] = 268923386;
assign addr[59292] = 287884725;
assign addr[59293] = 306823237;
assign addr[59294] = 325737419;
assign addr[59295] = 344625773;
assign addr[59296] = 363486799;
assign addr[59297] = 382319004;
assign addr[59298] = 401120892;
assign addr[59299] = 419890975;
assign addr[59300] = 438627762;
assign addr[59301] = 457329769;
assign addr[59302] = 475995513;
assign addr[59303] = 494623513;
assign addr[59304] = 513212292;
assign addr[59305] = 531760377;
assign addr[59306] = 550266296;
assign addr[59307] = 568728583;
assign addr[59308] = 587145773;
assign addr[59309] = 605516406;
assign addr[59310] = 623839025;
assign addr[59311] = 642112178;
assign addr[59312] = 660334415;
assign addr[59313] = 678504291;
assign addr[59314] = 696620367;
assign addr[59315] = 714681204;
assign addr[59316] = 732685372;
assign addr[59317] = 750631442;
assign addr[59318] = 768517992;
assign addr[59319] = 786343603;
assign addr[59320] = 804106861;
assign addr[59321] = 821806359;
assign addr[59322] = 839440693;
assign addr[59323] = 857008464;
assign addr[59324] = 874508280;
assign addr[59325] = 891938752;
assign addr[59326] = 909298500;
assign addr[59327] = 926586145;
assign addr[59328] = 943800318;
assign addr[59329] = 960939653;
assign addr[59330] = 978002791;
assign addr[59331] = 994988380;
assign addr[59332] = 1011895073;
assign addr[59333] = 1028721528;
assign addr[59334] = 1045466412;
assign addr[59335] = 1062128397;
assign addr[59336] = 1078706161;
assign addr[59337] = 1095198391;
assign addr[59338] = 1111603778;
assign addr[59339] = 1127921022;
assign addr[59340] = 1144148829;
assign addr[59341] = 1160285911;
assign addr[59342] = 1176330990;
assign addr[59343] = 1192282793;
assign addr[59344] = 1208140056;
assign addr[59345] = 1223901520;
assign addr[59346] = 1239565936;
assign addr[59347] = 1255132063;
assign addr[59348] = 1270598665;
assign addr[59349] = 1285964516;
assign addr[59350] = 1301228398;
assign addr[59351] = 1316389101;
assign addr[59352] = 1331445422;
assign addr[59353] = 1346396168;
assign addr[59354] = 1361240152;
assign addr[59355] = 1375976199;
assign addr[59356] = 1390603139;
assign addr[59357] = 1405119813;
assign addr[59358] = 1419525069;
assign addr[59359] = 1433817766;
assign addr[59360] = 1447996770;
assign addr[59361] = 1462060956;
assign addr[59362] = 1476009210;
assign addr[59363] = 1489840425;
assign addr[59364] = 1503553506;
assign addr[59365] = 1517147363;
assign addr[59366] = 1530620920;
assign addr[59367] = 1543973108;
assign addr[59368] = 1557202869;
assign addr[59369] = 1570309153;
assign addr[59370] = 1583290921;
assign addr[59371] = 1596147143;
assign addr[59372] = 1608876801;
assign addr[59373] = 1621478885;
assign addr[59374] = 1633952396;
assign addr[59375] = 1646296344;
assign addr[59376] = 1658509750;
assign addr[59377] = 1670591647;
assign addr[59378] = 1682541077;
assign addr[59379] = 1694357091;
assign addr[59380] = 1706038753;
assign addr[59381] = 1717585136;
assign addr[59382] = 1728995326;
assign addr[59383] = 1740268417;
assign addr[59384] = 1751403515;
assign addr[59385] = 1762399737;
assign addr[59386] = 1773256212;
assign addr[59387] = 1783972079;
assign addr[59388] = 1794546487;
assign addr[59389] = 1804978599;
assign addr[59390] = 1815267588;
assign addr[59391] = 1825412636;
assign addr[59392] = 1835412941;
assign addr[59393] = 1845267708;
assign addr[59394] = 1854976157;
assign addr[59395] = 1864537518;
assign addr[59396] = 1873951032;
assign addr[59397] = 1883215953;
assign addr[59398] = 1892331547;
assign addr[59399] = 1901297091;
assign addr[59400] = 1910111873;
assign addr[59401] = 1918775195;
assign addr[59402] = 1927286370;
assign addr[59403] = 1935644723;
assign addr[59404] = 1943849591;
assign addr[59405] = 1951900324;
assign addr[59406] = 1959796283;
assign addr[59407] = 1967536842;
assign addr[59408] = 1975121388;
assign addr[59409] = 1982549318;
assign addr[59410] = 1989820044;
assign addr[59411] = 1996932990;
assign addr[59412] = 2003887591;
assign addr[59413] = 2010683297;
assign addr[59414] = 2017319567;
assign addr[59415] = 2023795876;
assign addr[59416] = 2030111710;
assign addr[59417] = 2036266570;
assign addr[59418] = 2042259965;
assign addr[59419] = 2048091422;
assign addr[59420] = 2053760478;
assign addr[59421] = 2059266683;
assign addr[59422] = 2064609600;
assign addr[59423] = 2069788807;
assign addr[59424] = 2074803892;
assign addr[59425] = 2079654458;
assign addr[59426] = 2084340120;
assign addr[59427] = 2088860507;
assign addr[59428] = 2093215260;
assign addr[59429] = 2097404033;
assign addr[59430] = 2101426496;
assign addr[59431] = 2105282327;
assign addr[59432] = 2108971223;
assign addr[59433] = 2112492891;
assign addr[59434] = 2115847050;
assign addr[59435] = 2119033436;
assign addr[59436] = 2122051796;
assign addr[59437] = 2124901890;
assign addr[59438] = 2127583492;
assign addr[59439] = 2130096389;
assign addr[59440] = 2132440383;
assign addr[59441] = 2134615288;
assign addr[59442] = 2136620930;
assign addr[59443] = 2138457152;
assign addr[59444] = 2140123807;
assign addr[59445] = 2141620763;
assign addr[59446] = 2142947902;
assign addr[59447] = 2144105118;
assign addr[59448] = 2145092320;
assign addr[59449] = 2145909429;
assign addr[59450] = 2146556380;
assign addr[59451] = 2147033123;
assign addr[59452] = 2147339619;
assign addr[59453] = 2147475844;
assign addr[59454] = 2147441787;
assign addr[59455] = 2147237452;
assign addr[59456] = 2146862854;
assign addr[59457] = 2146318022;
assign addr[59458] = 2145603001;
assign addr[59459] = 2144717846;
assign addr[59460] = 2143662628;
assign addr[59461] = 2142437431;
assign addr[59462] = 2141042352;
assign addr[59463] = 2139477502;
assign addr[59464] = 2137743003;
assign addr[59465] = 2135838995;
assign addr[59466] = 2133765628;
assign addr[59467] = 2131523066;
assign addr[59468] = 2129111488;
assign addr[59469] = 2126531084;
assign addr[59470] = 2123782059;
assign addr[59471] = 2120864631;
assign addr[59472] = 2117779031;
assign addr[59473] = 2114525505;
assign addr[59474] = 2111104309;
assign addr[59475] = 2107515716;
assign addr[59476] = 2103760010;
assign addr[59477] = 2099837489;
assign addr[59478] = 2095748463;
assign addr[59479] = 2091493257;
assign addr[59480] = 2087072209;
assign addr[59481] = 2082485668;
assign addr[59482] = 2077733999;
assign addr[59483] = 2072817579;
assign addr[59484] = 2067736796;
assign addr[59485] = 2062492055;
assign addr[59486] = 2057083771;
assign addr[59487] = 2051512372;
assign addr[59488] = 2045778302;
assign addr[59489] = 2039882013;
assign addr[59490] = 2033823974;
assign addr[59491] = 2027604666;
assign addr[59492] = 2021224581;
assign addr[59493] = 2014684225;
assign addr[59494] = 2007984117;
assign addr[59495] = 2001124788;
assign addr[59496] = 1994106782;
assign addr[59497] = 1986930656;
assign addr[59498] = 1979596978;
assign addr[59499] = 1972106330;
assign addr[59500] = 1964459306;
assign addr[59501] = 1956656513;
assign addr[59502] = 1948698568;
assign addr[59503] = 1940586104;
assign addr[59504] = 1932319763;
assign addr[59505] = 1923900201;
assign addr[59506] = 1915328086;
assign addr[59507] = 1906604097;
assign addr[59508] = 1897728925;
assign addr[59509] = 1888703276;
assign addr[59510] = 1879527863;
assign addr[59511] = 1870203416;
assign addr[59512] = 1860730673;
assign addr[59513] = 1851110385;
assign addr[59514] = 1841343316;
assign addr[59515] = 1831430239;
assign addr[59516] = 1821371941;
assign addr[59517] = 1811169220;
assign addr[59518] = 1800822883;
assign addr[59519] = 1790333753;
assign addr[59520] = 1779702660;
assign addr[59521] = 1768930447;
assign addr[59522] = 1758017969;
assign addr[59523] = 1746966091;
assign addr[59524] = 1735775690;
assign addr[59525] = 1724447652;
assign addr[59526] = 1712982875;
assign addr[59527] = 1701382270;
assign addr[59528] = 1689646755;
assign addr[59529] = 1677777262;
assign addr[59530] = 1665774731;
assign addr[59531] = 1653640115;
assign addr[59532] = 1641374375;
assign addr[59533] = 1628978484;
assign addr[59534] = 1616453425;
assign addr[59535] = 1603800191;
assign addr[59536] = 1591019785;
assign addr[59537] = 1578113222;
assign addr[59538] = 1565081523;
assign addr[59539] = 1551925723;
assign addr[59540] = 1538646865;
assign addr[59541] = 1525246002;
assign addr[59542] = 1511724196;
assign addr[59543] = 1498082520;
assign addr[59544] = 1484322054;
assign addr[59545] = 1470443891;
assign addr[59546] = 1456449131;
assign addr[59547] = 1442338884;
assign addr[59548] = 1428114267;
assign addr[59549] = 1413776410;
assign addr[59550] = 1399326449;
assign addr[59551] = 1384765530;
assign addr[59552] = 1370094808;
assign addr[59553] = 1355315445;
assign addr[59554] = 1340428615;
assign addr[59555] = 1325435496;
assign addr[59556] = 1310337279;
assign addr[59557] = 1295135159;
assign addr[59558] = 1279830344;
assign addr[59559] = 1264424045;
assign addr[59560] = 1248917486;
assign addr[59561] = 1233311895;
assign addr[59562] = 1217608510;
assign addr[59563] = 1201808576;
assign addr[59564] = 1185913346;
assign addr[59565] = 1169924081;
assign addr[59566] = 1153842047;
assign addr[59567] = 1137668521;
assign addr[59568] = 1121404785;
assign addr[59569] = 1105052128;
assign addr[59570] = 1088611847;
assign addr[59571] = 1072085246;
assign addr[59572] = 1055473635;
assign addr[59573] = 1038778332;
assign addr[59574] = 1022000660;
assign addr[59575] = 1005141949;
assign addr[59576] = 988203537;
assign addr[59577] = 971186766;
assign addr[59578] = 954092986;
assign addr[59579] = 936923553;
assign addr[59580] = 919679827;
assign addr[59581] = 902363176;
assign addr[59582] = 884974973;
assign addr[59583] = 867516597;
assign addr[59584] = 849989433;
assign addr[59585] = 832394869;
assign addr[59586] = 814734301;
assign addr[59587] = 797009130;
assign addr[59588] = 779220762;
assign addr[59589] = 761370605;
assign addr[59590] = 743460077;
assign addr[59591] = 725490597;
assign addr[59592] = 707463589;
assign addr[59593] = 689380485;
assign addr[59594] = 671242716;
assign addr[59595] = 653051723;
assign addr[59596] = 634808946;
assign addr[59597] = 616515832;
assign addr[59598] = 598173833;
assign addr[59599] = 579784402;
assign addr[59600] = 561348998;
assign addr[59601] = 542869083;
assign addr[59602] = 524346121;
assign addr[59603] = 505781581;
assign addr[59604] = 487176937;
assign addr[59605] = 468533662;
assign addr[59606] = 449853235;
assign addr[59607] = 431137138;
assign addr[59608] = 412386854;
assign addr[59609] = 393603870;
assign addr[59610] = 374789676;
assign addr[59611] = 355945764;
assign addr[59612] = 337073627;
assign addr[59613] = 318174762;
assign addr[59614] = 299250668;
assign addr[59615] = 280302845;
assign addr[59616] = 261332796;
assign addr[59617] = 242342025;
assign addr[59618] = 223332037;
assign addr[59619] = 204304341;
assign addr[59620] = 185260444;
assign addr[59621] = 166201858;
assign addr[59622] = 147130093;
assign addr[59623] = 128046661;
assign addr[59624] = 108953076;
assign addr[59625] = 89850852;
assign addr[59626] = 70741503;
assign addr[59627] = 51626544;
assign addr[59628] = 32507492;
assign addr[59629] = 13385863;
assign addr[59630] = -5736829;
assign addr[59631] = -24859065;
assign addr[59632] = -43979330;
assign addr[59633] = -63096108;
assign addr[59634] = -82207882;
assign addr[59635] = -101313138;
assign addr[59636] = -120410361;
assign addr[59637] = -139498035;
assign addr[59638] = -158574649;
assign addr[59639] = -177638688;
assign addr[59640] = -196688642;
assign addr[59641] = -215722999;
assign addr[59642] = -234740251;
assign addr[59643] = -253738890;
assign addr[59644] = -272717408;
assign addr[59645] = -291674302;
assign addr[59646] = -310608068;
assign addr[59647] = -329517204;
assign addr[59648] = -348400212;
assign addr[59649] = -367255594;
assign addr[59650] = -386081854;
assign addr[59651] = -404877501;
assign addr[59652] = -423641043;
assign addr[59653] = -442370993;
assign addr[59654] = -461065866;
assign addr[59655] = -479724180;
assign addr[59656] = -498344454;
assign addr[59657] = -516925212;
assign addr[59658] = -535464981;
assign addr[59659] = -553962291;
assign addr[59660] = -572415676;
assign addr[59661] = -590823671;
assign addr[59662] = -609184818;
assign addr[59663] = -627497660;
assign addr[59664] = -645760745;
assign addr[59665] = -663972625;
assign addr[59666] = -682131857;
assign addr[59667] = -700236999;
assign addr[59668] = -718286617;
assign addr[59669] = -736279279;
assign addr[59670] = -754213559;
assign addr[59671] = -772088034;
assign addr[59672] = -789901288;
assign addr[59673] = -807651907;
assign addr[59674] = -825338484;
assign addr[59675] = -842959617;
assign addr[59676] = -860513908;
assign addr[59677] = -877999966;
assign addr[59678] = -895416404;
assign addr[59679] = -912761841;
assign addr[59680] = -930034901;
assign addr[59681] = -947234215;
assign addr[59682] = -964358420;
assign addr[59683] = -981406156;
assign addr[59684] = -998376073;
assign addr[59685] = -1015266825;
assign addr[59686] = -1032077073;
assign addr[59687] = -1048805483;
assign addr[59688] = -1065450729;
assign addr[59689] = -1082011492;
assign addr[59690] = -1098486458;
assign addr[59691] = -1114874320;
assign addr[59692] = -1131173780;
assign addr[59693] = -1147383544;
assign addr[59694] = -1163502328;
assign addr[59695] = -1179528853;
assign addr[59696] = -1195461849;
assign addr[59697] = -1211300053;
assign addr[59698] = -1227042207;
assign addr[59699] = -1242687064;
assign addr[59700] = -1258233384;
assign addr[59701] = -1273679934;
assign addr[59702] = -1289025489;
assign addr[59703] = -1304268832;
assign addr[59704] = -1319408754;
assign addr[59705] = -1334444055;
assign addr[59706] = -1349373543;
assign addr[59707] = -1364196034;
assign addr[59708] = -1378910353;
assign addr[59709] = -1393515332;
assign addr[59710] = -1408009814;
assign addr[59711] = -1422392650;
assign addr[59712] = -1436662698;
assign addr[59713] = -1450818828;
assign addr[59714] = -1464859917;
assign addr[59715] = -1478784851;
assign addr[59716] = -1492592527;
assign addr[59717] = -1506281850;
assign addr[59718] = -1519851733;
assign addr[59719] = -1533301101;
assign addr[59720] = -1546628888;
assign addr[59721] = -1559834037;
assign addr[59722] = -1572915501;
assign addr[59723] = -1585872242;
assign addr[59724] = -1598703233;
assign addr[59725] = -1611407456;
assign addr[59726] = -1623983905;
assign addr[59727] = -1636431582;
assign addr[59728] = -1648749499;
assign addr[59729] = -1660936681;
assign addr[59730] = -1672992161;
assign addr[59731] = -1684914983;
assign addr[59732] = -1696704201;
assign addr[59733] = -1708358881;
assign addr[59734] = -1719878099;
assign addr[59735] = -1731260941;
assign addr[59736] = -1742506504;
assign addr[59737] = -1753613897;
assign addr[59738] = -1764582240;
assign addr[59739] = -1775410662;
assign addr[59740] = -1786098304;
assign addr[59741] = -1796644320;
assign addr[59742] = -1807047873;
assign addr[59743] = -1817308138;
assign addr[59744] = -1827424302;
assign addr[59745] = -1837395562;
assign addr[59746] = -1847221128;
assign addr[59747] = -1856900221;
assign addr[59748] = -1866432072;
assign addr[59749] = -1875815927;
assign addr[59750] = -1885051042;
assign addr[59751] = -1894136683;
assign addr[59752] = -1903072131;
assign addr[59753] = -1911856677;
assign addr[59754] = -1920489624;
assign addr[59755] = -1928970288;
assign addr[59756] = -1937297997;
assign addr[59757] = -1945472089;
assign addr[59758] = -1953491918;
assign addr[59759] = -1961356847;
assign addr[59760] = -1969066252;
assign addr[59761] = -1976619522;
assign addr[59762] = -1984016058;
assign addr[59763] = -1991255274;
assign addr[59764] = -1998336596;
assign addr[59765] = -2005259462;
assign addr[59766] = -2012023322;
assign addr[59767] = -2018627642;
assign addr[59768] = -2025071897;
assign addr[59769] = -2031355576;
assign addr[59770] = -2037478181;
assign addr[59771] = -2043439226;
assign addr[59772] = -2049238240;
assign addr[59773] = -2054874761;
assign addr[59774] = -2060348343;
assign addr[59775] = -2065658552;
assign addr[59776] = -2070804967;
assign addr[59777] = -2075787180;
assign addr[59778] = -2080604795;
assign addr[59779] = -2085257431;
assign addr[59780] = -2089744719;
assign addr[59781] = -2094066304;
assign addr[59782] = -2098221841;
assign addr[59783] = -2102211002;
assign addr[59784] = -2106033471;
assign addr[59785] = -2109688944;
assign addr[59786] = -2113177132;
assign addr[59787] = -2116497758;
assign addr[59788] = -2119650558;
assign addr[59789] = -2122635283;
assign addr[59790] = -2125451696;
assign addr[59791] = -2128099574;
assign addr[59792] = -2130578706;
assign addr[59793] = -2132888897;
assign addr[59794] = -2135029962;
assign addr[59795] = -2137001733;
assign addr[59796] = -2138804053;
assign addr[59797] = -2140436778;
assign addr[59798] = -2141899780;
assign addr[59799] = -2143192942;
assign addr[59800] = -2144316162;
assign addr[59801] = -2145269351;
assign addr[59802] = -2146052433;
assign addr[59803] = -2146665347;
assign addr[59804] = -2147108043;
assign addr[59805] = -2147380486;
assign addr[59806] = -2147482655;
assign addr[59807] = -2147414542;
assign addr[59808] = -2147176152;
assign addr[59809] = -2146767505;
assign addr[59810] = -2146188631;
assign addr[59811] = -2145439578;
assign addr[59812] = -2144520405;
assign addr[59813] = -2143431184;
assign addr[59814] = -2142172003;
assign addr[59815] = -2140742960;
assign addr[59816] = -2139144169;
assign addr[59817] = -2137375758;
assign addr[59818] = -2135437865;
assign addr[59819] = -2133330646;
assign addr[59820] = -2131054266;
assign addr[59821] = -2128608907;
assign addr[59822] = -2125994762;
assign addr[59823] = -2123212038;
assign addr[59824] = -2120260957;
assign addr[59825] = -2117141752;
assign addr[59826] = -2113854671;
assign addr[59827] = -2110399974;
assign addr[59828] = -2106777935;
assign addr[59829] = -2102988841;
assign addr[59830] = -2099032994;
assign addr[59831] = -2094910706;
assign addr[59832] = -2090622304;
assign addr[59833] = -2086168128;
assign addr[59834] = -2081548533;
assign addr[59835] = -2076763883;
assign addr[59836] = -2071814558;
assign addr[59837] = -2066700952;
assign addr[59838] = -2061423468;
assign addr[59839] = -2055982526;
assign addr[59840] = -2050378558;
assign addr[59841] = -2044612007;
assign addr[59842] = -2038683330;
assign addr[59843] = -2032592999;
assign addr[59844] = -2026341495;
assign addr[59845] = -2019929315;
assign addr[59846] = -2013356967;
assign addr[59847] = -2006624971;
assign addr[59848] = -1999733863;
assign addr[59849] = -1992684188;
assign addr[59850] = -1985476506;
assign addr[59851] = -1978111387;
assign addr[59852] = -1970589416;
assign addr[59853] = -1962911189;
assign addr[59854] = -1955077316;
assign addr[59855] = -1947088417;
assign addr[59856] = -1938945125;
assign addr[59857] = -1930648088;
assign addr[59858] = -1922197961;
assign addr[59859] = -1913595416;
assign addr[59860] = -1904841135;
assign addr[59861] = -1895935811;
assign addr[59862] = -1886880151;
assign addr[59863] = -1877674873;
assign addr[59864] = -1868320707;
assign addr[59865] = -1858818395;
assign addr[59866] = -1849168689;
assign addr[59867] = -1839372356;
assign addr[59868] = -1829430172;
assign addr[59869] = -1819342925;
assign addr[59870] = -1809111415;
assign addr[59871] = -1798736454;
assign addr[59872] = -1788218865;
assign addr[59873] = -1777559480;
assign addr[59874] = -1766759146;
assign addr[59875] = -1755818718;
assign addr[59876] = -1744739065;
assign addr[59877] = -1733521064;
assign addr[59878] = -1722165606;
assign addr[59879] = -1710673591;
assign addr[59880] = -1699045930;
assign addr[59881] = -1687283545;
assign addr[59882] = -1675387369;
assign addr[59883] = -1663358344;
assign addr[59884] = -1651197426;
assign addr[59885] = -1638905577;
assign addr[59886] = -1626483774;
assign addr[59887] = -1613933000;
assign addr[59888] = -1601254251;
assign addr[59889] = -1588448533;
assign addr[59890] = -1575516860;
assign addr[59891] = -1562460258;
assign addr[59892] = -1549279763;
assign addr[59893] = -1535976419;
assign addr[59894] = -1522551282;
assign addr[59895] = -1509005416;
assign addr[59896] = -1495339895;
assign addr[59897] = -1481555802;
assign addr[59898] = -1467654232;
assign addr[59899] = -1453636285;
assign addr[59900] = -1439503074;
assign addr[59901] = -1425255719;
assign addr[59902] = -1410895350;
assign addr[59903] = -1396423105;
assign addr[59904] = -1381840133;
assign addr[59905] = -1367147589;
assign addr[59906] = -1352346639;
assign addr[59907] = -1337438456;
assign addr[59908] = -1322424222;
assign addr[59909] = -1307305128;
assign addr[59910] = -1292082373;
assign addr[59911] = -1276757164;
assign addr[59912] = -1261330715;
assign addr[59913] = -1245804251;
assign addr[59914] = -1230179002;
assign addr[59915] = -1214456207;
assign addr[59916] = -1198637114;
assign addr[59917] = -1182722976;
assign addr[59918] = -1166715055;
assign addr[59919] = -1150614620;
assign addr[59920] = -1134422949;
assign addr[59921] = -1118141326;
assign addr[59922] = -1101771040;
assign addr[59923] = -1085313391;
assign addr[59924] = -1068769683;
assign addr[59925] = -1052141228;
assign addr[59926] = -1035429345;
assign addr[59927] = -1018635358;
assign addr[59928] = -1001760600;
assign addr[59929] = -984806408;
assign addr[59930] = -967774128;
assign addr[59931] = -950665109;
assign addr[59932] = -933480707;
assign addr[59933] = -916222287;
assign addr[59934] = -898891215;
assign addr[59935] = -881488868;
assign addr[59936] = -864016623;
assign addr[59937] = -846475867;
assign addr[59938] = -828867991;
assign addr[59939] = -811194391;
assign addr[59940] = -793456467;
assign addr[59941] = -775655628;
assign addr[59942] = -757793284;
assign addr[59943] = -739870851;
assign addr[59944] = -721889752;
assign addr[59945] = -703851410;
assign addr[59946] = -685757258;
assign addr[59947] = -667608730;
assign addr[59948] = -649407264;
assign addr[59949] = -631154304;
assign addr[59950] = -612851297;
assign addr[59951] = -594499695;
assign addr[59952] = -576100953;
assign addr[59953] = -557656529;
assign addr[59954] = -539167887;
assign addr[59955] = -520636492;
assign addr[59956] = -502063814;
assign addr[59957] = -483451325;
assign addr[59958] = -464800501;
assign addr[59959] = -446112822;
assign addr[59960] = -427389768;
assign addr[59961] = -408632825;
assign addr[59962] = -389843480;
assign addr[59963] = -371023223;
assign addr[59964] = -352173546;
assign addr[59965] = -333295944;
assign addr[59966] = -314391913;
assign addr[59967] = -295462954;
assign addr[59968] = -276510565;
assign addr[59969] = -257536251;
assign addr[59970] = -238541516;
assign addr[59971] = -219527866;
assign addr[59972] = -200496809;
assign addr[59973] = -181449854;
assign addr[59974] = -162388511;
assign addr[59975] = -143314291;
assign addr[59976] = -124228708;
assign addr[59977] = -105133274;
assign addr[59978] = -86029503;
assign addr[59979] = -66918911;
assign addr[59980] = -47803013;
assign addr[59981] = -28683324;
assign addr[59982] = -9561361;
assign addr[59983] = 9561361;
assign addr[59984] = 28683324;
assign addr[59985] = 47803013;
assign addr[59986] = 66918911;
assign addr[59987] = 86029503;
assign addr[59988] = 105133274;
assign addr[59989] = 124228708;
assign addr[59990] = 143314291;
assign addr[59991] = 162388511;
assign addr[59992] = 181449854;
assign addr[59993] = 200496809;
assign addr[59994] = 219527866;
assign addr[59995] = 238541516;
assign addr[59996] = 257536251;
assign addr[59997] = 276510565;
assign addr[59998] = 295462953;
assign addr[59999] = 314391913;
assign addr[60000] = 333295944;
assign addr[60001] = 352173546;
assign addr[60002] = 371023223;
assign addr[60003] = 389843480;
assign addr[60004] = 408632825;
assign addr[60005] = 427389768;
assign addr[60006] = 446112822;
assign addr[60007] = 464800501;
assign addr[60008] = 483451325;
assign addr[60009] = 502063814;
assign addr[60010] = 520636492;
assign addr[60011] = 539167887;
assign addr[60012] = 557656529;
assign addr[60013] = 576100953;
assign addr[60014] = 594499695;
assign addr[60015] = 612851297;
assign addr[60016] = 631154304;
assign addr[60017] = 649407264;
assign addr[60018] = 667608730;
assign addr[60019] = 685757258;
assign addr[60020] = 703851410;
assign addr[60021] = 721889752;
assign addr[60022] = 739870851;
assign addr[60023] = 757793284;
assign addr[60024] = 775655628;
assign addr[60025] = 793456467;
assign addr[60026] = 811194391;
assign addr[60027] = 828867991;
assign addr[60028] = 846475867;
assign addr[60029] = 864016623;
assign addr[60030] = 881488868;
assign addr[60031] = 898891215;
assign addr[60032] = 916222287;
assign addr[60033] = 933480707;
assign addr[60034] = 950665109;
assign addr[60035] = 967774128;
assign addr[60036] = 984806408;
assign addr[60037] = 1001760600;
assign addr[60038] = 1018635358;
assign addr[60039] = 1035429345;
assign addr[60040] = 1052141228;
assign addr[60041] = 1068769683;
assign addr[60042] = 1085313391;
assign addr[60043] = 1101771040;
assign addr[60044] = 1118141326;
assign addr[60045] = 1134422949;
assign addr[60046] = 1150614620;
assign addr[60047] = 1166715055;
assign addr[60048] = 1182722976;
assign addr[60049] = 1198637114;
assign addr[60050] = 1214456207;
assign addr[60051] = 1230179002;
assign addr[60052] = 1245804251;
assign addr[60053] = 1261330715;
assign addr[60054] = 1276757164;
assign addr[60055] = 1292082373;
assign addr[60056] = 1307305128;
assign addr[60057] = 1322424222;
assign addr[60058] = 1337438456;
assign addr[60059] = 1352346639;
assign addr[60060] = 1367147589;
assign addr[60061] = 1381840133;
assign addr[60062] = 1396423105;
assign addr[60063] = 1410895350;
assign addr[60064] = 1425255719;
assign addr[60065] = 1439503074;
assign addr[60066] = 1453636285;
assign addr[60067] = 1467654232;
assign addr[60068] = 1481555802;
assign addr[60069] = 1495339895;
assign addr[60070] = 1509005416;
assign addr[60071] = 1522551282;
assign addr[60072] = 1535976419;
assign addr[60073] = 1549279763;
assign addr[60074] = 1562460258;
assign addr[60075] = 1575516860;
assign addr[60076] = 1588448533;
assign addr[60077] = 1601254251;
assign addr[60078] = 1613933000;
assign addr[60079] = 1626483774;
assign addr[60080] = 1638905577;
assign addr[60081] = 1651197426;
assign addr[60082] = 1663358344;
assign addr[60083] = 1675387369;
assign addr[60084] = 1687283545;
assign addr[60085] = 1699045930;
assign addr[60086] = 1710673591;
assign addr[60087] = 1722165606;
assign addr[60088] = 1733521064;
assign addr[60089] = 1744739065;
assign addr[60090] = 1755818718;
assign addr[60091] = 1766759146;
assign addr[60092] = 1777559480;
assign addr[60093] = 1788218865;
assign addr[60094] = 1798736454;
assign addr[60095] = 1809111415;
assign addr[60096] = 1819342925;
assign addr[60097] = 1829430172;
assign addr[60098] = 1839372356;
assign addr[60099] = 1849168689;
assign addr[60100] = 1858818395;
assign addr[60101] = 1868320707;
assign addr[60102] = 1877674873;
assign addr[60103] = 1886880151;
assign addr[60104] = 1895935811;
assign addr[60105] = 1904841135;
assign addr[60106] = 1913595416;
assign addr[60107] = 1922197961;
assign addr[60108] = 1930648088;
assign addr[60109] = 1938945125;
assign addr[60110] = 1947088417;
assign addr[60111] = 1955077316;
assign addr[60112] = 1962911189;
assign addr[60113] = 1970589416;
assign addr[60114] = 1978111387;
assign addr[60115] = 1985476506;
assign addr[60116] = 1992684188;
assign addr[60117] = 1999733863;
assign addr[60118] = 2006624971;
assign addr[60119] = 2013356967;
assign addr[60120] = 2019929315;
assign addr[60121] = 2026341495;
assign addr[60122] = 2032592999;
assign addr[60123] = 2038683330;
assign addr[60124] = 2044612007;
assign addr[60125] = 2050378558;
assign addr[60126] = 2055982526;
assign addr[60127] = 2061423468;
assign addr[60128] = 2066700952;
assign addr[60129] = 2071814558;
assign addr[60130] = 2076763883;
assign addr[60131] = 2081548533;
assign addr[60132] = 2086168128;
assign addr[60133] = 2090622304;
assign addr[60134] = 2094910706;
assign addr[60135] = 2099032994;
assign addr[60136] = 2102988841;
assign addr[60137] = 2106777935;
assign addr[60138] = 2110399974;
assign addr[60139] = 2113854671;
assign addr[60140] = 2117141752;
assign addr[60141] = 2120260957;
assign addr[60142] = 2123212038;
assign addr[60143] = 2125994762;
assign addr[60144] = 2128608907;
assign addr[60145] = 2131054266;
assign addr[60146] = 2133330646;
assign addr[60147] = 2135437865;
assign addr[60148] = 2137375758;
assign addr[60149] = 2139144169;
assign addr[60150] = 2140742960;
assign addr[60151] = 2142172003;
assign addr[60152] = 2143431184;
assign addr[60153] = 2144520405;
assign addr[60154] = 2145439578;
assign addr[60155] = 2146188631;
assign addr[60156] = 2146767505;
assign addr[60157] = 2147176152;
assign addr[60158] = 2147414542;
assign addr[60159] = 2147482655;
assign addr[60160] = 2147380486;
assign addr[60161] = 2147108043;
assign addr[60162] = 2146665347;
assign addr[60163] = 2146052433;
assign addr[60164] = 2145269351;
assign addr[60165] = 2144316162;
assign addr[60166] = 2143192942;
assign addr[60167] = 2141899780;
assign addr[60168] = 2140436778;
assign addr[60169] = 2138804053;
assign addr[60170] = 2137001733;
assign addr[60171] = 2135029962;
assign addr[60172] = 2132888897;
assign addr[60173] = 2130578706;
assign addr[60174] = 2128099574;
assign addr[60175] = 2125451696;
assign addr[60176] = 2122635283;
assign addr[60177] = 2119650558;
assign addr[60178] = 2116497758;
assign addr[60179] = 2113177132;
assign addr[60180] = 2109688944;
assign addr[60181] = 2106033471;
assign addr[60182] = 2102211002;
assign addr[60183] = 2098221841;
assign addr[60184] = 2094066304;
assign addr[60185] = 2089744719;
assign addr[60186] = 2085257431;
assign addr[60187] = 2080604795;
assign addr[60188] = 2075787180;
assign addr[60189] = 2070804967;
assign addr[60190] = 2065658552;
assign addr[60191] = 2060348343;
assign addr[60192] = 2054874761;
assign addr[60193] = 2049238240;
assign addr[60194] = 2043439226;
assign addr[60195] = 2037478181;
assign addr[60196] = 2031355576;
assign addr[60197] = 2025071897;
assign addr[60198] = 2018627642;
assign addr[60199] = 2012023322;
assign addr[60200] = 2005259462;
assign addr[60201] = 1998336596;
assign addr[60202] = 1991255274;
assign addr[60203] = 1984016058;
assign addr[60204] = 1976619522;
assign addr[60205] = 1969066252;
assign addr[60206] = 1961356847;
assign addr[60207] = 1953491918;
assign addr[60208] = 1945472089;
assign addr[60209] = 1937297997;
assign addr[60210] = 1928970288;
assign addr[60211] = 1920489624;
assign addr[60212] = 1911856677;
assign addr[60213] = 1903072131;
assign addr[60214] = 1894136683;
assign addr[60215] = 1885051042;
assign addr[60216] = 1875815927;
assign addr[60217] = 1866432072;
assign addr[60218] = 1856900221;
assign addr[60219] = 1847221128;
assign addr[60220] = 1837395562;
assign addr[60221] = 1827424302;
assign addr[60222] = 1817308138;
assign addr[60223] = 1807047873;
assign addr[60224] = 1796644320;
assign addr[60225] = 1786098304;
assign addr[60226] = 1775410662;
assign addr[60227] = 1764582240;
assign addr[60228] = 1753613897;
assign addr[60229] = 1742506504;
assign addr[60230] = 1731260941;
assign addr[60231] = 1719878099;
assign addr[60232] = 1708358881;
assign addr[60233] = 1696704201;
assign addr[60234] = 1684914983;
assign addr[60235] = 1672992161;
assign addr[60236] = 1660936681;
assign addr[60237] = 1648749499;
assign addr[60238] = 1636431582;
assign addr[60239] = 1623983905;
assign addr[60240] = 1611407456;
assign addr[60241] = 1598703233;
assign addr[60242] = 1585872242;
assign addr[60243] = 1572915501;
assign addr[60244] = 1559834037;
assign addr[60245] = 1546628888;
assign addr[60246] = 1533301101;
assign addr[60247] = 1519851733;
assign addr[60248] = 1506281850;
assign addr[60249] = 1492592527;
assign addr[60250] = 1478784851;
assign addr[60251] = 1464859917;
assign addr[60252] = 1450818828;
assign addr[60253] = 1436662698;
assign addr[60254] = 1422392650;
assign addr[60255] = 1408009814;
assign addr[60256] = 1393515332;
assign addr[60257] = 1378910353;
assign addr[60258] = 1364196034;
assign addr[60259] = 1349373543;
assign addr[60260] = 1334444055;
assign addr[60261] = 1319408754;
assign addr[60262] = 1304268832;
assign addr[60263] = 1289025489;
assign addr[60264] = 1273679934;
assign addr[60265] = 1258233384;
assign addr[60266] = 1242687064;
assign addr[60267] = 1227042207;
assign addr[60268] = 1211300053;
assign addr[60269] = 1195461849;
assign addr[60270] = 1179528853;
assign addr[60271] = 1163502328;
assign addr[60272] = 1147383544;
assign addr[60273] = 1131173780;
assign addr[60274] = 1114874320;
assign addr[60275] = 1098486458;
assign addr[60276] = 1082011492;
assign addr[60277] = 1065450729;
assign addr[60278] = 1048805483;
assign addr[60279] = 1032077073;
assign addr[60280] = 1015266825;
assign addr[60281] = 998376073;
assign addr[60282] = 981406156;
assign addr[60283] = 964358420;
assign addr[60284] = 947234215;
assign addr[60285] = 930034901;
assign addr[60286] = 912761841;
assign addr[60287] = 895416404;
assign addr[60288] = 877999966;
assign addr[60289] = 860513908;
assign addr[60290] = 842959617;
assign addr[60291] = 825338484;
assign addr[60292] = 807651907;
assign addr[60293] = 789901288;
assign addr[60294] = 772088034;
assign addr[60295] = 754213559;
assign addr[60296] = 736279279;
assign addr[60297] = 718286617;
assign addr[60298] = 700236999;
assign addr[60299] = 682131857;
assign addr[60300] = 663972625;
assign addr[60301] = 645760745;
assign addr[60302] = 627497660;
assign addr[60303] = 609184818;
assign addr[60304] = 590823671;
assign addr[60305] = 572415676;
assign addr[60306] = 553962291;
assign addr[60307] = 535464981;
assign addr[60308] = 516925212;
assign addr[60309] = 498344454;
assign addr[60310] = 479724180;
assign addr[60311] = 461065866;
assign addr[60312] = 442370993;
assign addr[60313] = 423641043;
assign addr[60314] = 404877501;
assign addr[60315] = 386081854;
assign addr[60316] = 367255594;
assign addr[60317] = 348400212;
assign addr[60318] = 329517204;
assign addr[60319] = 310608068;
assign addr[60320] = 291674302;
assign addr[60321] = 272717408;
assign addr[60322] = 253738890;
assign addr[60323] = 234740251;
assign addr[60324] = 215722999;
assign addr[60325] = 196688642;
assign addr[60326] = 177638688;
assign addr[60327] = 158574649;
assign addr[60328] = 139498035;
assign addr[60329] = 120410361;
assign addr[60330] = 101313138;
assign addr[60331] = 82207882;
assign addr[60332] = 63096108;
assign addr[60333] = 43979330;
assign addr[60334] = 24859065;
assign addr[60335] = 5736829;
assign addr[60336] = -13385863;
assign addr[60337] = -32507492;
assign addr[60338] = -51626544;
assign addr[60339] = -70741503;
assign addr[60340] = -89850852;
assign addr[60341] = -108953076;
assign addr[60342] = -128046661;
assign addr[60343] = -147130093;
assign addr[60344] = -166201858;
assign addr[60345] = -185260444;
assign addr[60346] = -204304341;
assign addr[60347] = -223332037;
assign addr[60348] = -242342025;
assign addr[60349] = -261332796;
assign addr[60350] = -280302845;
assign addr[60351] = -299250668;
assign addr[60352] = -318174762;
assign addr[60353] = -337073627;
assign addr[60354] = -355945764;
assign addr[60355] = -374789676;
assign addr[60356] = -393603870;
assign addr[60357] = -412386854;
assign addr[60358] = -431137138;
assign addr[60359] = -449853235;
assign addr[60360] = -468533662;
assign addr[60361] = -487176937;
assign addr[60362] = -505781581;
assign addr[60363] = -524346121;
assign addr[60364] = -542869083;
assign addr[60365] = -561348998;
assign addr[60366] = -579784402;
assign addr[60367] = -598173833;
assign addr[60368] = -616515832;
assign addr[60369] = -634808946;
assign addr[60370] = -653051723;
assign addr[60371] = -671242716;
assign addr[60372] = -689380485;
assign addr[60373] = -707463589;
assign addr[60374] = -725490597;
assign addr[60375] = -743460077;
assign addr[60376] = -761370605;
assign addr[60377] = -779220762;
assign addr[60378] = -797009130;
assign addr[60379] = -814734301;
assign addr[60380] = -832394869;
assign addr[60381] = -849989433;
assign addr[60382] = -867516597;
assign addr[60383] = -884974973;
assign addr[60384] = -902363176;
assign addr[60385] = -919679827;
assign addr[60386] = -936923553;
assign addr[60387] = -954092986;
assign addr[60388] = -971186766;
assign addr[60389] = -988203537;
assign addr[60390] = -1005141949;
assign addr[60391] = -1022000660;
assign addr[60392] = -1038778332;
assign addr[60393] = -1055473635;
assign addr[60394] = -1072085246;
assign addr[60395] = -1088611847;
assign addr[60396] = -1105052128;
assign addr[60397] = -1121404785;
assign addr[60398] = -1137668521;
assign addr[60399] = -1153842047;
assign addr[60400] = -1169924081;
assign addr[60401] = -1185913346;
assign addr[60402] = -1201808576;
assign addr[60403] = -1217608510;
assign addr[60404] = -1233311895;
assign addr[60405] = -1248917486;
assign addr[60406] = -1264424045;
assign addr[60407] = -1279830344;
assign addr[60408] = -1295135159;
assign addr[60409] = -1310337279;
assign addr[60410] = -1325435496;
assign addr[60411] = -1340428615;
assign addr[60412] = -1355315445;
assign addr[60413] = -1370094808;
assign addr[60414] = -1384765530;
assign addr[60415] = -1399326449;
assign addr[60416] = -1413776410;
assign addr[60417] = -1428114267;
assign addr[60418] = -1442338884;
assign addr[60419] = -1456449131;
assign addr[60420] = -1470443891;
assign addr[60421] = -1484322054;
assign addr[60422] = -1498082520;
assign addr[60423] = -1511724196;
assign addr[60424] = -1525246002;
assign addr[60425] = -1538646865;
assign addr[60426] = -1551925723;
assign addr[60427] = -1565081523;
assign addr[60428] = -1578113222;
assign addr[60429] = -1591019785;
assign addr[60430] = -1603800191;
assign addr[60431] = -1616453425;
assign addr[60432] = -1628978484;
assign addr[60433] = -1641374375;
assign addr[60434] = -1653640115;
assign addr[60435] = -1665774731;
assign addr[60436] = -1677777262;
assign addr[60437] = -1689646755;
assign addr[60438] = -1701382270;
assign addr[60439] = -1712982875;
assign addr[60440] = -1724447652;
assign addr[60441] = -1735775690;
assign addr[60442] = -1746966091;
assign addr[60443] = -1758017969;
assign addr[60444] = -1768930447;
assign addr[60445] = -1779702660;
assign addr[60446] = -1790333753;
assign addr[60447] = -1800822883;
assign addr[60448] = -1811169220;
assign addr[60449] = -1821371941;
assign addr[60450] = -1831430239;
assign addr[60451] = -1841343316;
assign addr[60452] = -1851110385;
assign addr[60453] = -1860730673;
assign addr[60454] = -1870203416;
assign addr[60455] = -1879527863;
assign addr[60456] = -1888703276;
assign addr[60457] = -1897728925;
assign addr[60458] = -1906604097;
assign addr[60459] = -1915328086;
assign addr[60460] = -1923900201;
assign addr[60461] = -1932319763;
assign addr[60462] = -1940586104;
assign addr[60463] = -1948698568;
assign addr[60464] = -1956656513;
assign addr[60465] = -1964459306;
assign addr[60466] = -1972106330;
assign addr[60467] = -1979596978;
assign addr[60468] = -1986930656;
assign addr[60469] = -1994106782;
assign addr[60470] = -2001124788;
assign addr[60471] = -2007984117;
assign addr[60472] = -2014684225;
assign addr[60473] = -2021224581;
assign addr[60474] = -2027604666;
assign addr[60475] = -2033823974;
assign addr[60476] = -2039882013;
assign addr[60477] = -2045778302;
assign addr[60478] = -2051512372;
assign addr[60479] = -2057083771;
assign addr[60480] = -2062492055;
assign addr[60481] = -2067736796;
assign addr[60482] = -2072817579;
assign addr[60483] = -2077733999;
assign addr[60484] = -2082485668;
assign addr[60485] = -2087072209;
assign addr[60486] = -2091493257;
assign addr[60487] = -2095748463;
assign addr[60488] = -2099837489;
assign addr[60489] = -2103760010;
assign addr[60490] = -2107515716;
assign addr[60491] = -2111104309;
assign addr[60492] = -2114525505;
assign addr[60493] = -2117779031;
assign addr[60494] = -2120864631;
assign addr[60495] = -2123782059;
assign addr[60496] = -2126531084;
assign addr[60497] = -2129111488;
assign addr[60498] = -2131523066;
assign addr[60499] = -2133765628;
assign addr[60500] = -2135838995;
assign addr[60501] = -2137743003;
assign addr[60502] = -2139477502;
assign addr[60503] = -2141042352;
assign addr[60504] = -2142437431;
assign addr[60505] = -2143662628;
assign addr[60506] = -2144717846;
assign addr[60507] = -2145603001;
assign addr[60508] = -2146318022;
assign addr[60509] = -2146862854;
assign addr[60510] = -2147237452;
assign addr[60511] = -2147441787;
assign addr[60512] = -2147475844;
assign addr[60513] = -2147339619;
assign addr[60514] = -2147033123;
assign addr[60515] = -2146556380;
assign addr[60516] = -2145909429;
assign addr[60517] = -2145092320;
assign addr[60518] = -2144105118;
assign addr[60519] = -2142947902;
assign addr[60520] = -2141620763;
assign addr[60521] = -2140123807;
assign addr[60522] = -2138457152;
assign addr[60523] = -2136620930;
assign addr[60524] = -2134615288;
assign addr[60525] = -2132440383;
assign addr[60526] = -2130096389;
assign addr[60527] = -2127583492;
assign addr[60528] = -2124901890;
assign addr[60529] = -2122051796;
assign addr[60530] = -2119033436;
assign addr[60531] = -2115847050;
assign addr[60532] = -2112492891;
assign addr[60533] = -2108971223;
assign addr[60534] = -2105282327;
assign addr[60535] = -2101426496;
assign addr[60536] = -2097404033;
assign addr[60537] = -2093215260;
assign addr[60538] = -2088860507;
assign addr[60539] = -2084340120;
assign addr[60540] = -2079654458;
assign addr[60541] = -2074803892;
assign addr[60542] = -2069788807;
assign addr[60543] = -2064609600;
assign addr[60544] = -2059266683;
assign addr[60545] = -2053760478;
assign addr[60546] = -2048091422;
assign addr[60547] = -2042259965;
assign addr[60548] = -2036266570;
assign addr[60549] = -2030111710;
assign addr[60550] = -2023795876;
assign addr[60551] = -2017319567;
assign addr[60552] = -2010683297;
assign addr[60553] = -2003887591;
assign addr[60554] = -1996932990;
assign addr[60555] = -1989820044;
assign addr[60556] = -1982549318;
assign addr[60557] = -1975121388;
assign addr[60558] = -1967536842;
assign addr[60559] = -1959796283;
assign addr[60560] = -1951900324;
assign addr[60561] = -1943849591;
assign addr[60562] = -1935644723;
assign addr[60563] = -1927286370;
assign addr[60564] = -1918775195;
assign addr[60565] = -1910111873;
assign addr[60566] = -1901297091;
assign addr[60567] = -1892331547;
assign addr[60568] = -1883215953;
assign addr[60569] = -1873951032;
assign addr[60570] = -1864537518;
assign addr[60571] = -1854976157;
assign addr[60572] = -1845267708;
assign addr[60573] = -1835412941;
assign addr[60574] = -1825412636;
assign addr[60575] = -1815267588;
assign addr[60576] = -1804978599;
assign addr[60577] = -1794546487;
assign addr[60578] = -1783972079;
assign addr[60579] = -1773256212;
assign addr[60580] = -1762399737;
assign addr[60581] = -1751403515;
assign addr[60582] = -1740268417;
assign addr[60583] = -1728995326;
assign addr[60584] = -1717585136;
assign addr[60585] = -1706038753;
assign addr[60586] = -1694357091;
assign addr[60587] = -1682541077;
assign addr[60588] = -1670591647;
assign addr[60589] = -1658509750;
assign addr[60590] = -1646296344;
assign addr[60591] = -1633952396;
assign addr[60592] = -1621478885;
assign addr[60593] = -1608876801;
assign addr[60594] = -1596147143;
assign addr[60595] = -1583290921;
assign addr[60596] = -1570309153;
assign addr[60597] = -1557202869;
assign addr[60598] = -1543973108;
assign addr[60599] = -1530620920;
assign addr[60600] = -1517147363;
assign addr[60601] = -1503553506;
assign addr[60602] = -1489840425;
assign addr[60603] = -1476009210;
assign addr[60604] = -1462060956;
assign addr[60605] = -1447996770;
assign addr[60606] = -1433817766;
assign addr[60607] = -1419525069;
assign addr[60608] = -1405119813;
assign addr[60609] = -1390603139;
assign addr[60610] = -1375976199;
assign addr[60611] = -1361240152;
assign addr[60612] = -1346396168;
assign addr[60613] = -1331445422;
assign addr[60614] = -1316389101;
assign addr[60615] = -1301228398;
assign addr[60616] = -1285964516;
assign addr[60617] = -1270598665;
assign addr[60618] = -1255132063;
assign addr[60619] = -1239565936;
assign addr[60620] = -1223901520;
assign addr[60621] = -1208140056;
assign addr[60622] = -1192282793;
assign addr[60623] = -1176330990;
assign addr[60624] = -1160285911;
assign addr[60625] = -1144148829;
assign addr[60626] = -1127921022;
assign addr[60627] = -1111603778;
assign addr[60628] = -1095198391;
assign addr[60629] = -1078706161;
assign addr[60630] = -1062128397;
assign addr[60631] = -1045466412;
assign addr[60632] = -1028721528;
assign addr[60633] = -1011895073;
assign addr[60634] = -994988380;
assign addr[60635] = -978002791;
assign addr[60636] = -960939653;
assign addr[60637] = -943800318;
assign addr[60638] = -926586145;
assign addr[60639] = -909298500;
assign addr[60640] = -891938752;
assign addr[60641] = -874508280;
assign addr[60642] = -857008464;
assign addr[60643] = -839440693;
assign addr[60644] = -821806359;
assign addr[60645] = -804106861;
assign addr[60646] = -786343603;
assign addr[60647] = -768517992;
assign addr[60648] = -750631442;
assign addr[60649] = -732685372;
assign addr[60650] = -714681204;
assign addr[60651] = -696620367;
assign addr[60652] = -678504291;
assign addr[60653] = -660334415;
assign addr[60654] = -642112178;
assign addr[60655] = -623839025;
assign addr[60656] = -605516406;
assign addr[60657] = -587145773;
assign addr[60658] = -568728583;
assign addr[60659] = -550266296;
assign addr[60660] = -531760377;
assign addr[60661] = -513212292;
assign addr[60662] = -494623513;
assign addr[60663] = -475995513;
assign addr[60664] = -457329769;
assign addr[60665] = -438627762;
assign addr[60666] = -419890975;
assign addr[60667] = -401120892;
assign addr[60668] = -382319004;
assign addr[60669] = -363486799;
assign addr[60670] = -344625773;
assign addr[60671] = -325737419;
assign addr[60672] = -306823237;
assign addr[60673] = -287884725;
assign addr[60674] = -268923386;
assign addr[60675] = -249940723;
assign addr[60676] = -230938242;
assign addr[60677] = -211917448;
assign addr[60678] = -192879850;
assign addr[60679] = -173826959;
assign addr[60680] = -154760284;
assign addr[60681] = -135681337;
assign addr[60682] = -116591632;
assign addr[60683] = -97492681;
assign addr[60684] = -78386000;
assign addr[60685] = -59273104;
assign addr[60686] = -40155507;
assign addr[60687] = -21034727;
assign addr[60688] = -1912278;
assign addr[60689] = 17210322;
assign addr[60690] = 36331557;
assign addr[60691] = 55449912;
assign addr[60692] = 74563870;
assign addr[60693] = 93671915;
assign addr[60694] = 112772533;
assign addr[60695] = 131864208;
assign addr[60696] = 150945428;
assign addr[60697] = 170014678;
assign addr[60698] = 189070447;
assign addr[60699] = 208111224;
assign addr[60700] = 227135500;
assign addr[60701] = 246141764;
assign addr[60702] = 265128512;
assign addr[60703] = 284094236;
assign addr[60704] = 303037433;
assign addr[60705] = 321956601;
assign addr[60706] = 340850240;
assign addr[60707] = 359716852;
assign addr[60708] = 378554940;
assign addr[60709] = 397363011;
assign addr[60710] = 416139574;
assign addr[60711] = 434883140;
assign addr[60712] = 453592221;
assign addr[60713] = 472265336;
assign addr[60714] = 490901003;
assign addr[60715] = 509497745;
assign addr[60716] = 528054086;
assign addr[60717] = 546568556;
assign addr[60718] = 565039687;
assign addr[60719] = 583466013;
assign addr[60720] = 601846074;
assign addr[60721] = 620178412;
assign addr[60722] = 638461574;
assign addr[60723] = 656694110;
assign addr[60724] = 674874574;
assign addr[60725] = 693001525;
assign addr[60726] = 711073524;
assign addr[60727] = 729089140;
assign addr[60728] = 747046944;
assign addr[60729] = 764945512;
assign addr[60730] = 782783424;
assign addr[60731] = 800559266;
assign addr[60732] = 818271628;
assign addr[60733] = 835919107;
assign addr[60734] = 853500302;
assign addr[60735] = 871013820;
assign addr[60736] = 888458272;
assign addr[60737] = 905832274;
assign addr[60738] = 923134450;
assign addr[60739] = 940363427;
assign addr[60740] = 957517838;
assign addr[60741] = 974596324;
assign addr[60742] = 991597531;
assign addr[60743] = 1008520110;
assign addr[60744] = 1025362720;
assign addr[60745] = 1042124025;
assign addr[60746] = 1058802695;
assign addr[60747] = 1075397409;
assign addr[60748] = 1091906851;
assign addr[60749] = 1108329711;
assign addr[60750] = 1124664687;
assign addr[60751] = 1140910484;
assign addr[60752] = 1157065814;
assign addr[60753] = 1173129396;
assign addr[60754] = 1189099956;
assign addr[60755] = 1204976227;
assign addr[60756] = 1220756951;
assign addr[60757] = 1236440877;
assign addr[60758] = 1252026760;
assign addr[60759] = 1267513365;
assign addr[60760] = 1282899464;
assign addr[60761] = 1298183838;
assign addr[60762] = 1313365273;
assign addr[60763] = 1328442566;
assign addr[60764] = 1343414522;
assign addr[60765] = 1358279953;
assign addr[60766] = 1373037681;
assign addr[60767] = 1387686535;
assign addr[60768] = 1402225355;
assign addr[60769] = 1416652986;
assign addr[60770] = 1430968286;
assign addr[60771] = 1445170118;
assign addr[60772] = 1459257358;
assign addr[60773] = 1473228887;
assign addr[60774] = 1487083598;
assign addr[60775] = 1500820393;
assign addr[60776] = 1514438181;
assign addr[60777] = 1527935884;
assign addr[60778] = 1541312431;
assign addr[60779] = 1554566762;
assign addr[60780] = 1567697824;
assign addr[60781] = 1580704578;
assign addr[60782] = 1593585992;
assign addr[60783] = 1606341043;
assign addr[60784] = 1618968722;
assign addr[60785] = 1631468027;
assign addr[60786] = 1643837966;
assign addr[60787] = 1656077559;
assign addr[60788] = 1668185835;
assign addr[60789] = 1680161834;
assign addr[60790] = 1692004606;
assign addr[60791] = 1703713213;
assign addr[60792] = 1715286726;
assign addr[60793] = 1726724227;
assign addr[60794] = 1738024810;
assign addr[60795] = 1749187577;
assign addr[60796] = 1760211645;
assign addr[60797] = 1771096139;
assign addr[60798] = 1781840195;
assign addr[60799] = 1792442963;
assign addr[60800] = 1802903601;
assign addr[60801] = 1813221279;
assign addr[60802] = 1823395180;
assign addr[60803] = 1833424497;
assign addr[60804] = 1843308435;
assign addr[60805] = 1853046210;
assign addr[60806] = 1862637049;
assign addr[60807] = 1872080193;
assign addr[60808] = 1881374892;
assign addr[60809] = 1890520410;
assign addr[60810] = 1899516021;
assign addr[60811] = 1908361011;
assign addr[60812] = 1917054681;
assign addr[60813] = 1925596340;
assign addr[60814] = 1933985310;
assign addr[60815] = 1942220928;
assign addr[60816] = 1950302539;
assign addr[60817] = 1958229503;
assign addr[60818] = 1966001192;
assign addr[60819] = 1973616989;
assign addr[60820] = 1981076290;
assign addr[60821] = 1988378503;
assign addr[60822] = 1995523051;
assign addr[60823] = 2002509365;
assign addr[60824] = 2009336893;
assign addr[60825] = 2016005093;
assign addr[60826] = 2022513436;
assign addr[60827] = 2028861406;
assign addr[60828] = 2035048499;
assign addr[60829] = 2041074226;
assign addr[60830] = 2046938108;
assign addr[60831] = 2052639680;
assign addr[60832] = 2058178491;
assign addr[60833] = 2063554100;
assign addr[60834] = 2068766083;
assign addr[60835] = 2073814024;
assign addr[60836] = 2078697525;
assign addr[60837] = 2083416198;
assign addr[60838] = 2087969669;
assign addr[60839] = 2092357577;
assign addr[60840] = 2096579573;
assign addr[60841] = 2100635323;
assign addr[60842] = 2104524506;
assign addr[60843] = 2108246813;
assign addr[60844] = 2111801949;
assign addr[60845] = 2115189632;
assign addr[60846] = 2118409593;
assign addr[60847] = 2121461578;
assign addr[60848] = 2124345343;
assign addr[60849] = 2127060661;
assign addr[60850] = 2129607316;
assign addr[60851] = 2131985106;
assign addr[60852] = 2134193842;
assign addr[60853] = 2136233350;
assign addr[60854] = 2138103468;
assign addr[60855] = 2139804048;
assign addr[60856] = 2141334954;
assign addr[60857] = 2142696065;
assign addr[60858] = 2143887273;
assign addr[60859] = 2144908484;
assign addr[60860] = 2145759618;
assign addr[60861] = 2146440605;
assign addr[60862] = 2146951393;
assign addr[60863] = 2147291941;
assign addr[60864] = 2147462221;
assign addr[60865] = 2147462221;
assign addr[60866] = 2147291941;
assign addr[60867] = 2146951393;
assign addr[60868] = 2146440605;
assign addr[60869] = 2145759618;
assign addr[60870] = 2144908484;
assign addr[60871] = 2143887273;
assign addr[60872] = 2142696065;
assign addr[60873] = 2141334954;
assign addr[60874] = 2139804048;
assign addr[60875] = 2138103468;
assign addr[60876] = 2136233350;
assign addr[60877] = 2134193842;
assign addr[60878] = 2131985106;
assign addr[60879] = 2129607316;
assign addr[60880] = 2127060661;
assign addr[60881] = 2124345343;
assign addr[60882] = 2121461578;
assign addr[60883] = 2118409593;
assign addr[60884] = 2115189632;
assign addr[60885] = 2111801949;
assign addr[60886] = 2108246813;
assign addr[60887] = 2104524506;
assign addr[60888] = 2100635323;
assign addr[60889] = 2096579573;
assign addr[60890] = 2092357577;
assign addr[60891] = 2087969669;
assign addr[60892] = 2083416198;
assign addr[60893] = 2078697525;
assign addr[60894] = 2073814024;
assign addr[60895] = 2068766083;
assign addr[60896] = 2063554100;
assign addr[60897] = 2058178491;
assign addr[60898] = 2052639680;
assign addr[60899] = 2046938108;
assign addr[60900] = 2041074226;
assign addr[60901] = 2035048499;
assign addr[60902] = 2028861406;
assign addr[60903] = 2022513436;
assign addr[60904] = 2016005093;
assign addr[60905] = 2009336893;
assign addr[60906] = 2002509365;
assign addr[60907] = 1995523051;
assign addr[60908] = 1988378503;
assign addr[60909] = 1981076290;
assign addr[60910] = 1973616989;
assign addr[60911] = 1966001192;
assign addr[60912] = 1958229503;
assign addr[60913] = 1950302539;
assign addr[60914] = 1942220928;
assign addr[60915] = 1933985310;
assign addr[60916] = 1925596340;
assign addr[60917] = 1917054681;
assign addr[60918] = 1908361011;
assign addr[60919] = 1899516021;
assign addr[60920] = 1890520410;
assign addr[60921] = 1881374892;
assign addr[60922] = 1872080193;
assign addr[60923] = 1862637049;
assign addr[60924] = 1853046210;
assign addr[60925] = 1843308435;
assign addr[60926] = 1833424497;
assign addr[60927] = 1823395180;
assign addr[60928] = 1813221279;
assign addr[60929] = 1802903601;
assign addr[60930] = 1792442963;
assign addr[60931] = 1781840195;
assign addr[60932] = 1771096139;
assign addr[60933] = 1760211645;
assign addr[60934] = 1749187577;
assign addr[60935] = 1738024810;
assign addr[60936] = 1726724227;
assign addr[60937] = 1715286726;
assign addr[60938] = 1703713213;
assign addr[60939] = 1692004606;
assign addr[60940] = 1680161834;
assign addr[60941] = 1668185835;
assign addr[60942] = 1656077559;
assign addr[60943] = 1643837966;
assign addr[60944] = 1631468027;
assign addr[60945] = 1618968722;
assign addr[60946] = 1606341043;
assign addr[60947] = 1593585992;
assign addr[60948] = 1580704578;
assign addr[60949] = 1567697824;
assign addr[60950] = 1554566762;
assign addr[60951] = 1541312431;
assign addr[60952] = 1527935884;
assign addr[60953] = 1514438181;
assign addr[60954] = 1500820393;
assign addr[60955] = 1487083598;
assign addr[60956] = 1473228887;
assign addr[60957] = 1459257358;
assign addr[60958] = 1445170118;
assign addr[60959] = 1430968286;
assign addr[60960] = 1416652986;
assign addr[60961] = 1402225355;
assign addr[60962] = 1387686535;
assign addr[60963] = 1373037681;
assign addr[60964] = 1358279953;
assign addr[60965] = 1343414522;
assign addr[60966] = 1328442566;
assign addr[60967] = 1313365273;
assign addr[60968] = 1298183838;
assign addr[60969] = 1282899464;
assign addr[60970] = 1267513365;
assign addr[60971] = 1252026760;
assign addr[60972] = 1236440877;
assign addr[60973] = 1220756951;
assign addr[60974] = 1204976227;
assign addr[60975] = 1189099956;
assign addr[60976] = 1173129396;
assign addr[60977] = 1157065814;
assign addr[60978] = 1140910484;
assign addr[60979] = 1124664687;
assign addr[60980] = 1108329711;
assign addr[60981] = 1091906851;
assign addr[60982] = 1075397409;
assign addr[60983] = 1058802695;
assign addr[60984] = 1042124025;
assign addr[60985] = 1025362720;
assign addr[60986] = 1008520110;
assign addr[60987] = 991597531;
assign addr[60988] = 974596324;
assign addr[60989] = 957517838;
assign addr[60990] = 940363427;
assign addr[60991] = 923134450;
assign addr[60992] = 905832274;
assign addr[60993] = 888458272;
assign addr[60994] = 871013820;
assign addr[60995] = 853500302;
assign addr[60996] = 835919107;
assign addr[60997] = 818271628;
assign addr[60998] = 800559266;
assign addr[60999] = 782783424;
assign addr[61000] = 764945512;
assign addr[61001] = 747046944;
assign addr[61002] = 729089140;
assign addr[61003] = 711073524;
assign addr[61004] = 693001525;
assign addr[61005] = 674874574;
assign addr[61006] = 656694110;
assign addr[61007] = 638461574;
assign addr[61008] = 620178412;
assign addr[61009] = 601846074;
assign addr[61010] = 583466013;
assign addr[61011] = 565039687;
assign addr[61012] = 546568556;
assign addr[61013] = 528054086;
assign addr[61014] = 509497745;
assign addr[61015] = 490901003;
assign addr[61016] = 472265336;
assign addr[61017] = 453592221;
assign addr[61018] = 434883140;
assign addr[61019] = 416139574;
assign addr[61020] = 397363011;
assign addr[61021] = 378554940;
assign addr[61022] = 359716852;
assign addr[61023] = 340850240;
assign addr[61024] = 321956601;
assign addr[61025] = 303037433;
assign addr[61026] = 284094236;
assign addr[61027] = 265128512;
assign addr[61028] = 246141764;
assign addr[61029] = 227135500;
assign addr[61030] = 208111224;
assign addr[61031] = 189070447;
assign addr[61032] = 170014678;
assign addr[61033] = 150945428;
assign addr[61034] = 131864208;
assign addr[61035] = 112772533;
assign addr[61036] = 93671915;
assign addr[61037] = 74563870;
assign addr[61038] = 55449912;
assign addr[61039] = 36331557;
assign addr[61040] = 17210322;
assign addr[61041] = -1912278;
assign addr[61042] = -21034727;
assign addr[61043] = -40155507;
assign addr[61044] = -59273104;
assign addr[61045] = -78386000;
assign addr[61046] = -97492681;
assign addr[61047] = -116591632;
assign addr[61048] = -135681337;
assign addr[61049] = -154760284;
assign addr[61050] = -173826959;
assign addr[61051] = -192879850;
assign addr[61052] = -211917448;
assign addr[61053] = -230938242;
assign addr[61054] = -249940723;
assign addr[61055] = -268923386;
assign addr[61056] = -287884725;
assign addr[61057] = -306823237;
assign addr[61058] = -325737419;
assign addr[61059] = -344625773;
assign addr[61060] = -363486799;
assign addr[61061] = -382319004;
assign addr[61062] = -401120892;
assign addr[61063] = -419890975;
assign addr[61064] = -438627762;
assign addr[61065] = -457329769;
assign addr[61066] = -475995513;
assign addr[61067] = -494623513;
assign addr[61068] = -513212292;
assign addr[61069] = -531760377;
assign addr[61070] = -550266296;
assign addr[61071] = -568728583;
assign addr[61072] = -587145773;
assign addr[61073] = -605516406;
assign addr[61074] = -623839025;
assign addr[61075] = -642112178;
assign addr[61076] = -660334415;
assign addr[61077] = -678504291;
assign addr[61078] = -696620367;
assign addr[61079] = -714681204;
assign addr[61080] = -732685372;
assign addr[61081] = -750631442;
assign addr[61082] = -768517992;
assign addr[61083] = -786343603;
assign addr[61084] = -804106861;
assign addr[61085] = -821806359;
assign addr[61086] = -839440693;
assign addr[61087] = -857008464;
assign addr[61088] = -874508280;
assign addr[61089] = -891938752;
assign addr[61090] = -909298500;
assign addr[61091] = -926586145;
assign addr[61092] = -943800318;
assign addr[61093] = -960939653;
assign addr[61094] = -978002791;
assign addr[61095] = -994988380;
assign addr[61096] = -1011895073;
assign addr[61097] = -1028721528;
assign addr[61098] = -1045466412;
assign addr[61099] = -1062128397;
assign addr[61100] = -1078706161;
assign addr[61101] = -1095198391;
assign addr[61102] = -1111603778;
assign addr[61103] = -1127921022;
assign addr[61104] = -1144148829;
assign addr[61105] = -1160285911;
assign addr[61106] = -1176330990;
assign addr[61107] = -1192282793;
assign addr[61108] = -1208140056;
assign addr[61109] = -1223901520;
assign addr[61110] = -1239565936;
assign addr[61111] = -1255132063;
assign addr[61112] = -1270598665;
assign addr[61113] = -1285964516;
assign addr[61114] = -1301228398;
assign addr[61115] = -1316389101;
assign addr[61116] = -1331445422;
assign addr[61117] = -1346396168;
assign addr[61118] = -1361240152;
assign addr[61119] = -1375976199;
assign addr[61120] = -1390603139;
assign addr[61121] = -1405119813;
assign addr[61122] = -1419525069;
assign addr[61123] = -1433817766;
assign addr[61124] = -1447996770;
assign addr[61125] = -1462060956;
assign addr[61126] = -1476009210;
assign addr[61127] = -1489840425;
assign addr[61128] = -1503553506;
assign addr[61129] = -1517147363;
assign addr[61130] = -1530620920;
assign addr[61131] = -1543973108;
assign addr[61132] = -1557202869;
assign addr[61133] = -1570309153;
assign addr[61134] = -1583290921;
assign addr[61135] = -1596147143;
assign addr[61136] = -1608876801;
assign addr[61137] = -1621478885;
assign addr[61138] = -1633952396;
assign addr[61139] = -1646296344;
assign addr[61140] = -1658509750;
assign addr[61141] = -1670591647;
assign addr[61142] = -1682541077;
assign addr[61143] = -1694357091;
assign addr[61144] = -1706038753;
assign addr[61145] = -1717585136;
assign addr[61146] = -1728995326;
assign addr[61147] = -1740268417;
assign addr[61148] = -1751403515;
assign addr[61149] = -1762399737;
assign addr[61150] = -1773256212;
assign addr[61151] = -1783972079;
assign addr[61152] = -1794546487;
assign addr[61153] = -1804978599;
assign addr[61154] = -1815267588;
assign addr[61155] = -1825412636;
assign addr[61156] = -1835412941;
assign addr[61157] = -1845267708;
assign addr[61158] = -1854976157;
assign addr[61159] = -1864537518;
assign addr[61160] = -1873951032;
assign addr[61161] = -1883215953;
assign addr[61162] = -1892331547;
assign addr[61163] = -1901297091;
assign addr[61164] = -1910111873;
assign addr[61165] = -1918775195;
assign addr[61166] = -1927286370;
assign addr[61167] = -1935644723;
assign addr[61168] = -1943849591;
assign addr[61169] = -1951900324;
assign addr[61170] = -1959796283;
assign addr[61171] = -1967536842;
assign addr[61172] = -1975121388;
assign addr[61173] = -1982549318;
assign addr[61174] = -1989820044;
assign addr[61175] = -1996932990;
assign addr[61176] = -2003887591;
assign addr[61177] = -2010683297;
assign addr[61178] = -2017319567;
assign addr[61179] = -2023795876;
assign addr[61180] = -2030111710;
assign addr[61181] = -2036266570;
assign addr[61182] = -2042259965;
assign addr[61183] = -2048091422;
assign addr[61184] = -2053760478;
assign addr[61185] = -2059266683;
assign addr[61186] = -2064609600;
assign addr[61187] = -2069788807;
assign addr[61188] = -2074803892;
assign addr[61189] = -2079654458;
assign addr[61190] = -2084340120;
assign addr[61191] = -2088860507;
assign addr[61192] = -2093215260;
assign addr[61193] = -2097404033;
assign addr[61194] = -2101426496;
assign addr[61195] = -2105282327;
assign addr[61196] = -2108971223;
assign addr[61197] = -2112492891;
assign addr[61198] = -2115847050;
assign addr[61199] = -2119033436;
assign addr[61200] = -2122051796;
assign addr[61201] = -2124901890;
assign addr[61202] = -2127583492;
assign addr[61203] = -2130096389;
assign addr[61204] = -2132440383;
assign addr[61205] = -2134615288;
assign addr[61206] = -2136620930;
assign addr[61207] = -2138457152;
assign addr[61208] = -2140123807;
assign addr[61209] = -2141620763;
assign addr[61210] = -2142947902;
assign addr[61211] = -2144105118;
assign addr[61212] = -2145092320;
assign addr[61213] = -2145909429;
assign addr[61214] = -2146556380;
assign addr[61215] = -2147033123;
assign addr[61216] = -2147339619;
assign addr[61217] = -2147475844;
assign addr[61218] = -2147441787;
assign addr[61219] = -2147237452;
assign addr[61220] = -2146862854;
assign addr[61221] = -2146318022;
assign addr[61222] = -2145603001;
assign addr[61223] = -2144717846;
assign addr[61224] = -2143662628;
assign addr[61225] = -2142437431;
assign addr[61226] = -2141042352;
assign addr[61227] = -2139477502;
assign addr[61228] = -2137743003;
assign addr[61229] = -2135838995;
assign addr[61230] = -2133765628;
assign addr[61231] = -2131523066;
assign addr[61232] = -2129111488;
assign addr[61233] = -2126531084;
assign addr[61234] = -2123782059;
assign addr[61235] = -2120864631;
assign addr[61236] = -2117779031;
assign addr[61237] = -2114525505;
assign addr[61238] = -2111104309;
assign addr[61239] = -2107515716;
assign addr[61240] = -2103760010;
assign addr[61241] = -2099837489;
assign addr[61242] = -2095748463;
assign addr[61243] = -2091493257;
assign addr[61244] = -2087072209;
assign addr[61245] = -2082485668;
assign addr[61246] = -2077733999;
assign addr[61247] = -2072817579;
assign addr[61248] = -2067736796;
assign addr[61249] = -2062492055;
assign addr[61250] = -2057083771;
assign addr[61251] = -2051512372;
assign addr[61252] = -2045778302;
assign addr[61253] = -2039882013;
assign addr[61254] = -2033823974;
assign addr[61255] = -2027604666;
assign addr[61256] = -2021224581;
assign addr[61257] = -2014684225;
assign addr[61258] = -2007984117;
assign addr[61259] = -2001124788;
assign addr[61260] = -1994106782;
assign addr[61261] = -1986930656;
assign addr[61262] = -1979596978;
assign addr[61263] = -1972106330;
assign addr[61264] = -1964459306;
assign addr[61265] = -1956656513;
assign addr[61266] = -1948698568;
assign addr[61267] = -1940586104;
assign addr[61268] = -1932319763;
assign addr[61269] = -1923900201;
assign addr[61270] = -1915328086;
assign addr[61271] = -1906604097;
assign addr[61272] = -1897728925;
assign addr[61273] = -1888703276;
assign addr[61274] = -1879527863;
assign addr[61275] = -1870203416;
assign addr[61276] = -1860730673;
assign addr[61277] = -1851110385;
assign addr[61278] = -1841343316;
assign addr[61279] = -1831430239;
assign addr[61280] = -1821371941;
assign addr[61281] = -1811169220;
assign addr[61282] = -1800822883;
assign addr[61283] = -1790333753;
assign addr[61284] = -1779702660;
assign addr[61285] = -1768930447;
assign addr[61286] = -1758017969;
assign addr[61287] = -1746966091;
assign addr[61288] = -1735775690;
assign addr[61289] = -1724447652;
assign addr[61290] = -1712982875;
assign addr[61291] = -1701382270;
assign addr[61292] = -1689646755;
assign addr[61293] = -1677777262;
assign addr[61294] = -1665774731;
assign addr[61295] = -1653640115;
assign addr[61296] = -1641374375;
assign addr[61297] = -1628978484;
assign addr[61298] = -1616453425;
assign addr[61299] = -1603800191;
assign addr[61300] = -1591019785;
assign addr[61301] = -1578113222;
assign addr[61302] = -1565081523;
assign addr[61303] = -1551925723;
assign addr[61304] = -1538646865;
assign addr[61305] = -1525246002;
assign addr[61306] = -1511724196;
assign addr[61307] = -1498082520;
assign addr[61308] = -1484322054;
assign addr[61309] = -1470443891;
assign addr[61310] = -1456449131;
assign addr[61311] = -1442338884;
assign addr[61312] = -1428114267;
assign addr[61313] = -1413776410;
assign addr[61314] = -1399326449;
assign addr[61315] = -1384765530;
assign addr[61316] = -1370094808;
assign addr[61317] = -1355315445;
assign addr[61318] = -1340428615;
assign addr[61319] = -1325435496;
assign addr[61320] = -1310337279;
assign addr[61321] = -1295135159;
assign addr[61322] = -1279830344;
assign addr[61323] = -1264424045;
assign addr[61324] = -1248917486;
assign addr[61325] = -1233311895;
assign addr[61326] = -1217608510;
assign addr[61327] = -1201808576;
assign addr[61328] = -1185913346;
assign addr[61329] = -1169924081;
assign addr[61330] = -1153842047;
assign addr[61331] = -1137668521;
assign addr[61332] = -1121404785;
assign addr[61333] = -1105052128;
assign addr[61334] = -1088611847;
assign addr[61335] = -1072085246;
assign addr[61336] = -1055473635;
assign addr[61337] = -1038778332;
assign addr[61338] = -1022000660;
assign addr[61339] = -1005141949;
assign addr[61340] = -988203537;
assign addr[61341] = -971186766;
assign addr[61342] = -954092986;
assign addr[61343] = -936923553;
assign addr[61344] = -919679827;
assign addr[61345] = -902363176;
assign addr[61346] = -884974973;
assign addr[61347] = -867516597;
assign addr[61348] = -849989433;
assign addr[61349] = -832394869;
assign addr[61350] = -814734301;
assign addr[61351] = -797009130;
assign addr[61352] = -779220762;
assign addr[61353] = -761370605;
assign addr[61354] = -743460077;
assign addr[61355] = -725490597;
assign addr[61356] = -707463589;
assign addr[61357] = -689380485;
assign addr[61358] = -671242716;
assign addr[61359] = -653051723;
assign addr[61360] = -634808946;
assign addr[61361] = -616515832;
assign addr[61362] = -598173833;
assign addr[61363] = -579784402;
assign addr[61364] = -561348998;
assign addr[61365] = -542869083;
assign addr[61366] = -524346121;
assign addr[61367] = -505781581;
assign addr[61368] = -487176937;
assign addr[61369] = -468533662;
assign addr[61370] = -449853235;
assign addr[61371] = -431137138;
assign addr[61372] = -412386854;
assign addr[61373] = -393603870;
assign addr[61374] = -374789676;
assign addr[61375] = -355945764;
assign addr[61376] = -337073627;
assign addr[61377] = -318174762;
assign addr[61378] = -299250668;
assign addr[61379] = -280302845;
assign addr[61380] = -261332796;
assign addr[61381] = -242342025;
assign addr[61382] = -223332037;
assign addr[61383] = -204304341;
assign addr[61384] = -185260444;
assign addr[61385] = -166201858;
assign addr[61386] = -147130093;
assign addr[61387] = -128046661;
assign addr[61388] = -108953076;
assign addr[61389] = -89850852;
assign addr[61390] = -70741503;
assign addr[61391] = -51626544;
assign addr[61392] = -32507492;
assign addr[61393] = -13385863;
assign addr[61394] = 5736829;
assign addr[61395] = 24859065;
assign addr[61396] = 43979330;
assign addr[61397] = 63096108;
assign addr[61398] = 82207882;
assign addr[61399] = 101313138;
assign addr[61400] = 120410361;
assign addr[61401] = 139498035;
assign addr[61402] = 158574649;
assign addr[61403] = 177638688;
assign addr[61404] = 196688642;
assign addr[61405] = 215722999;
assign addr[61406] = 234740251;
assign addr[61407] = 253738890;
assign addr[61408] = 272717408;
assign addr[61409] = 291674302;
assign addr[61410] = 310608068;
assign addr[61411] = 329517204;
assign addr[61412] = 348400212;
assign addr[61413] = 367255594;
assign addr[61414] = 386081854;
assign addr[61415] = 404877501;
assign addr[61416] = 423641043;
assign addr[61417] = 442370993;
assign addr[61418] = 461065866;
assign addr[61419] = 479724180;
assign addr[61420] = 498344454;
assign addr[61421] = 516925212;
assign addr[61422] = 535464981;
assign addr[61423] = 553962291;
assign addr[61424] = 572415676;
assign addr[61425] = 590823671;
assign addr[61426] = 609184818;
assign addr[61427] = 627497660;
assign addr[61428] = 645760745;
assign addr[61429] = 663972625;
assign addr[61430] = 682131857;
assign addr[61431] = 700236999;
assign addr[61432] = 718286617;
assign addr[61433] = 736279279;
assign addr[61434] = 754213559;
assign addr[61435] = 772088034;
assign addr[61436] = 789901288;
assign addr[61437] = 807651907;
assign addr[61438] = 825338484;
assign addr[61439] = 842959617;
assign addr[61440] = 860513908;
assign addr[61441] = 877999966;
assign addr[61442] = 895416404;
assign addr[61443] = 912761841;
assign addr[61444] = 930034901;
assign addr[61445] = 947234215;
assign addr[61446] = 964358420;
assign addr[61447] = 981406156;
assign addr[61448] = 998376073;
assign addr[61449] = 1015266825;
assign addr[61450] = 1032077073;
assign addr[61451] = 1048805483;
assign addr[61452] = 1065450729;
assign addr[61453] = 1082011492;
assign addr[61454] = 1098486458;
assign addr[61455] = 1114874320;
assign addr[61456] = 1131173780;
assign addr[61457] = 1147383544;
assign addr[61458] = 1163502328;
assign addr[61459] = 1179528853;
assign addr[61460] = 1195461849;
assign addr[61461] = 1211300053;
assign addr[61462] = 1227042207;
assign addr[61463] = 1242687064;
assign addr[61464] = 1258233384;
assign addr[61465] = 1273679934;
assign addr[61466] = 1289025489;
assign addr[61467] = 1304268832;
assign addr[61468] = 1319408754;
assign addr[61469] = 1334444055;
assign addr[61470] = 1349373543;
assign addr[61471] = 1364196034;
assign addr[61472] = 1378910353;
assign addr[61473] = 1393515332;
assign addr[61474] = 1408009814;
assign addr[61475] = 1422392650;
assign addr[61476] = 1436662698;
assign addr[61477] = 1450818828;
assign addr[61478] = 1464859917;
assign addr[61479] = 1478784851;
assign addr[61480] = 1492592527;
assign addr[61481] = 1506281850;
assign addr[61482] = 1519851733;
assign addr[61483] = 1533301101;
assign addr[61484] = 1546628888;
assign addr[61485] = 1559834037;
assign addr[61486] = 1572915501;
assign addr[61487] = 1585872242;
assign addr[61488] = 1598703233;
assign addr[61489] = 1611407456;
assign addr[61490] = 1623983905;
assign addr[61491] = 1636431582;
assign addr[61492] = 1648749499;
assign addr[61493] = 1660936681;
assign addr[61494] = 1672992161;
assign addr[61495] = 1684914983;
assign addr[61496] = 1696704201;
assign addr[61497] = 1708358881;
assign addr[61498] = 1719878099;
assign addr[61499] = 1731260941;
assign addr[61500] = 1742506504;
assign addr[61501] = 1753613897;
assign addr[61502] = 1764582240;
assign addr[61503] = 1775410662;
assign addr[61504] = 1786098304;
assign addr[61505] = 1796644320;
assign addr[61506] = 1807047873;
assign addr[61507] = 1817308138;
assign addr[61508] = 1827424302;
assign addr[61509] = 1837395562;
assign addr[61510] = 1847221128;
assign addr[61511] = 1856900221;
assign addr[61512] = 1866432072;
assign addr[61513] = 1875815927;
assign addr[61514] = 1885051042;
assign addr[61515] = 1894136683;
assign addr[61516] = 1903072131;
assign addr[61517] = 1911856677;
assign addr[61518] = 1920489624;
assign addr[61519] = 1928970288;
assign addr[61520] = 1937297997;
assign addr[61521] = 1945472089;
assign addr[61522] = 1953491918;
assign addr[61523] = 1961356847;
assign addr[61524] = 1969066252;
assign addr[61525] = 1976619522;
assign addr[61526] = 1984016058;
assign addr[61527] = 1991255274;
assign addr[61528] = 1998336596;
assign addr[61529] = 2005259462;
assign addr[61530] = 2012023322;
assign addr[61531] = 2018627642;
assign addr[61532] = 2025071897;
assign addr[61533] = 2031355576;
assign addr[61534] = 2037478181;
assign addr[61535] = 2043439226;
assign addr[61536] = 2049238240;
assign addr[61537] = 2054874761;
assign addr[61538] = 2060348343;
assign addr[61539] = 2065658552;
assign addr[61540] = 2070804967;
assign addr[61541] = 2075787180;
assign addr[61542] = 2080604795;
assign addr[61543] = 2085257431;
assign addr[61544] = 2089744719;
assign addr[61545] = 2094066304;
assign addr[61546] = 2098221841;
assign addr[61547] = 2102211002;
assign addr[61548] = 2106033471;
assign addr[61549] = 2109688944;
assign addr[61550] = 2113177132;
assign addr[61551] = 2116497758;
assign addr[61552] = 2119650558;
assign addr[61553] = 2122635283;
assign addr[61554] = 2125451696;
assign addr[61555] = 2128099574;
assign addr[61556] = 2130578706;
assign addr[61557] = 2132888897;
assign addr[61558] = 2135029962;
assign addr[61559] = 2137001733;
assign addr[61560] = 2138804053;
assign addr[61561] = 2140436778;
assign addr[61562] = 2141899780;
assign addr[61563] = 2143192942;
assign addr[61564] = 2144316162;
assign addr[61565] = 2145269351;
assign addr[61566] = 2146052433;
assign addr[61567] = 2146665347;
assign addr[61568] = 2147108043;
assign addr[61569] = 2147380486;
assign addr[61570] = 2147482655;
assign addr[61571] = 2147414542;
assign addr[61572] = 2147176152;
assign addr[61573] = 2146767505;
assign addr[61574] = 2146188631;
assign addr[61575] = 2145439578;
assign addr[61576] = 2144520405;
assign addr[61577] = 2143431184;
assign addr[61578] = 2142172003;
assign addr[61579] = 2140742960;
assign addr[61580] = 2139144169;
assign addr[61581] = 2137375758;
assign addr[61582] = 2135437865;
assign addr[61583] = 2133330646;
assign addr[61584] = 2131054266;
assign addr[61585] = 2128608907;
assign addr[61586] = 2125994762;
assign addr[61587] = 2123212038;
assign addr[61588] = 2120260957;
assign addr[61589] = 2117141752;
assign addr[61590] = 2113854671;
assign addr[61591] = 2110399974;
assign addr[61592] = 2106777935;
assign addr[61593] = 2102988841;
assign addr[61594] = 2099032994;
assign addr[61595] = 2094910706;
assign addr[61596] = 2090622304;
assign addr[61597] = 2086168128;
assign addr[61598] = 2081548533;
assign addr[61599] = 2076763883;
assign addr[61600] = 2071814558;
assign addr[61601] = 2066700952;
assign addr[61602] = 2061423468;
assign addr[61603] = 2055982526;
assign addr[61604] = 2050378558;
assign addr[61605] = 2044612007;
assign addr[61606] = 2038683330;
assign addr[61607] = 2032592999;
assign addr[61608] = 2026341495;
assign addr[61609] = 2019929315;
assign addr[61610] = 2013356967;
assign addr[61611] = 2006624971;
assign addr[61612] = 1999733863;
assign addr[61613] = 1992684188;
assign addr[61614] = 1985476506;
assign addr[61615] = 1978111387;
assign addr[61616] = 1970589416;
assign addr[61617] = 1962911189;
assign addr[61618] = 1955077316;
assign addr[61619] = 1947088417;
assign addr[61620] = 1938945125;
assign addr[61621] = 1930648088;
assign addr[61622] = 1922197961;
assign addr[61623] = 1913595416;
assign addr[61624] = 1904841135;
assign addr[61625] = 1895935811;
assign addr[61626] = 1886880151;
assign addr[61627] = 1877674873;
assign addr[61628] = 1868320707;
assign addr[61629] = 1858818395;
assign addr[61630] = 1849168689;
assign addr[61631] = 1839372356;
assign addr[61632] = 1829430172;
assign addr[61633] = 1819342925;
assign addr[61634] = 1809111415;
assign addr[61635] = 1798736454;
assign addr[61636] = 1788218865;
assign addr[61637] = 1777559480;
assign addr[61638] = 1766759146;
assign addr[61639] = 1755818718;
assign addr[61640] = 1744739065;
assign addr[61641] = 1733521064;
assign addr[61642] = 1722165606;
assign addr[61643] = 1710673591;
assign addr[61644] = 1699045930;
assign addr[61645] = 1687283545;
assign addr[61646] = 1675387369;
assign addr[61647] = 1663358344;
assign addr[61648] = 1651197426;
assign addr[61649] = 1638905577;
assign addr[61650] = 1626483774;
assign addr[61651] = 1613933000;
assign addr[61652] = 1601254251;
assign addr[61653] = 1588448533;
assign addr[61654] = 1575516860;
assign addr[61655] = 1562460258;
assign addr[61656] = 1549279763;
assign addr[61657] = 1535976419;
assign addr[61658] = 1522551282;
assign addr[61659] = 1509005416;
assign addr[61660] = 1495339895;
assign addr[61661] = 1481555802;
assign addr[61662] = 1467654232;
assign addr[61663] = 1453636285;
assign addr[61664] = 1439503074;
assign addr[61665] = 1425255719;
assign addr[61666] = 1410895350;
assign addr[61667] = 1396423105;
assign addr[61668] = 1381840133;
assign addr[61669] = 1367147589;
assign addr[61670] = 1352346639;
assign addr[61671] = 1337438456;
assign addr[61672] = 1322424222;
assign addr[61673] = 1307305128;
assign addr[61674] = 1292082373;
assign addr[61675] = 1276757164;
assign addr[61676] = 1261330715;
assign addr[61677] = 1245804251;
assign addr[61678] = 1230179002;
assign addr[61679] = 1214456207;
assign addr[61680] = 1198637114;
assign addr[61681] = 1182722976;
assign addr[61682] = 1166715055;
assign addr[61683] = 1150614620;
assign addr[61684] = 1134422949;
assign addr[61685] = 1118141326;
assign addr[61686] = 1101771040;
assign addr[61687] = 1085313391;
assign addr[61688] = 1068769683;
assign addr[61689] = 1052141228;
assign addr[61690] = 1035429345;
assign addr[61691] = 1018635358;
assign addr[61692] = 1001760600;
assign addr[61693] = 984806408;
assign addr[61694] = 967774128;
assign addr[61695] = 950665109;
assign addr[61696] = 933480707;
assign addr[61697] = 916222287;
assign addr[61698] = 898891215;
assign addr[61699] = 881488868;
assign addr[61700] = 864016623;
assign addr[61701] = 846475867;
assign addr[61702] = 828867991;
assign addr[61703] = 811194391;
assign addr[61704] = 793456467;
assign addr[61705] = 775655628;
assign addr[61706] = 757793284;
assign addr[61707] = 739870851;
assign addr[61708] = 721889752;
assign addr[61709] = 703851410;
assign addr[61710] = 685757258;
assign addr[61711] = 667608730;
assign addr[61712] = 649407264;
assign addr[61713] = 631154304;
assign addr[61714] = 612851297;
assign addr[61715] = 594499695;
assign addr[61716] = 576100953;
assign addr[61717] = 557656529;
assign addr[61718] = 539167887;
assign addr[61719] = 520636492;
assign addr[61720] = 502063814;
assign addr[61721] = 483451325;
assign addr[61722] = 464800501;
assign addr[61723] = 446112822;
assign addr[61724] = 427389768;
assign addr[61725] = 408632825;
assign addr[61726] = 389843480;
assign addr[61727] = 371023223;
assign addr[61728] = 352173546;
assign addr[61729] = 333295944;
assign addr[61730] = 314391913;
assign addr[61731] = 295462954;
assign addr[61732] = 276510565;
assign addr[61733] = 257536251;
assign addr[61734] = 238541516;
assign addr[61735] = 219527866;
assign addr[61736] = 200496809;
assign addr[61737] = 181449854;
assign addr[61738] = 162388511;
assign addr[61739] = 143314291;
assign addr[61740] = 124228708;
assign addr[61741] = 105133274;
assign addr[61742] = 86029503;
assign addr[61743] = 66918911;
assign addr[61744] = 47803013;
assign addr[61745] = 28683324;
assign addr[61746] = 9561361;
assign addr[61747] = -9561361;
assign addr[61748] = -28683324;
assign addr[61749] = -47803013;
assign addr[61750] = -66918911;
assign addr[61751] = -86029503;
assign addr[61752] = -105133274;
assign addr[61753] = -124228708;
assign addr[61754] = -143314291;
assign addr[61755] = -162388511;
assign addr[61756] = -181449854;
assign addr[61757] = -200496809;
assign addr[61758] = -219527866;
assign addr[61759] = -238541516;
assign addr[61760] = -257536251;
assign addr[61761] = -276510565;
assign addr[61762] = -295462953;
assign addr[61763] = -314391913;
assign addr[61764] = -333295944;
assign addr[61765] = -352173546;
assign addr[61766] = -371023223;
assign addr[61767] = -389843480;
assign addr[61768] = -408632825;
assign addr[61769] = -427389768;
assign addr[61770] = -446112822;
assign addr[61771] = -464800501;
assign addr[61772] = -483451325;
assign addr[61773] = -502063814;
assign addr[61774] = -520636492;
assign addr[61775] = -539167887;
assign addr[61776] = -557656529;
assign addr[61777] = -576100953;
assign addr[61778] = -594499695;
assign addr[61779] = -612851297;
assign addr[61780] = -631154304;
assign addr[61781] = -649407264;
assign addr[61782] = -667608730;
assign addr[61783] = -685757258;
assign addr[61784] = -703851410;
assign addr[61785] = -721889752;
assign addr[61786] = -739870851;
assign addr[61787] = -757793284;
assign addr[61788] = -775655628;
assign addr[61789] = -793456467;
assign addr[61790] = -811194391;
assign addr[61791] = -828867991;
assign addr[61792] = -846475867;
assign addr[61793] = -864016623;
assign addr[61794] = -881488868;
assign addr[61795] = -898891215;
assign addr[61796] = -916222287;
assign addr[61797] = -933480707;
assign addr[61798] = -950665109;
assign addr[61799] = -967774128;
assign addr[61800] = -984806408;
assign addr[61801] = -1001760600;
assign addr[61802] = -1018635358;
assign addr[61803] = -1035429345;
assign addr[61804] = -1052141228;
assign addr[61805] = -1068769683;
assign addr[61806] = -1085313391;
assign addr[61807] = -1101771040;
assign addr[61808] = -1118141326;
assign addr[61809] = -1134422949;
assign addr[61810] = -1150614620;
assign addr[61811] = -1166715055;
assign addr[61812] = -1182722976;
assign addr[61813] = -1198637114;
assign addr[61814] = -1214456207;
assign addr[61815] = -1230179002;
assign addr[61816] = -1245804251;
assign addr[61817] = -1261330715;
assign addr[61818] = -1276757164;
assign addr[61819] = -1292082373;
assign addr[61820] = -1307305128;
assign addr[61821] = -1322424222;
assign addr[61822] = -1337438456;
assign addr[61823] = -1352346639;
assign addr[61824] = -1367147589;
assign addr[61825] = -1381840133;
assign addr[61826] = -1396423105;
assign addr[61827] = -1410895350;
assign addr[61828] = -1425255719;
assign addr[61829] = -1439503074;
assign addr[61830] = -1453636285;
assign addr[61831] = -1467654232;
assign addr[61832] = -1481555802;
assign addr[61833] = -1495339895;
assign addr[61834] = -1509005416;
assign addr[61835] = -1522551282;
assign addr[61836] = -1535976419;
assign addr[61837] = -1549279763;
assign addr[61838] = -1562460258;
assign addr[61839] = -1575516860;
assign addr[61840] = -1588448533;
assign addr[61841] = -1601254251;
assign addr[61842] = -1613933000;
assign addr[61843] = -1626483774;
assign addr[61844] = -1638905577;
assign addr[61845] = -1651197426;
assign addr[61846] = -1663358344;
assign addr[61847] = -1675387369;
assign addr[61848] = -1687283545;
assign addr[61849] = -1699045930;
assign addr[61850] = -1710673591;
assign addr[61851] = -1722165606;
assign addr[61852] = -1733521064;
assign addr[61853] = -1744739065;
assign addr[61854] = -1755818718;
assign addr[61855] = -1766759146;
assign addr[61856] = -1777559480;
assign addr[61857] = -1788218865;
assign addr[61858] = -1798736454;
assign addr[61859] = -1809111415;
assign addr[61860] = -1819342925;
assign addr[61861] = -1829430172;
assign addr[61862] = -1839372356;
assign addr[61863] = -1849168689;
assign addr[61864] = -1858818395;
assign addr[61865] = -1868320707;
assign addr[61866] = -1877674873;
assign addr[61867] = -1886880151;
assign addr[61868] = -1895935811;
assign addr[61869] = -1904841135;
assign addr[61870] = -1913595416;
assign addr[61871] = -1922197961;
assign addr[61872] = -1930648088;
assign addr[61873] = -1938945125;
assign addr[61874] = -1947088417;
assign addr[61875] = -1955077316;
assign addr[61876] = -1962911189;
assign addr[61877] = -1970589416;
assign addr[61878] = -1978111387;
assign addr[61879] = -1985476506;
assign addr[61880] = -1992684188;
assign addr[61881] = -1999733863;
assign addr[61882] = -2006624971;
assign addr[61883] = -2013356967;
assign addr[61884] = -2019929315;
assign addr[61885] = -2026341495;
assign addr[61886] = -2032592999;
assign addr[61887] = -2038683330;
assign addr[61888] = -2044612007;
assign addr[61889] = -2050378558;
assign addr[61890] = -2055982526;
assign addr[61891] = -2061423468;
assign addr[61892] = -2066700952;
assign addr[61893] = -2071814558;
assign addr[61894] = -2076763883;
assign addr[61895] = -2081548533;
assign addr[61896] = -2086168128;
assign addr[61897] = -2090622304;
assign addr[61898] = -2094910706;
assign addr[61899] = -2099032994;
assign addr[61900] = -2102988841;
assign addr[61901] = -2106777935;
assign addr[61902] = -2110399974;
assign addr[61903] = -2113854671;
assign addr[61904] = -2117141752;
assign addr[61905] = -2120260957;
assign addr[61906] = -2123212038;
assign addr[61907] = -2125994762;
assign addr[61908] = -2128608907;
assign addr[61909] = -2131054266;
assign addr[61910] = -2133330646;
assign addr[61911] = -2135437865;
assign addr[61912] = -2137375758;
assign addr[61913] = -2139144169;
assign addr[61914] = -2140742960;
assign addr[61915] = -2142172003;
assign addr[61916] = -2143431184;
assign addr[61917] = -2144520405;
assign addr[61918] = -2145439578;
assign addr[61919] = -2146188631;
assign addr[61920] = -2146767505;
assign addr[61921] = -2147176152;
assign addr[61922] = -2147414542;
assign addr[61923] = -2147482655;
assign addr[61924] = -2147380486;
assign addr[61925] = -2147108043;
assign addr[61926] = -2146665347;
assign addr[61927] = -2146052433;
assign addr[61928] = -2145269351;
assign addr[61929] = -2144316162;
assign addr[61930] = -2143192942;
assign addr[61931] = -2141899780;
assign addr[61932] = -2140436778;
assign addr[61933] = -2138804053;
assign addr[61934] = -2137001733;
assign addr[61935] = -2135029962;
assign addr[61936] = -2132888897;
assign addr[61937] = -2130578706;
assign addr[61938] = -2128099574;
assign addr[61939] = -2125451696;
assign addr[61940] = -2122635283;
assign addr[61941] = -2119650558;
assign addr[61942] = -2116497758;
assign addr[61943] = -2113177132;
assign addr[61944] = -2109688944;
assign addr[61945] = -2106033471;
assign addr[61946] = -2102211002;
assign addr[61947] = -2098221841;
assign addr[61948] = -2094066304;
assign addr[61949] = -2089744719;
assign addr[61950] = -2085257431;
assign addr[61951] = -2080604795;
assign addr[61952] = -2075787180;
assign addr[61953] = -2070804967;
assign addr[61954] = -2065658552;
assign addr[61955] = -2060348343;
assign addr[61956] = -2054874761;
assign addr[61957] = -2049238240;
assign addr[61958] = -2043439226;
assign addr[61959] = -2037478181;
assign addr[61960] = -2031355576;
assign addr[61961] = -2025071897;
assign addr[61962] = -2018627642;
assign addr[61963] = -2012023322;
assign addr[61964] = -2005259462;
assign addr[61965] = -1998336596;
assign addr[61966] = -1991255274;
assign addr[61967] = -1984016058;
assign addr[61968] = -1976619522;
assign addr[61969] = -1969066252;
assign addr[61970] = -1961356847;
assign addr[61971] = -1953491918;
assign addr[61972] = -1945472089;
assign addr[61973] = -1937297997;
assign addr[61974] = -1928970288;
assign addr[61975] = -1920489624;
assign addr[61976] = -1911856677;
assign addr[61977] = -1903072131;
assign addr[61978] = -1894136683;
assign addr[61979] = -1885051042;
assign addr[61980] = -1875815927;
assign addr[61981] = -1866432072;
assign addr[61982] = -1856900221;
assign addr[61983] = -1847221128;
assign addr[61984] = -1837395562;
assign addr[61985] = -1827424302;
assign addr[61986] = -1817308138;
assign addr[61987] = -1807047873;
assign addr[61988] = -1796644320;
assign addr[61989] = -1786098304;
assign addr[61990] = -1775410662;
assign addr[61991] = -1764582240;
assign addr[61992] = -1753613897;
assign addr[61993] = -1742506504;
assign addr[61994] = -1731260941;
assign addr[61995] = -1719878099;
assign addr[61996] = -1708358881;
assign addr[61997] = -1696704201;
assign addr[61998] = -1684914983;
assign addr[61999] = -1672992161;
assign addr[62000] = -1660936681;
assign addr[62001] = -1648749499;
assign addr[62002] = -1636431582;
assign addr[62003] = -1623983905;
assign addr[62004] = -1611407456;
assign addr[62005] = -1598703233;
assign addr[62006] = -1585872242;
assign addr[62007] = -1572915501;
assign addr[62008] = -1559834037;
assign addr[62009] = -1546628888;
assign addr[62010] = -1533301101;
assign addr[62011] = -1519851733;
assign addr[62012] = -1506281850;
assign addr[62013] = -1492592527;
assign addr[62014] = -1478784851;
assign addr[62015] = -1464859917;
assign addr[62016] = -1450818828;
assign addr[62017] = -1436662698;
assign addr[62018] = -1422392650;
assign addr[62019] = -1408009814;
assign addr[62020] = -1393515332;
assign addr[62021] = -1378910353;
assign addr[62022] = -1364196034;
assign addr[62023] = -1349373543;
assign addr[62024] = -1334444055;
assign addr[62025] = -1319408754;
assign addr[62026] = -1304268832;
assign addr[62027] = -1289025489;
assign addr[62028] = -1273679934;
assign addr[62029] = -1258233384;
assign addr[62030] = -1242687064;
assign addr[62031] = -1227042207;
assign addr[62032] = -1211300053;
assign addr[62033] = -1195461849;
assign addr[62034] = -1179528853;
assign addr[62035] = -1163502328;
assign addr[62036] = -1147383544;
assign addr[62037] = -1131173780;
assign addr[62038] = -1114874320;
assign addr[62039] = -1098486458;
assign addr[62040] = -1082011492;
assign addr[62041] = -1065450729;
assign addr[62042] = -1048805483;
assign addr[62043] = -1032077073;
assign addr[62044] = -1015266825;
assign addr[62045] = -998376073;
assign addr[62046] = -981406156;
assign addr[62047] = -964358420;
assign addr[62048] = -947234215;
assign addr[62049] = -930034901;
assign addr[62050] = -912761841;
assign addr[62051] = -895416404;
assign addr[62052] = -877999966;
assign addr[62053] = -860513908;
assign addr[62054] = -842959617;
assign addr[62055] = -825338484;
assign addr[62056] = -807651907;
assign addr[62057] = -789901288;
assign addr[62058] = -772088034;
assign addr[62059] = -754213559;
assign addr[62060] = -736279279;
assign addr[62061] = -718286617;
assign addr[62062] = -700236999;
assign addr[62063] = -682131857;
assign addr[62064] = -663972625;
assign addr[62065] = -645760745;
assign addr[62066] = -627497660;
assign addr[62067] = -609184818;
assign addr[62068] = -590823671;
assign addr[62069] = -572415676;
assign addr[62070] = -553962291;
assign addr[62071] = -535464981;
assign addr[62072] = -516925212;
assign addr[62073] = -498344454;
assign addr[62074] = -479724180;
assign addr[62075] = -461065866;
assign addr[62076] = -442370993;
assign addr[62077] = -423641043;
assign addr[62078] = -404877501;
assign addr[62079] = -386081854;
assign addr[62080] = -367255594;
assign addr[62081] = -348400212;
assign addr[62082] = -329517204;
assign addr[62083] = -310608068;
assign addr[62084] = -291674302;
assign addr[62085] = -272717408;
assign addr[62086] = -253738890;
assign addr[62087] = -234740251;
assign addr[62088] = -215722999;
assign addr[62089] = -196688642;
assign addr[62090] = -177638688;
assign addr[62091] = -158574649;
assign addr[62092] = -139498035;
assign addr[62093] = -120410361;
assign addr[62094] = -101313138;
assign addr[62095] = -82207882;
assign addr[62096] = -63096108;
assign addr[62097] = -43979330;
assign addr[62098] = -24859065;
assign addr[62099] = -5736829;
assign addr[62100] = 13385863;
assign addr[62101] = 32507492;
assign addr[62102] = 51626544;
assign addr[62103] = 70741503;
assign addr[62104] = 89850852;
assign addr[62105] = 108953076;
assign addr[62106] = 128046661;
assign addr[62107] = 147130093;
assign addr[62108] = 166201858;
assign addr[62109] = 185260444;
assign addr[62110] = 204304341;
assign addr[62111] = 223332037;
assign addr[62112] = 242342025;
assign addr[62113] = 261332796;
assign addr[62114] = 280302845;
assign addr[62115] = 299250668;
assign addr[62116] = 318174762;
assign addr[62117] = 337073627;
assign addr[62118] = 355945764;
assign addr[62119] = 374789676;
assign addr[62120] = 393603870;
assign addr[62121] = 412386854;
assign addr[62122] = 431137138;
assign addr[62123] = 449853235;
assign addr[62124] = 468533662;
assign addr[62125] = 487176937;
assign addr[62126] = 505781581;
assign addr[62127] = 524346121;
assign addr[62128] = 542869083;
assign addr[62129] = 561348998;
assign addr[62130] = 579784402;
assign addr[62131] = 598173833;
assign addr[62132] = 616515832;
assign addr[62133] = 634808946;
assign addr[62134] = 653051723;
assign addr[62135] = 671242716;
assign addr[62136] = 689380485;
assign addr[62137] = 707463589;
assign addr[62138] = 725490597;
assign addr[62139] = 743460077;
assign addr[62140] = 761370605;
assign addr[62141] = 779220762;
assign addr[62142] = 797009130;
assign addr[62143] = 814734301;
assign addr[62144] = 832394869;
assign addr[62145] = 849989433;
assign addr[62146] = 867516597;
assign addr[62147] = 884974973;
assign addr[62148] = 902363176;
assign addr[62149] = 919679827;
assign addr[62150] = 936923553;
assign addr[62151] = 954092986;
assign addr[62152] = 971186766;
assign addr[62153] = 988203537;
assign addr[62154] = 1005141949;
assign addr[62155] = 1022000660;
assign addr[62156] = 1038778332;
assign addr[62157] = 1055473635;
assign addr[62158] = 1072085246;
assign addr[62159] = 1088611847;
assign addr[62160] = 1105052128;
assign addr[62161] = 1121404785;
assign addr[62162] = 1137668521;
assign addr[62163] = 1153842047;
assign addr[62164] = 1169924081;
assign addr[62165] = 1185913346;
assign addr[62166] = 1201808576;
assign addr[62167] = 1217608510;
assign addr[62168] = 1233311895;
assign addr[62169] = 1248917486;
assign addr[62170] = 1264424045;
assign addr[62171] = 1279830344;
assign addr[62172] = 1295135159;
assign addr[62173] = 1310337279;
assign addr[62174] = 1325435496;
assign addr[62175] = 1340428615;
assign addr[62176] = 1355315445;
assign addr[62177] = 1370094808;
assign addr[62178] = 1384765530;
assign addr[62179] = 1399326449;
assign addr[62180] = 1413776410;
assign addr[62181] = 1428114267;
assign addr[62182] = 1442338884;
assign addr[62183] = 1456449131;
assign addr[62184] = 1470443891;
assign addr[62185] = 1484322054;
assign addr[62186] = 1498082520;
assign addr[62187] = 1511724196;
assign addr[62188] = 1525246002;
assign addr[62189] = 1538646865;
assign addr[62190] = 1551925723;
assign addr[62191] = 1565081523;
assign addr[62192] = 1578113222;
assign addr[62193] = 1591019785;
assign addr[62194] = 1603800191;
assign addr[62195] = 1616453425;
assign addr[62196] = 1628978484;
assign addr[62197] = 1641374375;
assign addr[62198] = 1653640115;
assign addr[62199] = 1665774731;
assign addr[62200] = 1677777262;
assign addr[62201] = 1689646755;
assign addr[62202] = 1701382270;
assign addr[62203] = 1712982875;
assign addr[62204] = 1724447652;
assign addr[62205] = 1735775690;
assign addr[62206] = 1746966091;
assign addr[62207] = 1758017969;
assign addr[62208] = 1768930447;
assign addr[62209] = 1779702660;
assign addr[62210] = 1790333753;
assign addr[62211] = 1800822883;
assign addr[62212] = 1811169220;
assign addr[62213] = 1821371941;
assign addr[62214] = 1831430239;
assign addr[62215] = 1841343316;
assign addr[62216] = 1851110385;
assign addr[62217] = 1860730673;
assign addr[62218] = 1870203416;
assign addr[62219] = 1879527863;
assign addr[62220] = 1888703276;
assign addr[62221] = 1897728925;
assign addr[62222] = 1906604097;
assign addr[62223] = 1915328086;
assign addr[62224] = 1923900201;
assign addr[62225] = 1932319763;
assign addr[62226] = 1940586104;
assign addr[62227] = 1948698568;
assign addr[62228] = 1956656513;
assign addr[62229] = 1964459306;
assign addr[62230] = 1972106330;
assign addr[62231] = 1979596978;
assign addr[62232] = 1986930656;
assign addr[62233] = 1994106782;
assign addr[62234] = 2001124788;
assign addr[62235] = 2007984117;
assign addr[62236] = 2014684225;
assign addr[62237] = 2021224581;
assign addr[62238] = 2027604666;
assign addr[62239] = 2033823974;
assign addr[62240] = 2039882013;
assign addr[62241] = 2045778302;
assign addr[62242] = 2051512372;
assign addr[62243] = 2057083771;
assign addr[62244] = 2062492055;
assign addr[62245] = 2067736796;
assign addr[62246] = 2072817579;
assign addr[62247] = 2077733999;
assign addr[62248] = 2082485668;
assign addr[62249] = 2087072209;
assign addr[62250] = 2091493257;
assign addr[62251] = 2095748463;
assign addr[62252] = 2099837489;
assign addr[62253] = 2103760010;
assign addr[62254] = 2107515716;
assign addr[62255] = 2111104309;
assign addr[62256] = 2114525505;
assign addr[62257] = 2117779031;
assign addr[62258] = 2120864631;
assign addr[62259] = 2123782059;
assign addr[62260] = 2126531084;
assign addr[62261] = 2129111488;
assign addr[62262] = 2131523066;
assign addr[62263] = 2133765628;
assign addr[62264] = 2135838995;
assign addr[62265] = 2137743003;
assign addr[62266] = 2139477502;
assign addr[62267] = 2141042352;
assign addr[62268] = 2142437431;
assign addr[62269] = 2143662628;
assign addr[62270] = 2144717846;
assign addr[62271] = 2145603001;
assign addr[62272] = 2146318022;
assign addr[62273] = 2146862854;
assign addr[62274] = 2147237452;
assign addr[62275] = 2147441787;
assign addr[62276] = 2147475844;
assign addr[62277] = 2147339619;
assign addr[62278] = 2147033123;
assign addr[62279] = 2146556380;
assign addr[62280] = 2145909429;
assign addr[62281] = 2145092320;
assign addr[62282] = 2144105118;
assign addr[62283] = 2142947902;
assign addr[62284] = 2141620763;
assign addr[62285] = 2140123807;
assign addr[62286] = 2138457152;
assign addr[62287] = 2136620930;
assign addr[62288] = 2134615288;
assign addr[62289] = 2132440383;
assign addr[62290] = 2130096389;
assign addr[62291] = 2127583492;
assign addr[62292] = 2124901890;
assign addr[62293] = 2122051796;
assign addr[62294] = 2119033436;
assign addr[62295] = 2115847050;
assign addr[62296] = 2112492891;
assign addr[62297] = 2108971223;
assign addr[62298] = 2105282327;
assign addr[62299] = 2101426496;
assign addr[62300] = 2097404033;
assign addr[62301] = 2093215260;
assign addr[62302] = 2088860507;
assign addr[62303] = 2084340120;
assign addr[62304] = 2079654458;
assign addr[62305] = 2074803892;
assign addr[62306] = 2069788807;
assign addr[62307] = 2064609600;
assign addr[62308] = 2059266683;
assign addr[62309] = 2053760478;
assign addr[62310] = 2048091422;
assign addr[62311] = 2042259965;
assign addr[62312] = 2036266570;
assign addr[62313] = 2030111710;
assign addr[62314] = 2023795876;
assign addr[62315] = 2017319567;
assign addr[62316] = 2010683297;
assign addr[62317] = 2003887591;
assign addr[62318] = 1996932990;
assign addr[62319] = 1989820044;
assign addr[62320] = 1982549318;
assign addr[62321] = 1975121388;
assign addr[62322] = 1967536842;
assign addr[62323] = 1959796283;
assign addr[62324] = 1951900324;
assign addr[62325] = 1943849591;
assign addr[62326] = 1935644723;
assign addr[62327] = 1927286370;
assign addr[62328] = 1918775195;
assign addr[62329] = 1910111873;
assign addr[62330] = 1901297091;
assign addr[62331] = 1892331547;
assign addr[62332] = 1883215953;
assign addr[62333] = 1873951032;
assign addr[62334] = 1864537518;
assign addr[62335] = 1854976157;
assign addr[62336] = 1845267708;
assign addr[62337] = 1835412941;
assign addr[62338] = 1825412636;
assign addr[62339] = 1815267588;
assign addr[62340] = 1804978599;
assign addr[62341] = 1794546487;
assign addr[62342] = 1783972079;
assign addr[62343] = 1773256212;
assign addr[62344] = 1762399737;
assign addr[62345] = 1751403515;
assign addr[62346] = 1740268417;
assign addr[62347] = 1728995326;
assign addr[62348] = 1717585136;
assign addr[62349] = 1706038753;
assign addr[62350] = 1694357091;
assign addr[62351] = 1682541077;
assign addr[62352] = 1670591647;
assign addr[62353] = 1658509750;
assign addr[62354] = 1646296344;
assign addr[62355] = 1633952396;
assign addr[62356] = 1621478885;
assign addr[62357] = 1608876801;
assign addr[62358] = 1596147143;
assign addr[62359] = 1583290921;
assign addr[62360] = 1570309153;
assign addr[62361] = 1557202869;
assign addr[62362] = 1543973108;
assign addr[62363] = 1530620920;
assign addr[62364] = 1517147363;
assign addr[62365] = 1503553506;
assign addr[62366] = 1489840425;
assign addr[62367] = 1476009210;
assign addr[62368] = 1462060956;
assign addr[62369] = 1447996770;
assign addr[62370] = 1433817766;
assign addr[62371] = 1419525069;
assign addr[62372] = 1405119813;
assign addr[62373] = 1390603139;
assign addr[62374] = 1375976199;
assign addr[62375] = 1361240152;
assign addr[62376] = 1346396168;
assign addr[62377] = 1331445422;
assign addr[62378] = 1316389101;
assign addr[62379] = 1301228398;
assign addr[62380] = 1285964516;
assign addr[62381] = 1270598665;
assign addr[62382] = 1255132063;
assign addr[62383] = 1239565936;
assign addr[62384] = 1223901520;
assign addr[62385] = 1208140056;
assign addr[62386] = 1192282793;
assign addr[62387] = 1176330990;
assign addr[62388] = 1160285911;
assign addr[62389] = 1144148829;
assign addr[62390] = 1127921022;
assign addr[62391] = 1111603778;
assign addr[62392] = 1095198391;
assign addr[62393] = 1078706161;
assign addr[62394] = 1062128397;
assign addr[62395] = 1045466412;
assign addr[62396] = 1028721528;
assign addr[62397] = 1011895073;
assign addr[62398] = 994988380;
assign addr[62399] = 978002791;
assign addr[62400] = 960939653;
assign addr[62401] = 943800318;
assign addr[62402] = 926586145;
assign addr[62403] = 909298500;
assign addr[62404] = 891938752;
assign addr[62405] = 874508280;
assign addr[62406] = 857008464;
assign addr[62407] = 839440693;
assign addr[62408] = 821806359;
assign addr[62409] = 804106861;
assign addr[62410] = 786343603;
assign addr[62411] = 768517992;
assign addr[62412] = 750631442;
assign addr[62413] = 732685372;
assign addr[62414] = 714681204;
assign addr[62415] = 696620367;
assign addr[62416] = 678504291;
assign addr[62417] = 660334415;
assign addr[62418] = 642112178;
assign addr[62419] = 623839025;
assign addr[62420] = 605516406;
assign addr[62421] = 587145773;
assign addr[62422] = 568728583;
assign addr[62423] = 550266296;
assign addr[62424] = 531760377;
assign addr[62425] = 513212292;
assign addr[62426] = 494623513;
assign addr[62427] = 475995513;
assign addr[62428] = 457329769;
assign addr[62429] = 438627762;
assign addr[62430] = 419890975;
assign addr[62431] = 401120892;
assign addr[62432] = 382319004;
assign addr[62433] = 363486799;
assign addr[62434] = 344625773;
assign addr[62435] = 325737419;
assign addr[62436] = 306823237;
assign addr[62437] = 287884725;
assign addr[62438] = 268923386;
assign addr[62439] = 249940723;
assign addr[62440] = 230938242;
assign addr[62441] = 211917448;
assign addr[62442] = 192879850;
assign addr[62443] = 173826959;
assign addr[62444] = 154760284;
assign addr[62445] = 135681337;
assign addr[62446] = 116591632;
assign addr[62447] = 97492681;
assign addr[62448] = 78386000;
assign addr[62449] = 59273104;
assign addr[62450] = 40155507;
assign addr[62451] = 21034727;
assign addr[62452] = 1912278;
assign addr[62453] = -17210322;
assign addr[62454] = -36331557;
assign addr[62455] = -55449912;
assign addr[62456] = -74563870;
assign addr[62457] = -93671915;
assign addr[62458] = -112772533;
assign addr[62459] = -131864208;
assign addr[62460] = -150945428;
assign addr[62461] = -170014678;
assign addr[62462] = -189070447;
assign addr[62463] = -208111224;
assign addr[62464] = -227135500;
assign addr[62465] = -246141764;
assign addr[62466] = -265128512;
assign addr[62467] = -284094236;
assign addr[62468] = -303037433;
assign addr[62469] = -321956601;
assign addr[62470] = -340850240;
assign addr[62471] = -359716852;
assign addr[62472] = -378554940;
assign addr[62473] = -397363011;
assign addr[62474] = -416139574;
assign addr[62475] = -434883140;
assign addr[62476] = -453592221;
assign addr[62477] = -472265336;
assign addr[62478] = -490901003;
assign addr[62479] = -509497745;
assign addr[62480] = -528054086;
assign addr[62481] = -546568556;
assign addr[62482] = -565039687;
assign addr[62483] = -583466013;
assign addr[62484] = -601846074;
assign addr[62485] = -620178412;
assign addr[62486] = -638461574;
assign addr[62487] = -656694110;
assign addr[62488] = -674874574;
assign addr[62489] = -693001525;
assign addr[62490] = -711073524;
assign addr[62491] = -729089140;
assign addr[62492] = -747046944;
assign addr[62493] = -764945512;
assign addr[62494] = -782783424;
assign addr[62495] = -800559266;
assign addr[62496] = -818271628;
assign addr[62497] = -835919107;
assign addr[62498] = -853500302;
assign addr[62499] = -871013820;
assign addr[62500] = -888458272;
assign addr[62501] = -905832274;
assign addr[62502] = -923134450;
assign addr[62503] = -940363427;
assign addr[62504] = -957517838;
assign addr[62505] = -974596324;
assign addr[62506] = -991597531;
assign addr[62507] = -1008520110;
assign addr[62508] = -1025362720;
assign addr[62509] = -1042124025;
assign addr[62510] = -1058802695;
assign addr[62511] = -1075397409;
assign addr[62512] = -1091906851;
assign addr[62513] = -1108329711;
assign addr[62514] = -1124664687;
assign addr[62515] = -1140910484;
assign addr[62516] = -1157065814;
assign addr[62517] = -1173129396;
assign addr[62518] = -1189099956;
assign addr[62519] = -1204976227;
assign addr[62520] = -1220756951;
assign addr[62521] = -1236440877;
assign addr[62522] = -1252026760;
assign addr[62523] = -1267513365;
assign addr[62524] = -1282899464;
assign addr[62525] = -1298183838;
assign addr[62526] = -1313365273;
assign addr[62527] = -1328442566;
assign addr[62528] = -1343414522;
assign addr[62529] = -1358279953;
assign addr[62530] = -1373037681;
assign addr[62531] = -1387686535;
assign addr[62532] = -1402225355;
assign addr[62533] = -1416652986;
assign addr[62534] = -1430968286;
assign addr[62535] = -1445170118;
assign addr[62536] = -1459257358;
assign addr[62537] = -1473228887;
assign addr[62538] = -1487083598;
assign addr[62539] = -1500820393;
assign addr[62540] = -1514438181;
assign addr[62541] = -1527935884;
assign addr[62542] = -1541312431;
assign addr[62543] = -1554566762;
assign addr[62544] = -1567697824;
assign addr[62545] = -1580704578;
assign addr[62546] = -1593585992;
assign addr[62547] = -1606341043;
assign addr[62548] = -1618968722;
assign addr[62549] = -1631468027;
assign addr[62550] = -1643837966;
assign addr[62551] = -1656077559;
assign addr[62552] = -1668185835;
assign addr[62553] = -1680161834;
assign addr[62554] = -1692004606;
assign addr[62555] = -1703713213;
assign addr[62556] = -1715286726;
assign addr[62557] = -1726724227;
assign addr[62558] = -1738024810;
assign addr[62559] = -1749187577;
assign addr[62560] = -1760211645;
assign addr[62561] = -1771096139;
assign addr[62562] = -1781840195;
assign addr[62563] = -1792442963;
assign addr[62564] = -1802903601;
assign addr[62565] = -1813221279;
assign addr[62566] = -1823395180;
assign addr[62567] = -1833424497;
assign addr[62568] = -1843308435;
assign addr[62569] = -1853046210;
assign addr[62570] = -1862637049;
assign addr[62571] = -1872080193;
assign addr[62572] = -1881374892;
assign addr[62573] = -1890520410;
assign addr[62574] = -1899516021;
assign addr[62575] = -1908361011;
assign addr[62576] = -1917054681;
assign addr[62577] = -1925596340;
assign addr[62578] = -1933985310;
assign addr[62579] = -1942220928;
assign addr[62580] = -1950302539;
assign addr[62581] = -1958229503;
assign addr[62582] = -1966001192;
assign addr[62583] = -1973616989;
assign addr[62584] = -1981076290;
assign addr[62585] = -1988378503;
assign addr[62586] = -1995523051;
assign addr[62587] = -2002509365;
assign addr[62588] = -2009336893;
assign addr[62589] = -2016005093;
assign addr[62590] = -2022513436;
assign addr[62591] = -2028861406;
assign addr[62592] = -2035048499;
assign addr[62593] = -2041074226;
assign addr[62594] = -2046938108;
assign addr[62595] = -2052639680;
assign addr[62596] = -2058178491;
assign addr[62597] = -2063554100;
assign addr[62598] = -2068766083;
assign addr[62599] = -2073814024;
assign addr[62600] = -2078697525;
assign addr[62601] = -2083416198;
assign addr[62602] = -2087969669;
assign addr[62603] = -2092357577;
assign addr[62604] = -2096579573;
assign addr[62605] = -2100635323;
assign addr[62606] = -2104524506;
assign addr[62607] = -2108246813;
assign addr[62608] = -2111801949;
assign addr[62609] = -2115189632;
assign addr[62610] = -2118409593;
assign addr[62611] = -2121461578;
assign addr[62612] = -2124345343;
assign addr[62613] = -2127060661;
assign addr[62614] = -2129607316;
assign addr[62615] = -2131985106;
assign addr[62616] = -2134193842;
assign addr[62617] = -2136233350;
assign addr[62618] = -2138103468;
assign addr[62619] = -2139804048;
assign addr[62620] = -2141334954;
assign addr[62621] = -2142696065;
assign addr[62622] = -2143887273;
assign addr[62623] = -2144908484;
assign addr[62624] = -2145759618;
assign addr[62625] = -2146440605;
assign addr[62626] = -2146951393;
assign addr[62627] = -2147291941;
assign addr[62628] = -2147462221;
assign addr[62629] = -2147462221;
assign addr[62630] = -2147291941;
assign addr[62631] = -2146951393;
assign addr[62632] = -2146440605;
assign addr[62633] = -2145759618;
assign addr[62634] = -2144908484;
assign addr[62635] = -2143887273;
assign addr[62636] = -2142696065;
assign addr[62637] = -2141334954;
assign addr[62638] = -2139804048;
assign addr[62639] = -2138103468;
assign addr[62640] = -2136233350;
assign addr[62641] = -2134193842;
assign addr[62642] = -2131985106;
assign addr[62643] = -2129607316;
assign addr[62644] = -2127060661;
assign addr[62645] = -2124345343;
assign addr[62646] = -2121461578;
assign addr[62647] = -2118409593;
assign addr[62648] = -2115189632;
assign addr[62649] = -2111801949;
assign addr[62650] = -2108246813;
assign addr[62651] = -2104524506;
assign addr[62652] = -2100635323;
assign addr[62653] = -2096579573;
assign addr[62654] = -2092357577;
assign addr[62655] = -2087969669;
assign addr[62656] = -2083416198;
assign addr[62657] = -2078697525;
assign addr[62658] = -2073814024;
assign addr[62659] = -2068766083;
assign addr[62660] = -2063554100;
assign addr[62661] = -2058178491;
assign addr[62662] = -2052639680;
assign addr[62663] = -2046938108;
assign addr[62664] = -2041074226;
assign addr[62665] = -2035048499;
assign addr[62666] = -2028861406;
assign addr[62667] = -2022513436;
assign addr[62668] = -2016005093;
assign addr[62669] = -2009336893;
assign addr[62670] = -2002509365;
assign addr[62671] = -1995523051;
assign addr[62672] = -1988378503;
assign addr[62673] = -1981076290;
assign addr[62674] = -1973616989;
assign addr[62675] = -1966001192;
assign addr[62676] = -1958229503;
assign addr[62677] = -1950302539;
assign addr[62678] = -1942220928;
assign addr[62679] = -1933985310;
assign addr[62680] = -1925596340;
assign addr[62681] = -1917054681;
assign addr[62682] = -1908361011;
assign addr[62683] = -1899516021;
assign addr[62684] = -1890520410;
assign addr[62685] = -1881374892;
assign addr[62686] = -1872080193;
assign addr[62687] = -1862637049;
assign addr[62688] = -1853046210;
assign addr[62689] = -1843308435;
assign addr[62690] = -1833424497;
assign addr[62691] = -1823395180;
assign addr[62692] = -1813221279;
assign addr[62693] = -1802903601;
assign addr[62694] = -1792442963;
assign addr[62695] = -1781840195;
assign addr[62696] = -1771096139;
assign addr[62697] = -1760211645;
assign addr[62698] = -1749187577;
assign addr[62699] = -1738024810;
assign addr[62700] = -1726724227;
assign addr[62701] = -1715286726;
assign addr[62702] = -1703713213;
assign addr[62703] = -1692004606;
assign addr[62704] = -1680161834;
assign addr[62705] = -1668185835;
assign addr[62706] = -1656077559;
assign addr[62707] = -1643837966;
assign addr[62708] = -1631468027;
assign addr[62709] = -1618968722;
assign addr[62710] = -1606341043;
assign addr[62711] = -1593585992;
assign addr[62712] = -1580704578;
assign addr[62713] = -1567697824;
assign addr[62714] = -1554566762;
assign addr[62715] = -1541312431;
assign addr[62716] = -1527935884;
assign addr[62717] = -1514438181;
assign addr[62718] = -1500820393;
assign addr[62719] = -1487083598;
assign addr[62720] = -1473228887;
assign addr[62721] = -1459257358;
assign addr[62722] = -1445170118;
assign addr[62723] = -1430968286;
assign addr[62724] = -1416652986;
assign addr[62725] = -1402225355;
assign addr[62726] = -1387686535;
assign addr[62727] = -1373037681;
assign addr[62728] = -1358279953;
assign addr[62729] = -1343414522;
assign addr[62730] = -1328442566;
assign addr[62731] = -1313365273;
assign addr[62732] = -1298183838;
assign addr[62733] = -1282899464;
assign addr[62734] = -1267513365;
assign addr[62735] = -1252026760;
assign addr[62736] = -1236440877;
assign addr[62737] = -1220756951;
assign addr[62738] = -1204976227;
assign addr[62739] = -1189099956;
assign addr[62740] = -1173129396;
assign addr[62741] = -1157065814;
assign addr[62742] = -1140910484;
assign addr[62743] = -1124664687;
assign addr[62744] = -1108329711;
assign addr[62745] = -1091906851;
assign addr[62746] = -1075397409;
assign addr[62747] = -1058802695;
assign addr[62748] = -1042124025;
assign addr[62749] = -1025362720;
assign addr[62750] = -1008520110;
assign addr[62751] = -991597531;
assign addr[62752] = -974596324;
assign addr[62753] = -957517838;
assign addr[62754] = -940363427;
assign addr[62755] = -923134450;
assign addr[62756] = -905832274;
assign addr[62757] = -888458272;
assign addr[62758] = -871013820;
assign addr[62759] = -853500302;
assign addr[62760] = -835919107;
assign addr[62761] = -818271628;
assign addr[62762] = -800559266;
assign addr[62763] = -782783424;
assign addr[62764] = -764945512;
assign addr[62765] = -747046944;
assign addr[62766] = -729089140;
assign addr[62767] = -711073525;
assign addr[62768] = -693001525;
assign addr[62769] = -674874574;
assign addr[62770] = -656694110;
assign addr[62771] = -638461574;
assign addr[62772] = -620178412;
assign addr[62773] = -601846074;
assign addr[62774] = -583466013;
assign addr[62775] = -565039687;
assign addr[62776] = -546568556;
assign addr[62777] = -528054086;
assign addr[62778] = -509497745;
assign addr[62779] = -490901003;
assign addr[62780] = -472265336;
assign addr[62781] = -453592221;
assign addr[62782] = -434883140;
assign addr[62783] = -416139574;
assign addr[62784] = -397363011;
assign addr[62785] = -378554940;
assign addr[62786] = -359716852;
assign addr[62787] = -340850240;
assign addr[62788] = -321956601;
assign addr[62789] = -303037433;
assign addr[62790] = -284094236;
assign addr[62791] = -265128512;
assign addr[62792] = -246141764;
assign addr[62793] = -227135500;
assign addr[62794] = -208111224;
assign addr[62795] = -189070447;
assign addr[62796] = -170014678;
assign addr[62797] = -150945428;
assign addr[62798] = -131864208;
assign addr[62799] = -112772533;
assign addr[62800] = -93671915;
assign addr[62801] = -74563870;
assign addr[62802] = -55449912;
assign addr[62803] = -36331557;
assign addr[62804] = -17210322;
assign addr[62805] = 1912278;
assign addr[62806] = 21034727;
assign addr[62807] = 40155507;
assign addr[62808] = 59273104;
assign addr[62809] = 78386000;
assign addr[62810] = 97492681;
assign addr[62811] = 116591632;
assign addr[62812] = 135681337;
assign addr[62813] = 154760284;
assign addr[62814] = 173826959;
assign addr[62815] = 192879850;
assign addr[62816] = 211917448;
assign addr[62817] = 230938242;
assign addr[62818] = 249940723;
assign addr[62819] = 268923386;
assign addr[62820] = 287884725;
assign addr[62821] = 306823237;
assign addr[62822] = 325737419;
assign addr[62823] = 344625773;
assign addr[62824] = 363486799;
assign addr[62825] = 382319004;
assign addr[62826] = 401120892;
assign addr[62827] = 419890975;
assign addr[62828] = 438627762;
assign addr[62829] = 457329769;
assign addr[62830] = 475995513;
assign addr[62831] = 494623513;
assign addr[62832] = 513212292;
assign addr[62833] = 531760377;
assign addr[62834] = 550266296;
assign addr[62835] = 568728583;
assign addr[62836] = 587145773;
assign addr[62837] = 605516406;
assign addr[62838] = 623839025;
assign addr[62839] = 642112178;
assign addr[62840] = 660334415;
assign addr[62841] = 678504291;
assign addr[62842] = 696620367;
assign addr[62843] = 714681204;
assign addr[62844] = 732685372;
assign addr[62845] = 750631442;
assign addr[62846] = 768517992;
assign addr[62847] = 786343603;
assign addr[62848] = 804106861;
assign addr[62849] = 821806359;
assign addr[62850] = 839440693;
assign addr[62851] = 857008464;
assign addr[62852] = 874508280;
assign addr[62853] = 891938752;
assign addr[62854] = 909298500;
assign addr[62855] = 926586145;
assign addr[62856] = 943800318;
assign addr[62857] = 960939653;
assign addr[62858] = 978002791;
assign addr[62859] = 994988380;
assign addr[62860] = 1011895073;
assign addr[62861] = 1028721528;
assign addr[62862] = 1045466412;
assign addr[62863] = 1062128397;
assign addr[62864] = 1078706161;
assign addr[62865] = 1095198391;
assign addr[62866] = 1111603778;
assign addr[62867] = 1127921022;
assign addr[62868] = 1144148829;
assign addr[62869] = 1160285911;
assign addr[62870] = 1176330990;
assign addr[62871] = 1192282793;
assign addr[62872] = 1208140056;
assign addr[62873] = 1223901520;
assign addr[62874] = 1239565936;
assign addr[62875] = 1255132063;
assign addr[62876] = 1270598665;
assign addr[62877] = 1285964516;
assign addr[62878] = 1301228398;
assign addr[62879] = 1316389101;
assign addr[62880] = 1331445422;
assign addr[62881] = 1346396168;
assign addr[62882] = 1361240152;
assign addr[62883] = 1375976199;
assign addr[62884] = 1390603139;
assign addr[62885] = 1405119813;
assign addr[62886] = 1419525069;
assign addr[62887] = 1433817766;
assign addr[62888] = 1447996770;
assign addr[62889] = 1462060956;
assign addr[62890] = 1476009210;
assign addr[62891] = 1489840425;
assign addr[62892] = 1503553506;
assign addr[62893] = 1517147363;
assign addr[62894] = 1530620920;
assign addr[62895] = 1543973108;
assign addr[62896] = 1557202869;
assign addr[62897] = 1570309153;
assign addr[62898] = 1583290921;
assign addr[62899] = 1596147143;
assign addr[62900] = 1608876801;
assign addr[62901] = 1621478885;
assign addr[62902] = 1633952396;
assign addr[62903] = 1646296344;
assign addr[62904] = 1658509750;
assign addr[62905] = 1670591647;
assign addr[62906] = 1682541077;
assign addr[62907] = 1694357091;
assign addr[62908] = 1706038753;
assign addr[62909] = 1717585136;
assign addr[62910] = 1728995326;
assign addr[62911] = 1740268417;
assign addr[62912] = 1751403515;
assign addr[62913] = 1762399737;
assign addr[62914] = 1773256212;
assign addr[62915] = 1783972079;
assign addr[62916] = 1794546487;
assign addr[62917] = 1804978599;
assign addr[62918] = 1815267588;
assign addr[62919] = 1825412636;
assign addr[62920] = 1835412941;
assign addr[62921] = 1845267708;
assign addr[62922] = 1854976157;
assign addr[62923] = 1864537518;
assign addr[62924] = 1873951032;
assign addr[62925] = 1883215953;
assign addr[62926] = 1892331547;
assign addr[62927] = 1901297091;
assign addr[62928] = 1910111873;
assign addr[62929] = 1918775195;
assign addr[62930] = 1927286370;
assign addr[62931] = 1935644723;
assign addr[62932] = 1943849591;
assign addr[62933] = 1951900324;
assign addr[62934] = 1959796283;
assign addr[62935] = 1967536842;
assign addr[62936] = 1975121388;
assign addr[62937] = 1982549318;
assign addr[62938] = 1989820044;
assign addr[62939] = 1996932990;
assign addr[62940] = 2003887591;
assign addr[62941] = 2010683297;
assign addr[62942] = 2017319567;
assign addr[62943] = 2023795876;
assign addr[62944] = 2030111710;
assign addr[62945] = 2036266570;
assign addr[62946] = 2042259965;
assign addr[62947] = 2048091422;
assign addr[62948] = 2053760478;
assign addr[62949] = 2059266683;
assign addr[62950] = 2064609600;
assign addr[62951] = 2069788807;
assign addr[62952] = 2074803892;
assign addr[62953] = 2079654458;
assign addr[62954] = 2084340120;
assign addr[62955] = 2088860507;
assign addr[62956] = 2093215260;
assign addr[62957] = 2097404033;
assign addr[62958] = 2101426496;
assign addr[62959] = 2105282327;
assign addr[62960] = 2108971223;
assign addr[62961] = 2112492891;
assign addr[62962] = 2115847050;
assign addr[62963] = 2119033436;
assign addr[62964] = 2122051796;
assign addr[62965] = 2124901890;
assign addr[62966] = 2127583492;
assign addr[62967] = 2130096389;
assign addr[62968] = 2132440383;
assign addr[62969] = 2134615288;
assign addr[62970] = 2136620930;
assign addr[62971] = 2138457152;
assign addr[62972] = 2140123807;
assign addr[62973] = 2141620763;
assign addr[62974] = 2142947902;
assign addr[62975] = 2144105118;
assign addr[62976] = 2145092320;
assign addr[62977] = 2145909429;
assign addr[62978] = 2146556380;
assign addr[62979] = 2147033123;
assign addr[62980] = 2147339619;
assign addr[62981] = 2147475844;
assign addr[62982] = 2147441787;
assign addr[62983] = 2147237452;
assign addr[62984] = 2146862854;
assign addr[62985] = 2146318022;
assign addr[62986] = 2145603001;
assign addr[62987] = 2144717846;
assign addr[62988] = 2143662628;
assign addr[62989] = 2142437431;
assign addr[62990] = 2141042352;
assign addr[62991] = 2139477502;
assign addr[62992] = 2137743003;
assign addr[62993] = 2135838995;
assign addr[62994] = 2133765628;
assign addr[62995] = 2131523066;
assign addr[62996] = 2129111488;
assign addr[62997] = 2126531084;
assign addr[62998] = 2123782059;
assign addr[62999] = 2120864631;
assign addr[63000] = 2117779031;
assign addr[63001] = 2114525505;
assign addr[63002] = 2111104309;
assign addr[63003] = 2107515716;
assign addr[63004] = 2103760010;
assign addr[63005] = 2099837489;
assign addr[63006] = 2095748463;
assign addr[63007] = 2091493257;
assign addr[63008] = 2087072209;
assign addr[63009] = 2082485668;
assign addr[63010] = 2077733999;
assign addr[63011] = 2072817579;
assign addr[63012] = 2067736796;
assign addr[63013] = 2062492055;
assign addr[63014] = 2057083771;
assign addr[63015] = 2051512372;
assign addr[63016] = 2045778302;
assign addr[63017] = 2039882013;
assign addr[63018] = 2033823974;
assign addr[63019] = 2027604666;
assign addr[63020] = 2021224581;
assign addr[63021] = 2014684225;
assign addr[63022] = 2007984117;
assign addr[63023] = 2001124788;
assign addr[63024] = 1994106782;
assign addr[63025] = 1986930656;
assign addr[63026] = 1979596978;
assign addr[63027] = 1972106330;
assign addr[63028] = 1964459306;
assign addr[63029] = 1956656513;
assign addr[63030] = 1948698568;
assign addr[63031] = 1940586104;
assign addr[63032] = 1932319763;
assign addr[63033] = 1923900201;
assign addr[63034] = 1915328086;
assign addr[63035] = 1906604097;
assign addr[63036] = 1897728925;
assign addr[63037] = 1888703276;
assign addr[63038] = 1879527863;
assign addr[63039] = 1870203416;
assign addr[63040] = 1860730673;
assign addr[63041] = 1851110385;
assign addr[63042] = 1841343316;
assign addr[63043] = 1831430239;
assign addr[63044] = 1821371941;
assign addr[63045] = 1811169220;
assign addr[63046] = 1800822883;
assign addr[63047] = 1790333753;
assign addr[63048] = 1779702660;
assign addr[63049] = 1768930447;
assign addr[63050] = 1758017969;
assign addr[63051] = 1746966091;
assign addr[63052] = 1735775690;
assign addr[63053] = 1724447652;
assign addr[63054] = 1712982875;
assign addr[63055] = 1701382270;
assign addr[63056] = 1689646755;
assign addr[63057] = 1677777262;
assign addr[63058] = 1665774731;
assign addr[63059] = 1653640115;
assign addr[63060] = 1641374375;
assign addr[63061] = 1628978484;
assign addr[63062] = 1616453425;
assign addr[63063] = 1603800191;
assign addr[63064] = 1591019785;
assign addr[63065] = 1578113222;
assign addr[63066] = 1565081523;
assign addr[63067] = 1551925723;
assign addr[63068] = 1538646865;
assign addr[63069] = 1525246002;
assign addr[63070] = 1511724196;
assign addr[63071] = 1498082520;
assign addr[63072] = 1484322054;
assign addr[63073] = 1470443891;
assign addr[63074] = 1456449131;
assign addr[63075] = 1442338884;
assign addr[63076] = 1428114267;
assign addr[63077] = 1413776410;
assign addr[63078] = 1399326449;
assign addr[63079] = 1384765530;
assign addr[63080] = 1370094808;
assign addr[63081] = 1355315445;
assign addr[63082] = 1340428615;
assign addr[63083] = 1325435496;
assign addr[63084] = 1310337279;
assign addr[63085] = 1295135159;
assign addr[63086] = 1279830344;
assign addr[63087] = 1264424045;
assign addr[63088] = 1248917486;
assign addr[63089] = 1233311895;
assign addr[63090] = 1217608510;
assign addr[63091] = 1201808576;
assign addr[63092] = 1185913346;
assign addr[63093] = 1169924081;
assign addr[63094] = 1153842047;
assign addr[63095] = 1137668521;
assign addr[63096] = 1121404785;
assign addr[63097] = 1105052128;
assign addr[63098] = 1088611847;
assign addr[63099] = 1072085246;
assign addr[63100] = 1055473635;
assign addr[63101] = 1038778332;
assign addr[63102] = 1022000660;
assign addr[63103] = 1005141949;
assign addr[63104] = 988203537;
assign addr[63105] = 971186766;
assign addr[63106] = 954092986;
assign addr[63107] = 936923553;
assign addr[63108] = 919679827;
assign addr[63109] = 902363176;
assign addr[63110] = 884974973;
assign addr[63111] = 867516597;
assign addr[63112] = 849989433;
assign addr[63113] = 832394869;
assign addr[63114] = 814734301;
assign addr[63115] = 797009130;
assign addr[63116] = 779220762;
assign addr[63117] = 761370605;
assign addr[63118] = 743460077;
assign addr[63119] = 725490597;
assign addr[63120] = 707463589;
assign addr[63121] = 689380485;
assign addr[63122] = 671242716;
assign addr[63123] = 653051723;
assign addr[63124] = 634808946;
assign addr[63125] = 616515832;
assign addr[63126] = 598173833;
assign addr[63127] = 579784402;
assign addr[63128] = 561348998;
assign addr[63129] = 542869083;
assign addr[63130] = 524346121;
assign addr[63131] = 505781581;
assign addr[63132] = 487176937;
assign addr[63133] = 468533662;
assign addr[63134] = 449853235;
assign addr[63135] = 431137138;
assign addr[63136] = 412386854;
assign addr[63137] = 393603870;
assign addr[63138] = 374789676;
assign addr[63139] = 355945764;
assign addr[63140] = 337073627;
assign addr[63141] = 318174762;
assign addr[63142] = 299250668;
assign addr[63143] = 280302845;
assign addr[63144] = 261332796;
assign addr[63145] = 242342025;
assign addr[63146] = 223332037;
assign addr[63147] = 204304341;
assign addr[63148] = 185260444;
assign addr[63149] = 166201858;
assign addr[63150] = 147130093;
assign addr[63151] = 128046661;
assign addr[63152] = 108953076;
assign addr[63153] = 89850852;
assign addr[63154] = 70741503;
assign addr[63155] = 51626544;
assign addr[63156] = 32507492;
assign addr[63157] = 13385863;
assign addr[63158] = -5736829;
assign addr[63159] = -24859065;
assign addr[63160] = -43979330;
assign addr[63161] = -63096108;
assign addr[63162] = -82207882;
assign addr[63163] = -101313138;
assign addr[63164] = -120410361;
assign addr[63165] = -139498035;
assign addr[63166] = -158574649;
assign addr[63167] = -177638688;
assign addr[63168] = -196688642;
assign addr[63169] = -215722999;
assign addr[63170] = -234740251;
assign addr[63171] = -253738890;
assign addr[63172] = -272717408;
assign addr[63173] = -291674302;
assign addr[63174] = -310608068;
assign addr[63175] = -329517204;
assign addr[63176] = -348400212;
assign addr[63177] = -367255594;
assign addr[63178] = -386081854;
assign addr[63179] = -404877501;
assign addr[63180] = -423641043;
assign addr[63181] = -442370993;
assign addr[63182] = -461065866;
assign addr[63183] = -479724180;
assign addr[63184] = -498344454;
assign addr[63185] = -516925212;
assign addr[63186] = -535464981;
assign addr[63187] = -553962291;
assign addr[63188] = -572415676;
assign addr[63189] = -590823671;
assign addr[63190] = -609184818;
assign addr[63191] = -627497660;
assign addr[63192] = -645760745;
assign addr[63193] = -663972625;
assign addr[63194] = -682131857;
assign addr[63195] = -700236999;
assign addr[63196] = -718286617;
assign addr[63197] = -736279279;
assign addr[63198] = -754213559;
assign addr[63199] = -772088034;
assign addr[63200] = -789901288;
assign addr[63201] = -807651907;
assign addr[63202] = -825338484;
assign addr[63203] = -842959617;
assign addr[63204] = -860513908;
assign addr[63205] = -877999966;
assign addr[63206] = -895416404;
assign addr[63207] = -912761841;
assign addr[63208] = -930034901;
assign addr[63209] = -947234215;
assign addr[63210] = -964358420;
assign addr[63211] = -981406156;
assign addr[63212] = -998376073;
assign addr[63213] = -1015266825;
assign addr[63214] = -1032077073;
assign addr[63215] = -1048805483;
assign addr[63216] = -1065450729;
assign addr[63217] = -1082011492;
assign addr[63218] = -1098486458;
assign addr[63219] = -1114874320;
assign addr[63220] = -1131173780;
assign addr[63221] = -1147383544;
assign addr[63222] = -1163502328;
assign addr[63223] = -1179528853;
assign addr[63224] = -1195461849;
assign addr[63225] = -1211300053;
assign addr[63226] = -1227042207;
assign addr[63227] = -1242687064;
assign addr[63228] = -1258233384;
assign addr[63229] = -1273679934;
assign addr[63230] = -1289025489;
assign addr[63231] = -1304268832;
assign addr[63232] = -1319408754;
assign addr[63233] = -1334444055;
assign addr[63234] = -1349373543;
assign addr[63235] = -1364196034;
assign addr[63236] = -1378910353;
assign addr[63237] = -1393515332;
assign addr[63238] = -1408009814;
assign addr[63239] = -1422392650;
assign addr[63240] = -1436662698;
assign addr[63241] = -1450818828;
assign addr[63242] = -1464859917;
assign addr[63243] = -1478784851;
assign addr[63244] = -1492592527;
assign addr[63245] = -1506281850;
assign addr[63246] = -1519851733;
assign addr[63247] = -1533301101;
assign addr[63248] = -1546628888;
assign addr[63249] = -1559834037;
assign addr[63250] = -1572915501;
assign addr[63251] = -1585872242;
assign addr[63252] = -1598703233;
assign addr[63253] = -1611407456;
assign addr[63254] = -1623983905;
assign addr[63255] = -1636431582;
assign addr[63256] = -1648749499;
assign addr[63257] = -1660936681;
assign addr[63258] = -1672992161;
assign addr[63259] = -1684914983;
assign addr[63260] = -1696704201;
assign addr[63261] = -1708358881;
assign addr[63262] = -1719878099;
assign addr[63263] = -1731260941;
assign addr[63264] = -1742506504;
assign addr[63265] = -1753613897;
assign addr[63266] = -1764582240;
assign addr[63267] = -1775410662;
assign addr[63268] = -1786098304;
assign addr[63269] = -1796644320;
assign addr[63270] = -1807047873;
assign addr[63271] = -1817308138;
assign addr[63272] = -1827424302;
assign addr[63273] = -1837395562;
assign addr[63274] = -1847221128;
assign addr[63275] = -1856900221;
assign addr[63276] = -1866432072;
assign addr[63277] = -1875815927;
assign addr[63278] = -1885051042;
assign addr[63279] = -1894136683;
assign addr[63280] = -1903072131;
assign addr[63281] = -1911856677;
assign addr[63282] = -1920489624;
assign addr[63283] = -1928970288;
assign addr[63284] = -1937297997;
assign addr[63285] = -1945472089;
assign addr[63286] = -1953491918;
assign addr[63287] = -1961356847;
assign addr[63288] = -1969066252;
assign addr[63289] = -1976619522;
assign addr[63290] = -1984016058;
assign addr[63291] = -1991255274;
assign addr[63292] = -1998336596;
assign addr[63293] = -2005259462;
assign addr[63294] = -2012023322;
assign addr[63295] = -2018627642;
assign addr[63296] = -2025071897;
assign addr[63297] = -2031355576;
assign addr[63298] = -2037478181;
assign addr[63299] = -2043439226;
assign addr[63300] = -2049238240;
assign addr[63301] = -2054874761;
assign addr[63302] = -2060348343;
assign addr[63303] = -2065658552;
assign addr[63304] = -2070804967;
assign addr[63305] = -2075787180;
assign addr[63306] = -2080604795;
assign addr[63307] = -2085257431;
assign addr[63308] = -2089744719;
assign addr[63309] = -2094066304;
assign addr[63310] = -2098221841;
assign addr[63311] = -2102211002;
assign addr[63312] = -2106033471;
assign addr[63313] = -2109688944;
assign addr[63314] = -2113177132;
assign addr[63315] = -2116497758;
assign addr[63316] = -2119650558;
assign addr[63317] = -2122635283;
assign addr[63318] = -2125451696;
assign addr[63319] = -2128099574;
assign addr[63320] = -2130578706;
assign addr[63321] = -2132888897;
assign addr[63322] = -2135029962;
assign addr[63323] = -2137001733;
assign addr[63324] = -2138804053;
assign addr[63325] = -2140436778;
assign addr[63326] = -2141899780;
assign addr[63327] = -2143192942;
assign addr[63328] = -2144316162;
assign addr[63329] = -2145269351;
assign addr[63330] = -2146052433;
assign addr[63331] = -2146665347;
assign addr[63332] = -2147108043;
assign addr[63333] = -2147380486;
assign addr[63334] = -2147482655;
assign addr[63335] = -2147414542;
assign addr[63336] = -2147176152;
assign addr[63337] = -2146767505;
assign addr[63338] = -2146188631;
assign addr[63339] = -2145439578;
assign addr[63340] = -2144520405;
assign addr[63341] = -2143431184;
assign addr[63342] = -2142172003;
assign addr[63343] = -2140742960;
assign addr[63344] = -2139144169;
assign addr[63345] = -2137375758;
assign addr[63346] = -2135437865;
assign addr[63347] = -2133330646;
assign addr[63348] = -2131054266;
assign addr[63349] = -2128608907;
assign addr[63350] = -2125994762;
assign addr[63351] = -2123212038;
assign addr[63352] = -2120260957;
assign addr[63353] = -2117141752;
assign addr[63354] = -2113854671;
assign addr[63355] = -2110399974;
assign addr[63356] = -2106777935;
assign addr[63357] = -2102988841;
assign addr[63358] = -2099032994;
assign addr[63359] = -2094910706;
assign addr[63360] = -2090622304;
assign addr[63361] = -2086168128;
assign addr[63362] = -2081548533;
assign addr[63363] = -2076763883;
assign addr[63364] = -2071814558;
assign addr[63365] = -2066700952;
assign addr[63366] = -2061423468;
assign addr[63367] = -2055982526;
assign addr[63368] = -2050378558;
assign addr[63369] = -2044612007;
assign addr[63370] = -2038683330;
assign addr[63371] = -2032592999;
assign addr[63372] = -2026341495;
assign addr[63373] = -2019929315;
assign addr[63374] = -2013356967;
assign addr[63375] = -2006624971;
assign addr[63376] = -1999733863;
assign addr[63377] = -1992684188;
assign addr[63378] = -1985476506;
assign addr[63379] = -1978111387;
assign addr[63380] = -1970589416;
assign addr[63381] = -1962911189;
assign addr[63382] = -1955077316;
assign addr[63383] = -1947088417;
assign addr[63384] = -1938945125;
assign addr[63385] = -1930648088;
assign addr[63386] = -1922197961;
assign addr[63387] = -1913595416;
assign addr[63388] = -1904841135;
assign addr[63389] = -1895935811;
assign addr[63390] = -1886880151;
assign addr[63391] = -1877674873;
assign addr[63392] = -1868320707;
assign addr[63393] = -1858818395;
assign addr[63394] = -1849168689;
assign addr[63395] = -1839372356;
assign addr[63396] = -1829430172;
assign addr[63397] = -1819342925;
assign addr[63398] = -1809111415;
assign addr[63399] = -1798736454;
assign addr[63400] = -1788218865;
assign addr[63401] = -1777559480;
assign addr[63402] = -1766759146;
assign addr[63403] = -1755818718;
assign addr[63404] = -1744739065;
assign addr[63405] = -1733521064;
assign addr[63406] = -1722165606;
assign addr[63407] = -1710673591;
assign addr[63408] = -1699045930;
assign addr[63409] = -1687283545;
assign addr[63410] = -1675387369;
assign addr[63411] = -1663358344;
assign addr[63412] = -1651197426;
assign addr[63413] = -1638905577;
assign addr[63414] = -1626483774;
assign addr[63415] = -1613933000;
assign addr[63416] = -1601254251;
assign addr[63417] = -1588448533;
assign addr[63418] = -1575516860;
assign addr[63419] = -1562460258;
assign addr[63420] = -1549279763;
assign addr[63421] = -1535976419;
assign addr[63422] = -1522551282;
assign addr[63423] = -1509005416;
assign addr[63424] = -1495339895;
assign addr[63425] = -1481555802;
assign addr[63426] = -1467654232;
assign addr[63427] = -1453636285;
assign addr[63428] = -1439503074;
assign addr[63429] = -1425255719;
assign addr[63430] = -1410895350;
assign addr[63431] = -1396423105;
assign addr[63432] = -1381840133;
assign addr[63433] = -1367147589;
assign addr[63434] = -1352346639;
assign addr[63435] = -1337438456;
assign addr[63436] = -1322424222;
assign addr[63437] = -1307305128;
assign addr[63438] = -1292082373;
assign addr[63439] = -1276757164;
assign addr[63440] = -1261330715;
assign addr[63441] = -1245804251;
assign addr[63442] = -1230179002;
assign addr[63443] = -1214456207;
assign addr[63444] = -1198637114;
assign addr[63445] = -1182722976;
assign addr[63446] = -1166715055;
assign addr[63447] = -1150614620;
assign addr[63448] = -1134422949;
assign addr[63449] = -1118141326;
assign addr[63450] = -1101771040;
assign addr[63451] = -1085313391;
assign addr[63452] = -1068769683;
assign addr[63453] = -1052141228;
assign addr[63454] = -1035429345;
assign addr[63455] = -1018635358;
assign addr[63456] = -1001760600;
assign addr[63457] = -984806408;
assign addr[63458] = -967774128;
assign addr[63459] = -950665109;
assign addr[63460] = -933480707;
assign addr[63461] = -916222287;
assign addr[63462] = -898891215;
assign addr[63463] = -881488868;
assign addr[63464] = -864016623;
assign addr[63465] = -846475867;
assign addr[63466] = -828867991;
assign addr[63467] = -811194391;
assign addr[63468] = -793456467;
assign addr[63469] = -775655628;
assign addr[63470] = -757793284;
assign addr[63471] = -739870851;
assign addr[63472] = -721889752;
assign addr[63473] = -703851410;
assign addr[63474] = -685757258;
assign addr[63475] = -667608730;
assign addr[63476] = -649407264;
assign addr[63477] = -631154304;
assign addr[63478] = -612851297;
assign addr[63479] = -594499695;
assign addr[63480] = -576100953;
assign addr[63481] = -557656529;
assign addr[63482] = -539167887;
assign addr[63483] = -520636492;
assign addr[63484] = -502063814;
assign addr[63485] = -483451325;
assign addr[63486] = -464800501;
assign addr[63487] = -446112822;
assign addr[63488] = -427389768;
assign addr[63489] = -408632825;
assign addr[63490] = -389843480;
assign addr[63491] = -371023223;
assign addr[63492] = -352173546;
assign addr[63493] = -333295944;
assign addr[63494] = -314391913;
assign addr[63495] = -295462954;
assign addr[63496] = -276510565;
assign addr[63497] = -257536251;
assign addr[63498] = -238541516;
assign addr[63499] = -219527866;
assign addr[63500] = -200496809;
assign addr[63501] = -181449854;
assign addr[63502] = -162388511;
assign addr[63503] = -143314291;
assign addr[63504] = -124228708;
assign addr[63505] = -105133274;
assign addr[63506] = -86029503;
assign addr[63507] = -66918911;
assign addr[63508] = -47803013;
assign addr[63509] = -28683324;
assign addr[63510] = -9561361;
assign addr[63511] = 9561361;
assign addr[63512] = 28683324;
assign addr[63513] = 47803013;
assign addr[63514] = 66918911;
assign addr[63515] = 86029503;
assign addr[63516] = 105133274;
assign addr[63517] = 124228708;
assign addr[63518] = 143314291;
assign addr[63519] = 162388511;
assign addr[63520] = 181449854;
assign addr[63521] = 200496809;
assign addr[63522] = 219527866;
assign addr[63523] = 238541516;
assign addr[63524] = 257536251;
assign addr[63525] = 276510565;
assign addr[63526] = 295462953;
assign addr[63527] = 314391913;
assign addr[63528] = 333295944;
assign addr[63529] = 352173546;
assign addr[63530] = 371023223;
assign addr[63531] = 389843480;
assign addr[63532] = 408632825;
assign addr[63533] = 427389768;
assign addr[63534] = 446112822;
assign addr[63535] = 464800501;
assign addr[63536] = 483451325;
assign addr[63537] = 502063814;
assign addr[63538] = 520636492;
assign addr[63539] = 539167887;
assign addr[63540] = 557656529;
assign addr[63541] = 576100953;
assign addr[63542] = 594499695;
assign addr[63543] = 612851297;
assign addr[63544] = 631154304;
assign addr[63545] = 649407264;
assign addr[63546] = 667608730;
assign addr[63547] = 685757258;
assign addr[63548] = 703851410;
assign addr[63549] = 721889752;
assign addr[63550] = 739870851;
assign addr[63551] = 757793284;
assign addr[63552] = 775655628;
assign addr[63553] = 793456467;
assign addr[63554] = 811194391;
assign addr[63555] = 828867991;
assign addr[63556] = 846475867;
assign addr[63557] = 864016623;
assign addr[63558] = 881488868;
assign addr[63559] = 898891215;
assign addr[63560] = 916222287;
assign addr[63561] = 933480707;
assign addr[63562] = 950665109;
assign addr[63563] = 967774128;
assign addr[63564] = 984806408;
assign addr[63565] = 1001760600;
assign addr[63566] = 1018635358;
assign addr[63567] = 1035429345;
assign addr[63568] = 1052141228;
assign addr[63569] = 1068769683;
assign addr[63570] = 1085313391;
assign addr[63571] = 1101771040;
assign addr[63572] = 1118141326;
assign addr[63573] = 1134422949;
assign addr[63574] = 1150614620;
assign addr[63575] = 1166715055;
assign addr[63576] = 1182722976;
assign addr[63577] = 1198637114;
assign addr[63578] = 1214456207;
assign addr[63579] = 1230179002;
assign addr[63580] = 1245804251;
assign addr[63581] = 1261330715;
assign addr[63582] = 1276757164;
assign addr[63583] = 1292082373;
assign addr[63584] = 1307305128;
assign addr[63585] = 1322424222;
assign addr[63586] = 1337438456;
assign addr[63587] = 1352346639;
assign addr[63588] = 1367147589;
assign addr[63589] = 1381840133;
assign addr[63590] = 1396423105;
assign addr[63591] = 1410895350;
assign addr[63592] = 1425255719;
assign addr[63593] = 1439503074;
assign addr[63594] = 1453636285;
assign addr[63595] = 1467654232;
assign addr[63596] = 1481555802;
assign addr[63597] = 1495339895;
assign addr[63598] = 1509005416;
assign addr[63599] = 1522551282;
assign addr[63600] = 1535976419;
assign addr[63601] = 1549279763;
assign addr[63602] = 1562460258;
assign addr[63603] = 1575516860;
assign addr[63604] = 1588448533;
assign addr[63605] = 1601254251;
assign addr[63606] = 1613933000;
assign addr[63607] = 1626483774;
assign addr[63608] = 1638905577;
assign addr[63609] = 1651197426;
assign addr[63610] = 1663358344;
assign addr[63611] = 1675387369;
assign addr[63612] = 1687283545;
assign addr[63613] = 1699045930;
assign addr[63614] = 1710673591;
assign addr[63615] = 1722165606;
assign addr[63616] = 1733521064;
assign addr[63617] = 1744739065;
assign addr[63618] = 1755818718;
assign addr[63619] = 1766759146;
assign addr[63620] = 1777559480;
assign addr[63621] = 1788218865;
assign addr[63622] = 1798736454;
assign addr[63623] = 1809111415;
assign addr[63624] = 1819342925;
assign addr[63625] = 1829430172;
assign addr[63626] = 1839372356;
assign addr[63627] = 1849168689;
assign addr[63628] = 1858818395;
assign addr[63629] = 1868320707;
assign addr[63630] = 1877674873;
assign addr[63631] = 1886880151;
assign addr[63632] = 1895935811;
assign addr[63633] = 1904841135;
assign addr[63634] = 1913595416;
assign addr[63635] = 1922197961;
assign addr[63636] = 1930648088;
assign addr[63637] = 1938945125;
assign addr[63638] = 1947088417;
assign addr[63639] = 1955077316;
assign addr[63640] = 1962911189;
assign addr[63641] = 1970589416;
assign addr[63642] = 1978111387;
assign addr[63643] = 1985476506;
assign addr[63644] = 1992684188;
assign addr[63645] = 1999733863;
assign addr[63646] = 2006624971;
assign addr[63647] = 2013356967;
assign addr[63648] = 2019929315;
assign addr[63649] = 2026341495;
assign addr[63650] = 2032592999;
assign addr[63651] = 2038683330;
assign addr[63652] = 2044612007;
assign addr[63653] = 2050378558;
assign addr[63654] = 2055982526;
assign addr[63655] = 2061423468;
assign addr[63656] = 2066700952;
assign addr[63657] = 2071814558;
assign addr[63658] = 2076763883;
assign addr[63659] = 2081548533;
assign addr[63660] = 2086168128;
assign addr[63661] = 2090622304;
assign addr[63662] = 2094910706;
assign addr[63663] = 2099032994;
assign addr[63664] = 2102988841;
assign addr[63665] = 2106777935;
assign addr[63666] = 2110399974;
assign addr[63667] = 2113854671;
assign addr[63668] = 2117141752;
assign addr[63669] = 2120260957;
assign addr[63670] = 2123212038;
assign addr[63671] = 2125994762;
assign addr[63672] = 2128608907;
assign addr[63673] = 2131054266;
assign addr[63674] = 2133330646;
assign addr[63675] = 2135437865;
assign addr[63676] = 2137375758;
assign addr[63677] = 2139144169;
assign addr[63678] = 2140742960;
assign addr[63679] = 2142172003;
assign addr[63680] = 2143431184;
assign addr[63681] = 2144520405;
assign addr[63682] = 2145439578;
assign addr[63683] = 2146188631;
assign addr[63684] = 2146767505;
assign addr[63685] = 2147176152;
assign addr[63686] = 2147414542;
assign addr[63687] = 2147482655;
assign addr[63688] = 2147380486;
assign addr[63689] = 2147108043;
assign addr[63690] = 2146665347;
assign addr[63691] = 2146052433;
assign addr[63692] = 2145269351;
assign addr[63693] = 2144316162;
assign addr[63694] = 2143192942;
assign addr[63695] = 2141899780;
assign addr[63696] = 2140436778;
assign addr[63697] = 2138804053;
assign addr[63698] = 2137001733;
assign addr[63699] = 2135029962;
assign addr[63700] = 2132888897;
assign addr[63701] = 2130578706;
assign addr[63702] = 2128099574;
assign addr[63703] = 2125451696;
assign addr[63704] = 2122635283;
assign addr[63705] = 2119650558;
assign addr[63706] = 2116497758;
assign addr[63707] = 2113177132;
assign addr[63708] = 2109688944;
assign addr[63709] = 2106033471;
assign addr[63710] = 2102211002;
assign addr[63711] = 2098221841;
assign addr[63712] = 2094066304;
assign addr[63713] = 2089744719;
assign addr[63714] = 2085257431;
assign addr[63715] = 2080604795;
assign addr[63716] = 2075787180;
assign addr[63717] = 2070804967;
assign addr[63718] = 2065658552;
assign addr[63719] = 2060348343;
assign addr[63720] = 2054874761;
assign addr[63721] = 2049238240;
assign addr[63722] = 2043439226;
assign addr[63723] = 2037478181;
assign addr[63724] = 2031355576;
assign addr[63725] = 2025071897;
assign addr[63726] = 2018627642;
assign addr[63727] = 2012023322;
assign addr[63728] = 2005259462;
assign addr[63729] = 1998336596;
assign addr[63730] = 1991255274;
assign addr[63731] = 1984016058;
assign addr[63732] = 1976619522;
assign addr[63733] = 1969066252;
assign addr[63734] = 1961356847;
assign addr[63735] = 1953491918;
assign addr[63736] = 1945472089;
assign addr[63737] = 1937297997;
assign addr[63738] = 1928970288;
assign addr[63739] = 1920489624;
assign addr[63740] = 1911856677;
assign addr[63741] = 1903072131;
assign addr[63742] = 1894136683;
assign addr[63743] = 1885051042;
assign addr[63744] = 1875815927;
assign addr[63745] = 1866432072;
assign addr[63746] = 1856900221;
assign addr[63747] = 1847221128;
assign addr[63748] = 1837395562;
assign addr[63749] = 1827424302;
assign addr[63750] = 1817308138;
assign addr[63751] = 1807047873;
assign addr[63752] = 1796644320;
assign addr[63753] = 1786098304;
assign addr[63754] = 1775410662;
assign addr[63755] = 1764582240;
assign addr[63756] = 1753613897;
assign addr[63757] = 1742506504;
assign addr[63758] = 1731260941;
assign addr[63759] = 1719878099;
assign addr[63760] = 1708358881;
assign addr[63761] = 1696704201;
assign addr[63762] = 1684914983;
assign addr[63763] = 1672992161;
assign addr[63764] = 1660936681;
assign addr[63765] = 1648749499;
assign addr[63766] = 1636431582;
assign addr[63767] = 1623983905;
assign addr[63768] = 1611407456;
assign addr[63769] = 1598703233;
assign addr[63770] = 1585872242;
assign addr[63771] = 1572915501;
assign addr[63772] = 1559834037;
assign addr[63773] = 1546628888;
assign addr[63774] = 1533301101;
assign addr[63775] = 1519851733;
assign addr[63776] = 1506281850;
assign addr[63777] = 1492592527;
assign addr[63778] = 1478784851;
assign addr[63779] = 1464859917;
assign addr[63780] = 1450818828;
assign addr[63781] = 1436662698;
assign addr[63782] = 1422392650;
assign addr[63783] = 1408009814;
assign addr[63784] = 1393515332;
assign addr[63785] = 1378910353;
assign addr[63786] = 1364196034;
assign addr[63787] = 1349373543;
assign addr[63788] = 1334444055;
assign addr[63789] = 1319408754;
assign addr[63790] = 1304268832;
assign addr[63791] = 1289025489;
assign addr[63792] = 1273679934;
assign addr[63793] = 1258233384;
assign addr[63794] = 1242687064;
assign addr[63795] = 1227042207;
assign addr[63796] = 1211300053;
assign addr[63797] = 1195461849;
assign addr[63798] = 1179528853;
assign addr[63799] = 1163502328;
assign addr[63800] = 1147383544;
assign addr[63801] = 1131173780;
assign addr[63802] = 1114874320;
assign addr[63803] = 1098486458;
assign addr[63804] = 1082011492;
assign addr[63805] = 1065450729;
assign addr[63806] = 1048805483;
assign addr[63807] = 1032077073;
assign addr[63808] = 1015266825;
assign addr[63809] = 998376073;
assign addr[63810] = 981406156;
assign addr[63811] = 964358420;
assign addr[63812] = 947234215;
assign addr[63813] = 930034901;
assign addr[63814] = 912761841;
assign addr[63815] = 895416404;
assign addr[63816] = 877999966;
assign addr[63817] = 860513908;
assign addr[63818] = 842959617;
assign addr[63819] = 825338484;
assign addr[63820] = 807651907;
assign addr[63821] = 789901288;
assign addr[63822] = 772088034;
assign addr[63823] = 754213559;
assign addr[63824] = 736279279;
assign addr[63825] = 718286617;
assign addr[63826] = 700236999;
assign addr[63827] = 682131857;
assign addr[63828] = 663972625;
assign addr[63829] = 645760745;
assign addr[63830] = 627497660;
assign addr[63831] = 609184818;
assign addr[63832] = 590823671;
assign addr[63833] = 572415676;
assign addr[63834] = 553962291;
assign addr[63835] = 535464981;
assign addr[63836] = 516925212;
assign addr[63837] = 498344454;
assign addr[63838] = 479724180;
assign addr[63839] = 461065866;
assign addr[63840] = 442370993;
assign addr[63841] = 423641043;
assign addr[63842] = 404877501;
assign addr[63843] = 386081854;
assign addr[63844] = 367255594;
assign addr[63845] = 348400212;
assign addr[63846] = 329517204;
assign addr[63847] = 310608068;
assign addr[63848] = 291674302;
assign addr[63849] = 272717408;
assign addr[63850] = 253738890;
assign addr[63851] = 234740251;
assign addr[63852] = 215722999;
assign addr[63853] = 196688642;
assign addr[63854] = 177638688;
assign addr[63855] = 158574649;
assign addr[63856] = 139498035;
assign addr[63857] = 120410361;
assign addr[63858] = 101313138;
assign addr[63859] = 82207882;
assign addr[63860] = 63096108;
assign addr[63861] = 43979330;
assign addr[63862] = 24859065;
assign addr[63863] = 5736829;
assign addr[63864] = -13385863;
assign addr[63865] = -32507492;
assign addr[63866] = -51626544;
assign addr[63867] = -70741503;
assign addr[63868] = -89850852;
assign addr[63869] = -108953076;
assign addr[63870] = -128046661;
assign addr[63871] = -147130093;
assign addr[63872] = -166201858;
assign addr[63873] = -185260444;
assign addr[63874] = -204304341;
assign addr[63875] = -223332037;
assign addr[63876] = -242342025;
assign addr[63877] = -261332796;
assign addr[63878] = -280302845;
assign addr[63879] = -299250668;
assign addr[63880] = -318174762;
assign addr[63881] = -337073627;
assign addr[63882] = -355945764;
assign addr[63883] = -374789676;
assign addr[63884] = -393603870;
assign addr[63885] = -412386854;
assign addr[63886] = -431137138;
assign addr[63887] = -449853235;
assign addr[63888] = -468533662;
assign addr[63889] = -487176937;
assign addr[63890] = -505781581;
assign addr[63891] = -524346121;
assign addr[63892] = -542869083;
assign addr[63893] = -561348998;
assign addr[63894] = -579784402;
assign addr[63895] = -598173833;
assign addr[63896] = -616515832;
assign addr[63897] = -634808946;
assign addr[63898] = -653051723;
assign addr[63899] = -671242716;
assign addr[63900] = -689380485;
assign addr[63901] = -707463589;
assign addr[63902] = -725490597;
assign addr[63903] = -743460077;
assign addr[63904] = -761370605;
assign addr[63905] = -779220762;
assign addr[63906] = -797009130;
assign addr[63907] = -814734301;
assign addr[63908] = -832394869;
assign addr[63909] = -849989433;
assign addr[63910] = -867516597;
assign addr[63911] = -884974973;
assign addr[63912] = -902363176;
assign addr[63913] = -919679827;
assign addr[63914] = -936923553;
assign addr[63915] = -954092986;
assign addr[63916] = -971186766;
assign addr[63917] = -988203537;
assign addr[63918] = -1005141949;
assign addr[63919] = -1022000660;
assign addr[63920] = -1038778332;
assign addr[63921] = -1055473635;
assign addr[63922] = -1072085246;
assign addr[63923] = -1088611847;
assign addr[63924] = -1105052128;
assign addr[63925] = -1121404785;
assign addr[63926] = -1137668521;
assign addr[63927] = -1153842047;
assign addr[63928] = -1169924081;
assign addr[63929] = -1185913346;
assign addr[63930] = -1201808576;
assign addr[63931] = -1217608510;
assign addr[63932] = -1233311895;
assign addr[63933] = -1248917486;
assign addr[63934] = -1264424045;
assign addr[63935] = -1279830344;
assign addr[63936] = -1295135159;
assign addr[63937] = -1310337279;
assign addr[63938] = -1325435496;
assign addr[63939] = -1340428615;
assign addr[63940] = -1355315445;
assign addr[63941] = -1370094808;
assign addr[63942] = -1384765530;
assign addr[63943] = -1399326449;
assign addr[63944] = -1413776410;
assign addr[63945] = -1428114267;
assign addr[63946] = -1442338884;
assign addr[63947] = -1456449131;
assign addr[63948] = -1470443891;
assign addr[63949] = -1484322054;
assign addr[63950] = -1498082520;
assign addr[63951] = -1511724196;
assign addr[63952] = -1525246002;
assign addr[63953] = -1538646865;
assign addr[63954] = -1551925723;
assign addr[63955] = -1565081523;
assign addr[63956] = -1578113222;
assign addr[63957] = -1591019785;
assign addr[63958] = -1603800191;
assign addr[63959] = -1616453425;
assign addr[63960] = -1628978484;
assign addr[63961] = -1641374375;
assign addr[63962] = -1653640115;
assign addr[63963] = -1665774731;
assign addr[63964] = -1677777262;
assign addr[63965] = -1689646755;
assign addr[63966] = -1701382270;
assign addr[63967] = -1712982875;
assign addr[63968] = -1724447652;
assign addr[63969] = -1735775690;
assign addr[63970] = -1746966091;
assign addr[63971] = -1758017969;
assign addr[63972] = -1768930447;
assign addr[63973] = -1779702660;
assign addr[63974] = -1790333753;
assign addr[63975] = -1800822883;
assign addr[63976] = -1811169220;
assign addr[63977] = -1821371941;
assign addr[63978] = -1831430239;
assign addr[63979] = -1841343316;
assign addr[63980] = -1851110385;
assign addr[63981] = -1860730673;
assign addr[63982] = -1870203416;
assign addr[63983] = -1879527863;
assign addr[63984] = -1888703276;
assign addr[63985] = -1897728925;
assign addr[63986] = -1906604097;
assign addr[63987] = -1915328086;
assign addr[63988] = -1923900201;
assign addr[63989] = -1932319763;
assign addr[63990] = -1940586104;
assign addr[63991] = -1948698568;
assign addr[63992] = -1956656513;
assign addr[63993] = -1964459306;
assign addr[63994] = -1972106330;
assign addr[63995] = -1979596978;
assign addr[63996] = -1986930656;
assign addr[63997] = -1994106782;
assign addr[63998] = -2001124788;
assign addr[63999] = -2007984117;
assign addr[64000] = -2014684225;
assign addr[64001] = -2021224581;
assign addr[64002] = -2027604666;
assign addr[64003] = -2033823974;
assign addr[64004] = -2039882013;
assign addr[64005] = -2045778302;
assign addr[64006] = -2051512372;
assign addr[64007] = -2057083771;
assign addr[64008] = -2062492055;
assign addr[64009] = -2067736796;
assign addr[64010] = -2072817579;
assign addr[64011] = -2077733999;
assign addr[64012] = -2082485668;
assign addr[64013] = -2087072209;
assign addr[64014] = -2091493257;
assign addr[64015] = -2095748463;
assign addr[64016] = -2099837489;
assign addr[64017] = -2103760010;
assign addr[64018] = -2107515716;
assign addr[64019] = -2111104309;
assign addr[64020] = -2114525505;
assign addr[64021] = -2117779031;
assign addr[64022] = -2120864631;
assign addr[64023] = -2123782059;
assign addr[64024] = -2126531084;
assign addr[64025] = -2129111488;
assign addr[64026] = -2131523066;
assign addr[64027] = -2133765628;
assign addr[64028] = -2135838995;
assign addr[64029] = -2137743003;
assign addr[64030] = -2139477502;
assign addr[64031] = -2141042352;
assign addr[64032] = -2142437431;
assign addr[64033] = -2143662628;
assign addr[64034] = -2144717846;
assign addr[64035] = -2145603001;
assign addr[64036] = -2146318022;
assign addr[64037] = -2146862854;
assign addr[64038] = -2147237452;
assign addr[64039] = -2147441787;
assign addr[64040] = -2147475844;
assign addr[64041] = -2147339619;
assign addr[64042] = -2147033123;
assign addr[64043] = -2146556380;
assign addr[64044] = -2145909429;
assign addr[64045] = -2145092320;
assign addr[64046] = -2144105118;
assign addr[64047] = -2142947902;
assign addr[64048] = -2141620763;
assign addr[64049] = -2140123807;
assign addr[64050] = -2138457152;
assign addr[64051] = -2136620930;
assign addr[64052] = -2134615288;
assign addr[64053] = -2132440383;
assign addr[64054] = -2130096389;
assign addr[64055] = -2127583492;
assign addr[64056] = -2124901890;
assign addr[64057] = -2122051796;
assign addr[64058] = -2119033436;
assign addr[64059] = -2115847050;
assign addr[64060] = -2112492891;
assign addr[64061] = -2108971223;
assign addr[64062] = -2105282327;
assign addr[64063] = -2101426496;
assign addr[64064] = -2097404033;
assign addr[64065] = -2093215260;
assign addr[64066] = -2088860507;
assign addr[64067] = -2084340120;
assign addr[64068] = -2079654458;
assign addr[64069] = -2074803892;
assign addr[64070] = -2069788807;
assign addr[64071] = -2064609600;
assign addr[64072] = -2059266683;
assign addr[64073] = -2053760478;
assign addr[64074] = -2048091422;
assign addr[64075] = -2042259965;
assign addr[64076] = -2036266570;
assign addr[64077] = -2030111710;
assign addr[64078] = -2023795876;
assign addr[64079] = -2017319567;
assign addr[64080] = -2010683297;
assign addr[64081] = -2003887591;
assign addr[64082] = -1996932990;
assign addr[64083] = -1989820044;
assign addr[64084] = -1982549318;
assign addr[64085] = -1975121388;
assign addr[64086] = -1967536842;
assign addr[64087] = -1959796283;
assign addr[64088] = -1951900324;
assign addr[64089] = -1943849591;
assign addr[64090] = -1935644723;
assign addr[64091] = -1927286370;
assign addr[64092] = -1918775195;
assign addr[64093] = -1910111873;
assign addr[64094] = -1901297091;
assign addr[64095] = -1892331547;
assign addr[64096] = -1883215953;
assign addr[64097] = -1873951032;
assign addr[64098] = -1864537518;
assign addr[64099] = -1854976157;
assign addr[64100] = -1845267708;
assign addr[64101] = -1835412941;
assign addr[64102] = -1825412636;
assign addr[64103] = -1815267588;
assign addr[64104] = -1804978599;
assign addr[64105] = -1794546487;
assign addr[64106] = -1783972079;
assign addr[64107] = -1773256212;
assign addr[64108] = -1762399737;
assign addr[64109] = -1751403515;
assign addr[64110] = -1740268417;
assign addr[64111] = -1728995326;
assign addr[64112] = -1717585136;
assign addr[64113] = -1706038753;
assign addr[64114] = -1694357091;
assign addr[64115] = -1682541077;
assign addr[64116] = -1670591647;
assign addr[64117] = -1658509750;
assign addr[64118] = -1646296344;
assign addr[64119] = -1633952396;
assign addr[64120] = -1621478885;
assign addr[64121] = -1608876801;
assign addr[64122] = -1596147143;
assign addr[64123] = -1583290921;
assign addr[64124] = -1570309153;
assign addr[64125] = -1557202869;
assign addr[64126] = -1543973108;
assign addr[64127] = -1530620920;
assign addr[64128] = -1517147363;
assign addr[64129] = -1503553506;
assign addr[64130] = -1489840425;
assign addr[64131] = -1476009210;
assign addr[64132] = -1462060956;
assign addr[64133] = -1447996770;
assign addr[64134] = -1433817766;
assign addr[64135] = -1419525069;
assign addr[64136] = -1405119813;
assign addr[64137] = -1390603139;
assign addr[64138] = -1375976199;
assign addr[64139] = -1361240152;
assign addr[64140] = -1346396168;
assign addr[64141] = -1331445422;
assign addr[64142] = -1316389101;
assign addr[64143] = -1301228398;
assign addr[64144] = -1285964516;
assign addr[64145] = -1270598665;
assign addr[64146] = -1255132063;
assign addr[64147] = -1239565936;
assign addr[64148] = -1223901520;
assign addr[64149] = -1208140056;
assign addr[64150] = -1192282793;
assign addr[64151] = -1176330990;
assign addr[64152] = -1160285911;
assign addr[64153] = -1144148829;
assign addr[64154] = -1127921022;
assign addr[64155] = -1111603778;
assign addr[64156] = -1095198391;
assign addr[64157] = -1078706161;
assign addr[64158] = -1062128397;
assign addr[64159] = -1045466412;
assign addr[64160] = -1028721528;
assign addr[64161] = -1011895073;
assign addr[64162] = -994988380;
assign addr[64163] = -978002791;
assign addr[64164] = -960939653;
assign addr[64165] = -943800318;
assign addr[64166] = -926586145;
assign addr[64167] = -909298500;
assign addr[64168] = -891938752;
assign addr[64169] = -874508280;
assign addr[64170] = -857008464;
assign addr[64171] = -839440693;
assign addr[64172] = -821806359;
assign addr[64173] = -804106861;
assign addr[64174] = -786343603;
assign addr[64175] = -768517992;
assign addr[64176] = -750631442;
assign addr[64177] = -732685372;
assign addr[64178] = -714681204;
assign addr[64179] = -696620367;
assign addr[64180] = -678504291;
assign addr[64181] = -660334415;
assign addr[64182] = -642112178;
assign addr[64183] = -623839025;
assign addr[64184] = -605516406;
assign addr[64185] = -587145773;
assign addr[64186] = -568728583;
assign addr[64187] = -550266296;
assign addr[64188] = -531760377;
assign addr[64189] = -513212292;
assign addr[64190] = -494623513;
assign addr[64191] = -475995513;
assign addr[64192] = -457329769;
assign addr[64193] = -438627762;
assign addr[64194] = -419890975;
assign addr[64195] = -401120892;
assign addr[64196] = -382319004;
assign addr[64197] = -363486799;
assign addr[64198] = -344625773;
assign addr[64199] = -325737419;
assign addr[64200] = -306823237;
assign addr[64201] = -287884725;
assign addr[64202] = -268923386;
assign addr[64203] = -249940723;
assign addr[64204] = -230938242;
assign addr[64205] = -211917448;
assign addr[64206] = -192879850;
assign addr[64207] = -173826959;
assign addr[64208] = -154760284;
assign addr[64209] = -135681337;
assign addr[64210] = -116591632;
assign addr[64211] = -97492681;
assign addr[64212] = -78386000;
assign addr[64213] = -59273104;
assign addr[64214] = -40155507;
assign addr[64215] = -21034727;
assign addr[64216] = -1912278;
assign addr[64217] = 17210322;
assign addr[64218] = 36331557;
assign addr[64219] = 55449912;
assign addr[64220] = 74563870;
assign addr[64221] = 93671915;
assign addr[64222] = 112772533;
assign addr[64223] = 131864208;
assign addr[64224] = 150945428;
assign addr[64225] = 170014678;
assign addr[64226] = 189070447;
assign addr[64227] = 208111224;
assign addr[64228] = 227135500;
assign addr[64229] = 246141764;
assign addr[64230] = 265128512;
assign addr[64231] = 284094236;
assign addr[64232] = 303037433;
assign addr[64233] = 321956601;
assign addr[64234] = 340850240;
assign addr[64235] = 359716852;
assign addr[64236] = 378554940;
assign addr[64237] = 397363011;
assign addr[64238] = 416139574;
assign addr[64239] = 434883140;
assign addr[64240] = 453592221;
assign addr[64241] = 472265336;
assign addr[64242] = 490901003;
assign addr[64243] = 509497745;
assign addr[64244] = 528054086;
assign addr[64245] = 546568556;
assign addr[64246] = 565039687;
assign addr[64247] = 583466013;
assign addr[64248] = 601846074;
assign addr[64249] = 620178412;
assign addr[64250] = 638461574;
assign addr[64251] = 656694110;
assign addr[64252] = 674874574;
assign addr[64253] = 693001525;
assign addr[64254] = 711073524;
assign addr[64255] = 729089140;
assign addr[64256] = 747046944;
assign addr[64257] = 764945512;
assign addr[64258] = 782783424;
assign addr[64259] = 800559266;
assign addr[64260] = 818271628;
assign addr[64261] = 835919107;
assign addr[64262] = 853500302;
assign addr[64263] = 871013820;
assign addr[64264] = 888458272;
assign addr[64265] = 905832274;
assign addr[64266] = 923134450;
assign addr[64267] = 940363427;
assign addr[64268] = 957517838;
assign addr[64269] = 974596324;
assign addr[64270] = 991597531;
assign addr[64271] = 1008520110;
assign addr[64272] = 1025362720;
assign addr[64273] = 1042124025;
assign addr[64274] = 1058802695;
assign addr[64275] = 1075397409;
assign addr[64276] = 1091906851;
assign addr[64277] = 1108329711;
assign addr[64278] = 1124664687;
assign addr[64279] = 1140910484;
assign addr[64280] = 1157065814;
assign addr[64281] = 1173129396;
assign addr[64282] = 1189099956;
assign addr[64283] = 1204976227;
assign addr[64284] = 1220756951;
assign addr[64285] = 1236440877;
assign addr[64286] = 1252026760;
assign addr[64287] = 1267513365;
assign addr[64288] = 1282899464;
assign addr[64289] = 1298183838;
assign addr[64290] = 1313365273;
assign addr[64291] = 1328442566;
assign addr[64292] = 1343414522;
assign addr[64293] = 1358279953;
assign addr[64294] = 1373037681;
assign addr[64295] = 1387686535;
assign addr[64296] = 1402225355;
assign addr[64297] = 1416652986;
assign addr[64298] = 1430968286;
assign addr[64299] = 1445170118;
assign addr[64300] = 1459257358;
assign addr[64301] = 1473228887;
assign addr[64302] = 1487083598;
assign addr[64303] = 1500820393;
assign addr[64304] = 1514438181;
assign addr[64305] = 1527935884;
assign addr[64306] = 1541312431;
assign addr[64307] = 1554566762;
assign addr[64308] = 1567697824;
assign addr[64309] = 1580704578;
assign addr[64310] = 1593585992;
assign addr[64311] = 1606341043;
assign addr[64312] = 1618968722;
assign addr[64313] = 1631468027;
assign addr[64314] = 1643837966;
assign addr[64315] = 1656077559;
assign addr[64316] = 1668185835;
assign addr[64317] = 1680161834;
assign addr[64318] = 1692004606;
assign addr[64319] = 1703713213;
assign addr[64320] = 1715286726;
assign addr[64321] = 1726724227;
assign addr[64322] = 1738024810;
assign addr[64323] = 1749187577;
assign addr[64324] = 1760211645;
assign addr[64325] = 1771096139;
assign addr[64326] = 1781840195;
assign addr[64327] = 1792442963;
assign addr[64328] = 1802903601;
assign addr[64329] = 1813221279;
assign addr[64330] = 1823395180;
assign addr[64331] = 1833424497;
assign addr[64332] = 1843308435;
assign addr[64333] = 1853046210;
assign addr[64334] = 1862637049;
assign addr[64335] = 1872080193;
assign addr[64336] = 1881374892;
assign addr[64337] = 1890520410;
assign addr[64338] = 1899516021;
assign addr[64339] = 1908361011;
assign addr[64340] = 1917054681;
assign addr[64341] = 1925596340;
assign addr[64342] = 1933985310;
assign addr[64343] = 1942220928;
assign addr[64344] = 1950302539;
assign addr[64345] = 1958229503;
assign addr[64346] = 1966001192;
assign addr[64347] = 1973616989;
assign addr[64348] = 1981076290;
assign addr[64349] = 1988378503;
assign addr[64350] = 1995523051;
assign addr[64351] = 2002509365;
assign addr[64352] = 2009336893;
assign addr[64353] = 2016005093;
assign addr[64354] = 2022513436;
assign addr[64355] = 2028861406;
assign addr[64356] = 2035048499;
assign addr[64357] = 2041074226;
assign addr[64358] = 2046938108;
assign addr[64359] = 2052639680;
assign addr[64360] = 2058178491;
assign addr[64361] = 2063554100;
assign addr[64362] = 2068766083;
assign addr[64363] = 2073814024;
assign addr[64364] = 2078697525;
assign addr[64365] = 2083416198;
assign addr[64366] = 2087969669;
assign addr[64367] = 2092357577;
assign addr[64368] = 2096579573;
assign addr[64369] = 2100635323;
assign addr[64370] = 2104524506;
assign addr[64371] = 2108246813;
assign addr[64372] = 2111801949;
assign addr[64373] = 2115189632;
assign addr[64374] = 2118409593;
assign addr[64375] = 2121461578;
assign addr[64376] = 2124345343;
assign addr[64377] = 2127060661;
assign addr[64378] = 2129607316;
assign addr[64379] = 2131985106;
assign addr[64380] = 2134193842;
assign addr[64381] = 2136233350;
assign addr[64382] = 2138103468;
assign addr[64383] = 2139804048;
assign addr[64384] = 2141334954;
assign addr[64385] = 2142696065;
assign addr[64386] = 2143887273;
assign addr[64387] = 2144908484;
assign addr[64388] = 2145759618;
assign addr[64389] = 2146440605;
assign addr[64390] = 2146951393;
assign addr[64391] = 2147291941;
assign addr[64392] = 2147462221;
assign addr[64393] = 2147462221;
assign addr[64394] = 2147291941;
assign addr[64395] = 2146951393;
assign addr[64396] = 2146440605;
assign addr[64397] = 2145759618;
assign addr[64398] = 2144908484;
assign addr[64399] = 2143887273;
assign addr[64400] = 2142696065;
assign addr[64401] = 2141334954;
assign addr[64402] = 2139804048;
assign addr[64403] = 2138103468;
assign addr[64404] = 2136233350;
assign addr[64405] = 2134193842;
assign addr[64406] = 2131985106;
assign addr[64407] = 2129607316;
assign addr[64408] = 2127060661;
assign addr[64409] = 2124345343;
assign addr[64410] = 2121461578;
assign addr[64411] = 2118409593;
assign addr[64412] = 2115189632;
assign addr[64413] = 2111801949;
assign addr[64414] = 2108246813;
assign addr[64415] = 2104524506;
assign addr[64416] = 2100635323;
assign addr[64417] = 2096579573;
assign addr[64418] = 2092357577;
assign addr[64419] = 2087969669;
assign addr[64420] = 2083416198;
assign addr[64421] = 2078697525;
assign addr[64422] = 2073814024;
assign addr[64423] = 2068766083;
assign addr[64424] = 2063554100;
assign addr[64425] = 2058178491;
assign addr[64426] = 2052639680;
assign addr[64427] = 2046938108;
assign addr[64428] = 2041074226;
assign addr[64429] = 2035048499;
assign addr[64430] = 2028861406;
assign addr[64431] = 2022513436;
assign addr[64432] = 2016005093;
assign addr[64433] = 2009336893;
assign addr[64434] = 2002509365;
assign addr[64435] = 1995523051;
assign addr[64436] = 1988378503;
assign addr[64437] = 1981076290;
assign addr[64438] = 1973616989;
assign addr[64439] = 1966001192;
assign addr[64440] = 1958229503;
assign addr[64441] = 1950302539;
assign addr[64442] = 1942220928;
assign addr[64443] = 1933985310;
assign addr[64444] = 1925596340;
assign addr[64445] = 1917054681;
assign addr[64446] = 1908361011;
assign addr[64447] = 1899516021;
assign addr[64448] = 1890520410;
assign addr[64449] = 1881374892;
assign addr[64450] = 1872080193;
assign addr[64451] = 1862637049;
assign addr[64452] = 1853046210;
assign addr[64453] = 1843308435;
assign addr[64454] = 1833424497;
assign addr[64455] = 1823395180;
assign addr[64456] = 1813221279;
assign addr[64457] = 1802903601;
assign addr[64458] = 1792442963;
assign addr[64459] = 1781840195;
assign addr[64460] = 1771096139;
assign addr[64461] = 1760211645;
assign addr[64462] = 1749187577;
assign addr[64463] = 1738024810;
assign addr[64464] = 1726724227;
assign addr[64465] = 1715286726;
assign addr[64466] = 1703713213;
assign addr[64467] = 1692004606;
assign addr[64468] = 1680161834;
assign addr[64469] = 1668185835;
assign addr[64470] = 1656077559;
assign addr[64471] = 1643837966;
assign addr[64472] = 1631468027;
assign addr[64473] = 1618968722;
assign addr[64474] = 1606341043;
assign addr[64475] = 1593585992;
assign addr[64476] = 1580704578;
assign addr[64477] = 1567697824;
assign addr[64478] = 1554566762;
assign addr[64479] = 1541312431;
assign addr[64480] = 1527935884;
assign addr[64481] = 1514438181;
assign addr[64482] = 1500820393;
assign addr[64483] = 1487083598;
assign addr[64484] = 1473228887;
assign addr[64485] = 1459257358;
assign addr[64486] = 1445170118;
assign addr[64487] = 1430968286;
assign addr[64488] = 1416652986;
assign addr[64489] = 1402225355;
assign addr[64490] = 1387686535;
assign addr[64491] = 1373037681;
assign addr[64492] = 1358279953;
assign addr[64493] = 1343414522;
assign addr[64494] = 1328442566;
assign addr[64495] = 1313365273;
assign addr[64496] = 1298183838;
assign addr[64497] = 1282899464;
assign addr[64498] = 1267513365;
assign addr[64499] = 1252026760;
assign addr[64500] = 1236440877;
assign addr[64501] = 1220756951;
assign addr[64502] = 1204976227;
assign addr[64503] = 1189099956;
assign addr[64504] = 1173129396;
assign addr[64505] = 1157065814;
assign addr[64506] = 1140910484;
assign addr[64507] = 1124664687;
assign addr[64508] = 1108329711;
assign addr[64509] = 1091906851;
assign addr[64510] = 1075397409;
assign addr[64511] = 1058802695;
assign addr[64512] = 1042124025;
assign addr[64513] = 1025362720;
assign addr[64514] = 1008520110;
assign addr[64515] = 991597531;
assign addr[64516] = 974596324;
assign addr[64517] = 957517838;
assign addr[64518] = 940363427;
assign addr[64519] = 923134450;
assign addr[64520] = 905832274;
assign addr[64521] = 888458272;
assign addr[64522] = 871013820;
assign addr[64523] = 853500302;
assign addr[64524] = 835919107;
assign addr[64525] = 818271628;
assign addr[64526] = 800559266;
assign addr[64527] = 782783424;
assign addr[64528] = 764945512;
assign addr[64529] = 747046944;
assign addr[64530] = 729089140;
assign addr[64531] = 711073525;
assign addr[64532] = 693001525;
assign addr[64533] = 674874574;
assign addr[64534] = 656694110;
assign addr[64535] = 638461574;
assign addr[64536] = 620178412;
assign addr[64537] = 601846074;
assign addr[64538] = 583466013;
assign addr[64539] = 565039687;
assign addr[64540] = 546568556;
assign addr[64541] = 528054086;
assign addr[64542] = 509497745;
assign addr[64543] = 490901003;
assign addr[64544] = 472265336;
assign addr[64545] = 453592221;
assign addr[64546] = 434883140;
assign addr[64547] = 416139574;
assign addr[64548] = 397363011;
assign addr[64549] = 378554940;
assign addr[64550] = 359716852;
assign addr[64551] = 340850240;
assign addr[64552] = 321956601;
assign addr[64553] = 303037433;
assign addr[64554] = 284094236;
assign addr[64555] = 265128512;
assign addr[64556] = 246141764;
assign addr[64557] = 227135500;
assign addr[64558] = 208111224;
assign addr[64559] = 189070447;
assign addr[64560] = 170014678;
assign addr[64561] = 150945428;
assign addr[64562] = 131864208;
assign addr[64563] = 112772533;
assign addr[64564] = 93671915;
assign addr[64565] = 74563870;
assign addr[64566] = 55449912;
assign addr[64567] = 36331557;
assign addr[64568] = 17210322;
assign addr[64569] = -1912278;
assign addr[64570] = -21034727;
assign addr[64571] = -40155507;
assign addr[64572] = -59273104;
assign addr[64573] = -78386000;
assign addr[64574] = -97492681;
assign addr[64575] = -116591632;
assign addr[64576] = -135681337;
assign addr[64577] = -154760284;
assign addr[64578] = -173826959;
assign addr[64579] = -192879850;
assign addr[64580] = -211917448;
assign addr[64581] = -230938242;
assign addr[64582] = -249940723;
assign addr[64583] = -268923386;
assign addr[64584] = -287884725;
assign addr[64585] = -306823237;
assign addr[64586] = -325737419;
assign addr[64587] = -344625773;
assign addr[64588] = -363486799;
assign addr[64589] = -382319004;
assign addr[64590] = -401120892;
assign addr[64591] = -419890975;
assign addr[64592] = -438627762;
assign addr[64593] = -457329769;
assign addr[64594] = -475995513;
assign addr[64595] = -494623513;
assign addr[64596] = -513212292;
assign addr[64597] = -531760377;
assign addr[64598] = -550266296;
assign addr[64599] = -568728583;
assign addr[64600] = -587145773;
assign addr[64601] = -605516406;
assign addr[64602] = -623839025;
assign addr[64603] = -642112178;
assign addr[64604] = -660334415;
assign addr[64605] = -678504291;
assign addr[64606] = -696620367;
assign addr[64607] = -714681204;
assign addr[64608] = -732685372;
assign addr[64609] = -750631442;
assign addr[64610] = -768517992;
assign addr[64611] = -786343603;
assign addr[64612] = -804106861;
assign addr[64613] = -821806359;
assign addr[64614] = -839440693;
assign addr[64615] = -857008464;
assign addr[64616] = -874508280;
assign addr[64617] = -891938752;
assign addr[64618] = -909298500;
assign addr[64619] = -926586145;
assign addr[64620] = -943800318;
assign addr[64621] = -960939653;
assign addr[64622] = -978002791;
assign addr[64623] = -994988380;
assign addr[64624] = -1011895073;
assign addr[64625] = -1028721528;
assign addr[64626] = -1045466412;
assign addr[64627] = -1062128397;
assign addr[64628] = -1078706161;
assign addr[64629] = -1095198391;
assign addr[64630] = -1111603778;
assign addr[64631] = -1127921022;
assign addr[64632] = -1144148829;
assign addr[64633] = -1160285911;
assign addr[64634] = -1176330990;
assign addr[64635] = -1192282793;
assign addr[64636] = -1208140056;
assign addr[64637] = -1223901520;
assign addr[64638] = -1239565936;
assign addr[64639] = -1255132063;
assign addr[64640] = -1270598665;
assign addr[64641] = -1285964516;
assign addr[64642] = -1301228398;
assign addr[64643] = -1316389101;
assign addr[64644] = -1331445422;
assign addr[64645] = -1346396168;
assign addr[64646] = -1361240152;
assign addr[64647] = -1375976199;
assign addr[64648] = -1390603139;
assign addr[64649] = -1405119813;
assign addr[64650] = -1419525069;
assign addr[64651] = -1433817766;
assign addr[64652] = -1447996770;
assign addr[64653] = -1462060956;
assign addr[64654] = -1476009210;
assign addr[64655] = -1489840425;
assign addr[64656] = -1503553506;
assign addr[64657] = -1517147363;
assign addr[64658] = -1530620920;
assign addr[64659] = -1543973108;
assign addr[64660] = -1557202869;
assign addr[64661] = -1570309153;
assign addr[64662] = -1583290921;
assign addr[64663] = -1596147143;
assign addr[64664] = -1608876801;
assign addr[64665] = -1621478885;
assign addr[64666] = -1633952396;
assign addr[64667] = -1646296344;
assign addr[64668] = -1658509750;
assign addr[64669] = -1670591647;
assign addr[64670] = -1682541077;
assign addr[64671] = -1694357091;
assign addr[64672] = -1706038753;
assign addr[64673] = -1717585136;
assign addr[64674] = -1728995326;
assign addr[64675] = -1740268417;
assign addr[64676] = -1751403515;
assign addr[64677] = -1762399737;
assign addr[64678] = -1773256212;
assign addr[64679] = -1783972079;
assign addr[64680] = -1794546487;
assign addr[64681] = -1804978599;
assign addr[64682] = -1815267588;
assign addr[64683] = -1825412636;
assign addr[64684] = -1835412941;
assign addr[64685] = -1845267708;
assign addr[64686] = -1854976157;
assign addr[64687] = -1864537518;
assign addr[64688] = -1873951032;
assign addr[64689] = -1883215953;
assign addr[64690] = -1892331547;
assign addr[64691] = -1901297091;
assign addr[64692] = -1910111873;
assign addr[64693] = -1918775195;
assign addr[64694] = -1927286370;
assign addr[64695] = -1935644723;
assign addr[64696] = -1943849591;
assign addr[64697] = -1951900324;
assign addr[64698] = -1959796283;
assign addr[64699] = -1967536842;
assign addr[64700] = -1975121388;
assign addr[64701] = -1982549318;
assign addr[64702] = -1989820044;
assign addr[64703] = -1996932990;
assign addr[64704] = -2003887591;
assign addr[64705] = -2010683297;
assign addr[64706] = -2017319567;
assign addr[64707] = -2023795876;
assign addr[64708] = -2030111710;
assign addr[64709] = -2036266570;
assign addr[64710] = -2042259965;
assign addr[64711] = -2048091422;
assign addr[64712] = -2053760478;
assign addr[64713] = -2059266683;
assign addr[64714] = -2064609600;
assign addr[64715] = -2069788807;
assign addr[64716] = -2074803892;
assign addr[64717] = -2079654458;
assign addr[64718] = -2084340120;
assign addr[64719] = -2088860507;
assign addr[64720] = -2093215260;
assign addr[64721] = -2097404033;
assign addr[64722] = -2101426496;
assign addr[64723] = -2105282327;
assign addr[64724] = -2108971223;
assign addr[64725] = -2112492891;
assign addr[64726] = -2115847050;
assign addr[64727] = -2119033436;
assign addr[64728] = -2122051796;
assign addr[64729] = -2124901890;
assign addr[64730] = -2127583492;
assign addr[64731] = -2130096389;
assign addr[64732] = -2132440383;
assign addr[64733] = -2134615288;
assign addr[64734] = -2136620930;
assign addr[64735] = -2138457152;
assign addr[64736] = -2140123807;
assign addr[64737] = -2141620763;
assign addr[64738] = -2142947902;
assign addr[64739] = -2144105118;
assign addr[64740] = -2145092320;
assign addr[64741] = -2145909429;
assign addr[64742] = -2146556380;
assign addr[64743] = -2147033123;
assign addr[64744] = -2147339619;
assign addr[64745] = -2147475844;
assign addr[64746] = -2147441787;
assign addr[64747] = -2147237452;
assign addr[64748] = -2146862854;
assign addr[64749] = -2146318022;
assign addr[64750] = -2145603001;
assign addr[64751] = -2144717846;
assign addr[64752] = -2143662628;
assign addr[64753] = -2142437431;
assign addr[64754] = -2141042352;
assign addr[64755] = -2139477502;
assign addr[64756] = -2137743003;
assign addr[64757] = -2135838995;
assign addr[64758] = -2133765628;
assign addr[64759] = -2131523066;
assign addr[64760] = -2129111488;
assign addr[64761] = -2126531084;
assign addr[64762] = -2123782059;
assign addr[64763] = -2120864631;
assign addr[64764] = -2117779031;
assign addr[64765] = -2114525505;
assign addr[64766] = -2111104309;
assign addr[64767] = -2107515716;
assign addr[64768] = -2103760010;
assign addr[64769] = -2099837489;
assign addr[64770] = -2095748463;
assign addr[64771] = -2091493257;
assign addr[64772] = -2087072209;
assign addr[64773] = -2082485668;
assign addr[64774] = -2077733999;
assign addr[64775] = -2072817579;
assign addr[64776] = -2067736796;
assign addr[64777] = -2062492055;
assign addr[64778] = -2057083771;
assign addr[64779] = -2051512372;
assign addr[64780] = -2045778302;
assign addr[64781] = -2039882013;
assign addr[64782] = -2033823974;
assign addr[64783] = -2027604666;
assign addr[64784] = -2021224581;
assign addr[64785] = -2014684225;
assign addr[64786] = -2007984117;
assign addr[64787] = -2001124788;
assign addr[64788] = -1994106782;
assign addr[64789] = -1986930656;
assign addr[64790] = -1979596978;
assign addr[64791] = -1972106330;
assign addr[64792] = -1964459306;
assign addr[64793] = -1956656513;
assign addr[64794] = -1948698568;
assign addr[64795] = -1940586104;
assign addr[64796] = -1932319763;
assign addr[64797] = -1923900201;
assign addr[64798] = -1915328086;
assign addr[64799] = -1906604097;
assign addr[64800] = -1897728925;
assign addr[64801] = -1888703276;
assign addr[64802] = -1879527863;
assign addr[64803] = -1870203416;
assign addr[64804] = -1860730673;
assign addr[64805] = -1851110385;
assign addr[64806] = -1841343316;
assign addr[64807] = -1831430239;
assign addr[64808] = -1821371941;
assign addr[64809] = -1811169220;
assign addr[64810] = -1800822883;
assign addr[64811] = -1790333753;
assign addr[64812] = -1779702660;
assign addr[64813] = -1768930447;
assign addr[64814] = -1758017969;
assign addr[64815] = -1746966091;
assign addr[64816] = -1735775690;
assign addr[64817] = -1724447652;
assign addr[64818] = -1712982875;
assign addr[64819] = -1701382270;
assign addr[64820] = -1689646755;
assign addr[64821] = -1677777262;
assign addr[64822] = -1665774731;
assign addr[64823] = -1653640115;
assign addr[64824] = -1641374375;
assign addr[64825] = -1628978484;
assign addr[64826] = -1616453425;
assign addr[64827] = -1603800191;
assign addr[64828] = -1591019785;
assign addr[64829] = -1578113222;
assign addr[64830] = -1565081523;
assign addr[64831] = -1551925723;
assign addr[64832] = -1538646865;
assign addr[64833] = -1525246002;
assign addr[64834] = -1511724196;
assign addr[64835] = -1498082520;
assign addr[64836] = -1484322054;
assign addr[64837] = -1470443891;
assign addr[64838] = -1456449131;
assign addr[64839] = -1442338884;
assign addr[64840] = -1428114267;
assign addr[64841] = -1413776410;
assign addr[64842] = -1399326449;
assign addr[64843] = -1384765530;
assign addr[64844] = -1370094808;
assign addr[64845] = -1355315445;
assign addr[64846] = -1340428615;
assign addr[64847] = -1325435496;
assign addr[64848] = -1310337279;
assign addr[64849] = -1295135159;
assign addr[64850] = -1279830344;
assign addr[64851] = -1264424045;
assign addr[64852] = -1248917486;
assign addr[64853] = -1233311895;
assign addr[64854] = -1217608510;
assign addr[64855] = -1201808576;
assign addr[64856] = -1185913346;
assign addr[64857] = -1169924081;
assign addr[64858] = -1153842047;
assign addr[64859] = -1137668521;
assign addr[64860] = -1121404785;
assign addr[64861] = -1105052128;
assign addr[64862] = -1088611847;
assign addr[64863] = -1072085246;
assign addr[64864] = -1055473635;
assign addr[64865] = -1038778332;
assign addr[64866] = -1022000660;
assign addr[64867] = -1005141949;
assign addr[64868] = -988203537;
assign addr[64869] = -971186766;
assign addr[64870] = -954092986;
assign addr[64871] = -936923553;
assign addr[64872] = -919679827;
assign addr[64873] = -902363176;
assign addr[64874] = -884974973;
assign addr[64875] = -867516597;
assign addr[64876] = -849989433;
assign addr[64877] = -832394869;
assign addr[64878] = -814734301;
assign addr[64879] = -797009130;
assign addr[64880] = -779220762;
assign addr[64881] = -761370605;
assign addr[64882] = -743460077;
assign addr[64883] = -725490597;
assign addr[64884] = -707463589;
assign addr[64885] = -689380485;
assign addr[64886] = -671242716;
assign addr[64887] = -653051723;
assign addr[64888] = -634808946;
assign addr[64889] = -616515832;
assign addr[64890] = -598173833;
assign addr[64891] = -579784402;
assign addr[64892] = -561348998;
assign addr[64893] = -542869083;
assign addr[64894] = -524346121;
assign addr[64895] = -505781581;
assign addr[64896] = -487176937;
assign addr[64897] = -468533662;
assign addr[64898] = -449853235;
assign addr[64899] = -431137138;
assign addr[64900] = -412386854;
assign addr[64901] = -393603870;
assign addr[64902] = -374789676;
assign addr[64903] = -355945764;
assign addr[64904] = -337073627;
assign addr[64905] = -318174762;
assign addr[64906] = -299250668;
assign addr[64907] = -280302845;
assign addr[64908] = -261332796;
assign addr[64909] = -242342025;
assign addr[64910] = -223332037;
assign addr[64911] = -204304341;
assign addr[64912] = -185260444;
assign addr[64913] = -166201858;
assign addr[64914] = -147130093;
assign addr[64915] = -128046661;
assign addr[64916] = -108953076;
assign addr[64917] = -89850852;
assign addr[64918] = -70741503;
assign addr[64919] = -51626544;
assign addr[64920] = -32507492;
assign addr[64921] = -13385863;
assign addr[64922] = 5736829;
assign addr[64923] = 24859065;
assign addr[64924] = 43979330;
assign addr[64925] = 63096108;
assign addr[64926] = 82207882;
assign addr[64927] = 101313138;
assign addr[64928] = 120410361;
assign addr[64929] = 139498035;
assign addr[64930] = 158574649;
assign addr[64931] = 177638688;
assign addr[64932] = 196688642;
assign addr[64933] = 215722999;
assign addr[64934] = 234740251;
assign addr[64935] = 253738890;
assign addr[64936] = 272717408;
assign addr[64937] = 291674302;
assign addr[64938] = 310608068;
assign addr[64939] = 329517204;
assign addr[64940] = 348400212;
assign addr[64941] = 367255594;
assign addr[64942] = 386081854;
assign addr[64943] = 404877501;
assign addr[64944] = 423641043;
assign addr[64945] = 442370993;
assign addr[64946] = 461065866;
assign addr[64947] = 479724180;
assign addr[64948] = 498344454;
assign addr[64949] = 516925212;
assign addr[64950] = 535464981;
assign addr[64951] = 553962291;
assign addr[64952] = 572415676;
assign addr[64953] = 590823671;
assign addr[64954] = 609184818;
assign addr[64955] = 627497660;
assign addr[64956] = 645760745;
assign addr[64957] = 663972625;
assign addr[64958] = 682131857;
assign addr[64959] = 700236999;
assign addr[64960] = 718286617;
assign addr[64961] = 736279279;
assign addr[64962] = 754213559;
assign addr[64963] = 772088034;
assign addr[64964] = 789901288;
assign addr[64965] = 807651907;
assign addr[64966] = 825338484;
assign addr[64967] = 842959617;
assign addr[64968] = 860513908;
assign addr[64969] = 877999966;
assign addr[64970] = 895416404;
assign addr[64971] = 912761841;
assign addr[64972] = 930034901;
assign addr[64973] = 947234215;
assign addr[64974] = 964358420;
assign addr[64975] = 981406156;
assign addr[64976] = 998376073;
assign addr[64977] = 1015266825;
assign addr[64978] = 1032077073;
assign addr[64979] = 1048805483;
assign addr[64980] = 1065450729;
assign addr[64981] = 1082011492;
assign addr[64982] = 1098486458;
assign addr[64983] = 1114874320;
assign addr[64984] = 1131173780;
assign addr[64985] = 1147383544;
assign addr[64986] = 1163502328;
assign addr[64987] = 1179528853;
assign addr[64988] = 1195461849;
assign addr[64989] = 1211300053;
assign addr[64990] = 1227042207;
assign addr[64991] = 1242687064;
assign addr[64992] = 1258233384;
assign addr[64993] = 1273679934;
assign addr[64994] = 1289025489;
assign addr[64995] = 1304268832;
assign addr[64996] = 1319408754;
assign addr[64997] = 1334444055;
assign addr[64998] = 1349373543;
assign addr[64999] = 1364196034;
assign addr[65000] = 1378910353;
assign addr[65001] = 1393515332;
assign addr[65002] = 1408009814;
assign addr[65003] = 1422392650;
assign addr[65004] = 1436662698;
assign addr[65005] = 1450818828;
assign addr[65006] = 1464859917;
assign addr[65007] = 1478784851;
assign addr[65008] = 1492592527;
assign addr[65009] = 1506281850;
assign addr[65010] = 1519851733;
assign addr[65011] = 1533301101;
assign addr[65012] = 1546628888;
assign addr[65013] = 1559834037;
assign addr[65014] = 1572915501;
assign addr[65015] = 1585872242;
assign addr[65016] = 1598703233;
assign addr[65017] = 1611407456;
assign addr[65018] = 1623983905;
assign addr[65019] = 1636431582;
assign addr[65020] = 1648749499;
assign addr[65021] = 1660936681;
assign addr[65022] = 1672992161;
assign addr[65023] = 1684914983;
assign addr[65024] = 1696704201;
assign addr[65025] = 1708358881;
assign addr[65026] = 1719878099;
assign addr[65027] = 1731260941;
assign addr[65028] = 1742506504;
assign addr[65029] = 1753613897;
assign addr[65030] = 1764582240;
assign addr[65031] = 1775410662;
assign addr[65032] = 1786098304;
assign addr[65033] = 1796644320;
assign addr[65034] = 1807047873;
assign addr[65035] = 1817308138;
assign addr[65036] = 1827424302;
assign addr[65037] = 1837395562;
assign addr[65038] = 1847221128;
assign addr[65039] = 1856900221;
assign addr[65040] = 1866432072;
assign addr[65041] = 1875815927;
assign addr[65042] = 1885051042;
assign addr[65043] = 1894136683;
assign addr[65044] = 1903072131;
assign addr[65045] = 1911856677;
assign addr[65046] = 1920489624;
assign addr[65047] = 1928970288;
assign addr[65048] = 1937297997;
assign addr[65049] = 1945472089;
assign addr[65050] = 1953491918;
assign addr[65051] = 1961356847;
assign addr[65052] = 1969066252;
assign addr[65053] = 1976619522;
assign addr[65054] = 1984016058;
assign addr[65055] = 1991255274;
assign addr[65056] = 1998336596;
assign addr[65057] = 2005259462;
assign addr[65058] = 2012023322;
assign addr[65059] = 2018627642;
assign addr[65060] = 2025071897;
assign addr[65061] = 2031355576;
assign addr[65062] = 2037478181;
assign addr[65063] = 2043439226;
assign addr[65064] = 2049238240;
assign addr[65065] = 2054874761;
assign addr[65066] = 2060348343;
assign addr[65067] = 2065658552;
assign addr[65068] = 2070804967;
assign addr[65069] = 2075787180;
assign addr[65070] = 2080604795;
assign addr[65071] = 2085257431;
assign addr[65072] = 2089744719;
assign addr[65073] = 2094066304;
assign addr[65074] = 2098221841;
assign addr[65075] = 2102211002;
assign addr[65076] = 2106033471;
assign addr[65077] = 2109688944;
assign addr[65078] = 2113177132;
assign addr[65079] = 2116497758;
assign addr[65080] = 2119650558;
assign addr[65081] = 2122635283;
assign addr[65082] = 2125451696;
assign addr[65083] = 2128099574;
assign addr[65084] = 2130578706;
assign addr[65085] = 2132888897;
assign addr[65086] = 2135029962;
assign addr[65087] = 2137001733;
assign addr[65088] = 2138804053;
assign addr[65089] = 2140436778;
assign addr[65090] = 2141899780;
assign addr[65091] = 2143192942;
assign addr[65092] = 2144316162;
assign addr[65093] = 2145269351;
assign addr[65094] = 2146052433;
assign addr[65095] = 2146665347;
assign addr[65096] = 2147108043;
assign addr[65097] = 2147380486;
assign addr[65098] = 2147482655;
assign addr[65099] = 2147414542;
assign addr[65100] = 2147176152;
assign addr[65101] = 2146767505;
assign addr[65102] = 2146188631;
assign addr[65103] = 2145439578;
assign addr[65104] = 2144520405;
assign addr[65105] = 2143431184;
assign addr[65106] = 2142172003;
assign addr[65107] = 2140742960;
assign addr[65108] = 2139144169;
assign addr[65109] = 2137375758;
assign addr[65110] = 2135437865;
assign addr[65111] = 2133330646;
assign addr[65112] = 2131054266;
assign addr[65113] = 2128608907;
assign addr[65114] = 2125994762;
assign addr[65115] = 2123212038;
assign addr[65116] = 2120260957;
assign addr[65117] = 2117141752;
assign addr[65118] = 2113854671;
assign addr[65119] = 2110399974;
assign addr[65120] = 2106777935;
assign addr[65121] = 2102988841;
assign addr[65122] = 2099032994;
assign addr[65123] = 2094910706;
assign addr[65124] = 2090622304;
assign addr[65125] = 2086168128;
assign addr[65126] = 2081548533;
assign addr[65127] = 2076763883;
assign addr[65128] = 2071814558;
assign addr[65129] = 2066700952;
assign addr[65130] = 2061423468;
assign addr[65131] = 2055982526;
assign addr[65132] = 2050378558;
assign addr[65133] = 2044612007;
assign addr[65134] = 2038683330;
assign addr[65135] = 2032592999;
assign addr[65136] = 2026341495;
assign addr[65137] = 2019929315;
assign addr[65138] = 2013356967;
assign addr[65139] = 2006624971;
assign addr[65140] = 1999733863;
assign addr[65141] = 1992684188;
assign addr[65142] = 1985476506;
assign addr[65143] = 1978111387;
assign addr[65144] = 1970589416;
assign addr[65145] = 1962911189;
assign addr[65146] = 1955077316;
assign addr[65147] = 1947088417;
assign addr[65148] = 1938945125;
assign addr[65149] = 1930648088;
assign addr[65150] = 1922197961;
assign addr[65151] = 1913595416;
assign addr[65152] = 1904841135;
assign addr[65153] = 1895935811;
assign addr[65154] = 1886880151;
assign addr[65155] = 1877674873;
assign addr[65156] = 1868320707;
assign addr[65157] = 1858818395;
assign addr[65158] = 1849168689;
assign addr[65159] = 1839372356;
assign addr[65160] = 1829430172;
assign addr[65161] = 1819342925;
assign addr[65162] = 1809111415;
assign addr[65163] = 1798736454;
assign addr[65164] = 1788218865;
assign addr[65165] = 1777559480;
assign addr[65166] = 1766759146;
assign addr[65167] = 1755818718;
assign addr[65168] = 1744739065;
assign addr[65169] = 1733521064;
assign addr[65170] = 1722165606;
assign addr[65171] = 1710673591;
assign addr[65172] = 1699045930;
assign addr[65173] = 1687283545;
assign addr[65174] = 1675387369;
assign addr[65175] = 1663358344;
assign addr[65176] = 1651197426;
assign addr[65177] = 1638905577;
assign addr[65178] = 1626483774;
assign addr[65179] = 1613933000;
assign addr[65180] = 1601254251;
assign addr[65181] = 1588448533;
assign addr[65182] = 1575516860;
assign addr[65183] = 1562460258;
assign addr[65184] = 1549279763;
assign addr[65185] = 1535976419;
assign addr[65186] = 1522551282;
assign addr[65187] = 1509005416;
assign addr[65188] = 1495339895;
assign addr[65189] = 1481555802;
assign addr[65190] = 1467654232;
assign addr[65191] = 1453636285;
assign addr[65192] = 1439503074;
assign addr[65193] = 1425255719;
assign addr[65194] = 1410895350;
assign addr[65195] = 1396423105;
assign addr[65196] = 1381840133;
assign addr[65197] = 1367147589;
assign addr[65198] = 1352346639;
assign addr[65199] = 1337438456;
assign addr[65200] = 1322424222;
assign addr[65201] = 1307305128;
assign addr[65202] = 1292082373;
assign addr[65203] = 1276757164;
assign addr[65204] = 1261330715;
assign addr[65205] = 1245804251;
assign addr[65206] = 1230179002;
assign addr[65207] = 1214456207;
assign addr[65208] = 1198637114;
assign addr[65209] = 1182722976;
assign addr[65210] = 1166715055;
assign addr[65211] = 1150614620;
assign addr[65212] = 1134422949;
assign addr[65213] = 1118141326;
assign addr[65214] = 1101771040;
assign addr[65215] = 1085313391;
assign addr[65216] = 1068769683;
assign addr[65217] = 1052141228;
assign addr[65218] = 1035429345;
assign addr[65219] = 1018635358;
assign addr[65220] = 1001760600;
assign addr[65221] = 984806408;
assign addr[65222] = 967774128;
assign addr[65223] = 950665109;
assign addr[65224] = 933480707;
assign addr[65225] = 916222287;
assign addr[65226] = 898891215;
assign addr[65227] = 881488868;
assign addr[65228] = 864016623;
assign addr[65229] = 846475867;
assign addr[65230] = 828867991;
assign addr[65231] = 811194391;
assign addr[65232] = 793456467;
assign addr[65233] = 775655628;
assign addr[65234] = 757793284;
assign addr[65235] = 739870851;
assign addr[65236] = 721889752;
assign addr[65237] = 703851410;
assign addr[65238] = 685757258;
assign addr[65239] = 667608730;
assign addr[65240] = 649407264;
assign addr[65241] = 631154304;
assign addr[65242] = 612851297;
assign addr[65243] = 594499695;
assign addr[65244] = 576100953;
assign addr[65245] = 557656529;
assign addr[65246] = 539167887;
assign addr[65247] = 520636492;
assign addr[65248] = 502063814;
assign addr[65249] = 483451325;
assign addr[65250] = 464800501;
assign addr[65251] = 446112822;
assign addr[65252] = 427389768;
assign addr[65253] = 408632825;
assign addr[65254] = 389843480;
assign addr[65255] = 371023223;
assign addr[65256] = 352173546;
assign addr[65257] = 333295944;
assign addr[65258] = 314391913;
assign addr[65259] = 295462954;
assign addr[65260] = 276510565;
assign addr[65261] = 257536251;
assign addr[65262] = 238541516;
assign addr[65263] = 219527866;
assign addr[65264] = 200496809;
assign addr[65265] = 181449854;
assign addr[65266] = 162388511;
assign addr[65267] = 143314291;
assign addr[65268] = 124228708;
assign addr[65269] = 105133274;
assign addr[65270] = 86029503;
assign addr[65271] = 66918911;
assign addr[65272] = 47803013;
assign addr[65273] = 28683324;
assign addr[65274] = 9561361;
assign addr[65275] = -9561361;
assign addr[65276] = -28683324;
assign addr[65277] = -47803013;
assign addr[65278] = -66918911;
assign addr[65279] = -86029503;
assign addr[65280] = -105133274;
assign addr[65281] = -124228708;
assign addr[65282] = -143314291;
assign addr[65283] = -162388511;
assign addr[65284] = -181449854;
assign addr[65285] = -200496809;
assign addr[65286] = -219527866;
assign addr[65287] = -238541516;
assign addr[65288] = -257536251;
assign addr[65289] = -276510565;
assign addr[65290] = -295462953;
assign addr[65291] = -314391913;
assign addr[65292] = -333295944;
assign addr[65293] = -352173546;
assign addr[65294] = -371023223;
assign addr[65295] = -389843480;
assign addr[65296] = -408632825;
assign addr[65297] = -427389768;
assign addr[65298] = -446112822;
assign addr[65299] = -464800501;
assign addr[65300] = -483451325;
assign addr[65301] = -502063814;
assign addr[65302] = -520636492;
assign addr[65303] = -539167887;
assign addr[65304] = -557656529;
assign addr[65305] = -576100953;
assign addr[65306] = -594499695;
assign addr[65307] = -612851297;
assign addr[65308] = -631154304;
assign addr[65309] = -649407264;
assign addr[65310] = -667608730;
assign addr[65311] = -685757258;
assign addr[65312] = -703851410;
assign addr[65313] = -721889752;
assign addr[65314] = -739870851;
assign addr[65315] = -757793284;
assign addr[65316] = -775655628;
assign addr[65317] = -793456467;
assign addr[65318] = -811194391;
assign addr[65319] = -828867991;
assign addr[65320] = -846475867;
assign addr[65321] = -864016623;
assign addr[65322] = -881488868;
assign addr[65323] = -898891215;
assign addr[65324] = -916222287;
assign addr[65325] = -933480707;
assign addr[65326] = -950665109;
assign addr[65327] = -967774128;
assign addr[65328] = -984806408;
assign addr[65329] = -1001760600;
assign addr[65330] = -1018635358;
assign addr[65331] = -1035429345;
assign addr[65332] = -1052141228;
assign addr[65333] = -1068769683;
assign addr[65334] = -1085313391;
assign addr[65335] = -1101771040;
assign addr[65336] = -1118141326;
assign addr[65337] = -1134422949;
assign addr[65338] = -1150614620;
assign addr[65339] = -1166715055;
assign addr[65340] = -1182722976;
assign addr[65341] = -1198637114;
assign addr[65342] = -1214456207;
assign addr[65343] = -1230179002;
assign addr[65344] = -1245804251;
assign addr[65345] = -1261330715;
assign addr[65346] = -1276757164;
assign addr[65347] = -1292082373;
assign addr[65348] = -1307305128;
assign addr[65349] = -1322424222;
assign addr[65350] = -1337438456;
assign addr[65351] = -1352346639;
assign addr[65352] = -1367147589;
assign addr[65353] = -1381840133;
assign addr[65354] = -1396423105;
assign addr[65355] = -1410895350;
assign addr[65356] = -1425255719;
assign addr[65357] = -1439503074;
assign addr[65358] = -1453636285;
assign addr[65359] = -1467654232;
assign addr[65360] = -1481555802;
assign addr[65361] = -1495339895;
assign addr[65362] = -1509005416;
assign addr[65363] = -1522551282;
assign addr[65364] = -1535976419;
assign addr[65365] = -1549279763;
assign addr[65366] = -1562460258;
assign addr[65367] = -1575516860;
assign addr[65368] = -1588448533;
assign addr[65369] = -1601254251;
assign addr[65370] = -1613933000;
assign addr[65371] = -1626483774;
assign addr[65372] = -1638905577;
assign addr[65373] = -1651197426;
assign addr[65374] = -1663358344;
assign addr[65375] = -1675387369;
assign addr[65376] = -1687283545;
assign addr[65377] = -1699045930;
assign addr[65378] = -1710673591;
assign addr[65379] = -1722165606;
assign addr[65380] = -1733521064;
assign addr[65381] = -1744739065;
assign addr[65382] = -1755818718;
assign addr[65383] = -1766759146;
assign addr[65384] = -1777559480;
assign addr[65385] = -1788218865;
assign addr[65386] = -1798736454;
assign addr[65387] = -1809111415;
assign addr[65388] = -1819342925;
assign addr[65389] = -1829430172;
assign addr[65390] = -1839372356;
assign addr[65391] = -1849168689;
assign addr[65392] = -1858818395;
assign addr[65393] = -1868320707;
assign addr[65394] = -1877674873;
assign addr[65395] = -1886880151;
assign addr[65396] = -1895935811;
assign addr[65397] = -1904841135;
assign addr[65398] = -1913595416;
assign addr[65399] = -1922197961;
assign addr[65400] = -1930648088;
assign addr[65401] = -1938945125;
assign addr[65402] = -1947088417;
assign addr[65403] = -1955077316;
assign addr[65404] = -1962911189;
assign addr[65405] = -1970589416;
assign addr[65406] = -1978111387;
assign addr[65407] = -1985476506;
assign addr[65408] = -1992684188;
assign addr[65409] = -1999733863;
assign addr[65410] = -2006624971;
assign addr[65411] = -2013356967;
assign addr[65412] = -2019929315;
assign addr[65413] = -2026341495;
assign addr[65414] = -2032592999;
assign addr[65415] = -2038683330;
assign addr[65416] = -2044612007;
assign addr[65417] = -2050378558;
assign addr[65418] = -2055982526;
assign addr[65419] = -2061423468;
assign addr[65420] = -2066700952;
assign addr[65421] = -2071814558;
assign addr[65422] = -2076763883;
assign addr[65423] = -2081548533;
assign addr[65424] = -2086168128;
assign addr[65425] = -2090622304;
assign addr[65426] = -2094910706;
assign addr[65427] = -2099032994;
assign addr[65428] = -2102988841;
assign addr[65429] = -2106777935;
assign addr[65430] = -2110399974;
assign addr[65431] = -2113854671;
assign addr[65432] = -2117141752;
assign addr[65433] = -2120260957;
assign addr[65434] = -2123212038;
assign addr[65435] = -2125994762;
assign addr[65436] = -2128608907;
assign addr[65437] = -2131054266;
assign addr[65438] = -2133330646;
assign addr[65439] = -2135437865;
assign addr[65440] = -2137375758;
assign addr[65441] = -2139144169;
assign addr[65442] = -2140742960;
assign addr[65443] = -2142172003;
assign addr[65444] = -2143431184;
assign addr[65445] = -2144520405;
assign addr[65446] = -2145439578;
assign addr[65447] = -2146188631;
assign addr[65448] = -2146767505;
assign addr[65449] = -2147176152;
assign addr[65450] = -2147414542;
assign addr[65451] = -2147482655;
assign addr[65452] = -2147380486;
assign addr[65453] = -2147108043;
assign addr[65454] = -2146665347;
assign addr[65455] = -2146052433;
assign addr[65456] = -2145269351;
assign addr[65457] = -2144316162;
assign addr[65458] = -2143192942;
assign addr[65459] = -2141899780;
assign addr[65460] = -2140436778;
assign addr[65461] = -2138804053;
assign addr[65462] = -2137001733;
assign addr[65463] = -2135029962;
assign addr[65464] = -2132888897;
assign addr[65465] = -2130578706;
assign addr[65466] = -2128099574;
assign addr[65467] = -2125451696;
assign addr[65468] = -2122635283;
assign addr[65469] = -2119650558;
assign addr[65470] = -2116497758;
assign addr[65471] = -2113177132;
assign addr[65472] = -2109688944;
assign addr[65473] = -2106033471;
assign addr[65474] = -2102211002;
assign addr[65475] = -2098221841;
assign addr[65476] = -2094066304;
assign addr[65477] = -2089744719;
assign addr[65478] = -2085257431;
assign addr[65479] = -2080604795;
assign addr[65480] = -2075787180;
assign addr[65481] = -2070804967;
assign addr[65482] = -2065658552;
assign addr[65483] = -2060348343;
assign addr[65484] = -2054874761;
assign addr[65485] = -2049238240;
assign addr[65486] = -2043439226;
assign addr[65487] = -2037478181;
assign addr[65488] = -2031355576;
assign addr[65489] = -2025071897;
assign addr[65490] = -2018627642;
assign addr[65491] = -2012023322;
assign addr[65492] = -2005259462;
assign addr[65493] = -1998336596;
assign addr[65494] = -1991255274;
assign addr[65495] = -1984016058;
assign addr[65496] = -1976619522;
assign addr[65497] = -1969066252;
assign addr[65498] = -1961356847;
assign addr[65499] = -1953491918;
assign addr[65500] = -1945472089;
assign addr[65501] = -1937297997;
assign addr[65502] = -1928970288;
assign addr[65503] = -1920489624;
assign addr[65504] = -1911856677;
assign addr[65505] = -1903072131;
assign addr[65506] = -1894136683;
assign addr[65507] = -1885051042;
assign addr[65508] = -1875815927;
assign addr[65509] = -1866432072;
assign addr[65510] = -1856900221;
assign addr[65511] = -1847221128;
assign addr[65512] = -1837395562;
assign addr[65513] = -1827424302;
assign addr[65514] = -1817308138;
assign addr[65515] = -1807047873;
assign addr[65516] = -1796644320;
assign addr[65517] = -1786098304;
assign addr[65518] = -1775410662;
assign addr[65519] = -1764582240;
assign addr[65520] = -1753613897;
assign addr[65521] = -1742506504;
assign addr[65522] = -1731260941;
assign addr[65523] = -1719878099;
assign addr[65524] = -1708358881;
assign addr[65525] = -1696704201;
assign addr[65526] = -1684914983;
assign addr[65527] = -1672992161;
assign addr[65528] = -1660936681;
assign addr[65529] = -1648749499;
assign addr[65530] = -1636431582;
assign addr[65531] = -1623983905;
assign addr[65532] = -1611407456;
assign addr[65533] = -1598703233;
assign addr[65534] = -1585872242;
assign addr[65535] = -1572915501;
endmodule