module rompcm44(
	input clk,//45m
	input reset_n,
	output signed [31:0]addrout
);

wire signed [31:0]addr[0:65535];
reg [9:0]k;
wire lrck;
always @(posedge clk or negedge reset_n)begin
	if(reset_n ==0) 
	k = 0;
	
	else
	k <= k+1;

end
assign lrck = k[9];
reg [15:0]i;
always @(posedge lrck or negedge reset_n)begin
	if(reset_n ==0)begin
		i <= 0;
	//	addrout <= 32'd0;
		end
	
	else begin
		i <= i+1;
	//	addrout <= addr[i];
		end
end

assign addrout = addr[i];

assign addr[0]= 0;
assign addr[1]= 304930476;
assign addr[2]= 603681519;
assign addr[3]= 890198924;
assign addr[4]= 1158676398;
assign addr[5]= 1403673233;
assign addr[6]= 1620224553;
assign addr[7]= 1803941934;
assign addr[8]= 1951102334;
assign addr[9]= 2058723538;
assign addr[10]= 2124624598;
assign addr[11]= 2147470025;
assign addr[12]= 2126796855;
assign addr[13]= 2063024031;
assign addr[14]= 1957443913;
assign addr[15]= 1812196087;
assign addr[16]= 1630224009;
assign addr[17]= 1415215352;
assign addr[18]= 1171527280;
assign addr[19]= 904098143;
assign addr[20]= 618347408;
assign addr[21]= 320065829;
assign addr[22]= 15298099;
assign addr[23]= -289779648;
assign addr[24]= -588984994;
assign addr[25]= -876254528;
assign addr[26]= -1145766716;
assign addr[27]= -1392059879;
assign addr[28]= -1610142873;
assign addr[29]= -1795596234;
assign addr[30]= -1944661739;
assign addr[31]= -2054318569;
assign addr[32]= -2122344521;
assign addr[33]= -2147361045;
assign addr[34]= -2128861181;
assign addr[35]= -2067219829;
assign addr[36]= -1963686155;
assign addr[37]= -1820358275;
assign addr[38]= -1640140734;
assign addr[39]= -1426685652;
assign addr[40]= -1184318708;
assign addr[41]= -917951481;
assign addr[42]= -632981917;
assign addr[43]= -335184940;
assign addr[44]= -30595422;
assign addr[45]= 274614114;
assign addr[46]= 574258580;
assign addr[47]= 862265664;
assign addr[48]= 1132798888;
assign addr[49]= 1380375881;
assign addr[50]= 1599979481;
assign addr[51]= 1787159411;
assign addr[52]= 1938122457;
assign addr[53]= 2049809346;
assign addr[54]= 2119956737;
assign addr[55]= 2147143090;
assign addr[56]= 2130817471;
assign addr[57]= 2071310720;
assign addr[58]= 1969828744;
assign addr[59]= 1828428082;
assign addr[60]= 1649974225;
assign addr[61]= 1438083551;
assign addr[62]= 1197050035;
assign addr[63]= 931758235;
assign addr[64]= 647584304;
assign addr[65]= 350287041;
assign addr[66]= 45891193;
assign addr[67]= -259434643;
assign addr[68]= -559503022;
assign addr[69]= -848233042;
assign addr[70]= -1119773573;
assign addr[71]= -1368621831;
assign addr[72]= -1589734894;
assign addr[73]= -1778631892;
assign addr[74]= -1931484818;
assign addr[75]= -2045196100;
assign addr[76]= -2117461370;
assign addr[77]= -2146816171;
assign addr[78]= -2132665626;
assign addr[79]= -2075296495;
assign addr[80]= -1975871368;
assign addr[81]= -1836405100;
assign addr[82]= -1659723983;
assign addr[83]= -1449408469;
assign addr[84]= -1209720613;
assign addr[85]= -945517704;
assign addr[86]= -662153826;
assign addr[87]= -365371365;
assign addr[88]= -61184634;
assign addr[89]= 244242007;
assign addr[90]= 544719071;
assign addr[91]= 834157373;
assign addr[92]= 1106691431;
assign addr[93]= 1356798326;
assign addr[94]= 1579409630;
assign addr[95]= 1770014111;
assign addr[96]= 1924749160;
assign addr[97]= 2040479063;
assign addr[98]= 2114858546;
assign addr[99]= 2146380306;
assign addr[100]= 2134405552;
assign addr[101]= 2079176953;
assign addr[102]= 1981813720;
assign addr[103]= 1844288924;
assign addr[104]= 1669389513;
assign addr[105]= 1460659832;
assign addr[106]= 1222329801;
assign addr[107]= 959229189;
assign addr[108]= 676689746;
assign addr[109]= 380437148;
assign addr[110]= 76474970;
assign addr[111]= -229036977;
assign addr[112]= -529907477;
assign addr[113]= -820039373;
assign addr[114]= -1093553126;
assign addr[115]= -1344905966;
assign addr[116]= -1569004214;
assign addr[117]= -1761306505;
assign addr[118]= -1917915825;
assign addr[119]= -2035658475;
assign addr[120]= -2112148396;
assign addr[121]= -2145835515;
assign addr[122]= -2136037160;
assign addr[123]= -2082951896;
assign addr[124]= -1987655498;
assign addr[125]= -1852079154;
assign addr[126]= -1678970324;
assign addr[127]= -1471837070;
assign addr[128]= -1234876957;
assign addr[129]= -972891995;
assign addr[130]= -691191324;
assign addr[131]= -395483624;
assign addr[132]= -91761426;
assign addr[133]= 213820322;
assign addr[134]= 515068990;
assign addr[135]= 805879757;
assign addr[136]= 1080359326;
assign addr[137]= 1332945355;
assign addr[138]= 1558519173;
assign addr[139]= 1752509516;
assign addr[140]= 1910985158;
assign addr[141]= 2030734582;
assign addr[142]= 2109331059;
assign addr[143]= 2145181827;
assign addr[144]= 2137560369;
assign addr[145]= 2086621133;
assign addr[146]= 1993396407;
assign addr[147]= 1859775393;
assign addr[148]= 1688465931;
assign addr[149]= 1482939614;
assign addr[150]= 1247361445;
assign addr[151]= 986505429;
assign addr[152]= 705657826;
assign addr[153]= 410510029;
assign addr[154]= 107043224;
assign addr[155]= -198592817;
assign addr[156]= -500204365;
assign addr[157]= -791679244;
assign addr[158]= -1067110699;
assign addr[159]= -1320917099;
assign addr[160]= -1547955041;
assign addr[161]= -1743623590;
assign addr[162]= -1903957513;
assign addr[163]= -2025707632;
assign addr[164]= -2106406677;
assign addr[165]= -2144419275;
assign addr[166]= -2138975100;
assign addr[167]= -2090184478;
assign addr[168]= -1999036154;
assign addr[169]= -1867377253;
assign addr[170]= -1697875851;
assign addr[171]= -1493966902;
assign addr[172]= -1259782632;
assign addr[173]= -1000068799;
assign addr[174]= -720088517;
assign addr[175]= -425515602;
assign addr[176]= -122319591;
assign addr[177]= 183355234;
assign addr[178]= 485314355;
assign addr[179]= 777438554;
assign addr[180]= 1053807919;
assign addr[181]= 1308821808;
assign addr[182]= 1537312353;
assign addr[183]= 1734649179;
assign addr[184]= 1896833245;
assign addr[185]= 2020577882;
assign addr[186]= 2103375398;
assign addr[187]= 2143547897;
assign addr[188]= 2140281282;
assign addr[189]= 2093641749;
assign addr[190]= 2004574453;
assign addr[191]= 1874884346;
assign addr[192]= 1707199606;
assign addr[193]= 1504918373;
assign addr[194]= 1272139887;
assign addr[195]= 1013581418;
assign addr[196]= 734482665;
assign addr[197]= 440499581;
assign addr[198]= 137589750;
assign addr[199]= -168108346;
assign addr[200]= -470399716;
assign addr[201]= -763158411;
assign addr[202]= -1040451659;
assign addr[203]= -1296660098;
assign addr[204]= -1526591649;
assign addr[205]= -1725586737;
assign addr[206]= -1889612716;
assign addr[207]= -2015345591;
assign addr[208]= -2100237377;
assign addr[209]= -2142567738;
assign addr[210]= -2141478848;
assign addr[211]= -2096992772;
assign addr[212]= -2010011024;
assign addr[213]= -1882296293;
assign addr[214]= -1716436725;
assign addr[215]= -1515793473;
assign addr[216]= -1284432584;
assign addr[217]= -1027042599;
assign addr[218]= -748839539;
assign addr[219]= -455461206;
assign addr[220]= -152852926;
assign addr[221]= 152852926;
assign addr[222]= 455461206;
assign addr[223]= 748839539;
assign addr[224]= 1027042599;
assign addr[225]= 1284432584;
assign addr[226]= 1515793473;
assign addr[227]= 1716436725;
assign addr[228]= 1882296293;
assign addr[229]= 2010011024;
assign addr[230]= 2096992772;
assign addr[231]= 2141478848;
assign addr[232]= 2142567738;
assign addr[233]= 2100237377;
assign addr[234]= 2015345591;
assign addr[235]= 1889612716;
assign addr[236]= 1725586737;
assign addr[237]= 1526591649;
assign addr[238]= 1296660098;
assign addr[239]= 1040451659;
assign addr[240]= 763158411;
assign addr[241]= 470399716;
assign addr[242]= 168108346;
assign addr[243]= -137589750;
assign addr[244]= -440499581;
assign addr[245]= -734482665;
assign addr[246]= -1013581418;
assign addr[247]= -1272139887;
assign addr[248]= -1504918373;
assign addr[249]= -1707199606;
assign addr[250]= -1874884346;
assign addr[251]= -2004574453;
assign addr[252]= -2093641749;
assign addr[253]= -2140281282;
assign addr[254]= -2143547897;
assign addr[255]= -2103375398;
assign addr[256]= -2020577882;
assign addr[257]= -1896833245;
assign addr[258]= -1734649179;
assign addr[259]= -1537312353;
assign addr[260]= -1308821808;
assign addr[261]= -1053807919;
assign addr[262]= -777438554;
assign addr[263]= -485314355;
assign addr[264]= -183355234;
assign addr[265]= 122319591;
assign addr[266]= 425515602;
assign addr[267]= 720088517;
assign addr[268]= 1000068799;
assign addr[269]= 1259782632;
assign addr[270]= 1493966902;
assign addr[271]= 1697875851;
assign addr[272]= 1867377253;
assign addr[273]= 1999036154;
assign addr[274]= 2090184478;
assign addr[275]= 2138975100;
assign addr[276]= 2144419275;
assign addr[277]= 2106406677;
assign addr[278]= 2025707632;
assign addr[279]= 1903957513;
assign addr[280]= 1743623590;
assign addr[281]= 1547955041;
assign addr[282]= 1320917099;
assign addr[283]= 1067110699;
assign addr[284]= 791679244;
assign addr[285]= 500204365;
assign addr[286]= 198592817;
assign addr[287]= -107043224;
assign addr[288]= -410510029;
assign addr[289]= -705657826;
assign addr[290]= -986505429;
assign addr[291]= -1247361445;
assign addr[292]= -1482939614;
assign addr[293]= -1688465931;
assign addr[294]= -1859775393;
assign addr[295]= -1993396407;
assign addr[296]= -2086621133;
assign addr[297]= -2137560369;
assign addr[298]= -2145181827;
assign addr[299]= -2109331059;
assign addr[300]= -2030734582;
assign addr[301]= -1910985158;
assign addr[302]= -1752509516;
assign addr[303]= -1558519173;
assign addr[304]= -1332945355;
assign addr[305]= -1080359326;
assign addr[306]= -805879757;
assign addr[307]= -515068990;
assign addr[308]= -213820322;
assign addr[309]= 91761426;
assign addr[310]= 395483624;
assign addr[311]= 691191324;
assign addr[312]= 972891995;
assign addr[313]= 1234876957;
assign addr[314]= 1471837070;
assign addr[315]= 1678970324;
assign addr[316]= 1852079154;
assign addr[317]= 1987655498;
assign addr[318]= 2082951896;
assign addr[319]= 2136037160;
assign addr[320]= 2145835515;
assign addr[321]= 2112148396;
assign addr[322]= 2035658475;
assign addr[323]= 1917915825;
assign addr[324]= 1761306505;
assign addr[325]= 1569004214;
assign addr[326]= 1344905966;
assign addr[327]= 1093553126;
assign addr[328]= 820039373;
assign addr[329]= 529907477;
assign addr[330]= 229036977;
assign addr[331]= -76474970;
assign addr[332]= -380437148;
assign addr[333]= -676689746;
assign addr[334]= -959229189;
assign addr[335]= -1222329801;
assign addr[336]= -1460659832;
assign addr[337]= -1669389513;
assign addr[338]= -1844288924;
assign addr[339]= -1981813720;
assign addr[340]= -2079176953;
assign addr[341]= -2134405552;
assign addr[342]= -2146380306;
assign addr[343]= -2114858546;
assign addr[344]= -2040479063;
assign addr[345]= -1924749160;
assign addr[346]= -1770014111;
assign addr[347]= -1579409630;
assign addr[348]= -1356798326;
assign addr[349]= -1106691431;
assign addr[350]= -834157373;
assign addr[351]= -544719071;
assign addr[352]= -244242007;
assign addr[353]= 61184634;
assign addr[354]= 365371365;
assign addr[355]= 662153826;
assign addr[356]= 945517704;
assign addr[357]= 1209720613;
assign addr[358]= 1449408469;
assign addr[359]= 1659723983;
assign addr[360]= 1836405100;
assign addr[361]= 1975871368;
assign addr[362]= 2075296495;
assign addr[363]= 2132665626;
assign addr[364]= 2146816171;
assign addr[365]= 2117461370;
assign addr[366]= 2045196100;
assign addr[367]= 1931484818;
assign addr[368]= 1778631892;
assign addr[369]= 1589734894;
assign addr[370]= 1368621831;
assign addr[371]= 1119773573;
assign addr[372]= 848233042;
assign addr[373]= 559503022;
assign addr[374]= 259434643;
assign addr[375]= -45891193;
assign addr[376]= -350287041;
assign addr[377]= -647584304;
assign addr[378]= -931758235;
assign addr[379]= -1197050035;
assign addr[380]= -1438083551;
assign addr[381]= -1649974225;
assign addr[382]= -1828428082;
assign addr[383]= -1969828744;
assign addr[384]= -2071310720;
assign addr[385]= -2130817471;
assign addr[386]= -2147143090;
assign addr[387]= -2119956737;
assign addr[388]= -2049809346;
assign addr[389]= -1938122457;
assign addr[390]= -1787159411;
assign addr[391]= -1599979481;
assign addr[392]= -1380375881;
assign addr[393]= -1132798888;
assign addr[394]= -862265664;
assign addr[395]= -574258580;
assign addr[396]= -274614114;
assign addr[397]= 30595422;
assign addr[398]= 335184940;
assign addr[399]= 632981917;
assign addr[400]= 917951481;
assign addr[401]= 1184318708;
assign addr[402]= 1426685652;
assign addr[403]= 1640140734;
assign addr[404]= 1820358275;
assign addr[405]= 1963686155;
assign addr[406]= 2067219829;
assign addr[407]= 2128861181;
assign addr[408]= 2147361045;
assign addr[409]= 2122344521;
assign addr[410]= 2054318569;
assign addr[411]= 1944661739;
assign addr[412]= 1795596234;
assign addr[413]= 1610142873;
assign addr[414]= 1392059879;
assign addr[415]= 1145766716;
assign addr[416]= 876254528;
assign addr[417]= 588984994;
assign addr[418]= 289779648;
assign addr[419]= -15298099;
assign addr[420]= -320065829;
assign addr[421]= -618347408;
assign addr[422]= -904098143;
assign addr[423]= -1171527280;
assign addr[424]= -1415215352;
assign addr[425]= -1630224009;
assign addr[426]= -1812196087;
assign addr[427]= -1957443913;
assign addr[428]= -2063024031;
assign addr[429]= -2126796855;
assign addr[430]= -2147470025;
assign addr[431]= -2124624598;
assign addr[432]= -2058723538;
assign addr[433]= -1951102334;
assign addr[434]= -1803941934;
assign addr[435]= -1620224553;
assign addr[436]= -1403673233;
assign addr[437]= -1158676398;
assign addr[438]= -890198924;
assign addr[439]= -603681519;
assign addr[440]= -304930476;
assign addr[441]= 0;
assign addr[442]= 304930476;
assign addr[443]= 603681519;
assign addr[444]= 890198924;
assign addr[445]= 1158676398;
assign addr[446]= 1403673233;
assign addr[447]= 1620224553;
assign addr[448]= 1803941934;
assign addr[449]= 1951102334;
assign addr[450]= 2058723538;
assign addr[451]= 2124624598;
assign addr[452]= 2147470025;
assign addr[453]= 2126796855;
assign addr[454]= 2063024031;
assign addr[455]= 1957443913;
assign addr[456]= 1812196087;
assign addr[457]= 1630224009;
assign addr[458]= 1415215352;
assign addr[459]= 1171527280;
assign addr[460]= 904098143;
assign addr[461]= 618347408;
assign addr[462]= 320065829;
assign addr[463]= 15298099;
assign addr[464]= -289779648;
assign addr[465]= -588984994;
assign addr[466]= -876254528;
assign addr[467]= -1145766716;
assign addr[468]= -1392059879;
assign addr[469]= -1610142873;
assign addr[470]= -1795596234;
assign addr[471]= -1944661739;
assign addr[472]= -2054318569;
assign addr[473]= -2122344521;
assign addr[474]= -2147361045;
assign addr[475]= -2128861181;
assign addr[476]= -2067219829;
assign addr[477]= -1963686155;
assign addr[478]= -1820358275;
assign addr[479]= -1640140734;
assign addr[480]= -1426685652;
assign addr[481]= -1184318708;
assign addr[482]= -917951481;
assign addr[483]= -632981917;
assign addr[484]= -335184940;
assign addr[485]= -30595422;
assign addr[486]= 274614114;
assign addr[487]= 574258580;
assign addr[488]= 862265664;
assign addr[489]= 1132798888;
assign addr[490]= 1380375881;
assign addr[491]= 1599979481;
assign addr[492]= 1787159411;
assign addr[493]= 1938122457;
assign addr[494]= 2049809346;
assign addr[495]= 2119956737;
assign addr[496]= 2147143090;
assign addr[497]= 2130817471;
assign addr[498]= 2071310720;
assign addr[499]= 1969828744;
assign addr[500]= 1828428082;
assign addr[501]= 1649974225;
assign addr[502]= 1438083551;
assign addr[503]= 1197050035;
assign addr[504]= 931758235;
assign addr[505]= 647584304;
assign addr[506]= 350287041;
assign addr[507]= 45891193;
assign addr[508]= -259434643;
assign addr[509]= -559503022;
assign addr[510]= -848233042;
assign addr[511]= -1119773573;
assign addr[512]= -1368621831;
assign addr[513]= -1589734894;
assign addr[514]= -1778631892;
assign addr[515]= -1931484818;
assign addr[516]= -2045196100;
assign addr[517]= -2117461370;
assign addr[518]= -2146816171;
assign addr[519]= -2132665626;
assign addr[520]= -2075296495;
assign addr[521]= -1975871368;
assign addr[522]= -1836405100;
assign addr[523]= -1659723983;
assign addr[524]= -1449408469;
assign addr[525]= -1209720613;
assign addr[526]= -945517704;
assign addr[527]= -662153826;
assign addr[528]= -365371365;
assign addr[529]= -61184634;
assign addr[530]= 244242007;
assign addr[531]= 544719071;
assign addr[532]= 834157373;
assign addr[533]= 1106691431;
assign addr[534]= 1356798326;
assign addr[535]= 1579409630;
assign addr[536]= 1770014111;
assign addr[537]= 1924749160;
assign addr[538]= 2040479063;
assign addr[539]= 2114858546;
assign addr[540]= 2146380306;
assign addr[541]= 2134405552;
assign addr[542]= 2079176953;
assign addr[543]= 1981813720;
assign addr[544]= 1844288924;
assign addr[545]= 1669389513;
assign addr[546]= 1460659832;
assign addr[547]= 1222329801;
assign addr[548]= 959229189;
assign addr[549]= 676689746;
assign addr[550]= 380437148;
assign addr[551]= 76474970;
assign addr[552]= -229036977;
assign addr[553]= -529907477;
assign addr[554]= -820039373;
assign addr[555]= -1093553126;
assign addr[556]= -1344905966;
assign addr[557]= -1569004214;
assign addr[558]= -1761306505;
assign addr[559]= -1917915825;
assign addr[560]= -2035658475;
assign addr[561]= -2112148396;
assign addr[562]= -2145835515;
assign addr[563]= -2136037160;
assign addr[564]= -2082951896;
assign addr[565]= -1987655498;
assign addr[566]= -1852079154;
assign addr[567]= -1678970324;
assign addr[568]= -1471837070;
assign addr[569]= -1234876957;
assign addr[570]= -972891995;
assign addr[571]= -691191324;
assign addr[572]= -395483624;
assign addr[573]= -91761426;
assign addr[574]= 213820322;
assign addr[575]= 515068990;
assign addr[576]= 805879757;
assign addr[577]= 1080359326;
assign addr[578]= 1332945355;
assign addr[579]= 1558519173;
assign addr[580]= 1752509516;
assign addr[581]= 1910985158;
assign addr[582]= 2030734582;
assign addr[583]= 2109331059;
assign addr[584]= 2145181827;
assign addr[585]= 2137560369;
assign addr[586]= 2086621133;
assign addr[587]= 1993396407;
assign addr[588]= 1859775393;
assign addr[589]= 1688465931;
assign addr[590]= 1482939614;
assign addr[591]= 1247361445;
assign addr[592]= 986505429;
assign addr[593]= 705657826;
assign addr[594]= 410510029;
assign addr[595]= 107043224;
assign addr[596]= -198592817;
assign addr[597]= -500204365;
assign addr[598]= -791679244;
assign addr[599]= -1067110699;
assign addr[600]= -1320917099;
assign addr[601]= -1547955041;
assign addr[602]= -1743623590;
assign addr[603]= -1903957513;
assign addr[604]= -2025707632;
assign addr[605]= -2106406677;
assign addr[606]= -2144419275;
assign addr[607]= -2138975100;
assign addr[608]= -2090184478;
assign addr[609]= -1999036154;
assign addr[610]= -1867377253;
assign addr[611]= -1697875851;
assign addr[612]= -1493966902;
assign addr[613]= -1259782632;
assign addr[614]= -1000068799;
assign addr[615]= -720088517;
assign addr[616]= -425515602;
assign addr[617]= -122319591;
assign addr[618]= 183355234;
assign addr[619]= 485314355;
assign addr[620]= 777438554;
assign addr[621]= 1053807919;
assign addr[622]= 1308821808;
assign addr[623]= 1537312353;
assign addr[624]= 1734649179;
assign addr[625]= 1896833245;
assign addr[626]= 2020577882;
assign addr[627]= 2103375398;
assign addr[628]= 2143547897;
assign addr[629]= 2140281282;
assign addr[630]= 2093641749;
assign addr[631]= 2004574453;
assign addr[632]= 1874884346;
assign addr[633]= 1707199606;
assign addr[634]= 1504918373;
assign addr[635]= 1272139887;
assign addr[636]= 1013581418;
assign addr[637]= 734482665;
assign addr[638]= 440499581;
assign addr[639]= 137589750;
assign addr[640]= -168108346;
assign addr[641]= -470399716;
assign addr[642]= -763158411;
assign addr[643]= -1040451659;
assign addr[644]= -1296660098;
assign addr[645]= -1526591649;
assign addr[646]= -1725586737;
assign addr[647]= -1889612716;
assign addr[648]= -2015345591;
assign addr[649]= -2100237377;
assign addr[650]= -2142567738;
assign addr[651]= -2141478848;
assign addr[652]= -2096992772;
assign addr[653]= -2010011024;
assign addr[654]= -1882296293;
assign addr[655]= -1716436725;
assign addr[656]= -1515793473;
assign addr[657]= -1284432584;
assign addr[658]= -1027042599;
assign addr[659]= -748839539;
assign addr[660]= -455461206;
assign addr[661]= -152852926;
assign addr[662]= 152852926;
assign addr[663]= 455461206;
assign addr[664]= 748839539;
assign addr[665]= 1027042599;
assign addr[666]= 1284432584;
assign addr[667]= 1515793473;
assign addr[668]= 1716436725;
assign addr[669]= 1882296293;
assign addr[670]= 2010011024;
assign addr[671]= 2096992772;
assign addr[672]= 2141478848;
assign addr[673]= 2142567738;
assign addr[674]= 2100237377;
assign addr[675]= 2015345591;
assign addr[676]= 1889612716;
assign addr[677]= 1725586737;
assign addr[678]= 1526591649;
assign addr[679]= 1296660098;
assign addr[680]= 1040451659;
assign addr[681]= 763158411;
assign addr[682]= 470399716;
assign addr[683]= 168108346;
assign addr[684]= -137589750;
assign addr[685]= -440499581;
assign addr[686]= -734482665;
assign addr[687]= -1013581418;
assign addr[688]= -1272139887;
assign addr[689]= -1504918373;
assign addr[690]= -1707199606;
assign addr[691]= -1874884346;
assign addr[692]= -2004574453;
assign addr[693]= -2093641749;
assign addr[694]= -2140281282;
assign addr[695]= -2143547897;
assign addr[696]= -2103375398;
assign addr[697]= -2020577882;
assign addr[698]= -1896833245;
assign addr[699]= -1734649179;
assign addr[700]= -1537312353;
assign addr[701]= -1308821808;
assign addr[702]= -1053807919;
assign addr[703]= -777438554;
assign addr[704]= -485314355;
assign addr[705]= -183355234;
assign addr[706]= 122319591;
assign addr[707]= 425515602;
assign addr[708]= 720088517;
assign addr[709]= 1000068799;
assign addr[710]= 1259782632;
assign addr[711]= 1493966902;
assign addr[712]= 1697875851;
assign addr[713]= 1867377253;
assign addr[714]= 1999036154;
assign addr[715]= 2090184478;
assign addr[716]= 2138975100;
assign addr[717]= 2144419275;
assign addr[718]= 2106406677;
assign addr[719]= 2025707632;
assign addr[720]= 1903957513;
assign addr[721]= 1743623590;
assign addr[722]= 1547955041;
assign addr[723]= 1320917099;
assign addr[724]= 1067110699;
assign addr[725]= 791679244;
assign addr[726]= 500204365;
assign addr[727]= 198592817;
assign addr[728]= -107043224;
assign addr[729]= -410510029;
assign addr[730]= -705657826;
assign addr[731]= -986505429;
assign addr[732]= -1247361445;
assign addr[733]= -1482939614;
assign addr[734]= -1688465931;
assign addr[735]= -1859775393;
assign addr[736]= -1993396407;
assign addr[737]= -2086621133;
assign addr[738]= -2137560369;
assign addr[739]= -2145181827;
assign addr[740]= -2109331059;
assign addr[741]= -2030734582;
assign addr[742]= -1910985158;
assign addr[743]= -1752509516;
assign addr[744]= -1558519173;
assign addr[745]= -1332945355;
assign addr[746]= -1080359326;
assign addr[747]= -805879757;
assign addr[748]= -515068990;
assign addr[749]= -213820322;
assign addr[750]= 91761426;
assign addr[751]= 395483624;
assign addr[752]= 691191324;
assign addr[753]= 972891995;
assign addr[754]= 1234876957;
assign addr[755]= 1471837070;
assign addr[756]= 1678970324;
assign addr[757]= 1852079154;
assign addr[758]= 1987655498;
assign addr[759]= 2082951896;
assign addr[760]= 2136037160;
assign addr[761]= 2145835515;
assign addr[762]= 2112148396;
assign addr[763]= 2035658475;
assign addr[764]= 1917915825;
assign addr[765]= 1761306505;
assign addr[766]= 1569004214;
assign addr[767]= 1344905966;
assign addr[768]= 1093553126;
assign addr[769]= 820039373;
assign addr[770]= 529907477;
assign addr[771]= 229036977;
assign addr[772]= -76474970;
assign addr[773]= -380437148;
assign addr[774]= -676689746;
assign addr[775]= -959229189;
assign addr[776]= -1222329801;
assign addr[777]= -1460659832;
assign addr[778]= -1669389513;
assign addr[779]= -1844288924;
assign addr[780]= -1981813720;
assign addr[781]= -2079176953;
assign addr[782]= -2134405552;
assign addr[783]= -2146380306;
assign addr[784]= -2114858546;
assign addr[785]= -2040479063;
assign addr[786]= -1924749160;
assign addr[787]= -1770014111;
assign addr[788]= -1579409630;
assign addr[789]= -1356798326;
assign addr[790]= -1106691431;
assign addr[791]= -834157373;
assign addr[792]= -544719071;
assign addr[793]= -244242007;
assign addr[794]= 61184634;
assign addr[795]= 365371365;
assign addr[796]= 662153826;
assign addr[797]= 945517704;
assign addr[798]= 1209720613;
assign addr[799]= 1449408469;
assign addr[800]= 1659723983;
assign addr[801]= 1836405100;
assign addr[802]= 1975871368;
assign addr[803]= 2075296495;
assign addr[804]= 2132665626;
assign addr[805]= 2146816171;
assign addr[806]= 2117461370;
assign addr[807]= 2045196100;
assign addr[808]= 1931484818;
assign addr[809]= 1778631892;
assign addr[810]= 1589734894;
assign addr[811]= 1368621831;
assign addr[812]= 1119773573;
assign addr[813]= 848233042;
assign addr[814]= 559503022;
assign addr[815]= 259434643;
assign addr[816]= -45891193;
assign addr[817]= -350287041;
assign addr[818]= -647584304;
assign addr[819]= -931758235;
assign addr[820]= -1197050035;
assign addr[821]= -1438083551;
assign addr[822]= -1649974225;
assign addr[823]= -1828428082;
assign addr[824]= -1969828744;
assign addr[825]= -2071310720;
assign addr[826]= -2130817471;
assign addr[827]= -2147143090;
assign addr[828]= -2119956737;
assign addr[829]= -2049809346;
assign addr[830]= -1938122457;
assign addr[831]= -1787159411;
assign addr[832]= -1599979481;
assign addr[833]= -1380375881;
assign addr[834]= -1132798888;
assign addr[835]= -862265664;
assign addr[836]= -574258580;
assign addr[837]= -274614114;
assign addr[838]= 30595422;
assign addr[839]= 335184940;
assign addr[840]= 632981917;
assign addr[841]= 917951481;
assign addr[842]= 1184318708;
assign addr[843]= 1426685652;
assign addr[844]= 1640140734;
assign addr[845]= 1820358275;
assign addr[846]= 1963686155;
assign addr[847]= 2067219829;
assign addr[848]= 2128861181;
assign addr[849]= 2147361045;
assign addr[850]= 2122344521;
assign addr[851]= 2054318569;
assign addr[852]= 1944661739;
assign addr[853]= 1795596234;
assign addr[854]= 1610142873;
assign addr[855]= 1392059879;
assign addr[856]= 1145766716;
assign addr[857]= 876254528;
assign addr[858]= 588984994;
assign addr[859]= 289779648;
assign addr[860]= -15298099;
assign addr[861]= -320065829;
assign addr[862]= -618347408;
assign addr[863]= -904098143;
assign addr[864]= -1171527280;
assign addr[865]= -1415215352;
assign addr[866]= -1630224009;
assign addr[867]= -1812196087;
assign addr[868]= -1957443913;
assign addr[869]= -2063024031;
assign addr[870]= -2126796855;
assign addr[871]= -2147470025;
assign addr[872]= -2124624598;
assign addr[873]= -2058723538;
assign addr[874]= -1951102334;
assign addr[875]= -1803941934;
assign addr[876]= -1620224553;
assign addr[877]= -1403673233;
assign addr[878]= -1158676398;
assign addr[879]= -890198924;
assign addr[880]= -603681519;
assign addr[881]= -304930476;
assign addr[882]= 0;
assign addr[883]= 304930476;
assign addr[884]= 603681519;
assign addr[885]= 890198924;
assign addr[886]= 1158676398;
assign addr[887]= 1403673233;
assign addr[888]= 1620224553;
assign addr[889]= 1803941934;
assign addr[890]= 1951102334;
assign addr[891]= 2058723538;
assign addr[892]= 2124624598;
assign addr[893]= 2147470025;
assign addr[894]= 2126796855;
assign addr[895]= 2063024031;
assign addr[896]= 1957443913;
assign addr[897]= 1812196087;
assign addr[898]= 1630224009;
assign addr[899]= 1415215352;
assign addr[900]= 1171527280;
assign addr[901]= 904098143;
assign addr[902]= 618347408;
assign addr[903]= 320065829;
assign addr[904]= 15298099;
assign addr[905]= -289779648;
assign addr[906]= -588984994;
assign addr[907]= -876254528;
assign addr[908]= -1145766716;
assign addr[909]= -1392059879;
assign addr[910]= -1610142873;
assign addr[911]= -1795596234;
assign addr[912]= -1944661739;
assign addr[913]= -2054318569;
assign addr[914]= -2122344521;
assign addr[915]= -2147361045;
assign addr[916]= -2128861181;
assign addr[917]= -2067219829;
assign addr[918]= -1963686155;
assign addr[919]= -1820358275;
assign addr[920]= -1640140734;
assign addr[921]= -1426685652;
assign addr[922]= -1184318708;
assign addr[923]= -917951481;
assign addr[924]= -632981917;
assign addr[925]= -335184940;
assign addr[926]= -30595422;
assign addr[927]= 274614114;
assign addr[928]= 574258580;
assign addr[929]= 862265664;
assign addr[930]= 1132798888;
assign addr[931]= 1380375881;
assign addr[932]= 1599979481;
assign addr[933]= 1787159411;
assign addr[934]= 1938122457;
assign addr[935]= 2049809346;
assign addr[936]= 2119956737;
assign addr[937]= 2147143090;
assign addr[938]= 2130817471;
assign addr[939]= 2071310720;
assign addr[940]= 1969828744;
assign addr[941]= 1828428082;
assign addr[942]= 1649974225;
assign addr[943]= 1438083551;
assign addr[944]= 1197050035;
assign addr[945]= 931758235;
assign addr[946]= 647584304;
assign addr[947]= 350287041;
assign addr[948]= 45891193;
assign addr[949]= -259434643;
assign addr[950]= -559503022;
assign addr[951]= -848233042;
assign addr[952]= -1119773573;
assign addr[953]= -1368621831;
assign addr[954]= -1589734894;
assign addr[955]= -1778631892;
assign addr[956]= -1931484818;
assign addr[957]= -2045196100;
assign addr[958]= -2117461370;
assign addr[959]= -2146816171;
assign addr[960]= -2132665626;
assign addr[961]= -2075296495;
assign addr[962]= -1975871368;
assign addr[963]= -1836405100;
assign addr[964]= -1659723983;
assign addr[965]= -1449408469;
assign addr[966]= -1209720613;
assign addr[967]= -945517704;
assign addr[968]= -662153826;
assign addr[969]= -365371365;
assign addr[970]= -61184634;
assign addr[971]= 244242007;
assign addr[972]= 544719071;
assign addr[973]= 834157373;
assign addr[974]= 1106691431;
assign addr[975]= 1356798326;
assign addr[976]= 1579409630;
assign addr[977]= 1770014111;
assign addr[978]= 1924749160;
assign addr[979]= 2040479063;
assign addr[980]= 2114858546;
assign addr[981]= 2146380306;
assign addr[982]= 2134405552;
assign addr[983]= 2079176953;
assign addr[984]= 1981813720;
assign addr[985]= 1844288924;
assign addr[986]= 1669389513;
assign addr[987]= 1460659832;
assign addr[988]= 1222329801;
assign addr[989]= 959229189;
assign addr[990]= 676689746;
assign addr[991]= 380437148;
assign addr[992]= 76474970;
assign addr[993]= -229036977;
assign addr[994]= -529907477;
assign addr[995]= -820039373;
assign addr[996]= -1093553126;
assign addr[997]= -1344905966;
assign addr[998]= -1569004214;
assign addr[999]= -1761306505;
assign addr[1000]= -1917915825;
assign addr[1001]= -2035658475;
assign addr[1002]= -2112148396;
assign addr[1003]= -2145835515;
assign addr[1004]= -2136037160;
assign addr[1005]= -2082951896;
assign addr[1006]= -1987655498;
assign addr[1007]= -1852079154;
assign addr[1008]= -1678970324;
assign addr[1009]= -1471837070;
assign addr[1010]= -1234876957;
assign addr[1011]= -972891995;
assign addr[1012]= -691191324;
assign addr[1013]= -395483624;
assign addr[1014]= -91761426;
assign addr[1015]= 213820322;
assign addr[1016]= 515068990;
assign addr[1017]= 805879757;
assign addr[1018]= 1080359326;
assign addr[1019]= 1332945355;
assign addr[1020]= 1558519173;
assign addr[1021]= 1752509516;
assign addr[1022]= 1910985158;
assign addr[1023]= 2030734582;
assign addr[1024]= 2109331059;
assign addr[1025]= 2145181827;
assign addr[1026]= 2137560369;
assign addr[1027]= 2086621133;
assign addr[1028]= 1993396407;
assign addr[1029]= 1859775393;
assign addr[1030]= 1688465931;
assign addr[1031]= 1482939614;
assign addr[1032]= 1247361445;
assign addr[1033]= 986505429;
assign addr[1034]= 705657826;
assign addr[1035]= 410510029;
assign addr[1036]= 107043224;
assign addr[1037]= -198592817;
assign addr[1038]= -500204365;
assign addr[1039]= -791679244;
assign addr[1040]= -1067110699;
assign addr[1041]= -1320917099;
assign addr[1042]= -1547955041;
assign addr[1043]= -1743623590;
assign addr[1044]= -1903957513;
assign addr[1045]= -2025707632;
assign addr[1046]= -2106406677;
assign addr[1047]= -2144419275;
assign addr[1048]= -2138975100;
assign addr[1049]= -2090184478;
assign addr[1050]= -1999036154;
assign addr[1051]= -1867377253;
assign addr[1052]= -1697875851;
assign addr[1053]= -1493966902;
assign addr[1054]= -1259782632;
assign addr[1055]= -1000068799;
assign addr[1056]= -720088517;
assign addr[1057]= -425515602;
assign addr[1058]= -122319591;
assign addr[1059]= 183355234;
assign addr[1060]= 485314355;
assign addr[1061]= 777438554;
assign addr[1062]= 1053807919;
assign addr[1063]= 1308821808;
assign addr[1064]= 1537312353;
assign addr[1065]= 1734649179;
assign addr[1066]= 1896833245;
assign addr[1067]= 2020577882;
assign addr[1068]= 2103375398;
assign addr[1069]= 2143547897;
assign addr[1070]= 2140281282;
assign addr[1071]= 2093641749;
assign addr[1072]= 2004574453;
assign addr[1073]= 1874884346;
assign addr[1074]= 1707199606;
assign addr[1075]= 1504918373;
assign addr[1076]= 1272139887;
assign addr[1077]= 1013581418;
assign addr[1078]= 734482665;
assign addr[1079]= 440499581;
assign addr[1080]= 137589750;
assign addr[1081]= -168108346;
assign addr[1082]= -470399716;
assign addr[1083]= -763158411;
assign addr[1084]= -1040451659;
assign addr[1085]= -1296660098;
assign addr[1086]= -1526591649;
assign addr[1087]= -1725586737;
assign addr[1088]= -1889612716;
assign addr[1089]= -2015345591;
assign addr[1090]= -2100237377;
assign addr[1091]= -2142567738;
assign addr[1092]= -2141478848;
assign addr[1093]= -2096992772;
assign addr[1094]= -2010011024;
assign addr[1095]= -1882296293;
assign addr[1096]= -1716436725;
assign addr[1097]= -1515793473;
assign addr[1098]= -1284432584;
assign addr[1099]= -1027042599;
assign addr[1100]= -748839539;
assign addr[1101]= -455461206;
assign addr[1102]= -152852926;
assign addr[1103]= 152852926;
assign addr[1104]= 455461206;
assign addr[1105]= 748839539;
assign addr[1106]= 1027042599;
assign addr[1107]= 1284432584;
assign addr[1108]= 1515793473;
assign addr[1109]= 1716436725;
assign addr[1110]= 1882296293;
assign addr[1111]= 2010011024;
assign addr[1112]= 2096992772;
assign addr[1113]= 2141478848;
assign addr[1114]= 2142567738;
assign addr[1115]= 2100237377;
assign addr[1116]= 2015345591;
assign addr[1117]= 1889612716;
assign addr[1118]= 1725586737;
assign addr[1119]= 1526591649;
assign addr[1120]= 1296660098;
assign addr[1121]= 1040451659;
assign addr[1122]= 763158411;
assign addr[1123]= 470399716;
assign addr[1124]= 168108346;
assign addr[1125]= -137589750;
assign addr[1126]= -440499581;
assign addr[1127]= -734482665;
assign addr[1128]= -1013581418;
assign addr[1129]= -1272139887;
assign addr[1130]= -1504918373;
assign addr[1131]= -1707199606;
assign addr[1132]= -1874884346;
assign addr[1133]= -2004574453;
assign addr[1134]= -2093641749;
assign addr[1135]= -2140281282;
assign addr[1136]= -2143547897;
assign addr[1137]= -2103375398;
assign addr[1138]= -2020577882;
assign addr[1139]= -1896833245;
assign addr[1140]= -1734649179;
assign addr[1141]= -1537312353;
assign addr[1142]= -1308821808;
assign addr[1143]= -1053807919;
assign addr[1144]= -777438554;
assign addr[1145]= -485314355;
assign addr[1146]= -183355234;
assign addr[1147]= 122319591;
assign addr[1148]= 425515602;
assign addr[1149]= 720088517;
assign addr[1150]= 1000068799;
assign addr[1151]= 1259782632;
assign addr[1152]= 1493966902;
assign addr[1153]= 1697875851;
assign addr[1154]= 1867377253;
assign addr[1155]= 1999036154;
assign addr[1156]= 2090184478;
assign addr[1157]= 2138975100;
assign addr[1158]= 2144419275;
assign addr[1159]= 2106406677;
assign addr[1160]= 2025707632;
assign addr[1161]= 1903957513;
assign addr[1162]= 1743623590;
assign addr[1163]= 1547955041;
assign addr[1164]= 1320917099;
assign addr[1165]= 1067110699;
assign addr[1166]= 791679244;
assign addr[1167]= 500204365;
assign addr[1168]= 198592817;
assign addr[1169]= -107043224;
assign addr[1170]= -410510029;
assign addr[1171]= -705657826;
assign addr[1172]= -986505429;
assign addr[1173]= -1247361445;
assign addr[1174]= -1482939614;
assign addr[1175]= -1688465931;
assign addr[1176]= -1859775393;
assign addr[1177]= -1993396407;
assign addr[1178]= -2086621133;
assign addr[1179]= -2137560369;
assign addr[1180]= -2145181827;
assign addr[1181]= -2109331059;
assign addr[1182]= -2030734582;
assign addr[1183]= -1910985158;
assign addr[1184]= -1752509516;
assign addr[1185]= -1558519173;
assign addr[1186]= -1332945355;
assign addr[1187]= -1080359326;
assign addr[1188]= -805879757;
assign addr[1189]= -515068990;
assign addr[1190]= -213820322;
assign addr[1191]= 91761426;
assign addr[1192]= 395483624;
assign addr[1193]= 691191324;
assign addr[1194]= 972891995;
assign addr[1195]= 1234876957;
assign addr[1196]= 1471837070;
assign addr[1197]= 1678970324;
assign addr[1198]= 1852079154;
assign addr[1199]= 1987655498;
assign addr[1200]= 2082951896;
assign addr[1201]= 2136037160;
assign addr[1202]= 2145835515;
assign addr[1203]= 2112148396;
assign addr[1204]= 2035658475;
assign addr[1205]= 1917915825;
assign addr[1206]= 1761306505;
assign addr[1207]= 1569004214;
assign addr[1208]= 1344905966;
assign addr[1209]= 1093553126;
assign addr[1210]= 820039373;
assign addr[1211]= 529907477;
assign addr[1212]= 229036977;
assign addr[1213]= -76474970;
assign addr[1214]= -380437148;
assign addr[1215]= -676689746;
assign addr[1216]= -959229189;
assign addr[1217]= -1222329801;
assign addr[1218]= -1460659832;
assign addr[1219]= -1669389513;
assign addr[1220]= -1844288924;
assign addr[1221]= -1981813720;
assign addr[1222]= -2079176953;
assign addr[1223]= -2134405552;
assign addr[1224]= -2146380306;
assign addr[1225]= -2114858546;
assign addr[1226]= -2040479063;
assign addr[1227]= -1924749160;
assign addr[1228]= -1770014111;
assign addr[1229]= -1579409630;
assign addr[1230]= -1356798326;
assign addr[1231]= -1106691431;
assign addr[1232]= -834157373;
assign addr[1233]= -544719071;
assign addr[1234]= -244242007;
assign addr[1235]= 61184634;
assign addr[1236]= 365371365;
assign addr[1237]= 662153826;
assign addr[1238]= 945517704;
assign addr[1239]= 1209720613;
assign addr[1240]= 1449408469;
assign addr[1241]= 1659723983;
assign addr[1242]= 1836405100;
assign addr[1243]= 1975871368;
assign addr[1244]= 2075296495;
assign addr[1245]= 2132665626;
assign addr[1246]= 2146816171;
assign addr[1247]= 2117461370;
assign addr[1248]= 2045196100;
assign addr[1249]= 1931484818;
assign addr[1250]= 1778631892;
assign addr[1251]= 1589734894;
assign addr[1252]= 1368621831;
assign addr[1253]= 1119773573;
assign addr[1254]= 848233042;
assign addr[1255]= 559503022;
assign addr[1256]= 259434643;
assign addr[1257]= -45891193;
assign addr[1258]= -350287041;
assign addr[1259]= -647584304;
assign addr[1260]= -931758235;
assign addr[1261]= -1197050035;
assign addr[1262]= -1438083551;
assign addr[1263]= -1649974225;
assign addr[1264]= -1828428082;
assign addr[1265]= -1969828744;
assign addr[1266]= -2071310720;
assign addr[1267]= -2130817471;
assign addr[1268]= -2147143090;
assign addr[1269]= -2119956737;
assign addr[1270]= -2049809346;
assign addr[1271]= -1938122457;
assign addr[1272]= -1787159411;
assign addr[1273]= -1599979481;
assign addr[1274]= -1380375881;
assign addr[1275]= -1132798888;
assign addr[1276]= -862265664;
assign addr[1277]= -574258580;
assign addr[1278]= -274614114;
assign addr[1279]= 30595422;
assign addr[1280]= 335184940;
assign addr[1281]= 632981917;
assign addr[1282]= 917951481;
assign addr[1283]= 1184318708;
assign addr[1284]= 1426685652;
assign addr[1285]= 1640140734;
assign addr[1286]= 1820358275;
assign addr[1287]= 1963686155;
assign addr[1288]= 2067219829;
assign addr[1289]= 2128861181;
assign addr[1290]= 2147361045;
assign addr[1291]= 2122344521;
assign addr[1292]= 2054318569;
assign addr[1293]= 1944661739;
assign addr[1294]= 1795596234;
assign addr[1295]= 1610142873;
assign addr[1296]= 1392059879;
assign addr[1297]= 1145766716;
assign addr[1298]= 876254528;
assign addr[1299]= 588984994;
assign addr[1300]= 289779648;
assign addr[1301]= -15298099;
assign addr[1302]= -320065829;
assign addr[1303]= -618347408;
assign addr[1304]= -904098143;
assign addr[1305]= -1171527280;
assign addr[1306]= -1415215352;
assign addr[1307]= -1630224009;
assign addr[1308]= -1812196087;
assign addr[1309]= -1957443913;
assign addr[1310]= -2063024031;
assign addr[1311]= -2126796855;
assign addr[1312]= -2147470025;
assign addr[1313]= -2124624598;
assign addr[1314]= -2058723538;
assign addr[1315]= -1951102334;
assign addr[1316]= -1803941934;
assign addr[1317]= -1620224553;
assign addr[1318]= -1403673233;
assign addr[1319]= -1158676398;
assign addr[1320]= -890198924;
assign addr[1321]= -603681519;
assign addr[1322]= -304930476;
assign addr[1323]= 0;
assign addr[1324]= 304930476;
assign addr[1325]= 603681519;
assign addr[1326]= 890198924;
assign addr[1327]= 1158676398;
assign addr[1328]= 1403673233;
assign addr[1329]= 1620224553;
assign addr[1330]= 1803941934;
assign addr[1331]= 1951102334;
assign addr[1332]= 2058723538;
assign addr[1333]= 2124624598;
assign addr[1334]= 2147470025;
assign addr[1335]= 2126796855;
assign addr[1336]= 2063024031;
assign addr[1337]= 1957443913;
assign addr[1338]= 1812196087;
assign addr[1339]= 1630224009;
assign addr[1340]= 1415215352;
assign addr[1341]= 1171527280;
assign addr[1342]= 904098143;
assign addr[1343]= 618347408;
assign addr[1344]= 320065829;
assign addr[1345]= 15298099;
assign addr[1346]= -289779648;
assign addr[1347]= -588984994;
assign addr[1348]= -876254528;
assign addr[1349]= -1145766716;
assign addr[1350]= -1392059879;
assign addr[1351]= -1610142873;
assign addr[1352]= -1795596234;
assign addr[1353]= -1944661739;
assign addr[1354]= -2054318569;
assign addr[1355]= -2122344521;
assign addr[1356]= -2147361045;
assign addr[1357]= -2128861181;
assign addr[1358]= -2067219829;
assign addr[1359]= -1963686155;
assign addr[1360]= -1820358275;
assign addr[1361]= -1640140734;
assign addr[1362]= -1426685652;
assign addr[1363]= -1184318708;
assign addr[1364]= -917951481;
assign addr[1365]= -632981917;
assign addr[1366]= -335184940;
assign addr[1367]= -30595422;
assign addr[1368]= 274614114;
assign addr[1369]= 574258580;
assign addr[1370]= 862265664;
assign addr[1371]= 1132798888;
assign addr[1372]= 1380375881;
assign addr[1373]= 1599979481;
assign addr[1374]= 1787159411;
assign addr[1375]= 1938122457;
assign addr[1376]= 2049809346;
assign addr[1377]= 2119956737;
assign addr[1378]= 2147143090;
assign addr[1379]= 2130817471;
assign addr[1380]= 2071310720;
assign addr[1381]= 1969828744;
assign addr[1382]= 1828428082;
assign addr[1383]= 1649974225;
assign addr[1384]= 1438083551;
assign addr[1385]= 1197050035;
assign addr[1386]= 931758235;
assign addr[1387]= 647584304;
assign addr[1388]= 350287041;
assign addr[1389]= 45891193;
assign addr[1390]= -259434643;
assign addr[1391]= -559503022;
assign addr[1392]= -848233042;
assign addr[1393]= -1119773573;
assign addr[1394]= -1368621831;
assign addr[1395]= -1589734894;
assign addr[1396]= -1778631892;
assign addr[1397]= -1931484818;
assign addr[1398]= -2045196100;
assign addr[1399]= -2117461370;
assign addr[1400]= -2146816171;
assign addr[1401]= -2132665626;
assign addr[1402]= -2075296495;
assign addr[1403]= -1975871368;
assign addr[1404]= -1836405100;
assign addr[1405]= -1659723983;
assign addr[1406]= -1449408469;
assign addr[1407]= -1209720613;
assign addr[1408]= -945517704;
assign addr[1409]= -662153826;
assign addr[1410]= -365371365;
assign addr[1411]= -61184634;
assign addr[1412]= 244242007;
assign addr[1413]= 544719071;
assign addr[1414]= 834157373;
assign addr[1415]= 1106691431;
assign addr[1416]= 1356798326;
assign addr[1417]= 1579409630;
assign addr[1418]= 1770014111;
assign addr[1419]= 1924749160;
assign addr[1420]= 2040479063;
assign addr[1421]= 2114858546;
assign addr[1422]= 2146380306;
assign addr[1423]= 2134405552;
assign addr[1424]= 2079176953;
assign addr[1425]= 1981813720;
assign addr[1426]= 1844288924;
assign addr[1427]= 1669389513;
assign addr[1428]= 1460659832;
assign addr[1429]= 1222329801;
assign addr[1430]= 959229189;
assign addr[1431]= 676689746;
assign addr[1432]= 380437148;
assign addr[1433]= 76474970;
assign addr[1434]= -229036977;
assign addr[1435]= -529907477;
assign addr[1436]= -820039373;
assign addr[1437]= -1093553126;
assign addr[1438]= -1344905966;
assign addr[1439]= -1569004214;
assign addr[1440]= -1761306505;
assign addr[1441]= -1917915825;
assign addr[1442]= -2035658475;
assign addr[1443]= -2112148396;
assign addr[1444]= -2145835515;
assign addr[1445]= -2136037160;
assign addr[1446]= -2082951896;
assign addr[1447]= -1987655498;
assign addr[1448]= -1852079154;
assign addr[1449]= -1678970324;
assign addr[1450]= -1471837070;
assign addr[1451]= -1234876957;
assign addr[1452]= -972891995;
assign addr[1453]= -691191324;
assign addr[1454]= -395483624;
assign addr[1455]= -91761426;
assign addr[1456]= 213820322;
assign addr[1457]= 515068990;
assign addr[1458]= 805879757;
assign addr[1459]= 1080359326;
assign addr[1460]= 1332945355;
assign addr[1461]= 1558519173;
assign addr[1462]= 1752509516;
assign addr[1463]= 1910985158;
assign addr[1464]= 2030734582;
assign addr[1465]= 2109331059;
assign addr[1466]= 2145181827;
assign addr[1467]= 2137560369;
assign addr[1468]= 2086621133;
assign addr[1469]= 1993396407;
assign addr[1470]= 1859775393;
assign addr[1471]= 1688465931;
assign addr[1472]= 1482939614;
assign addr[1473]= 1247361445;
assign addr[1474]= 986505429;
assign addr[1475]= 705657826;
assign addr[1476]= 410510029;
assign addr[1477]= 107043224;
assign addr[1478]= -198592817;
assign addr[1479]= -500204365;
assign addr[1480]= -791679244;
assign addr[1481]= -1067110699;
assign addr[1482]= -1320917099;
assign addr[1483]= -1547955041;
assign addr[1484]= -1743623590;
assign addr[1485]= -1903957513;
assign addr[1486]= -2025707632;
assign addr[1487]= -2106406677;
assign addr[1488]= -2144419275;
assign addr[1489]= -2138975100;
assign addr[1490]= -2090184478;
assign addr[1491]= -1999036154;
assign addr[1492]= -1867377253;
assign addr[1493]= -1697875851;
assign addr[1494]= -1493966902;
assign addr[1495]= -1259782632;
assign addr[1496]= -1000068799;
assign addr[1497]= -720088517;
assign addr[1498]= -425515602;
assign addr[1499]= -122319591;
assign addr[1500]= 183355234;
assign addr[1501]= 485314355;
assign addr[1502]= 777438554;
assign addr[1503]= 1053807919;
assign addr[1504]= 1308821808;
assign addr[1505]= 1537312353;
assign addr[1506]= 1734649179;
assign addr[1507]= 1896833245;
assign addr[1508]= 2020577882;
assign addr[1509]= 2103375398;
assign addr[1510]= 2143547897;
assign addr[1511]= 2140281282;
assign addr[1512]= 2093641749;
assign addr[1513]= 2004574453;
assign addr[1514]= 1874884346;
assign addr[1515]= 1707199606;
assign addr[1516]= 1504918373;
assign addr[1517]= 1272139887;
assign addr[1518]= 1013581418;
assign addr[1519]= 734482665;
assign addr[1520]= 440499581;
assign addr[1521]= 137589750;
assign addr[1522]= -168108346;
assign addr[1523]= -470399716;
assign addr[1524]= -763158411;
assign addr[1525]= -1040451659;
assign addr[1526]= -1296660098;
assign addr[1527]= -1526591649;
assign addr[1528]= -1725586737;
assign addr[1529]= -1889612716;
assign addr[1530]= -2015345591;
assign addr[1531]= -2100237377;
assign addr[1532]= -2142567738;
assign addr[1533]= -2141478848;
assign addr[1534]= -2096992772;
assign addr[1535]= -2010011024;
assign addr[1536]= -1882296293;
assign addr[1537]= -1716436725;
assign addr[1538]= -1515793473;
assign addr[1539]= -1284432584;
assign addr[1540]= -1027042599;
assign addr[1541]= -748839539;
assign addr[1542]= -455461206;
assign addr[1543]= -152852926;
assign addr[1544]= 152852926;
assign addr[1545]= 455461206;
assign addr[1546]= 748839539;
assign addr[1547]= 1027042599;
assign addr[1548]= 1284432584;
assign addr[1549]= 1515793473;
assign addr[1550]= 1716436725;
assign addr[1551]= 1882296293;
assign addr[1552]= 2010011024;
assign addr[1553]= 2096992772;
assign addr[1554]= 2141478848;
assign addr[1555]= 2142567738;
assign addr[1556]= 2100237377;
assign addr[1557]= 2015345591;
assign addr[1558]= 1889612716;
assign addr[1559]= 1725586737;
assign addr[1560]= 1526591649;
assign addr[1561]= 1296660098;
assign addr[1562]= 1040451659;
assign addr[1563]= 763158411;
assign addr[1564]= 470399716;
assign addr[1565]= 168108346;
assign addr[1566]= -137589750;
assign addr[1567]= -440499581;
assign addr[1568]= -734482665;
assign addr[1569]= -1013581418;
assign addr[1570]= -1272139887;
assign addr[1571]= -1504918373;
assign addr[1572]= -1707199606;
assign addr[1573]= -1874884346;
assign addr[1574]= -2004574453;
assign addr[1575]= -2093641749;
assign addr[1576]= -2140281282;
assign addr[1577]= -2143547897;
assign addr[1578]= -2103375398;
assign addr[1579]= -2020577882;
assign addr[1580]= -1896833245;
assign addr[1581]= -1734649179;
assign addr[1582]= -1537312353;
assign addr[1583]= -1308821808;
assign addr[1584]= -1053807919;
assign addr[1585]= -777438554;
assign addr[1586]= -485314355;
assign addr[1587]= -183355234;
assign addr[1588]= 122319591;
assign addr[1589]= 425515602;
assign addr[1590]= 720088517;
assign addr[1591]= 1000068799;
assign addr[1592]= 1259782632;
assign addr[1593]= 1493966902;
assign addr[1594]= 1697875851;
assign addr[1595]= 1867377253;
assign addr[1596]= 1999036154;
assign addr[1597]= 2090184478;
assign addr[1598]= 2138975100;
assign addr[1599]= 2144419275;
assign addr[1600]= 2106406677;
assign addr[1601]= 2025707632;
assign addr[1602]= 1903957513;
assign addr[1603]= 1743623590;
assign addr[1604]= 1547955041;
assign addr[1605]= 1320917099;
assign addr[1606]= 1067110699;
assign addr[1607]= 791679244;
assign addr[1608]= 500204365;
assign addr[1609]= 198592817;
assign addr[1610]= -107043224;
assign addr[1611]= -410510029;
assign addr[1612]= -705657826;
assign addr[1613]= -986505429;
assign addr[1614]= -1247361445;
assign addr[1615]= -1482939614;
assign addr[1616]= -1688465931;
assign addr[1617]= -1859775393;
assign addr[1618]= -1993396407;
assign addr[1619]= -2086621133;
assign addr[1620]= -2137560369;
assign addr[1621]= -2145181827;
assign addr[1622]= -2109331059;
assign addr[1623]= -2030734582;
assign addr[1624]= -1910985158;
assign addr[1625]= -1752509516;
assign addr[1626]= -1558519173;
assign addr[1627]= -1332945355;
assign addr[1628]= -1080359326;
assign addr[1629]= -805879757;
assign addr[1630]= -515068990;
assign addr[1631]= -213820322;
assign addr[1632]= 91761426;
assign addr[1633]= 395483624;
assign addr[1634]= 691191324;
assign addr[1635]= 972891995;
assign addr[1636]= 1234876957;
assign addr[1637]= 1471837070;
assign addr[1638]= 1678970324;
assign addr[1639]= 1852079154;
assign addr[1640]= 1987655498;
assign addr[1641]= 2082951896;
assign addr[1642]= 2136037160;
assign addr[1643]= 2145835515;
assign addr[1644]= 2112148396;
assign addr[1645]= 2035658475;
assign addr[1646]= 1917915825;
assign addr[1647]= 1761306505;
assign addr[1648]= 1569004214;
assign addr[1649]= 1344905966;
assign addr[1650]= 1093553126;
assign addr[1651]= 820039373;
assign addr[1652]= 529907477;
assign addr[1653]= 229036977;
assign addr[1654]= -76474970;
assign addr[1655]= -380437148;
assign addr[1656]= -676689746;
assign addr[1657]= -959229189;
assign addr[1658]= -1222329801;
assign addr[1659]= -1460659832;
assign addr[1660]= -1669389513;
assign addr[1661]= -1844288924;
assign addr[1662]= -1981813720;
assign addr[1663]= -2079176953;
assign addr[1664]= -2134405552;
assign addr[1665]= -2146380306;
assign addr[1666]= -2114858546;
assign addr[1667]= -2040479063;
assign addr[1668]= -1924749160;
assign addr[1669]= -1770014111;
assign addr[1670]= -1579409630;
assign addr[1671]= -1356798326;
assign addr[1672]= -1106691431;
assign addr[1673]= -834157373;
assign addr[1674]= -544719071;
assign addr[1675]= -244242007;
assign addr[1676]= 61184634;
assign addr[1677]= 365371365;
assign addr[1678]= 662153826;
assign addr[1679]= 945517704;
assign addr[1680]= 1209720613;
assign addr[1681]= 1449408469;
assign addr[1682]= 1659723983;
assign addr[1683]= 1836405100;
assign addr[1684]= 1975871368;
assign addr[1685]= 2075296495;
assign addr[1686]= 2132665626;
assign addr[1687]= 2146816171;
assign addr[1688]= 2117461370;
assign addr[1689]= 2045196100;
assign addr[1690]= 1931484818;
assign addr[1691]= 1778631892;
assign addr[1692]= 1589734894;
assign addr[1693]= 1368621831;
assign addr[1694]= 1119773573;
assign addr[1695]= 848233042;
assign addr[1696]= 559503022;
assign addr[1697]= 259434643;
assign addr[1698]= -45891193;
assign addr[1699]= -350287041;
assign addr[1700]= -647584304;
assign addr[1701]= -931758235;
assign addr[1702]= -1197050035;
assign addr[1703]= -1438083551;
assign addr[1704]= -1649974225;
assign addr[1705]= -1828428082;
assign addr[1706]= -1969828744;
assign addr[1707]= -2071310720;
assign addr[1708]= -2130817471;
assign addr[1709]= -2147143090;
assign addr[1710]= -2119956737;
assign addr[1711]= -2049809346;
assign addr[1712]= -1938122457;
assign addr[1713]= -1787159411;
assign addr[1714]= -1599979481;
assign addr[1715]= -1380375881;
assign addr[1716]= -1132798888;
assign addr[1717]= -862265664;
assign addr[1718]= -574258580;
assign addr[1719]= -274614114;
assign addr[1720]= 30595422;
assign addr[1721]= 335184940;
assign addr[1722]= 632981917;
assign addr[1723]= 917951481;
assign addr[1724]= 1184318708;
assign addr[1725]= 1426685652;
assign addr[1726]= 1640140734;
assign addr[1727]= 1820358275;
assign addr[1728]= 1963686155;
assign addr[1729]= 2067219829;
assign addr[1730]= 2128861181;
assign addr[1731]= 2147361045;
assign addr[1732]= 2122344521;
assign addr[1733]= 2054318569;
assign addr[1734]= 1944661739;
assign addr[1735]= 1795596234;
assign addr[1736]= 1610142873;
assign addr[1737]= 1392059879;
assign addr[1738]= 1145766716;
assign addr[1739]= 876254528;
assign addr[1740]= 588984994;
assign addr[1741]= 289779648;
assign addr[1742]= -15298099;
assign addr[1743]= -320065829;
assign addr[1744]= -618347408;
assign addr[1745]= -904098143;
assign addr[1746]= -1171527280;
assign addr[1747]= -1415215352;
assign addr[1748]= -1630224009;
assign addr[1749]= -1812196087;
assign addr[1750]= -1957443913;
assign addr[1751]= -2063024031;
assign addr[1752]= -2126796855;
assign addr[1753]= -2147470025;
assign addr[1754]= -2124624598;
assign addr[1755]= -2058723538;
assign addr[1756]= -1951102334;
assign addr[1757]= -1803941934;
assign addr[1758]= -1620224553;
assign addr[1759]= -1403673233;
assign addr[1760]= -1158676398;
assign addr[1761]= -890198924;
assign addr[1762]= -603681519;
assign addr[1763]= -304930476;
assign addr[1764]= 0;
assign addr[1765]= 304930476;
assign addr[1766]= 603681519;
assign addr[1767]= 890198924;
assign addr[1768]= 1158676398;
assign addr[1769]= 1403673233;
assign addr[1770]= 1620224553;
assign addr[1771]= 1803941934;
assign addr[1772]= 1951102334;
assign addr[1773]= 2058723538;
assign addr[1774]= 2124624598;
assign addr[1775]= 2147470025;
assign addr[1776]= 2126796855;
assign addr[1777]= 2063024031;
assign addr[1778]= 1957443913;
assign addr[1779]= 1812196087;
assign addr[1780]= 1630224009;
assign addr[1781]= 1415215352;
assign addr[1782]= 1171527280;
assign addr[1783]= 904098143;
assign addr[1784]= 618347408;
assign addr[1785]= 320065829;
assign addr[1786]= 15298099;
assign addr[1787]= -289779648;
assign addr[1788]= -588984994;
assign addr[1789]= -876254528;
assign addr[1790]= -1145766716;
assign addr[1791]= -1392059879;
assign addr[1792]= -1610142873;
assign addr[1793]= -1795596234;
assign addr[1794]= -1944661739;
assign addr[1795]= -2054318569;
assign addr[1796]= -2122344521;
assign addr[1797]= -2147361045;
assign addr[1798]= -2128861181;
assign addr[1799]= -2067219829;
assign addr[1800]= -1963686155;
assign addr[1801]= -1820358275;
assign addr[1802]= -1640140734;
assign addr[1803]= -1426685652;
assign addr[1804]= -1184318708;
assign addr[1805]= -917951481;
assign addr[1806]= -632981917;
assign addr[1807]= -335184940;
assign addr[1808]= -30595422;
assign addr[1809]= 274614114;
assign addr[1810]= 574258580;
assign addr[1811]= 862265664;
assign addr[1812]= 1132798888;
assign addr[1813]= 1380375881;
assign addr[1814]= 1599979481;
assign addr[1815]= 1787159411;
assign addr[1816]= 1938122457;
assign addr[1817]= 2049809346;
assign addr[1818]= 2119956737;
assign addr[1819]= 2147143090;
assign addr[1820]= 2130817471;
assign addr[1821]= 2071310720;
assign addr[1822]= 1969828744;
assign addr[1823]= 1828428082;
assign addr[1824]= 1649974225;
assign addr[1825]= 1438083551;
assign addr[1826]= 1197050035;
assign addr[1827]= 931758235;
assign addr[1828]= 647584304;
assign addr[1829]= 350287041;
assign addr[1830]= 45891193;
assign addr[1831]= -259434643;
assign addr[1832]= -559503022;
assign addr[1833]= -848233042;
assign addr[1834]= -1119773573;
assign addr[1835]= -1368621831;
assign addr[1836]= -1589734894;
assign addr[1837]= -1778631892;
assign addr[1838]= -1931484818;
assign addr[1839]= -2045196100;
assign addr[1840]= -2117461370;
assign addr[1841]= -2146816171;
assign addr[1842]= -2132665626;
assign addr[1843]= -2075296495;
assign addr[1844]= -1975871368;
assign addr[1845]= -1836405100;
assign addr[1846]= -1659723983;
assign addr[1847]= -1449408469;
assign addr[1848]= -1209720613;
assign addr[1849]= -945517704;
assign addr[1850]= -662153826;
assign addr[1851]= -365371365;
assign addr[1852]= -61184634;
assign addr[1853]= 244242007;
assign addr[1854]= 544719071;
assign addr[1855]= 834157373;
assign addr[1856]= 1106691431;
assign addr[1857]= 1356798326;
assign addr[1858]= 1579409630;
assign addr[1859]= 1770014111;
assign addr[1860]= 1924749160;
assign addr[1861]= 2040479063;
assign addr[1862]= 2114858546;
assign addr[1863]= 2146380306;
assign addr[1864]= 2134405552;
assign addr[1865]= 2079176953;
assign addr[1866]= 1981813720;
assign addr[1867]= 1844288924;
assign addr[1868]= 1669389513;
assign addr[1869]= 1460659832;
assign addr[1870]= 1222329801;
assign addr[1871]= 959229189;
assign addr[1872]= 676689746;
assign addr[1873]= 380437148;
assign addr[1874]= 76474970;
assign addr[1875]= -229036977;
assign addr[1876]= -529907477;
assign addr[1877]= -820039373;
assign addr[1878]= -1093553126;
assign addr[1879]= -1344905966;
assign addr[1880]= -1569004214;
assign addr[1881]= -1761306505;
assign addr[1882]= -1917915825;
assign addr[1883]= -2035658475;
assign addr[1884]= -2112148396;
assign addr[1885]= -2145835515;
assign addr[1886]= -2136037160;
assign addr[1887]= -2082951896;
assign addr[1888]= -1987655498;
assign addr[1889]= -1852079154;
assign addr[1890]= -1678970324;
assign addr[1891]= -1471837070;
assign addr[1892]= -1234876957;
assign addr[1893]= -972891995;
assign addr[1894]= -691191324;
assign addr[1895]= -395483624;
assign addr[1896]= -91761426;
assign addr[1897]= 213820322;
assign addr[1898]= 515068990;
assign addr[1899]= 805879757;
assign addr[1900]= 1080359326;
assign addr[1901]= 1332945355;
assign addr[1902]= 1558519173;
assign addr[1903]= 1752509516;
assign addr[1904]= 1910985158;
assign addr[1905]= 2030734582;
assign addr[1906]= 2109331059;
assign addr[1907]= 2145181827;
assign addr[1908]= 2137560369;
assign addr[1909]= 2086621133;
assign addr[1910]= 1993396407;
assign addr[1911]= 1859775393;
assign addr[1912]= 1688465931;
assign addr[1913]= 1482939614;
assign addr[1914]= 1247361445;
assign addr[1915]= 986505429;
assign addr[1916]= 705657826;
assign addr[1917]= 410510029;
assign addr[1918]= 107043224;
assign addr[1919]= -198592817;
assign addr[1920]= -500204365;
assign addr[1921]= -791679244;
assign addr[1922]= -1067110699;
assign addr[1923]= -1320917099;
assign addr[1924]= -1547955041;
assign addr[1925]= -1743623590;
assign addr[1926]= -1903957513;
assign addr[1927]= -2025707632;
assign addr[1928]= -2106406677;
assign addr[1929]= -2144419275;
assign addr[1930]= -2138975100;
assign addr[1931]= -2090184478;
assign addr[1932]= -1999036154;
assign addr[1933]= -1867377253;
assign addr[1934]= -1697875851;
assign addr[1935]= -1493966902;
assign addr[1936]= -1259782632;
assign addr[1937]= -1000068799;
assign addr[1938]= -720088517;
assign addr[1939]= -425515602;
assign addr[1940]= -122319591;
assign addr[1941]= 183355234;
assign addr[1942]= 485314355;
assign addr[1943]= 777438554;
assign addr[1944]= 1053807919;
assign addr[1945]= 1308821808;
assign addr[1946]= 1537312353;
assign addr[1947]= 1734649179;
assign addr[1948]= 1896833245;
assign addr[1949]= 2020577882;
assign addr[1950]= 2103375398;
assign addr[1951]= 2143547897;
assign addr[1952]= 2140281282;
assign addr[1953]= 2093641749;
assign addr[1954]= 2004574453;
assign addr[1955]= 1874884346;
assign addr[1956]= 1707199606;
assign addr[1957]= 1504918373;
assign addr[1958]= 1272139887;
assign addr[1959]= 1013581418;
assign addr[1960]= 734482665;
assign addr[1961]= 440499581;
assign addr[1962]= 137589750;
assign addr[1963]= -168108346;
assign addr[1964]= -470399716;
assign addr[1965]= -763158411;
assign addr[1966]= -1040451659;
assign addr[1967]= -1296660098;
assign addr[1968]= -1526591649;
assign addr[1969]= -1725586737;
assign addr[1970]= -1889612716;
assign addr[1971]= -2015345591;
assign addr[1972]= -2100237377;
assign addr[1973]= -2142567738;
assign addr[1974]= -2141478848;
assign addr[1975]= -2096992772;
assign addr[1976]= -2010011024;
assign addr[1977]= -1882296293;
assign addr[1978]= -1716436725;
assign addr[1979]= -1515793473;
assign addr[1980]= -1284432584;
assign addr[1981]= -1027042599;
assign addr[1982]= -748839539;
assign addr[1983]= -455461206;
assign addr[1984]= -152852926;
assign addr[1985]= 152852926;
assign addr[1986]= 455461206;
assign addr[1987]= 748839539;
assign addr[1988]= 1027042599;
assign addr[1989]= 1284432584;
assign addr[1990]= 1515793473;
assign addr[1991]= 1716436725;
assign addr[1992]= 1882296293;
assign addr[1993]= 2010011024;
assign addr[1994]= 2096992772;
assign addr[1995]= 2141478848;
assign addr[1996]= 2142567738;
assign addr[1997]= 2100237377;
assign addr[1998]= 2015345591;
assign addr[1999]= 1889612716;
assign addr[2000]= 1725586737;
assign addr[2001]= 1526591649;
assign addr[2002]= 1296660098;
assign addr[2003]= 1040451659;
assign addr[2004]= 763158411;
assign addr[2005]= 470399716;
assign addr[2006]= 168108346;
assign addr[2007]= -137589750;
assign addr[2008]= -440499581;
assign addr[2009]= -734482665;
assign addr[2010]= -1013581418;
assign addr[2011]= -1272139887;
assign addr[2012]= -1504918373;
assign addr[2013]= -1707199606;
assign addr[2014]= -1874884346;
assign addr[2015]= -2004574453;
assign addr[2016]= -2093641749;
assign addr[2017]= -2140281282;
assign addr[2018]= -2143547897;
assign addr[2019]= -2103375398;
assign addr[2020]= -2020577882;
assign addr[2021]= -1896833245;
assign addr[2022]= -1734649179;
assign addr[2023]= -1537312353;
assign addr[2024]= -1308821808;
assign addr[2025]= -1053807919;
assign addr[2026]= -777438554;
assign addr[2027]= -485314355;
assign addr[2028]= -183355234;
assign addr[2029]= 122319591;
assign addr[2030]= 425515602;
assign addr[2031]= 720088517;
assign addr[2032]= 1000068799;
assign addr[2033]= 1259782632;
assign addr[2034]= 1493966902;
assign addr[2035]= 1697875851;
assign addr[2036]= 1867377253;
assign addr[2037]= 1999036154;
assign addr[2038]= 2090184478;
assign addr[2039]= 2138975100;
assign addr[2040]= 2144419275;
assign addr[2041]= 2106406677;
assign addr[2042]= 2025707632;
assign addr[2043]= 1903957513;
assign addr[2044]= 1743623590;
assign addr[2045]= 1547955041;
assign addr[2046]= 1320917099;
assign addr[2047]= 1067110699;
assign addr[2048]= 791679244;
assign addr[2049]= 500204365;
assign addr[2050]= 198592817;
assign addr[2051]= -107043224;
assign addr[2052]= -410510029;
assign addr[2053]= -705657826;
assign addr[2054]= -986505429;
assign addr[2055]= -1247361445;
assign addr[2056]= -1482939614;
assign addr[2057]= -1688465931;
assign addr[2058]= -1859775393;
assign addr[2059]= -1993396407;
assign addr[2060]= -2086621133;
assign addr[2061]= -2137560369;
assign addr[2062]= -2145181827;
assign addr[2063]= -2109331059;
assign addr[2064]= -2030734582;
assign addr[2065]= -1910985158;
assign addr[2066]= -1752509516;
assign addr[2067]= -1558519173;
assign addr[2068]= -1332945355;
assign addr[2069]= -1080359326;
assign addr[2070]= -805879757;
assign addr[2071]= -515068990;
assign addr[2072]= -213820322;
assign addr[2073]= 91761426;
assign addr[2074]= 395483624;
assign addr[2075]= 691191324;
assign addr[2076]= 972891995;
assign addr[2077]= 1234876957;
assign addr[2078]= 1471837070;
assign addr[2079]= 1678970324;
assign addr[2080]= 1852079154;
assign addr[2081]= 1987655498;
assign addr[2082]= 2082951896;
assign addr[2083]= 2136037160;
assign addr[2084]= 2145835515;
assign addr[2085]= 2112148396;
assign addr[2086]= 2035658475;
assign addr[2087]= 1917915825;
assign addr[2088]= 1761306505;
assign addr[2089]= 1569004214;
assign addr[2090]= 1344905966;
assign addr[2091]= 1093553126;
assign addr[2092]= 820039373;
assign addr[2093]= 529907477;
assign addr[2094]= 229036977;
assign addr[2095]= -76474970;
assign addr[2096]= -380437148;
assign addr[2097]= -676689746;
assign addr[2098]= -959229189;
assign addr[2099]= -1222329801;
assign addr[2100]= -1460659832;
assign addr[2101]= -1669389513;
assign addr[2102]= -1844288924;
assign addr[2103]= -1981813720;
assign addr[2104]= -2079176953;
assign addr[2105]= -2134405552;
assign addr[2106]= -2146380306;
assign addr[2107]= -2114858546;
assign addr[2108]= -2040479063;
assign addr[2109]= -1924749160;
assign addr[2110]= -1770014111;
assign addr[2111]= -1579409630;
assign addr[2112]= -1356798326;
assign addr[2113]= -1106691431;
assign addr[2114]= -834157373;
assign addr[2115]= -544719071;
assign addr[2116]= -244242007;
assign addr[2117]= 61184634;
assign addr[2118]= 365371365;
assign addr[2119]= 662153826;
assign addr[2120]= 945517704;
assign addr[2121]= 1209720613;
assign addr[2122]= 1449408469;
assign addr[2123]= 1659723983;
assign addr[2124]= 1836405100;
assign addr[2125]= 1975871368;
assign addr[2126]= 2075296495;
assign addr[2127]= 2132665626;
assign addr[2128]= 2146816171;
assign addr[2129]= 2117461370;
assign addr[2130]= 2045196100;
assign addr[2131]= 1931484818;
assign addr[2132]= 1778631892;
assign addr[2133]= 1589734894;
assign addr[2134]= 1368621831;
assign addr[2135]= 1119773573;
assign addr[2136]= 848233042;
assign addr[2137]= 559503022;
assign addr[2138]= 259434643;
assign addr[2139]= -45891193;
assign addr[2140]= -350287041;
assign addr[2141]= -647584304;
assign addr[2142]= -931758235;
assign addr[2143]= -1197050035;
assign addr[2144]= -1438083551;
assign addr[2145]= -1649974225;
assign addr[2146]= -1828428082;
assign addr[2147]= -1969828744;
assign addr[2148]= -2071310720;
assign addr[2149]= -2130817471;
assign addr[2150]= -2147143090;
assign addr[2151]= -2119956737;
assign addr[2152]= -2049809346;
assign addr[2153]= -1938122457;
assign addr[2154]= -1787159411;
assign addr[2155]= -1599979481;
assign addr[2156]= -1380375881;
assign addr[2157]= -1132798888;
assign addr[2158]= -862265664;
assign addr[2159]= -574258580;
assign addr[2160]= -274614114;
assign addr[2161]= 30595422;
assign addr[2162]= 335184940;
assign addr[2163]= 632981917;
assign addr[2164]= 917951481;
assign addr[2165]= 1184318708;
assign addr[2166]= 1426685652;
assign addr[2167]= 1640140734;
assign addr[2168]= 1820358275;
assign addr[2169]= 1963686155;
assign addr[2170]= 2067219829;
assign addr[2171]= 2128861181;
assign addr[2172]= 2147361045;
assign addr[2173]= 2122344521;
assign addr[2174]= 2054318569;
assign addr[2175]= 1944661739;
assign addr[2176]= 1795596234;
assign addr[2177]= 1610142873;
assign addr[2178]= 1392059879;
assign addr[2179]= 1145766716;
assign addr[2180]= 876254528;
assign addr[2181]= 588984994;
assign addr[2182]= 289779648;
assign addr[2183]= -15298099;
assign addr[2184]= -320065829;
assign addr[2185]= -618347408;
assign addr[2186]= -904098143;
assign addr[2187]= -1171527280;
assign addr[2188]= -1415215352;
assign addr[2189]= -1630224009;
assign addr[2190]= -1812196087;
assign addr[2191]= -1957443913;
assign addr[2192]= -2063024031;
assign addr[2193]= -2126796855;
assign addr[2194]= -2147470025;
assign addr[2195]= -2124624598;
assign addr[2196]= -2058723538;
assign addr[2197]= -1951102334;
assign addr[2198]= -1803941934;
assign addr[2199]= -1620224553;
assign addr[2200]= -1403673233;
assign addr[2201]= -1158676398;
assign addr[2202]= -890198924;
assign addr[2203]= -603681519;
assign addr[2204]= -304930476;
assign addr[2205]= 0;
assign addr[2206]= 304930476;
assign addr[2207]= 603681519;
assign addr[2208]= 890198924;
assign addr[2209]= 1158676398;
assign addr[2210]= 1403673233;
assign addr[2211]= 1620224553;
assign addr[2212]= 1803941934;
assign addr[2213]= 1951102334;
assign addr[2214]= 2058723538;
assign addr[2215]= 2124624598;
assign addr[2216]= 2147470025;
assign addr[2217]= 2126796855;
assign addr[2218]= 2063024031;
assign addr[2219]= 1957443913;
assign addr[2220]= 1812196087;
assign addr[2221]= 1630224009;
assign addr[2222]= 1415215352;
assign addr[2223]= 1171527280;
assign addr[2224]= 904098143;
assign addr[2225]= 618347408;
assign addr[2226]= 320065829;
assign addr[2227]= 15298099;
assign addr[2228]= -289779648;
assign addr[2229]= -588984994;
assign addr[2230]= -876254528;
assign addr[2231]= -1145766716;
assign addr[2232]= -1392059879;
assign addr[2233]= -1610142873;
assign addr[2234]= -1795596234;
assign addr[2235]= -1944661739;
assign addr[2236]= -2054318569;
assign addr[2237]= -2122344521;
assign addr[2238]= -2147361045;
assign addr[2239]= -2128861181;
assign addr[2240]= -2067219829;
assign addr[2241]= -1963686155;
assign addr[2242]= -1820358275;
assign addr[2243]= -1640140734;
assign addr[2244]= -1426685652;
assign addr[2245]= -1184318708;
assign addr[2246]= -917951481;
assign addr[2247]= -632981917;
assign addr[2248]= -335184940;
assign addr[2249]= -30595422;
assign addr[2250]= 274614114;
assign addr[2251]= 574258580;
assign addr[2252]= 862265664;
assign addr[2253]= 1132798888;
assign addr[2254]= 1380375881;
assign addr[2255]= 1599979481;
assign addr[2256]= 1787159411;
assign addr[2257]= 1938122457;
assign addr[2258]= 2049809346;
assign addr[2259]= 2119956737;
assign addr[2260]= 2147143090;
assign addr[2261]= 2130817471;
assign addr[2262]= 2071310720;
assign addr[2263]= 1969828744;
assign addr[2264]= 1828428082;
assign addr[2265]= 1649974225;
assign addr[2266]= 1438083551;
assign addr[2267]= 1197050035;
assign addr[2268]= 931758235;
assign addr[2269]= 647584304;
assign addr[2270]= 350287041;
assign addr[2271]= 45891193;
assign addr[2272]= -259434643;
assign addr[2273]= -559503022;
assign addr[2274]= -848233042;
assign addr[2275]= -1119773573;
assign addr[2276]= -1368621831;
assign addr[2277]= -1589734894;
assign addr[2278]= -1778631892;
assign addr[2279]= -1931484818;
assign addr[2280]= -2045196100;
assign addr[2281]= -2117461370;
assign addr[2282]= -2146816171;
assign addr[2283]= -2132665626;
assign addr[2284]= -2075296495;
assign addr[2285]= -1975871368;
assign addr[2286]= -1836405100;
assign addr[2287]= -1659723983;
assign addr[2288]= -1449408469;
assign addr[2289]= -1209720613;
assign addr[2290]= -945517704;
assign addr[2291]= -662153826;
assign addr[2292]= -365371365;
assign addr[2293]= -61184634;
assign addr[2294]= 244242007;
assign addr[2295]= 544719071;
assign addr[2296]= 834157373;
assign addr[2297]= 1106691431;
assign addr[2298]= 1356798326;
assign addr[2299]= 1579409630;
assign addr[2300]= 1770014111;
assign addr[2301]= 1924749160;
assign addr[2302]= 2040479063;
assign addr[2303]= 2114858546;
assign addr[2304]= 2146380306;
assign addr[2305]= 2134405552;
assign addr[2306]= 2079176953;
assign addr[2307]= 1981813720;
assign addr[2308]= 1844288924;
assign addr[2309]= 1669389513;
assign addr[2310]= 1460659832;
assign addr[2311]= 1222329801;
assign addr[2312]= 959229189;
assign addr[2313]= 676689746;
assign addr[2314]= 380437148;
assign addr[2315]= 76474970;
assign addr[2316]= -229036977;
assign addr[2317]= -529907477;
assign addr[2318]= -820039373;
assign addr[2319]= -1093553126;
assign addr[2320]= -1344905966;
assign addr[2321]= -1569004214;
assign addr[2322]= -1761306505;
assign addr[2323]= -1917915825;
assign addr[2324]= -2035658475;
assign addr[2325]= -2112148396;
assign addr[2326]= -2145835515;
assign addr[2327]= -2136037160;
assign addr[2328]= -2082951896;
assign addr[2329]= -1987655498;
assign addr[2330]= -1852079154;
assign addr[2331]= -1678970324;
assign addr[2332]= -1471837070;
assign addr[2333]= -1234876957;
assign addr[2334]= -972891995;
assign addr[2335]= -691191324;
assign addr[2336]= -395483624;
assign addr[2337]= -91761426;
assign addr[2338]= 213820322;
assign addr[2339]= 515068990;
assign addr[2340]= 805879757;
assign addr[2341]= 1080359326;
assign addr[2342]= 1332945355;
assign addr[2343]= 1558519173;
assign addr[2344]= 1752509516;
assign addr[2345]= 1910985158;
assign addr[2346]= 2030734582;
assign addr[2347]= 2109331059;
assign addr[2348]= 2145181827;
assign addr[2349]= 2137560369;
assign addr[2350]= 2086621133;
assign addr[2351]= 1993396407;
assign addr[2352]= 1859775393;
assign addr[2353]= 1688465931;
assign addr[2354]= 1482939614;
assign addr[2355]= 1247361445;
assign addr[2356]= 986505429;
assign addr[2357]= 705657826;
assign addr[2358]= 410510029;
assign addr[2359]= 107043224;
assign addr[2360]= -198592817;
assign addr[2361]= -500204365;
assign addr[2362]= -791679244;
assign addr[2363]= -1067110699;
assign addr[2364]= -1320917099;
assign addr[2365]= -1547955041;
assign addr[2366]= -1743623590;
assign addr[2367]= -1903957513;
assign addr[2368]= -2025707632;
assign addr[2369]= -2106406677;
assign addr[2370]= -2144419275;
assign addr[2371]= -2138975100;
assign addr[2372]= -2090184478;
assign addr[2373]= -1999036154;
assign addr[2374]= -1867377253;
assign addr[2375]= -1697875851;
assign addr[2376]= -1493966902;
assign addr[2377]= -1259782632;
assign addr[2378]= -1000068799;
assign addr[2379]= -720088517;
assign addr[2380]= -425515602;
assign addr[2381]= -122319591;
assign addr[2382]= 183355234;
assign addr[2383]= 485314355;
assign addr[2384]= 777438554;
assign addr[2385]= 1053807919;
assign addr[2386]= 1308821808;
assign addr[2387]= 1537312353;
assign addr[2388]= 1734649179;
assign addr[2389]= 1896833245;
assign addr[2390]= 2020577882;
assign addr[2391]= 2103375398;
assign addr[2392]= 2143547897;
assign addr[2393]= 2140281282;
assign addr[2394]= 2093641749;
assign addr[2395]= 2004574453;
assign addr[2396]= 1874884346;
assign addr[2397]= 1707199606;
assign addr[2398]= 1504918373;
assign addr[2399]= 1272139887;
assign addr[2400]= 1013581418;
assign addr[2401]= 734482665;
assign addr[2402]= 440499581;
assign addr[2403]= 137589750;
assign addr[2404]= -168108346;
assign addr[2405]= -470399716;
assign addr[2406]= -763158411;
assign addr[2407]= -1040451659;
assign addr[2408]= -1296660098;
assign addr[2409]= -1526591649;
assign addr[2410]= -1725586737;
assign addr[2411]= -1889612716;
assign addr[2412]= -2015345591;
assign addr[2413]= -2100237377;
assign addr[2414]= -2142567738;
assign addr[2415]= -2141478848;
assign addr[2416]= -2096992772;
assign addr[2417]= -2010011024;
assign addr[2418]= -1882296293;
assign addr[2419]= -1716436725;
assign addr[2420]= -1515793473;
assign addr[2421]= -1284432584;
assign addr[2422]= -1027042599;
assign addr[2423]= -748839539;
assign addr[2424]= -455461206;
assign addr[2425]= -152852926;
assign addr[2426]= 152852926;
assign addr[2427]= 455461206;
assign addr[2428]= 748839539;
assign addr[2429]= 1027042599;
assign addr[2430]= 1284432584;
assign addr[2431]= 1515793473;
assign addr[2432]= 1716436725;
assign addr[2433]= 1882296293;
assign addr[2434]= 2010011024;
assign addr[2435]= 2096992772;
assign addr[2436]= 2141478848;
assign addr[2437]= 2142567738;
assign addr[2438]= 2100237377;
assign addr[2439]= 2015345591;
assign addr[2440]= 1889612716;
assign addr[2441]= 1725586737;
assign addr[2442]= 1526591649;
assign addr[2443]= 1296660098;
assign addr[2444]= 1040451659;
assign addr[2445]= 763158411;
assign addr[2446]= 470399716;
assign addr[2447]= 168108346;
assign addr[2448]= -137589750;
assign addr[2449]= -440499581;
assign addr[2450]= -734482665;
assign addr[2451]= -1013581418;
assign addr[2452]= -1272139887;
assign addr[2453]= -1504918373;
assign addr[2454]= -1707199606;
assign addr[2455]= -1874884346;
assign addr[2456]= -2004574453;
assign addr[2457]= -2093641749;
assign addr[2458]= -2140281282;
assign addr[2459]= -2143547897;
assign addr[2460]= -2103375398;
assign addr[2461]= -2020577882;
assign addr[2462]= -1896833245;
assign addr[2463]= -1734649179;
assign addr[2464]= -1537312353;
assign addr[2465]= -1308821808;
assign addr[2466]= -1053807919;
assign addr[2467]= -777438554;
assign addr[2468]= -485314355;
assign addr[2469]= -183355234;
assign addr[2470]= 122319591;
assign addr[2471]= 425515602;
assign addr[2472]= 720088517;
assign addr[2473]= 1000068799;
assign addr[2474]= 1259782632;
assign addr[2475]= 1493966902;
assign addr[2476]= 1697875851;
assign addr[2477]= 1867377253;
assign addr[2478]= 1999036154;
assign addr[2479]= 2090184478;
assign addr[2480]= 2138975100;
assign addr[2481]= 2144419275;
assign addr[2482]= 2106406677;
assign addr[2483]= 2025707632;
assign addr[2484]= 1903957513;
assign addr[2485]= 1743623590;
assign addr[2486]= 1547955041;
assign addr[2487]= 1320917099;
assign addr[2488]= 1067110699;
assign addr[2489]= 791679244;
assign addr[2490]= 500204365;
assign addr[2491]= 198592817;
assign addr[2492]= -107043224;
assign addr[2493]= -410510029;
assign addr[2494]= -705657826;
assign addr[2495]= -986505429;
assign addr[2496]= -1247361445;
assign addr[2497]= -1482939614;
assign addr[2498]= -1688465931;
assign addr[2499]= -1859775393;
assign addr[2500]= -1993396407;
assign addr[2501]= -2086621133;
assign addr[2502]= -2137560369;
assign addr[2503]= -2145181827;
assign addr[2504]= -2109331059;
assign addr[2505]= -2030734582;
assign addr[2506]= -1910985158;
assign addr[2507]= -1752509516;
assign addr[2508]= -1558519173;
assign addr[2509]= -1332945355;
assign addr[2510]= -1080359326;
assign addr[2511]= -805879757;
assign addr[2512]= -515068990;
assign addr[2513]= -213820322;
assign addr[2514]= 91761426;
assign addr[2515]= 395483624;
assign addr[2516]= 691191324;
assign addr[2517]= 972891995;
assign addr[2518]= 1234876957;
assign addr[2519]= 1471837070;
assign addr[2520]= 1678970324;
assign addr[2521]= 1852079154;
assign addr[2522]= 1987655498;
assign addr[2523]= 2082951896;
assign addr[2524]= 2136037160;
assign addr[2525]= 2145835515;
assign addr[2526]= 2112148396;
assign addr[2527]= 2035658475;
assign addr[2528]= 1917915825;
assign addr[2529]= 1761306505;
assign addr[2530]= 1569004214;
assign addr[2531]= 1344905966;
assign addr[2532]= 1093553126;
assign addr[2533]= 820039373;
assign addr[2534]= 529907477;
assign addr[2535]= 229036977;
assign addr[2536]= -76474970;
assign addr[2537]= -380437148;
assign addr[2538]= -676689746;
assign addr[2539]= -959229189;
assign addr[2540]= -1222329801;
assign addr[2541]= -1460659832;
assign addr[2542]= -1669389513;
assign addr[2543]= -1844288924;
assign addr[2544]= -1981813720;
assign addr[2545]= -2079176953;
assign addr[2546]= -2134405552;
assign addr[2547]= -2146380306;
assign addr[2548]= -2114858546;
assign addr[2549]= -2040479063;
assign addr[2550]= -1924749160;
assign addr[2551]= -1770014111;
assign addr[2552]= -1579409630;
assign addr[2553]= -1356798326;
assign addr[2554]= -1106691431;
assign addr[2555]= -834157373;
assign addr[2556]= -544719071;
assign addr[2557]= -244242007;
assign addr[2558]= 61184634;
assign addr[2559]= 365371365;
assign addr[2560]= 662153826;
assign addr[2561]= 945517704;
assign addr[2562]= 1209720613;
assign addr[2563]= 1449408469;
assign addr[2564]= 1659723983;
assign addr[2565]= 1836405100;
assign addr[2566]= 1975871368;
assign addr[2567]= 2075296495;
assign addr[2568]= 2132665626;
assign addr[2569]= 2146816171;
assign addr[2570]= 2117461370;
assign addr[2571]= 2045196100;
assign addr[2572]= 1931484818;
assign addr[2573]= 1778631892;
assign addr[2574]= 1589734894;
assign addr[2575]= 1368621831;
assign addr[2576]= 1119773573;
assign addr[2577]= 848233042;
assign addr[2578]= 559503022;
assign addr[2579]= 259434643;
assign addr[2580]= -45891193;
assign addr[2581]= -350287041;
assign addr[2582]= -647584304;
assign addr[2583]= -931758235;
assign addr[2584]= -1197050035;
assign addr[2585]= -1438083551;
assign addr[2586]= -1649974225;
assign addr[2587]= -1828428082;
assign addr[2588]= -1969828744;
assign addr[2589]= -2071310720;
assign addr[2590]= -2130817471;
assign addr[2591]= -2147143090;
assign addr[2592]= -2119956737;
assign addr[2593]= -2049809346;
assign addr[2594]= -1938122457;
assign addr[2595]= -1787159411;
assign addr[2596]= -1599979481;
assign addr[2597]= -1380375881;
assign addr[2598]= -1132798888;
assign addr[2599]= -862265664;
assign addr[2600]= -574258580;
assign addr[2601]= -274614114;
assign addr[2602]= 30595422;
assign addr[2603]= 335184940;
assign addr[2604]= 632981917;
assign addr[2605]= 917951481;
assign addr[2606]= 1184318708;
assign addr[2607]= 1426685652;
assign addr[2608]= 1640140734;
assign addr[2609]= 1820358275;
assign addr[2610]= 1963686155;
assign addr[2611]= 2067219829;
assign addr[2612]= 2128861181;
assign addr[2613]= 2147361045;
assign addr[2614]= 2122344521;
assign addr[2615]= 2054318569;
assign addr[2616]= 1944661739;
assign addr[2617]= 1795596234;
assign addr[2618]= 1610142873;
assign addr[2619]= 1392059879;
assign addr[2620]= 1145766716;
assign addr[2621]= 876254528;
assign addr[2622]= 588984994;
assign addr[2623]= 289779648;
assign addr[2624]= -15298099;
assign addr[2625]= -320065829;
assign addr[2626]= -618347408;
assign addr[2627]= -904098143;
assign addr[2628]= -1171527280;
assign addr[2629]= -1415215352;
assign addr[2630]= -1630224009;
assign addr[2631]= -1812196087;
assign addr[2632]= -1957443913;
assign addr[2633]= -2063024031;
assign addr[2634]= -2126796855;
assign addr[2635]= -2147470025;
assign addr[2636]= -2124624598;
assign addr[2637]= -2058723538;
assign addr[2638]= -1951102334;
assign addr[2639]= -1803941934;
assign addr[2640]= -1620224553;
assign addr[2641]= -1403673233;
assign addr[2642]= -1158676398;
assign addr[2643]= -890198924;
assign addr[2644]= -603681519;
assign addr[2645]= -304930476;
assign addr[2646]= 0;
assign addr[2647]= 304930476;
assign addr[2648]= 603681519;
assign addr[2649]= 890198924;
assign addr[2650]= 1158676398;
assign addr[2651]= 1403673233;
assign addr[2652]= 1620224553;
assign addr[2653]= 1803941934;
assign addr[2654]= 1951102334;
assign addr[2655]= 2058723538;
assign addr[2656]= 2124624598;
assign addr[2657]= 2147470025;
assign addr[2658]= 2126796855;
assign addr[2659]= 2063024031;
assign addr[2660]= 1957443913;
assign addr[2661]= 1812196087;
assign addr[2662]= 1630224009;
assign addr[2663]= 1415215352;
assign addr[2664]= 1171527280;
assign addr[2665]= 904098143;
assign addr[2666]= 618347408;
assign addr[2667]= 320065829;
assign addr[2668]= 15298099;
assign addr[2669]= -289779648;
assign addr[2670]= -588984994;
assign addr[2671]= -876254528;
assign addr[2672]= -1145766716;
assign addr[2673]= -1392059879;
assign addr[2674]= -1610142873;
assign addr[2675]= -1795596234;
assign addr[2676]= -1944661739;
assign addr[2677]= -2054318569;
assign addr[2678]= -2122344521;
assign addr[2679]= -2147361045;
assign addr[2680]= -2128861181;
assign addr[2681]= -2067219829;
assign addr[2682]= -1963686155;
assign addr[2683]= -1820358275;
assign addr[2684]= -1640140734;
assign addr[2685]= -1426685652;
assign addr[2686]= -1184318708;
assign addr[2687]= -917951481;
assign addr[2688]= -632981917;
assign addr[2689]= -335184940;
assign addr[2690]= -30595422;
assign addr[2691]= 274614114;
assign addr[2692]= 574258580;
assign addr[2693]= 862265664;
assign addr[2694]= 1132798888;
assign addr[2695]= 1380375881;
assign addr[2696]= 1599979481;
assign addr[2697]= 1787159411;
assign addr[2698]= 1938122457;
assign addr[2699]= 2049809346;
assign addr[2700]= 2119956737;
assign addr[2701]= 2147143090;
assign addr[2702]= 2130817471;
assign addr[2703]= 2071310720;
assign addr[2704]= 1969828744;
assign addr[2705]= 1828428082;
assign addr[2706]= 1649974225;
assign addr[2707]= 1438083551;
assign addr[2708]= 1197050035;
assign addr[2709]= 931758235;
assign addr[2710]= 647584304;
assign addr[2711]= 350287041;
assign addr[2712]= 45891193;
assign addr[2713]= -259434643;
assign addr[2714]= -559503022;
assign addr[2715]= -848233042;
assign addr[2716]= -1119773573;
assign addr[2717]= -1368621831;
assign addr[2718]= -1589734894;
assign addr[2719]= -1778631892;
assign addr[2720]= -1931484818;
assign addr[2721]= -2045196100;
assign addr[2722]= -2117461370;
assign addr[2723]= -2146816171;
assign addr[2724]= -2132665626;
assign addr[2725]= -2075296495;
assign addr[2726]= -1975871368;
assign addr[2727]= -1836405100;
assign addr[2728]= -1659723983;
assign addr[2729]= -1449408469;
assign addr[2730]= -1209720613;
assign addr[2731]= -945517704;
assign addr[2732]= -662153826;
assign addr[2733]= -365371365;
assign addr[2734]= -61184634;
assign addr[2735]= 244242007;
assign addr[2736]= 544719071;
assign addr[2737]= 834157373;
assign addr[2738]= 1106691431;
assign addr[2739]= 1356798326;
assign addr[2740]= 1579409630;
assign addr[2741]= 1770014111;
assign addr[2742]= 1924749160;
assign addr[2743]= 2040479063;
assign addr[2744]= 2114858546;
assign addr[2745]= 2146380306;
assign addr[2746]= 2134405552;
assign addr[2747]= 2079176953;
assign addr[2748]= 1981813720;
assign addr[2749]= 1844288924;
assign addr[2750]= 1669389513;
assign addr[2751]= 1460659832;
assign addr[2752]= 1222329801;
assign addr[2753]= 959229189;
assign addr[2754]= 676689746;
assign addr[2755]= 380437148;
assign addr[2756]= 76474970;
assign addr[2757]= -229036977;
assign addr[2758]= -529907477;
assign addr[2759]= -820039373;
assign addr[2760]= -1093553126;
assign addr[2761]= -1344905966;
assign addr[2762]= -1569004214;
assign addr[2763]= -1761306505;
assign addr[2764]= -1917915825;
assign addr[2765]= -2035658475;
assign addr[2766]= -2112148396;
assign addr[2767]= -2145835515;
assign addr[2768]= -2136037160;
assign addr[2769]= -2082951896;
assign addr[2770]= -1987655498;
assign addr[2771]= -1852079154;
assign addr[2772]= -1678970324;
assign addr[2773]= -1471837070;
assign addr[2774]= -1234876957;
assign addr[2775]= -972891995;
assign addr[2776]= -691191324;
assign addr[2777]= -395483624;
assign addr[2778]= -91761426;
assign addr[2779]= 213820322;
assign addr[2780]= 515068990;
assign addr[2781]= 805879757;
assign addr[2782]= 1080359326;
assign addr[2783]= 1332945355;
assign addr[2784]= 1558519173;
assign addr[2785]= 1752509516;
assign addr[2786]= 1910985158;
assign addr[2787]= 2030734582;
assign addr[2788]= 2109331059;
assign addr[2789]= 2145181827;
assign addr[2790]= 2137560369;
assign addr[2791]= 2086621133;
assign addr[2792]= 1993396407;
assign addr[2793]= 1859775393;
assign addr[2794]= 1688465931;
assign addr[2795]= 1482939614;
assign addr[2796]= 1247361445;
assign addr[2797]= 986505429;
assign addr[2798]= 705657826;
assign addr[2799]= 410510029;
assign addr[2800]= 107043224;
assign addr[2801]= -198592817;
assign addr[2802]= -500204365;
assign addr[2803]= -791679244;
assign addr[2804]= -1067110699;
assign addr[2805]= -1320917099;
assign addr[2806]= -1547955041;
assign addr[2807]= -1743623590;
assign addr[2808]= -1903957513;
assign addr[2809]= -2025707632;
assign addr[2810]= -2106406677;
assign addr[2811]= -2144419275;
assign addr[2812]= -2138975100;
assign addr[2813]= -2090184478;
assign addr[2814]= -1999036154;
assign addr[2815]= -1867377253;
assign addr[2816]= -1697875851;
assign addr[2817]= -1493966902;
assign addr[2818]= -1259782632;
assign addr[2819]= -1000068799;
assign addr[2820]= -720088517;
assign addr[2821]= -425515602;
assign addr[2822]= -122319591;
assign addr[2823]= 183355234;
assign addr[2824]= 485314355;
assign addr[2825]= 777438554;
assign addr[2826]= 1053807919;
assign addr[2827]= 1308821808;
assign addr[2828]= 1537312353;
assign addr[2829]= 1734649179;
assign addr[2830]= 1896833245;
assign addr[2831]= 2020577882;
assign addr[2832]= 2103375398;
assign addr[2833]= 2143547897;
assign addr[2834]= 2140281282;
assign addr[2835]= 2093641749;
assign addr[2836]= 2004574453;
assign addr[2837]= 1874884346;
assign addr[2838]= 1707199606;
assign addr[2839]= 1504918373;
assign addr[2840]= 1272139887;
assign addr[2841]= 1013581418;
assign addr[2842]= 734482665;
assign addr[2843]= 440499581;
assign addr[2844]= 137589750;
assign addr[2845]= -168108346;
assign addr[2846]= -470399716;
assign addr[2847]= -763158411;
assign addr[2848]= -1040451659;
assign addr[2849]= -1296660098;
assign addr[2850]= -1526591649;
assign addr[2851]= -1725586737;
assign addr[2852]= -1889612716;
assign addr[2853]= -2015345591;
assign addr[2854]= -2100237377;
assign addr[2855]= -2142567738;
assign addr[2856]= -2141478848;
assign addr[2857]= -2096992772;
assign addr[2858]= -2010011024;
assign addr[2859]= -1882296293;
assign addr[2860]= -1716436725;
assign addr[2861]= -1515793473;
assign addr[2862]= -1284432584;
assign addr[2863]= -1027042599;
assign addr[2864]= -748839539;
assign addr[2865]= -455461206;
assign addr[2866]= -152852926;
assign addr[2867]= 152852926;
assign addr[2868]= 455461206;
assign addr[2869]= 748839539;
assign addr[2870]= 1027042599;
assign addr[2871]= 1284432584;
assign addr[2872]= 1515793473;
assign addr[2873]= 1716436725;
assign addr[2874]= 1882296293;
assign addr[2875]= 2010011024;
assign addr[2876]= 2096992772;
assign addr[2877]= 2141478848;
assign addr[2878]= 2142567738;
assign addr[2879]= 2100237377;
assign addr[2880]= 2015345591;
assign addr[2881]= 1889612716;
assign addr[2882]= 1725586737;
assign addr[2883]= 1526591649;
assign addr[2884]= 1296660098;
assign addr[2885]= 1040451659;
assign addr[2886]= 763158411;
assign addr[2887]= 470399716;
assign addr[2888]= 168108346;
assign addr[2889]= -137589750;
assign addr[2890]= -440499581;
assign addr[2891]= -734482665;
assign addr[2892]= -1013581418;
assign addr[2893]= -1272139887;
assign addr[2894]= -1504918373;
assign addr[2895]= -1707199606;
assign addr[2896]= -1874884346;
assign addr[2897]= -2004574453;
assign addr[2898]= -2093641749;
assign addr[2899]= -2140281282;
assign addr[2900]= -2143547897;
assign addr[2901]= -2103375398;
assign addr[2902]= -2020577882;
assign addr[2903]= -1896833245;
assign addr[2904]= -1734649179;
assign addr[2905]= -1537312353;
assign addr[2906]= -1308821808;
assign addr[2907]= -1053807919;
assign addr[2908]= -777438554;
assign addr[2909]= -485314355;
assign addr[2910]= -183355234;
assign addr[2911]= 122319591;
assign addr[2912]= 425515602;
assign addr[2913]= 720088517;
assign addr[2914]= 1000068799;
assign addr[2915]= 1259782632;
assign addr[2916]= 1493966902;
assign addr[2917]= 1697875851;
assign addr[2918]= 1867377253;
assign addr[2919]= 1999036154;
assign addr[2920]= 2090184478;
assign addr[2921]= 2138975100;
assign addr[2922]= 2144419275;
assign addr[2923]= 2106406677;
assign addr[2924]= 2025707632;
assign addr[2925]= 1903957513;
assign addr[2926]= 1743623590;
assign addr[2927]= 1547955041;
assign addr[2928]= 1320917099;
assign addr[2929]= 1067110699;
assign addr[2930]= 791679244;
assign addr[2931]= 500204365;
assign addr[2932]= 198592817;
assign addr[2933]= -107043224;
assign addr[2934]= -410510029;
assign addr[2935]= -705657826;
assign addr[2936]= -986505429;
assign addr[2937]= -1247361445;
assign addr[2938]= -1482939614;
assign addr[2939]= -1688465931;
assign addr[2940]= -1859775393;
assign addr[2941]= -1993396407;
assign addr[2942]= -2086621133;
assign addr[2943]= -2137560369;
assign addr[2944]= -2145181827;
assign addr[2945]= -2109331059;
assign addr[2946]= -2030734582;
assign addr[2947]= -1910985158;
assign addr[2948]= -1752509516;
assign addr[2949]= -1558519173;
assign addr[2950]= -1332945355;
assign addr[2951]= -1080359326;
assign addr[2952]= -805879757;
assign addr[2953]= -515068990;
assign addr[2954]= -213820322;
assign addr[2955]= 91761426;
assign addr[2956]= 395483624;
assign addr[2957]= 691191324;
assign addr[2958]= 972891995;
assign addr[2959]= 1234876957;
assign addr[2960]= 1471837070;
assign addr[2961]= 1678970324;
assign addr[2962]= 1852079154;
assign addr[2963]= 1987655498;
assign addr[2964]= 2082951896;
assign addr[2965]= 2136037160;
assign addr[2966]= 2145835515;
assign addr[2967]= 2112148396;
assign addr[2968]= 2035658475;
assign addr[2969]= 1917915825;
assign addr[2970]= 1761306505;
assign addr[2971]= 1569004214;
assign addr[2972]= 1344905966;
assign addr[2973]= 1093553126;
assign addr[2974]= 820039373;
assign addr[2975]= 529907477;
assign addr[2976]= 229036977;
assign addr[2977]= -76474970;
assign addr[2978]= -380437148;
assign addr[2979]= -676689746;
assign addr[2980]= -959229189;
assign addr[2981]= -1222329801;
assign addr[2982]= -1460659832;
assign addr[2983]= -1669389513;
assign addr[2984]= -1844288924;
assign addr[2985]= -1981813720;
assign addr[2986]= -2079176953;
assign addr[2987]= -2134405552;
assign addr[2988]= -2146380306;
assign addr[2989]= -2114858546;
assign addr[2990]= -2040479063;
assign addr[2991]= -1924749160;
assign addr[2992]= -1770014111;
assign addr[2993]= -1579409630;
assign addr[2994]= -1356798326;
assign addr[2995]= -1106691431;
assign addr[2996]= -834157373;
assign addr[2997]= -544719071;
assign addr[2998]= -244242007;
assign addr[2999]= 61184634;
assign addr[3000]= 365371365;
assign addr[3001]= 662153826;
assign addr[3002]= 945517704;
assign addr[3003]= 1209720613;
assign addr[3004]= 1449408469;
assign addr[3005]= 1659723983;
assign addr[3006]= 1836405100;
assign addr[3007]= 1975871368;
assign addr[3008]= 2075296495;
assign addr[3009]= 2132665626;
assign addr[3010]= 2146816171;
assign addr[3011]= 2117461370;
assign addr[3012]= 2045196100;
assign addr[3013]= 1931484818;
assign addr[3014]= 1778631892;
assign addr[3015]= 1589734894;
assign addr[3016]= 1368621831;
assign addr[3017]= 1119773573;
assign addr[3018]= 848233042;
assign addr[3019]= 559503022;
assign addr[3020]= 259434643;
assign addr[3021]= -45891193;
assign addr[3022]= -350287041;
assign addr[3023]= -647584304;
assign addr[3024]= -931758235;
assign addr[3025]= -1197050035;
assign addr[3026]= -1438083551;
assign addr[3027]= -1649974225;
assign addr[3028]= -1828428082;
assign addr[3029]= -1969828744;
assign addr[3030]= -2071310720;
assign addr[3031]= -2130817471;
assign addr[3032]= -2147143090;
assign addr[3033]= -2119956737;
assign addr[3034]= -2049809346;
assign addr[3035]= -1938122457;
assign addr[3036]= -1787159411;
assign addr[3037]= -1599979481;
assign addr[3038]= -1380375881;
assign addr[3039]= -1132798888;
assign addr[3040]= -862265664;
assign addr[3041]= -574258580;
assign addr[3042]= -274614114;
assign addr[3043]= 30595422;
assign addr[3044]= 335184940;
assign addr[3045]= 632981917;
assign addr[3046]= 917951481;
assign addr[3047]= 1184318708;
assign addr[3048]= 1426685652;
assign addr[3049]= 1640140734;
assign addr[3050]= 1820358275;
assign addr[3051]= 1963686155;
assign addr[3052]= 2067219829;
assign addr[3053]= 2128861181;
assign addr[3054]= 2147361045;
assign addr[3055]= 2122344521;
assign addr[3056]= 2054318569;
assign addr[3057]= 1944661739;
assign addr[3058]= 1795596234;
assign addr[3059]= 1610142873;
assign addr[3060]= 1392059879;
assign addr[3061]= 1145766716;
assign addr[3062]= 876254528;
assign addr[3063]= 588984994;
assign addr[3064]= 289779648;
assign addr[3065]= -15298099;
assign addr[3066]= -320065829;
assign addr[3067]= -618347408;
assign addr[3068]= -904098143;
assign addr[3069]= -1171527280;
assign addr[3070]= -1415215352;
assign addr[3071]= -1630224009;
assign addr[3072]= -1812196087;
assign addr[3073]= -1957443913;
assign addr[3074]= -2063024031;
assign addr[3075]= -2126796855;
assign addr[3076]= -2147470025;
assign addr[3077]= -2124624598;
assign addr[3078]= -2058723538;
assign addr[3079]= -1951102334;
assign addr[3080]= -1803941934;
assign addr[3081]= -1620224553;
assign addr[3082]= -1403673233;
assign addr[3083]= -1158676398;
assign addr[3084]= -890198924;
assign addr[3085]= -603681519;
assign addr[3086]= -304930476;
assign addr[3087]= 0;
assign addr[3088]= 304930476;
assign addr[3089]= 603681519;
assign addr[3090]= 890198924;
assign addr[3091]= 1158676398;
assign addr[3092]= 1403673233;
assign addr[3093]= 1620224553;
assign addr[3094]= 1803941934;
assign addr[3095]= 1951102334;
assign addr[3096]= 2058723538;
assign addr[3097]= 2124624598;
assign addr[3098]= 2147470025;
assign addr[3099]= 2126796855;
assign addr[3100]= 2063024031;
assign addr[3101]= 1957443913;
assign addr[3102]= 1812196087;
assign addr[3103]= 1630224009;
assign addr[3104]= 1415215352;
assign addr[3105]= 1171527280;
assign addr[3106]= 904098143;
assign addr[3107]= 618347408;
assign addr[3108]= 320065829;
assign addr[3109]= 15298099;
assign addr[3110]= -289779648;
assign addr[3111]= -588984994;
assign addr[3112]= -876254528;
assign addr[3113]= -1145766716;
assign addr[3114]= -1392059879;
assign addr[3115]= -1610142873;
assign addr[3116]= -1795596234;
assign addr[3117]= -1944661739;
assign addr[3118]= -2054318569;
assign addr[3119]= -2122344521;
assign addr[3120]= -2147361045;
assign addr[3121]= -2128861181;
assign addr[3122]= -2067219829;
assign addr[3123]= -1963686155;
assign addr[3124]= -1820358275;
assign addr[3125]= -1640140734;
assign addr[3126]= -1426685652;
assign addr[3127]= -1184318708;
assign addr[3128]= -917951481;
assign addr[3129]= -632981917;
assign addr[3130]= -335184940;
assign addr[3131]= -30595422;
assign addr[3132]= 274614114;
assign addr[3133]= 574258580;
assign addr[3134]= 862265664;
assign addr[3135]= 1132798888;
assign addr[3136]= 1380375881;
assign addr[3137]= 1599979481;
assign addr[3138]= 1787159411;
assign addr[3139]= 1938122457;
assign addr[3140]= 2049809346;
assign addr[3141]= 2119956737;
assign addr[3142]= 2147143090;
assign addr[3143]= 2130817471;
assign addr[3144]= 2071310720;
assign addr[3145]= 1969828744;
assign addr[3146]= 1828428082;
assign addr[3147]= 1649974225;
assign addr[3148]= 1438083551;
assign addr[3149]= 1197050035;
assign addr[3150]= 931758235;
assign addr[3151]= 647584304;
assign addr[3152]= 350287041;
assign addr[3153]= 45891193;
assign addr[3154]= -259434643;
assign addr[3155]= -559503022;
assign addr[3156]= -848233042;
assign addr[3157]= -1119773573;
assign addr[3158]= -1368621831;
assign addr[3159]= -1589734894;
assign addr[3160]= -1778631892;
assign addr[3161]= -1931484818;
assign addr[3162]= -2045196100;
assign addr[3163]= -2117461370;
assign addr[3164]= -2146816171;
assign addr[3165]= -2132665626;
assign addr[3166]= -2075296495;
assign addr[3167]= -1975871368;
assign addr[3168]= -1836405100;
assign addr[3169]= -1659723983;
assign addr[3170]= -1449408469;
assign addr[3171]= -1209720613;
assign addr[3172]= -945517704;
assign addr[3173]= -662153826;
assign addr[3174]= -365371365;
assign addr[3175]= -61184634;
assign addr[3176]= 244242007;
assign addr[3177]= 544719071;
assign addr[3178]= 834157373;
assign addr[3179]= 1106691431;
assign addr[3180]= 1356798326;
assign addr[3181]= 1579409630;
assign addr[3182]= 1770014111;
assign addr[3183]= 1924749160;
assign addr[3184]= 2040479063;
assign addr[3185]= 2114858546;
assign addr[3186]= 2146380306;
assign addr[3187]= 2134405552;
assign addr[3188]= 2079176953;
assign addr[3189]= 1981813720;
assign addr[3190]= 1844288924;
assign addr[3191]= 1669389513;
assign addr[3192]= 1460659832;
assign addr[3193]= 1222329801;
assign addr[3194]= 959229189;
assign addr[3195]= 676689746;
assign addr[3196]= 380437148;
assign addr[3197]= 76474970;
assign addr[3198]= -229036977;
assign addr[3199]= -529907477;
assign addr[3200]= -820039373;
assign addr[3201]= -1093553126;
assign addr[3202]= -1344905966;
assign addr[3203]= -1569004214;
assign addr[3204]= -1761306505;
assign addr[3205]= -1917915825;
assign addr[3206]= -2035658475;
assign addr[3207]= -2112148396;
assign addr[3208]= -2145835515;
assign addr[3209]= -2136037160;
assign addr[3210]= -2082951896;
assign addr[3211]= -1987655498;
assign addr[3212]= -1852079154;
assign addr[3213]= -1678970324;
assign addr[3214]= -1471837070;
assign addr[3215]= -1234876957;
assign addr[3216]= -972891995;
assign addr[3217]= -691191324;
assign addr[3218]= -395483624;
assign addr[3219]= -91761426;
assign addr[3220]= 213820322;
assign addr[3221]= 515068990;
assign addr[3222]= 805879757;
assign addr[3223]= 1080359326;
assign addr[3224]= 1332945355;
assign addr[3225]= 1558519173;
assign addr[3226]= 1752509516;
assign addr[3227]= 1910985158;
assign addr[3228]= 2030734582;
assign addr[3229]= 2109331059;
assign addr[3230]= 2145181827;
assign addr[3231]= 2137560369;
assign addr[3232]= 2086621133;
assign addr[3233]= 1993396407;
assign addr[3234]= 1859775393;
assign addr[3235]= 1688465931;
assign addr[3236]= 1482939614;
assign addr[3237]= 1247361445;
assign addr[3238]= 986505429;
assign addr[3239]= 705657826;
assign addr[3240]= 410510029;
assign addr[3241]= 107043224;
assign addr[3242]= -198592817;
assign addr[3243]= -500204365;
assign addr[3244]= -791679244;
assign addr[3245]= -1067110699;
assign addr[3246]= -1320917099;
assign addr[3247]= -1547955041;
assign addr[3248]= -1743623590;
assign addr[3249]= -1903957513;
assign addr[3250]= -2025707632;
assign addr[3251]= -2106406677;
assign addr[3252]= -2144419275;
assign addr[3253]= -2138975100;
assign addr[3254]= -2090184478;
assign addr[3255]= -1999036154;
assign addr[3256]= -1867377253;
assign addr[3257]= -1697875851;
assign addr[3258]= -1493966902;
assign addr[3259]= -1259782632;
assign addr[3260]= -1000068799;
assign addr[3261]= -720088517;
assign addr[3262]= -425515602;
assign addr[3263]= -122319591;
assign addr[3264]= 183355234;
assign addr[3265]= 485314355;
assign addr[3266]= 777438554;
assign addr[3267]= 1053807919;
assign addr[3268]= 1308821808;
assign addr[3269]= 1537312353;
assign addr[3270]= 1734649179;
assign addr[3271]= 1896833245;
assign addr[3272]= 2020577882;
assign addr[3273]= 2103375398;
assign addr[3274]= 2143547897;
assign addr[3275]= 2140281282;
assign addr[3276]= 2093641749;
assign addr[3277]= 2004574453;
assign addr[3278]= 1874884346;
assign addr[3279]= 1707199606;
assign addr[3280]= 1504918373;
assign addr[3281]= 1272139887;
assign addr[3282]= 1013581418;
assign addr[3283]= 734482665;
assign addr[3284]= 440499581;
assign addr[3285]= 137589750;
assign addr[3286]= -168108346;
assign addr[3287]= -470399716;
assign addr[3288]= -763158411;
assign addr[3289]= -1040451659;
assign addr[3290]= -1296660098;
assign addr[3291]= -1526591649;
assign addr[3292]= -1725586737;
assign addr[3293]= -1889612716;
assign addr[3294]= -2015345591;
assign addr[3295]= -2100237377;
assign addr[3296]= -2142567738;
assign addr[3297]= -2141478848;
assign addr[3298]= -2096992772;
assign addr[3299]= -2010011024;
assign addr[3300]= -1882296293;
assign addr[3301]= -1716436725;
assign addr[3302]= -1515793473;
assign addr[3303]= -1284432584;
assign addr[3304]= -1027042599;
assign addr[3305]= -748839539;
assign addr[3306]= -455461206;
assign addr[3307]= -152852926;
assign addr[3308]= 152852926;
assign addr[3309]= 455461206;
assign addr[3310]= 748839539;
assign addr[3311]= 1027042599;
assign addr[3312]= 1284432584;
assign addr[3313]= 1515793473;
assign addr[3314]= 1716436725;
assign addr[3315]= 1882296293;
assign addr[3316]= 2010011024;
assign addr[3317]= 2096992772;
assign addr[3318]= 2141478848;
assign addr[3319]= 2142567738;
assign addr[3320]= 2100237377;
assign addr[3321]= 2015345591;
assign addr[3322]= 1889612716;
assign addr[3323]= 1725586737;
assign addr[3324]= 1526591649;
assign addr[3325]= 1296660098;
assign addr[3326]= 1040451659;
assign addr[3327]= 763158411;
assign addr[3328]= 470399716;
assign addr[3329]= 168108346;
assign addr[3330]= -137589750;
assign addr[3331]= -440499581;
assign addr[3332]= -734482665;
assign addr[3333]= -1013581418;
assign addr[3334]= -1272139887;
assign addr[3335]= -1504918373;
assign addr[3336]= -1707199606;
assign addr[3337]= -1874884346;
assign addr[3338]= -2004574453;
assign addr[3339]= -2093641749;
assign addr[3340]= -2140281282;
assign addr[3341]= -2143547897;
assign addr[3342]= -2103375398;
assign addr[3343]= -2020577882;
assign addr[3344]= -1896833245;
assign addr[3345]= -1734649179;
assign addr[3346]= -1537312353;
assign addr[3347]= -1308821808;
assign addr[3348]= -1053807919;
assign addr[3349]= -777438554;
assign addr[3350]= -485314355;
assign addr[3351]= -183355234;
assign addr[3352]= 122319591;
assign addr[3353]= 425515602;
assign addr[3354]= 720088517;
assign addr[3355]= 1000068799;
assign addr[3356]= 1259782632;
assign addr[3357]= 1493966902;
assign addr[3358]= 1697875851;
assign addr[3359]= 1867377253;
assign addr[3360]= 1999036154;
assign addr[3361]= 2090184478;
assign addr[3362]= 2138975100;
assign addr[3363]= 2144419275;
assign addr[3364]= 2106406677;
assign addr[3365]= 2025707632;
assign addr[3366]= 1903957513;
assign addr[3367]= 1743623590;
assign addr[3368]= 1547955041;
assign addr[3369]= 1320917099;
assign addr[3370]= 1067110699;
assign addr[3371]= 791679244;
assign addr[3372]= 500204365;
assign addr[3373]= 198592817;
assign addr[3374]= -107043224;
assign addr[3375]= -410510029;
assign addr[3376]= -705657826;
assign addr[3377]= -986505429;
assign addr[3378]= -1247361445;
assign addr[3379]= -1482939614;
assign addr[3380]= -1688465931;
assign addr[3381]= -1859775393;
assign addr[3382]= -1993396407;
assign addr[3383]= -2086621133;
assign addr[3384]= -2137560369;
assign addr[3385]= -2145181827;
assign addr[3386]= -2109331059;
assign addr[3387]= -2030734582;
assign addr[3388]= -1910985158;
assign addr[3389]= -1752509516;
assign addr[3390]= -1558519173;
assign addr[3391]= -1332945355;
assign addr[3392]= -1080359326;
assign addr[3393]= -805879757;
assign addr[3394]= -515068990;
assign addr[3395]= -213820322;
assign addr[3396]= 91761426;
assign addr[3397]= 395483624;
assign addr[3398]= 691191324;
assign addr[3399]= 972891995;
assign addr[3400]= 1234876957;
assign addr[3401]= 1471837070;
assign addr[3402]= 1678970324;
assign addr[3403]= 1852079154;
assign addr[3404]= 1987655498;
assign addr[3405]= 2082951896;
assign addr[3406]= 2136037160;
assign addr[3407]= 2145835515;
assign addr[3408]= 2112148396;
assign addr[3409]= 2035658475;
assign addr[3410]= 1917915825;
assign addr[3411]= 1761306505;
assign addr[3412]= 1569004214;
assign addr[3413]= 1344905966;
assign addr[3414]= 1093553126;
assign addr[3415]= 820039373;
assign addr[3416]= 529907477;
assign addr[3417]= 229036977;
assign addr[3418]= -76474970;
assign addr[3419]= -380437148;
assign addr[3420]= -676689746;
assign addr[3421]= -959229189;
assign addr[3422]= -1222329801;
assign addr[3423]= -1460659832;
assign addr[3424]= -1669389513;
assign addr[3425]= -1844288924;
assign addr[3426]= -1981813720;
assign addr[3427]= -2079176953;
assign addr[3428]= -2134405552;
assign addr[3429]= -2146380306;
assign addr[3430]= -2114858546;
assign addr[3431]= -2040479063;
assign addr[3432]= -1924749160;
assign addr[3433]= -1770014111;
assign addr[3434]= -1579409630;
assign addr[3435]= -1356798326;
assign addr[3436]= -1106691431;
assign addr[3437]= -834157373;
assign addr[3438]= -544719071;
assign addr[3439]= -244242007;
assign addr[3440]= 61184634;
assign addr[3441]= 365371365;
assign addr[3442]= 662153826;
assign addr[3443]= 945517704;
assign addr[3444]= 1209720613;
assign addr[3445]= 1449408469;
assign addr[3446]= 1659723983;
assign addr[3447]= 1836405100;
assign addr[3448]= 1975871368;
assign addr[3449]= 2075296495;
assign addr[3450]= 2132665626;
assign addr[3451]= 2146816171;
assign addr[3452]= 2117461370;
assign addr[3453]= 2045196100;
assign addr[3454]= 1931484818;
assign addr[3455]= 1778631892;
assign addr[3456]= 1589734894;
assign addr[3457]= 1368621831;
assign addr[3458]= 1119773573;
assign addr[3459]= 848233042;
assign addr[3460]= 559503022;
assign addr[3461]= 259434643;
assign addr[3462]= -45891193;
assign addr[3463]= -350287041;
assign addr[3464]= -647584304;
assign addr[3465]= -931758235;
assign addr[3466]= -1197050035;
assign addr[3467]= -1438083551;
assign addr[3468]= -1649974225;
assign addr[3469]= -1828428082;
assign addr[3470]= -1969828744;
assign addr[3471]= -2071310720;
assign addr[3472]= -2130817471;
assign addr[3473]= -2147143090;
assign addr[3474]= -2119956737;
assign addr[3475]= -2049809346;
assign addr[3476]= -1938122457;
assign addr[3477]= -1787159411;
assign addr[3478]= -1599979481;
assign addr[3479]= -1380375881;
assign addr[3480]= -1132798888;
assign addr[3481]= -862265664;
assign addr[3482]= -574258580;
assign addr[3483]= -274614114;
assign addr[3484]= 30595422;
assign addr[3485]= 335184940;
assign addr[3486]= 632981917;
assign addr[3487]= 917951481;
assign addr[3488]= 1184318708;
assign addr[3489]= 1426685652;
assign addr[3490]= 1640140734;
assign addr[3491]= 1820358275;
assign addr[3492]= 1963686155;
assign addr[3493]= 2067219829;
assign addr[3494]= 2128861181;
assign addr[3495]= 2147361045;
assign addr[3496]= 2122344521;
assign addr[3497]= 2054318569;
assign addr[3498]= 1944661739;
assign addr[3499]= 1795596234;
assign addr[3500]= 1610142873;
assign addr[3501]= 1392059879;
assign addr[3502]= 1145766716;
assign addr[3503]= 876254528;
assign addr[3504]= 588984994;
assign addr[3505]= 289779648;
assign addr[3506]= -15298099;
assign addr[3507]= -320065829;
assign addr[3508]= -618347408;
assign addr[3509]= -904098143;
assign addr[3510]= -1171527280;
assign addr[3511]= -1415215352;
assign addr[3512]= -1630224009;
assign addr[3513]= -1812196087;
assign addr[3514]= -1957443913;
assign addr[3515]= -2063024031;
assign addr[3516]= -2126796855;
assign addr[3517]= -2147470025;
assign addr[3518]= -2124624598;
assign addr[3519]= -2058723538;
assign addr[3520]= -1951102334;
assign addr[3521]= -1803941934;
assign addr[3522]= -1620224553;
assign addr[3523]= -1403673233;
assign addr[3524]= -1158676398;
assign addr[3525]= -890198924;
assign addr[3526]= -603681519;
assign addr[3527]= -304930476;
assign addr[3528]= 0;
assign addr[3529]= 304930476;
assign addr[3530]= 603681519;
assign addr[3531]= 890198924;
assign addr[3532]= 1158676398;
assign addr[3533]= 1403673233;
assign addr[3534]= 1620224553;
assign addr[3535]= 1803941934;
assign addr[3536]= 1951102334;
assign addr[3537]= 2058723538;
assign addr[3538]= 2124624598;
assign addr[3539]= 2147470025;
assign addr[3540]= 2126796855;
assign addr[3541]= 2063024031;
assign addr[3542]= 1957443913;
assign addr[3543]= 1812196087;
assign addr[3544]= 1630224009;
assign addr[3545]= 1415215352;
assign addr[3546]= 1171527280;
assign addr[3547]= 904098143;
assign addr[3548]= 618347408;
assign addr[3549]= 320065829;
assign addr[3550]= 15298099;
assign addr[3551]= -289779648;
assign addr[3552]= -588984994;
assign addr[3553]= -876254528;
assign addr[3554]= -1145766716;
assign addr[3555]= -1392059879;
assign addr[3556]= -1610142873;
assign addr[3557]= -1795596234;
assign addr[3558]= -1944661739;
assign addr[3559]= -2054318569;
assign addr[3560]= -2122344521;
assign addr[3561]= -2147361045;
assign addr[3562]= -2128861181;
assign addr[3563]= -2067219829;
assign addr[3564]= -1963686155;
assign addr[3565]= -1820358275;
assign addr[3566]= -1640140734;
assign addr[3567]= -1426685652;
assign addr[3568]= -1184318708;
assign addr[3569]= -917951481;
assign addr[3570]= -632981917;
assign addr[3571]= -335184940;
assign addr[3572]= -30595422;
assign addr[3573]= 274614114;
assign addr[3574]= 574258580;
assign addr[3575]= 862265664;
assign addr[3576]= 1132798888;
assign addr[3577]= 1380375881;
assign addr[3578]= 1599979481;
assign addr[3579]= 1787159411;
assign addr[3580]= 1938122457;
assign addr[3581]= 2049809346;
assign addr[3582]= 2119956737;
assign addr[3583]= 2147143090;
assign addr[3584]= 2130817471;
assign addr[3585]= 2071310720;
assign addr[3586]= 1969828744;
assign addr[3587]= 1828428082;
assign addr[3588]= 1649974225;
assign addr[3589]= 1438083551;
assign addr[3590]= 1197050035;
assign addr[3591]= 931758235;
assign addr[3592]= 647584304;
assign addr[3593]= 350287041;
assign addr[3594]= 45891193;
assign addr[3595]= -259434643;
assign addr[3596]= -559503022;
assign addr[3597]= -848233042;
assign addr[3598]= -1119773573;
assign addr[3599]= -1368621831;
assign addr[3600]= -1589734894;
assign addr[3601]= -1778631892;
assign addr[3602]= -1931484818;
assign addr[3603]= -2045196100;
assign addr[3604]= -2117461370;
assign addr[3605]= -2146816171;
assign addr[3606]= -2132665626;
assign addr[3607]= -2075296495;
assign addr[3608]= -1975871368;
assign addr[3609]= -1836405100;
assign addr[3610]= -1659723983;
assign addr[3611]= -1449408469;
assign addr[3612]= -1209720613;
assign addr[3613]= -945517704;
assign addr[3614]= -662153826;
assign addr[3615]= -365371365;
assign addr[3616]= -61184634;
assign addr[3617]= 244242007;
assign addr[3618]= 544719071;
assign addr[3619]= 834157373;
assign addr[3620]= 1106691431;
assign addr[3621]= 1356798326;
assign addr[3622]= 1579409630;
assign addr[3623]= 1770014111;
assign addr[3624]= 1924749160;
assign addr[3625]= 2040479063;
assign addr[3626]= 2114858546;
assign addr[3627]= 2146380306;
assign addr[3628]= 2134405552;
assign addr[3629]= 2079176953;
assign addr[3630]= 1981813720;
assign addr[3631]= 1844288924;
assign addr[3632]= 1669389513;
assign addr[3633]= 1460659832;
assign addr[3634]= 1222329801;
assign addr[3635]= 959229189;
assign addr[3636]= 676689746;
assign addr[3637]= 380437148;
assign addr[3638]= 76474970;
assign addr[3639]= -229036977;
assign addr[3640]= -529907477;
assign addr[3641]= -820039373;
assign addr[3642]= -1093553126;
assign addr[3643]= -1344905966;
assign addr[3644]= -1569004214;
assign addr[3645]= -1761306505;
assign addr[3646]= -1917915825;
assign addr[3647]= -2035658475;
assign addr[3648]= -2112148396;
assign addr[3649]= -2145835515;
assign addr[3650]= -2136037160;
assign addr[3651]= -2082951896;
assign addr[3652]= -1987655498;
assign addr[3653]= -1852079154;
assign addr[3654]= -1678970324;
assign addr[3655]= -1471837070;
assign addr[3656]= -1234876957;
assign addr[3657]= -972891995;
assign addr[3658]= -691191324;
assign addr[3659]= -395483624;
assign addr[3660]= -91761426;
assign addr[3661]= 213820322;
assign addr[3662]= 515068990;
assign addr[3663]= 805879757;
assign addr[3664]= 1080359326;
assign addr[3665]= 1332945355;
assign addr[3666]= 1558519173;
assign addr[3667]= 1752509516;
assign addr[3668]= 1910985158;
assign addr[3669]= 2030734582;
assign addr[3670]= 2109331059;
assign addr[3671]= 2145181827;
assign addr[3672]= 2137560369;
assign addr[3673]= 2086621133;
assign addr[3674]= 1993396407;
assign addr[3675]= 1859775393;
assign addr[3676]= 1688465931;
assign addr[3677]= 1482939614;
assign addr[3678]= 1247361445;
assign addr[3679]= 986505429;
assign addr[3680]= 705657826;
assign addr[3681]= 410510029;
assign addr[3682]= 107043224;
assign addr[3683]= -198592817;
assign addr[3684]= -500204365;
assign addr[3685]= -791679244;
assign addr[3686]= -1067110699;
assign addr[3687]= -1320917099;
assign addr[3688]= -1547955041;
assign addr[3689]= -1743623590;
assign addr[3690]= -1903957513;
assign addr[3691]= -2025707632;
assign addr[3692]= -2106406677;
assign addr[3693]= -2144419275;
assign addr[3694]= -2138975100;
assign addr[3695]= -2090184478;
assign addr[3696]= -1999036154;
assign addr[3697]= -1867377253;
assign addr[3698]= -1697875851;
assign addr[3699]= -1493966902;
assign addr[3700]= -1259782632;
assign addr[3701]= -1000068799;
assign addr[3702]= -720088517;
assign addr[3703]= -425515602;
assign addr[3704]= -122319591;
assign addr[3705]= 183355234;
assign addr[3706]= 485314355;
assign addr[3707]= 777438554;
assign addr[3708]= 1053807919;
assign addr[3709]= 1308821808;
assign addr[3710]= 1537312353;
assign addr[3711]= 1734649179;
assign addr[3712]= 1896833245;
assign addr[3713]= 2020577882;
assign addr[3714]= 2103375398;
assign addr[3715]= 2143547897;
assign addr[3716]= 2140281282;
assign addr[3717]= 2093641749;
assign addr[3718]= 2004574453;
assign addr[3719]= 1874884346;
assign addr[3720]= 1707199606;
assign addr[3721]= 1504918373;
assign addr[3722]= 1272139887;
assign addr[3723]= 1013581418;
assign addr[3724]= 734482665;
assign addr[3725]= 440499581;
assign addr[3726]= 137589750;
assign addr[3727]= -168108346;
assign addr[3728]= -470399716;
assign addr[3729]= -763158411;
assign addr[3730]= -1040451659;
assign addr[3731]= -1296660098;
assign addr[3732]= -1526591649;
assign addr[3733]= -1725586737;
assign addr[3734]= -1889612716;
assign addr[3735]= -2015345591;
assign addr[3736]= -2100237377;
assign addr[3737]= -2142567738;
assign addr[3738]= -2141478848;
assign addr[3739]= -2096992772;
assign addr[3740]= -2010011024;
assign addr[3741]= -1882296293;
assign addr[3742]= -1716436725;
assign addr[3743]= -1515793473;
assign addr[3744]= -1284432584;
assign addr[3745]= -1027042599;
assign addr[3746]= -748839539;
assign addr[3747]= -455461206;
assign addr[3748]= -152852926;
assign addr[3749]= 152852926;
assign addr[3750]= 455461206;
assign addr[3751]= 748839539;
assign addr[3752]= 1027042599;
assign addr[3753]= 1284432584;
assign addr[3754]= 1515793473;
assign addr[3755]= 1716436725;
assign addr[3756]= 1882296293;
assign addr[3757]= 2010011024;
assign addr[3758]= 2096992772;
assign addr[3759]= 2141478848;
assign addr[3760]= 2142567738;
assign addr[3761]= 2100237377;
assign addr[3762]= 2015345591;
assign addr[3763]= 1889612716;
assign addr[3764]= 1725586737;
assign addr[3765]= 1526591649;
assign addr[3766]= 1296660098;
assign addr[3767]= 1040451659;
assign addr[3768]= 763158411;
assign addr[3769]= 470399716;
assign addr[3770]= 168108346;
assign addr[3771]= -137589750;
assign addr[3772]= -440499581;
assign addr[3773]= -734482665;
assign addr[3774]= -1013581418;
assign addr[3775]= -1272139887;
assign addr[3776]= -1504918373;
assign addr[3777]= -1707199606;
assign addr[3778]= -1874884346;
assign addr[3779]= -2004574453;
assign addr[3780]= -2093641749;
assign addr[3781]= -2140281282;
assign addr[3782]= -2143547897;
assign addr[3783]= -2103375398;
assign addr[3784]= -2020577882;
assign addr[3785]= -1896833245;
assign addr[3786]= -1734649179;
assign addr[3787]= -1537312353;
assign addr[3788]= -1308821808;
assign addr[3789]= -1053807919;
assign addr[3790]= -777438554;
assign addr[3791]= -485314355;
assign addr[3792]= -183355234;
assign addr[3793]= 122319591;
assign addr[3794]= 425515602;
assign addr[3795]= 720088517;
assign addr[3796]= 1000068799;
assign addr[3797]= 1259782632;
assign addr[3798]= 1493966902;
assign addr[3799]= 1697875851;
assign addr[3800]= 1867377253;
assign addr[3801]= 1999036154;
assign addr[3802]= 2090184478;
assign addr[3803]= 2138975100;
assign addr[3804]= 2144419275;
assign addr[3805]= 2106406677;
assign addr[3806]= 2025707632;
assign addr[3807]= 1903957513;
assign addr[3808]= 1743623590;
assign addr[3809]= 1547955041;
assign addr[3810]= 1320917099;
assign addr[3811]= 1067110699;
assign addr[3812]= 791679244;
assign addr[3813]= 500204365;
assign addr[3814]= 198592817;
assign addr[3815]= -107043224;
assign addr[3816]= -410510029;
assign addr[3817]= -705657826;
assign addr[3818]= -986505429;
assign addr[3819]= -1247361445;
assign addr[3820]= -1482939614;
assign addr[3821]= -1688465931;
assign addr[3822]= -1859775393;
assign addr[3823]= -1993396407;
assign addr[3824]= -2086621133;
assign addr[3825]= -2137560369;
assign addr[3826]= -2145181827;
assign addr[3827]= -2109331059;
assign addr[3828]= -2030734582;
assign addr[3829]= -1910985158;
assign addr[3830]= -1752509516;
assign addr[3831]= -1558519173;
assign addr[3832]= -1332945355;
assign addr[3833]= -1080359326;
assign addr[3834]= -805879757;
assign addr[3835]= -515068990;
assign addr[3836]= -213820322;
assign addr[3837]= 91761426;
assign addr[3838]= 395483624;
assign addr[3839]= 691191324;
assign addr[3840]= 972891995;
assign addr[3841]= 1234876957;
assign addr[3842]= 1471837070;
assign addr[3843]= 1678970324;
assign addr[3844]= 1852079154;
assign addr[3845]= 1987655498;
assign addr[3846]= 2082951896;
assign addr[3847]= 2136037160;
assign addr[3848]= 2145835515;
assign addr[3849]= 2112148396;
assign addr[3850]= 2035658475;
assign addr[3851]= 1917915825;
assign addr[3852]= 1761306505;
assign addr[3853]= 1569004214;
assign addr[3854]= 1344905966;
assign addr[3855]= 1093553126;
assign addr[3856]= 820039373;
assign addr[3857]= 529907477;
assign addr[3858]= 229036977;
assign addr[3859]= -76474970;
assign addr[3860]= -380437148;
assign addr[3861]= -676689746;
assign addr[3862]= -959229189;
assign addr[3863]= -1222329801;
assign addr[3864]= -1460659832;
assign addr[3865]= -1669389513;
assign addr[3866]= -1844288924;
assign addr[3867]= -1981813720;
assign addr[3868]= -2079176953;
assign addr[3869]= -2134405552;
assign addr[3870]= -2146380306;
assign addr[3871]= -2114858546;
assign addr[3872]= -2040479063;
assign addr[3873]= -1924749160;
assign addr[3874]= -1770014111;
assign addr[3875]= -1579409630;
assign addr[3876]= -1356798326;
assign addr[3877]= -1106691431;
assign addr[3878]= -834157373;
assign addr[3879]= -544719071;
assign addr[3880]= -244242007;
assign addr[3881]= 61184634;
assign addr[3882]= 365371365;
assign addr[3883]= 662153826;
assign addr[3884]= 945517704;
assign addr[3885]= 1209720613;
assign addr[3886]= 1449408469;
assign addr[3887]= 1659723983;
assign addr[3888]= 1836405100;
assign addr[3889]= 1975871368;
assign addr[3890]= 2075296495;
assign addr[3891]= 2132665626;
assign addr[3892]= 2146816171;
assign addr[3893]= 2117461370;
assign addr[3894]= 2045196100;
assign addr[3895]= 1931484818;
assign addr[3896]= 1778631892;
assign addr[3897]= 1589734894;
assign addr[3898]= 1368621831;
assign addr[3899]= 1119773573;
assign addr[3900]= 848233042;
assign addr[3901]= 559503022;
assign addr[3902]= 259434643;
assign addr[3903]= -45891193;
assign addr[3904]= -350287041;
assign addr[3905]= -647584304;
assign addr[3906]= -931758235;
assign addr[3907]= -1197050035;
assign addr[3908]= -1438083551;
assign addr[3909]= -1649974225;
assign addr[3910]= -1828428082;
assign addr[3911]= -1969828744;
assign addr[3912]= -2071310720;
assign addr[3913]= -2130817471;
assign addr[3914]= -2147143090;
assign addr[3915]= -2119956737;
assign addr[3916]= -2049809346;
assign addr[3917]= -1938122457;
assign addr[3918]= -1787159411;
assign addr[3919]= -1599979481;
assign addr[3920]= -1380375881;
assign addr[3921]= -1132798888;
assign addr[3922]= -862265664;
assign addr[3923]= -574258580;
assign addr[3924]= -274614114;
assign addr[3925]= 30595422;
assign addr[3926]= 335184940;
assign addr[3927]= 632981917;
assign addr[3928]= 917951481;
assign addr[3929]= 1184318708;
assign addr[3930]= 1426685652;
assign addr[3931]= 1640140734;
assign addr[3932]= 1820358275;
assign addr[3933]= 1963686155;
assign addr[3934]= 2067219829;
assign addr[3935]= 2128861181;
assign addr[3936]= 2147361045;
assign addr[3937]= 2122344521;
assign addr[3938]= 2054318569;
assign addr[3939]= 1944661739;
assign addr[3940]= 1795596234;
assign addr[3941]= 1610142873;
assign addr[3942]= 1392059879;
assign addr[3943]= 1145766716;
assign addr[3944]= 876254528;
assign addr[3945]= 588984994;
assign addr[3946]= 289779648;
assign addr[3947]= -15298099;
assign addr[3948]= -320065829;
assign addr[3949]= -618347408;
assign addr[3950]= -904098143;
assign addr[3951]= -1171527280;
assign addr[3952]= -1415215352;
assign addr[3953]= -1630224009;
assign addr[3954]= -1812196087;
assign addr[3955]= -1957443913;
assign addr[3956]= -2063024031;
assign addr[3957]= -2126796855;
assign addr[3958]= -2147470025;
assign addr[3959]= -2124624598;
assign addr[3960]= -2058723538;
assign addr[3961]= -1951102334;
assign addr[3962]= -1803941934;
assign addr[3963]= -1620224553;
assign addr[3964]= -1403673233;
assign addr[3965]= -1158676398;
assign addr[3966]= -890198924;
assign addr[3967]= -603681519;
assign addr[3968]= -304930476;
assign addr[3969]= 0;
assign addr[3970]= 304930476;
assign addr[3971]= 603681519;
assign addr[3972]= 890198924;
assign addr[3973]= 1158676398;
assign addr[3974]= 1403673233;
assign addr[3975]= 1620224553;
assign addr[3976]= 1803941934;
assign addr[3977]= 1951102334;
assign addr[3978]= 2058723538;
assign addr[3979]= 2124624598;
assign addr[3980]= 2147470025;
assign addr[3981]= 2126796855;
assign addr[3982]= 2063024031;
assign addr[3983]= 1957443913;
assign addr[3984]= 1812196087;
assign addr[3985]= 1630224009;
assign addr[3986]= 1415215352;
assign addr[3987]= 1171527280;
assign addr[3988]= 904098143;
assign addr[3989]= 618347408;
assign addr[3990]= 320065829;
assign addr[3991]= 15298099;
assign addr[3992]= -289779648;
assign addr[3993]= -588984994;
assign addr[3994]= -876254528;
assign addr[3995]= -1145766716;
assign addr[3996]= -1392059879;
assign addr[3997]= -1610142873;
assign addr[3998]= -1795596234;
assign addr[3999]= -1944661739;
assign addr[4000]= -2054318569;
assign addr[4001]= -2122344521;
assign addr[4002]= -2147361045;
assign addr[4003]= -2128861181;
assign addr[4004]= -2067219829;
assign addr[4005]= -1963686155;
assign addr[4006]= -1820358275;
assign addr[4007]= -1640140734;
assign addr[4008]= -1426685652;
assign addr[4009]= -1184318708;
assign addr[4010]= -917951481;
assign addr[4011]= -632981917;
assign addr[4012]= -335184940;
assign addr[4013]= -30595422;
assign addr[4014]= 274614114;
assign addr[4015]= 574258580;
assign addr[4016]= 862265664;
assign addr[4017]= 1132798888;
assign addr[4018]= 1380375881;
assign addr[4019]= 1599979481;
assign addr[4020]= 1787159411;
assign addr[4021]= 1938122457;
assign addr[4022]= 2049809346;
assign addr[4023]= 2119956737;
assign addr[4024]= 2147143090;
assign addr[4025]= 2130817471;
assign addr[4026]= 2071310720;
assign addr[4027]= 1969828744;
assign addr[4028]= 1828428082;
assign addr[4029]= 1649974225;
assign addr[4030]= 1438083551;
assign addr[4031]= 1197050035;
assign addr[4032]= 931758235;
assign addr[4033]= 647584304;
assign addr[4034]= 350287041;
assign addr[4035]= 45891193;
assign addr[4036]= -259434643;
assign addr[4037]= -559503022;
assign addr[4038]= -848233042;
assign addr[4039]= -1119773573;
assign addr[4040]= -1368621831;
assign addr[4041]= -1589734894;
assign addr[4042]= -1778631892;
assign addr[4043]= -1931484818;
assign addr[4044]= -2045196100;
assign addr[4045]= -2117461370;
assign addr[4046]= -2146816171;
assign addr[4047]= -2132665626;
assign addr[4048]= -2075296495;
assign addr[4049]= -1975871368;
assign addr[4050]= -1836405100;
assign addr[4051]= -1659723983;
assign addr[4052]= -1449408469;
assign addr[4053]= -1209720613;
assign addr[4054]= -945517704;
assign addr[4055]= -662153826;
assign addr[4056]= -365371365;
assign addr[4057]= -61184634;
assign addr[4058]= 244242007;
assign addr[4059]= 544719071;
assign addr[4060]= 834157373;
assign addr[4061]= 1106691431;
assign addr[4062]= 1356798326;
assign addr[4063]= 1579409630;
assign addr[4064]= 1770014111;
assign addr[4065]= 1924749160;
assign addr[4066]= 2040479063;
assign addr[4067]= 2114858546;
assign addr[4068]= 2146380306;
assign addr[4069]= 2134405552;
assign addr[4070]= 2079176953;
assign addr[4071]= 1981813720;
assign addr[4072]= 1844288924;
assign addr[4073]= 1669389513;
assign addr[4074]= 1460659832;
assign addr[4075]= 1222329801;
assign addr[4076]= 959229189;
assign addr[4077]= 676689746;
assign addr[4078]= 380437148;
assign addr[4079]= 76474970;
assign addr[4080]= -229036977;
assign addr[4081]= -529907477;
assign addr[4082]= -820039373;
assign addr[4083]= -1093553126;
assign addr[4084]= -1344905966;
assign addr[4085]= -1569004214;
assign addr[4086]= -1761306505;
assign addr[4087]= -1917915825;
assign addr[4088]= -2035658475;
assign addr[4089]= -2112148396;
assign addr[4090]= -2145835515;
assign addr[4091]= -2136037160;
assign addr[4092]= -2082951896;
assign addr[4093]= -1987655498;
assign addr[4094]= -1852079154;
assign addr[4095]= -1678970324;
assign addr[4096]= -1471837070;
assign addr[4097]= -1234876957;
assign addr[4098]= -972891995;
assign addr[4099]= -691191324;
assign addr[4100]= -395483624;
assign addr[4101]= -91761426;
assign addr[4102]= 213820322;
assign addr[4103]= 515068990;
assign addr[4104]= 805879757;
assign addr[4105]= 1080359326;
assign addr[4106]= 1332945355;
assign addr[4107]= 1558519173;
assign addr[4108]= 1752509516;
assign addr[4109]= 1910985158;
assign addr[4110]= 2030734582;
assign addr[4111]= 2109331059;
assign addr[4112]= 2145181827;
assign addr[4113]= 2137560369;
assign addr[4114]= 2086621133;
assign addr[4115]= 1993396407;
assign addr[4116]= 1859775393;
assign addr[4117]= 1688465931;
assign addr[4118]= 1482939614;
assign addr[4119]= 1247361445;
assign addr[4120]= 986505429;
assign addr[4121]= 705657826;
assign addr[4122]= 410510029;
assign addr[4123]= 107043224;
assign addr[4124]= -198592817;
assign addr[4125]= -500204365;
assign addr[4126]= -791679244;
assign addr[4127]= -1067110699;
assign addr[4128]= -1320917099;
assign addr[4129]= -1547955041;
assign addr[4130]= -1743623590;
assign addr[4131]= -1903957513;
assign addr[4132]= -2025707632;
assign addr[4133]= -2106406677;
assign addr[4134]= -2144419275;
assign addr[4135]= -2138975100;
assign addr[4136]= -2090184478;
assign addr[4137]= -1999036154;
assign addr[4138]= -1867377253;
assign addr[4139]= -1697875851;
assign addr[4140]= -1493966902;
assign addr[4141]= -1259782632;
assign addr[4142]= -1000068799;
assign addr[4143]= -720088517;
assign addr[4144]= -425515602;
assign addr[4145]= -122319591;
assign addr[4146]= 183355234;
assign addr[4147]= 485314355;
assign addr[4148]= 777438554;
assign addr[4149]= 1053807919;
assign addr[4150]= 1308821808;
assign addr[4151]= 1537312353;
assign addr[4152]= 1734649179;
assign addr[4153]= 1896833245;
assign addr[4154]= 2020577882;
assign addr[4155]= 2103375398;
assign addr[4156]= 2143547897;
assign addr[4157]= 2140281282;
assign addr[4158]= 2093641749;
assign addr[4159]= 2004574453;
assign addr[4160]= 1874884346;
assign addr[4161]= 1707199606;
assign addr[4162]= 1504918373;
assign addr[4163]= 1272139887;
assign addr[4164]= 1013581418;
assign addr[4165]= 734482665;
assign addr[4166]= 440499581;
assign addr[4167]= 137589750;
assign addr[4168]= -168108346;
assign addr[4169]= -470399716;
assign addr[4170]= -763158411;
assign addr[4171]= -1040451659;
assign addr[4172]= -1296660098;
assign addr[4173]= -1526591649;
assign addr[4174]= -1725586737;
assign addr[4175]= -1889612716;
assign addr[4176]= -2015345591;
assign addr[4177]= -2100237377;
assign addr[4178]= -2142567738;
assign addr[4179]= -2141478848;
assign addr[4180]= -2096992772;
assign addr[4181]= -2010011024;
assign addr[4182]= -1882296293;
assign addr[4183]= -1716436725;
assign addr[4184]= -1515793473;
assign addr[4185]= -1284432584;
assign addr[4186]= -1027042599;
assign addr[4187]= -748839539;
assign addr[4188]= -455461206;
assign addr[4189]= -152852926;
assign addr[4190]= 152852926;
assign addr[4191]= 455461206;
assign addr[4192]= 748839539;
assign addr[4193]= 1027042599;
assign addr[4194]= 1284432584;
assign addr[4195]= 1515793473;
assign addr[4196]= 1716436725;
assign addr[4197]= 1882296293;
assign addr[4198]= 2010011024;
assign addr[4199]= 2096992772;
assign addr[4200]= 2141478848;
assign addr[4201]= 2142567738;
assign addr[4202]= 2100237377;
assign addr[4203]= 2015345591;
assign addr[4204]= 1889612716;
assign addr[4205]= 1725586737;
assign addr[4206]= 1526591649;
assign addr[4207]= 1296660098;
assign addr[4208]= 1040451659;
assign addr[4209]= 763158411;
assign addr[4210]= 470399716;
assign addr[4211]= 168108346;
assign addr[4212]= -137589750;
assign addr[4213]= -440499581;
assign addr[4214]= -734482665;
assign addr[4215]= -1013581418;
assign addr[4216]= -1272139887;
assign addr[4217]= -1504918373;
assign addr[4218]= -1707199606;
assign addr[4219]= -1874884346;
assign addr[4220]= -2004574453;
assign addr[4221]= -2093641749;
assign addr[4222]= -2140281282;
assign addr[4223]= -2143547897;
assign addr[4224]= -2103375398;
assign addr[4225]= -2020577882;
assign addr[4226]= -1896833245;
assign addr[4227]= -1734649179;
assign addr[4228]= -1537312353;
assign addr[4229]= -1308821808;
assign addr[4230]= -1053807919;
assign addr[4231]= -777438554;
assign addr[4232]= -485314355;
assign addr[4233]= -183355234;
assign addr[4234]= 122319591;
assign addr[4235]= 425515602;
assign addr[4236]= 720088517;
assign addr[4237]= 1000068799;
assign addr[4238]= 1259782632;
assign addr[4239]= 1493966902;
assign addr[4240]= 1697875851;
assign addr[4241]= 1867377253;
assign addr[4242]= 1999036154;
assign addr[4243]= 2090184478;
assign addr[4244]= 2138975100;
assign addr[4245]= 2144419275;
assign addr[4246]= 2106406677;
assign addr[4247]= 2025707632;
assign addr[4248]= 1903957513;
assign addr[4249]= 1743623590;
assign addr[4250]= 1547955041;
assign addr[4251]= 1320917099;
assign addr[4252]= 1067110699;
assign addr[4253]= 791679244;
assign addr[4254]= 500204365;
assign addr[4255]= 198592817;
assign addr[4256]= -107043224;
assign addr[4257]= -410510029;
assign addr[4258]= -705657826;
assign addr[4259]= -986505429;
assign addr[4260]= -1247361445;
assign addr[4261]= -1482939614;
assign addr[4262]= -1688465931;
assign addr[4263]= -1859775393;
assign addr[4264]= -1993396407;
assign addr[4265]= -2086621133;
assign addr[4266]= -2137560369;
assign addr[4267]= -2145181827;
assign addr[4268]= -2109331059;
assign addr[4269]= -2030734582;
assign addr[4270]= -1910985158;
assign addr[4271]= -1752509516;
assign addr[4272]= -1558519173;
assign addr[4273]= -1332945355;
assign addr[4274]= -1080359326;
assign addr[4275]= -805879757;
assign addr[4276]= -515068990;
assign addr[4277]= -213820322;
assign addr[4278]= 91761426;
assign addr[4279]= 395483624;
assign addr[4280]= 691191324;
assign addr[4281]= 972891995;
assign addr[4282]= 1234876957;
assign addr[4283]= 1471837070;
assign addr[4284]= 1678970324;
assign addr[4285]= 1852079154;
assign addr[4286]= 1987655498;
assign addr[4287]= 2082951896;
assign addr[4288]= 2136037160;
assign addr[4289]= 2145835515;
assign addr[4290]= 2112148396;
assign addr[4291]= 2035658475;
assign addr[4292]= 1917915825;
assign addr[4293]= 1761306505;
assign addr[4294]= 1569004214;
assign addr[4295]= 1344905966;
assign addr[4296]= 1093553126;
assign addr[4297]= 820039373;
assign addr[4298]= 529907477;
assign addr[4299]= 229036977;
assign addr[4300]= -76474970;
assign addr[4301]= -380437148;
assign addr[4302]= -676689746;
assign addr[4303]= -959229189;
assign addr[4304]= -1222329801;
assign addr[4305]= -1460659832;
assign addr[4306]= -1669389513;
assign addr[4307]= -1844288924;
assign addr[4308]= -1981813720;
assign addr[4309]= -2079176953;
assign addr[4310]= -2134405552;
assign addr[4311]= -2146380306;
assign addr[4312]= -2114858546;
assign addr[4313]= -2040479063;
assign addr[4314]= -1924749160;
assign addr[4315]= -1770014111;
assign addr[4316]= -1579409630;
assign addr[4317]= -1356798326;
assign addr[4318]= -1106691431;
assign addr[4319]= -834157373;
assign addr[4320]= -544719071;
assign addr[4321]= -244242007;
assign addr[4322]= 61184634;
assign addr[4323]= 365371365;
assign addr[4324]= 662153826;
assign addr[4325]= 945517704;
assign addr[4326]= 1209720613;
assign addr[4327]= 1449408469;
assign addr[4328]= 1659723983;
assign addr[4329]= 1836405100;
assign addr[4330]= 1975871368;
assign addr[4331]= 2075296495;
assign addr[4332]= 2132665626;
assign addr[4333]= 2146816171;
assign addr[4334]= 2117461370;
assign addr[4335]= 2045196100;
assign addr[4336]= 1931484818;
assign addr[4337]= 1778631892;
assign addr[4338]= 1589734894;
assign addr[4339]= 1368621831;
assign addr[4340]= 1119773573;
assign addr[4341]= 848233042;
assign addr[4342]= 559503022;
assign addr[4343]= 259434643;
assign addr[4344]= -45891193;
assign addr[4345]= -350287041;
assign addr[4346]= -647584304;
assign addr[4347]= -931758235;
assign addr[4348]= -1197050035;
assign addr[4349]= -1438083551;
assign addr[4350]= -1649974225;
assign addr[4351]= -1828428082;
assign addr[4352]= -1969828744;
assign addr[4353]= -2071310720;
assign addr[4354]= -2130817471;
assign addr[4355]= -2147143090;
assign addr[4356]= -2119956737;
assign addr[4357]= -2049809346;
assign addr[4358]= -1938122457;
assign addr[4359]= -1787159411;
assign addr[4360]= -1599979481;
assign addr[4361]= -1380375881;
assign addr[4362]= -1132798888;
assign addr[4363]= -862265664;
assign addr[4364]= -574258580;
assign addr[4365]= -274614114;
assign addr[4366]= 30595422;
assign addr[4367]= 335184940;
assign addr[4368]= 632981917;
assign addr[4369]= 917951481;
assign addr[4370]= 1184318708;
assign addr[4371]= 1426685652;
assign addr[4372]= 1640140734;
assign addr[4373]= 1820358275;
assign addr[4374]= 1963686155;
assign addr[4375]= 2067219829;
assign addr[4376]= 2128861181;
assign addr[4377]= 2147361045;
assign addr[4378]= 2122344521;
assign addr[4379]= 2054318569;
assign addr[4380]= 1944661739;
assign addr[4381]= 1795596234;
assign addr[4382]= 1610142873;
assign addr[4383]= 1392059879;
assign addr[4384]= 1145766716;
assign addr[4385]= 876254528;
assign addr[4386]= 588984994;
assign addr[4387]= 289779648;
assign addr[4388]= -15298099;
assign addr[4389]= -320065829;
assign addr[4390]= -618347408;
assign addr[4391]= -904098143;
assign addr[4392]= -1171527280;
assign addr[4393]= -1415215352;
assign addr[4394]= -1630224009;
assign addr[4395]= -1812196087;
assign addr[4396]= -1957443913;
assign addr[4397]= -2063024031;
assign addr[4398]= -2126796855;
assign addr[4399]= -2147470025;
assign addr[4400]= -2124624598;
assign addr[4401]= -2058723538;
assign addr[4402]= -1951102334;
assign addr[4403]= -1803941934;
assign addr[4404]= -1620224553;
assign addr[4405]= -1403673233;
assign addr[4406]= -1158676398;
assign addr[4407]= -890198924;
assign addr[4408]= -603681519;
assign addr[4409]= -304930476;
assign addr[4410]= 0;
assign addr[4411]= 304930476;
assign addr[4412]= 603681519;
assign addr[4413]= 890198924;
assign addr[4414]= 1158676398;
assign addr[4415]= 1403673233;
assign addr[4416]= 1620224553;
assign addr[4417]= 1803941934;
assign addr[4418]= 1951102334;
assign addr[4419]= 2058723538;
assign addr[4420]= 2124624598;
assign addr[4421]= 2147470025;
assign addr[4422]= 2126796855;
assign addr[4423]= 2063024031;
assign addr[4424]= 1957443913;
assign addr[4425]= 1812196087;
assign addr[4426]= 1630224009;
assign addr[4427]= 1415215352;
assign addr[4428]= 1171527280;
assign addr[4429]= 904098143;
assign addr[4430]= 618347408;
assign addr[4431]= 320065829;
assign addr[4432]= 15298099;
assign addr[4433]= -289779648;
assign addr[4434]= -588984994;
assign addr[4435]= -876254528;
assign addr[4436]= -1145766716;
assign addr[4437]= -1392059879;
assign addr[4438]= -1610142873;
assign addr[4439]= -1795596234;
assign addr[4440]= -1944661739;
assign addr[4441]= -2054318569;
assign addr[4442]= -2122344521;
assign addr[4443]= -2147361045;
assign addr[4444]= -2128861181;
assign addr[4445]= -2067219829;
assign addr[4446]= -1963686155;
assign addr[4447]= -1820358275;
assign addr[4448]= -1640140734;
assign addr[4449]= -1426685652;
assign addr[4450]= -1184318708;
assign addr[4451]= -917951481;
assign addr[4452]= -632981917;
assign addr[4453]= -335184940;
assign addr[4454]= -30595422;
assign addr[4455]= 274614114;
assign addr[4456]= 574258580;
assign addr[4457]= 862265664;
assign addr[4458]= 1132798888;
assign addr[4459]= 1380375881;
assign addr[4460]= 1599979481;
assign addr[4461]= 1787159411;
assign addr[4462]= 1938122457;
assign addr[4463]= 2049809346;
assign addr[4464]= 2119956737;
assign addr[4465]= 2147143090;
assign addr[4466]= 2130817471;
assign addr[4467]= 2071310720;
assign addr[4468]= 1969828744;
assign addr[4469]= 1828428082;
assign addr[4470]= 1649974225;
assign addr[4471]= 1438083551;
assign addr[4472]= 1197050035;
assign addr[4473]= 931758235;
assign addr[4474]= 647584304;
assign addr[4475]= 350287041;
assign addr[4476]= 45891193;
assign addr[4477]= -259434643;
assign addr[4478]= -559503022;
assign addr[4479]= -848233042;
assign addr[4480]= -1119773573;
assign addr[4481]= -1368621831;
assign addr[4482]= -1589734894;
assign addr[4483]= -1778631892;
assign addr[4484]= -1931484818;
assign addr[4485]= -2045196100;
assign addr[4486]= -2117461370;
assign addr[4487]= -2146816171;
assign addr[4488]= -2132665626;
assign addr[4489]= -2075296495;
assign addr[4490]= -1975871368;
assign addr[4491]= -1836405100;
assign addr[4492]= -1659723983;
assign addr[4493]= -1449408469;
assign addr[4494]= -1209720613;
assign addr[4495]= -945517704;
assign addr[4496]= -662153826;
assign addr[4497]= -365371365;
assign addr[4498]= -61184634;
assign addr[4499]= 244242007;
assign addr[4500]= 544719071;
assign addr[4501]= 834157373;
assign addr[4502]= 1106691431;
assign addr[4503]= 1356798326;
assign addr[4504]= 1579409630;
assign addr[4505]= 1770014111;
assign addr[4506]= 1924749160;
assign addr[4507]= 2040479063;
assign addr[4508]= 2114858546;
assign addr[4509]= 2146380306;
assign addr[4510]= 2134405552;
assign addr[4511]= 2079176953;
assign addr[4512]= 1981813720;
assign addr[4513]= 1844288924;
assign addr[4514]= 1669389513;
assign addr[4515]= 1460659832;
assign addr[4516]= 1222329801;
assign addr[4517]= 959229189;
assign addr[4518]= 676689746;
assign addr[4519]= 380437148;
assign addr[4520]= 76474970;
assign addr[4521]= -229036977;
assign addr[4522]= -529907477;
assign addr[4523]= -820039373;
assign addr[4524]= -1093553126;
assign addr[4525]= -1344905966;
assign addr[4526]= -1569004214;
assign addr[4527]= -1761306505;
assign addr[4528]= -1917915825;
assign addr[4529]= -2035658475;
assign addr[4530]= -2112148396;
assign addr[4531]= -2145835515;
assign addr[4532]= -2136037160;
assign addr[4533]= -2082951896;
assign addr[4534]= -1987655498;
assign addr[4535]= -1852079154;
assign addr[4536]= -1678970324;
assign addr[4537]= -1471837070;
assign addr[4538]= -1234876957;
assign addr[4539]= -972891995;
assign addr[4540]= -691191324;
assign addr[4541]= -395483624;
assign addr[4542]= -91761426;
assign addr[4543]= 213820322;
assign addr[4544]= 515068990;
assign addr[4545]= 805879757;
assign addr[4546]= 1080359326;
assign addr[4547]= 1332945355;
assign addr[4548]= 1558519173;
assign addr[4549]= 1752509516;
assign addr[4550]= 1910985158;
assign addr[4551]= 2030734582;
assign addr[4552]= 2109331059;
assign addr[4553]= 2145181827;
assign addr[4554]= 2137560369;
assign addr[4555]= 2086621133;
assign addr[4556]= 1993396407;
assign addr[4557]= 1859775393;
assign addr[4558]= 1688465931;
assign addr[4559]= 1482939614;
assign addr[4560]= 1247361445;
assign addr[4561]= 986505429;
assign addr[4562]= 705657826;
assign addr[4563]= 410510029;
assign addr[4564]= 107043224;
assign addr[4565]= -198592817;
assign addr[4566]= -500204365;
assign addr[4567]= -791679244;
assign addr[4568]= -1067110699;
assign addr[4569]= -1320917099;
assign addr[4570]= -1547955041;
assign addr[4571]= -1743623590;
assign addr[4572]= -1903957513;
assign addr[4573]= -2025707632;
assign addr[4574]= -2106406677;
assign addr[4575]= -2144419275;
assign addr[4576]= -2138975100;
assign addr[4577]= -2090184478;
assign addr[4578]= -1999036154;
assign addr[4579]= -1867377253;
assign addr[4580]= -1697875851;
assign addr[4581]= -1493966902;
assign addr[4582]= -1259782632;
assign addr[4583]= -1000068799;
assign addr[4584]= -720088517;
assign addr[4585]= -425515602;
assign addr[4586]= -122319591;
assign addr[4587]= 183355234;
assign addr[4588]= 485314355;
assign addr[4589]= 777438554;
assign addr[4590]= 1053807919;
assign addr[4591]= 1308821808;
assign addr[4592]= 1537312353;
assign addr[4593]= 1734649179;
assign addr[4594]= 1896833245;
assign addr[4595]= 2020577882;
assign addr[4596]= 2103375398;
assign addr[4597]= 2143547897;
assign addr[4598]= 2140281282;
assign addr[4599]= 2093641749;
assign addr[4600]= 2004574453;
assign addr[4601]= 1874884346;
assign addr[4602]= 1707199606;
assign addr[4603]= 1504918373;
assign addr[4604]= 1272139887;
assign addr[4605]= 1013581418;
assign addr[4606]= 734482665;
assign addr[4607]= 440499581;
assign addr[4608]= 137589750;
assign addr[4609]= -168108346;
assign addr[4610]= -470399716;
assign addr[4611]= -763158411;
assign addr[4612]= -1040451659;
assign addr[4613]= -1296660098;
assign addr[4614]= -1526591649;
assign addr[4615]= -1725586737;
assign addr[4616]= -1889612716;
assign addr[4617]= -2015345591;
assign addr[4618]= -2100237377;
assign addr[4619]= -2142567738;
assign addr[4620]= -2141478848;
assign addr[4621]= -2096992772;
assign addr[4622]= -2010011024;
assign addr[4623]= -1882296293;
assign addr[4624]= -1716436725;
assign addr[4625]= -1515793473;
assign addr[4626]= -1284432584;
assign addr[4627]= -1027042599;
assign addr[4628]= -748839539;
assign addr[4629]= -455461206;
assign addr[4630]= -152852926;
assign addr[4631]= 152852926;
assign addr[4632]= 455461206;
assign addr[4633]= 748839539;
assign addr[4634]= 1027042599;
assign addr[4635]= 1284432584;
assign addr[4636]= 1515793473;
assign addr[4637]= 1716436725;
assign addr[4638]= 1882296293;
assign addr[4639]= 2010011024;
assign addr[4640]= 2096992772;
assign addr[4641]= 2141478848;
assign addr[4642]= 2142567738;
assign addr[4643]= 2100237377;
assign addr[4644]= 2015345591;
assign addr[4645]= 1889612716;
assign addr[4646]= 1725586737;
assign addr[4647]= 1526591649;
assign addr[4648]= 1296660098;
assign addr[4649]= 1040451659;
assign addr[4650]= 763158411;
assign addr[4651]= 470399716;
assign addr[4652]= 168108346;
assign addr[4653]= -137589750;
assign addr[4654]= -440499581;
assign addr[4655]= -734482665;
assign addr[4656]= -1013581418;
assign addr[4657]= -1272139887;
assign addr[4658]= -1504918373;
assign addr[4659]= -1707199606;
assign addr[4660]= -1874884346;
assign addr[4661]= -2004574453;
assign addr[4662]= -2093641749;
assign addr[4663]= -2140281282;
assign addr[4664]= -2143547897;
assign addr[4665]= -2103375398;
assign addr[4666]= -2020577882;
assign addr[4667]= -1896833245;
assign addr[4668]= -1734649179;
assign addr[4669]= -1537312353;
assign addr[4670]= -1308821808;
assign addr[4671]= -1053807919;
assign addr[4672]= -777438554;
assign addr[4673]= -485314355;
assign addr[4674]= -183355234;
assign addr[4675]= 122319591;
assign addr[4676]= 425515602;
assign addr[4677]= 720088517;
assign addr[4678]= 1000068799;
assign addr[4679]= 1259782632;
assign addr[4680]= 1493966902;
assign addr[4681]= 1697875851;
assign addr[4682]= 1867377253;
assign addr[4683]= 1999036154;
assign addr[4684]= 2090184478;
assign addr[4685]= 2138975100;
assign addr[4686]= 2144419275;
assign addr[4687]= 2106406677;
assign addr[4688]= 2025707632;
assign addr[4689]= 1903957513;
assign addr[4690]= 1743623590;
assign addr[4691]= 1547955041;
assign addr[4692]= 1320917099;
assign addr[4693]= 1067110699;
assign addr[4694]= 791679244;
assign addr[4695]= 500204365;
assign addr[4696]= 198592817;
assign addr[4697]= -107043224;
assign addr[4698]= -410510029;
assign addr[4699]= -705657826;
assign addr[4700]= -986505429;
assign addr[4701]= -1247361445;
assign addr[4702]= -1482939614;
assign addr[4703]= -1688465931;
assign addr[4704]= -1859775393;
assign addr[4705]= -1993396407;
assign addr[4706]= -2086621133;
assign addr[4707]= -2137560369;
assign addr[4708]= -2145181827;
assign addr[4709]= -2109331059;
assign addr[4710]= -2030734582;
assign addr[4711]= -1910985158;
assign addr[4712]= -1752509516;
assign addr[4713]= -1558519173;
assign addr[4714]= -1332945355;
assign addr[4715]= -1080359326;
assign addr[4716]= -805879757;
assign addr[4717]= -515068990;
assign addr[4718]= -213820322;
assign addr[4719]= 91761426;
assign addr[4720]= 395483624;
assign addr[4721]= 691191324;
assign addr[4722]= 972891995;
assign addr[4723]= 1234876957;
assign addr[4724]= 1471837070;
assign addr[4725]= 1678970324;
assign addr[4726]= 1852079154;
assign addr[4727]= 1987655498;
assign addr[4728]= 2082951896;
assign addr[4729]= 2136037160;
assign addr[4730]= 2145835515;
assign addr[4731]= 2112148396;
assign addr[4732]= 2035658475;
assign addr[4733]= 1917915825;
assign addr[4734]= 1761306505;
assign addr[4735]= 1569004214;
assign addr[4736]= 1344905966;
assign addr[4737]= 1093553126;
assign addr[4738]= 820039373;
assign addr[4739]= 529907477;
assign addr[4740]= 229036977;
assign addr[4741]= -76474970;
assign addr[4742]= -380437148;
assign addr[4743]= -676689746;
assign addr[4744]= -959229189;
assign addr[4745]= -1222329801;
assign addr[4746]= -1460659832;
assign addr[4747]= -1669389513;
assign addr[4748]= -1844288924;
assign addr[4749]= -1981813720;
assign addr[4750]= -2079176953;
assign addr[4751]= -2134405552;
assign addr[4752]= -2146380306;
assign addr[4753]= -2114858546;
assign addr[4754]= -2040479063;
assign addr[4755]= -1924749160;
assign addr[4756]= -1770014111;
assign addr[4757]= -1579409630;
assign addr[4758]= -1356798326;
assign addr[4759]= -1106691431;
assign addr[4760]= -834157373;
assign addr[4761]= -544719071;
assign addr[4762]= -244242007;
assign addr[4763]= 61184634;
assign addr[4764]= 365371365;
assign addr[4765]= 662153826;
assign addr[4766]= 945517704;
assign addr[4767]= 1209720613;
assign addr[4768]= 1449408469;
assign addr[4769]= 1659723983;
assign addr[4770]= 1836405100;
assign addr[4771]= 1975871368;
assign addr[4772]= 2075296495;
assign addr[4773]= 2132665626;
assign addr[4774]= 2146816171;
assign addr[4775]= 2117461370;
assign addr[4776]= 2045196100;
assign addr[4777]= 1931484818;
assign addr[4778]= 1778631892;
assign addr[4779]= 1589734894;
assign addr[4780]= 1368621831;
assign addr[4781]= 1119773573;
assign addr[4782]= 848233042;
assign addr[4783]= 559503022;
assign addr[4784]= 259434643;
assign addr[4785]= -45891193;
assign addr[4786]= -350287041;
assign addr[4787]= -647584304;
assign addr[4788]= -931758235;
assign addr[4789]= -1197050035;
assign addr[4790]= -1438083551;
assign addr[4791]= -1649974225;
assign addr[4792]= -1828428082;
assign addr[4793]= -1969828744;
assign addr[4794]= -2071310720;
assign addr[4795]= -2130817471;
assign addr[4796]= -2147143090;
assign addr[4797]= -2119956737;
assign addr[4798]= -2049809346;
assign addr[4799]= -1938122457;
assign addr[4800]= -1787159411;
assign addr[4801]= -1599979481;
assign addr[4802]= -1380375881;
assign addr[4803]= -1132798888;
assign addr[4804]= -862265664;
assign addr[4805]= -574258580;
assign addr[4806]= -274614114;
assign addr[4807]= 30595422;
assign addr[4808]= 335184940;
assign addr[4809]= 632981917;
assign addr[4810]= 917951481;
assign addr[4811]= 1184318708;
assign addr[4812]= 1426685652;
assign addr[4813]= 1640140734;
assign addr[4814]= 1820358275;
assign addr[4815]= 1963686155;
assign addr[4816]= 2067219829;
assign addr[4817]= 2128861181;
assign addr[4818]= 2147361045;
assign addr[4819]= 2122344521;
assign addr[4820]= 2054318569;
assign addr[4821]= 1944661739;
assign addr[4822]= 1795596234;
assign addr[4823]= 1610142873;
assign addr[4824]= 1392059879;
assign addr[4825]= 1145766716;
assign addr[4826]= 876254528;
assign addr[4827]= 588984994;
assign addr[4828]= 289779648;
assign addr[4829]= -15298099;
assign addr[4830]= -320065829;
assign addr[4831]= -618347408;
assign addr[4832]= -904098143;
assign addr[4833]= -1171527280;
assign addr[4834]= -1415215352;
assign addr[4835]= -1630224009;
assign addr[4836]= -1812196087;
assign addr[4837]= -1957443913;
assign addr[4838]= -2063024031;
assign addr[4839]= -2126796855;
assign addr[4840]= -2147470025;
assign addr[4841]= -2124624598;
assign addr[4842]= -2058723538;
assign addr[4843]= -1951102334;
assign addr[4844]= -1803941934;
assign addr[4845]= -1620224553;
assign addr[4846]= -1403673233;
assign addr[4847]= -1158676398;
assign addr[4848]= -890198924;
assign addr[4849]= -603681519;
assign addr[4850]= -304930476;
assign addr[4851]= 0;
assign addr[4852]= 304930476;
assign addr[4853]= 603681519;
assign addr[4854]= 890198924;
assign addr[4855]= 1158676398;
assign addr[4856]= 1403673233;
assign addr[4857]= 1620224553;
assign addr[4858]= 1803941934;
assign addr[4859]= 1951102334;
assign addr[4860]= 2058723538;
assign addr[4861]= 2124624598;
assign addr[4862]= 2147470025;
assign addr[4863]= 2126796855;
assign addr[4864]= 2063024031;
assign addr[4865]= 1957443913;
assign addr[4866]= 1812196087;
assign addr[4867]= 1630224009;
assign addr[4868]= 1415215352;
assign addr[4869]= 1171527280;
assign addr[4870]= 904098143;
assign addr[4871]= 618347408;
assign addr[4872]= 320065829;
assign addr[4873]= 15298099;
assign addr[4874]= -289779648;
assign addr[4875]= -588984994;
assign addr[4876]= -876254528;
assign addr[4877]= -1145766716;
assign addr[4878]= -1392059879;
assign addr[4879]= -1610142873;
assign addr[4880]= -1795596234;
assign addr[4881]= -1944661739;
assign addr[4882]= -2054318569;
assign addr[4883]= -2122344521;
assign addr[4884]= -2147361045;
assign addr[4885]= -2128861181;
assign addr[4886]= -2067219829;
assign addr[4887]= -1963686155;
assign addr[4888]= -1820358275;
assign addr[4889]= -1640140734;
assign addr[4890]= -1426685652;
assign addr[4891]= -1184318708;
assign addr[4892]= -917951481;
assign addr[4893]= -632981917;
assign addr[4894]= -335184940;
assign addr[4895]= -30595422;
assign addr[4896]= 274614114;
assign addr[4897]= 574258580;
assign addr[4898]= 862265664;
assign addr[4899]= 1132798888;
assign addr[4900]= 1380375881;
assign addr[4901]= 1599979481;
assign addr[4902]= 1787159411;
assign addr[4903]= 1938122457;
assign addr[4904]= 2049809346;
assign addr[4905]= 2119956737;
assign addr[4906]= 2147143090;
assign addr[4907]= 2130817471;
assign addr[4908]= 2071310720;
assign addr[4909]= 1969828744;
assign addr[4910]= 1828428082;
assign addr[4911]= 1649974225;
assign addr[4912]= 1438083551;
assign addr[4913]= 1197050035;
assign addr[4914]= 931758235;
assign addr[4915]= 647584304;
assign addr[4916]= 350287041;
assign addr[4917]= 45891193;
assign addr[4918]= -259434643;
assign addr[4919]= -559503022;
assign addr[4920]= -848233042;
assign addr[4921]= -1119773573;
assign addr[4922]= -1368621831;
assign addr[4923]= -1589734894;
assign addr[4924]= -1778631892;
assign addr[4925]= -1931484818;
assign addr[4926]= -2045196100;
assign addr[4927]= -2117461370;
assign addr[4928]= -2146816171;
assign addr[4929]= -2132665626;
assign addr[4930]= -2075296495;
assign addr[4931]= -1975871368;
assign addr[4932]= -1836405100;
assign addr[4933]= -1659723983;
assign addr[4934]= -1449408469;
assign addr[4935]= -1209720613;
assign addr[4936]= -945517704;
assign addr[4937]= -662153826;
assign addr[4938]= -365371365;
assign addr[4939]= -61184634;
assign addr[4940]= 244242007;
assign addr[4941]= 544719071;
assign addr[4942]= 834157373;
assign addr[4943]= 1106691431;
assign addr[4944]= 1356798326;
assign addr[4945]= 1579409630;
assign addr[4946]= 1770014111;
assign addr[4947]= 1924749160;
assign addr[4948]= 2040479063;
assign addr[4949]= 2114858546;
assign addr[4950]= 2146380306;
assign addr[4951]= 2134405552;
assign addr[4952]= 2079176953;
assign addr[4953]= 1981813720;
assign addr[4954]= 1844288924;
assign addr[4955]= 1669389513;
assign addr[4956]= 1460659832;
assign addr[4957]= 1222329801;
assign addr[4958]= 959229189;
assign addr[4959]= 676689746;
assign addr[4960]= 380437148;
assign addr[4961]= 76474970;
assign addr[4962]= -229036977;
assign addr[4963]= -529907477;
assign addr[4964]= -820039373;
assign addr[4965]= -1093553126;
assign addr[4966]= -1344905966;
assign addr[4967]= -1569004214;
assign addr[4968]= -1761306505;
assign addr[4969]= -1917915825;
assign addr[4970]= -2035658475;
assign addr[4971]= -2112148396;
assign addr[4972]= -2145835515;
assign addr[4973]= -2136037160;
assign addr[4974]= -2082951896;
assign addr[4975]= -1987655498;
assign addr[4976]= -1852079154;
assign addr[4977]= -1678970324;
assign addr[4978]= -1471837070;
assign addr[4979]= -1234876957;
assign addr[4980]= -972891995;
assign addr[4981]= -691191324;
assign addr[4982]= -395483624;
assign addr[4983]= -91761426;
assign addr[4984]= 213820322;
assign addr[4985]= 515068990;
assign addr[4986]= 805879757;
assign addr[4987]= 1080359326;
assign addr[4988]= 1332945355;
assign addr[4989]= 1558519173;
assign addr[4990]= 1752509516;
assign addr[4991]= 1910985158;
assign addr[4992]= 2030734582;
assign addr[4993]= 2109331059;
assign addr[4994]= 2145181827;
assign addr[4995]= 2137560369;
assign addr[4996]= 2086621133;
assign addr[4997]= 1993396407;
assign addr[4998]= 1859775393;
assign addr[4999]= 1688465931;
assign addr[5000]= 1482939614;
assign addr[5001]= 1247361445;
assign addr[5002]= 986505429;
assign addr[5003]= 705657826;
assign addr[5004]= 410510029;
assign addr[5005]= 107043224;
assign addr[5006]= -198592817;
assign addr[5007]= -500204365;
assign addr[5008]= -791679244;
assign addr[5009]= -1067110699;
assign addr[5010]= -1320917099;
assign addr[5011]= -1547955041;
assign addr[5012]= -1743623590;
assign addr[5013]= -1903957513;
assign addr[5014]= -2025707632;
assign addr[5015]= -2106406677;
assign addr[5016]= -2144419275;
assign addr[5017]= -2138975100;
assign addr[5018]= -2090184478;
assign addr[5019]= -1999036154;
assign addr[5020]= -1867377253;
assign addr[5021]= -1697875851;
assign addr[5022]= -1493966902;
assign addr[5023]= -1259782632;
assign addr[5024]= -1000068799;
assign addr[5025]= -720088517;
assign addr[5026]= -425515602;
assign addr[5027]= -122319591;
assign addr[5028]= 183355234;
assign addr[5029]= 485314355;
assign addr[5030]= 777438554;
assign addr[5031]= 1053807919;
assign addr[5032]= 1308821808;
assign addr[5033]= 1537312353;
assign addr[5034]= 1734649179;
assign addr[5035]= 1896833245;
assign addr[5036]= 2020577882;
assign addr[5037]= 2103375398;
assign addr[5038]= 2143547897;
assign addr[5039]= 2140281282;
assign addr[5040]= 2093641749;
assign addr[5041]= 2004574453;
assign addr[5042]= 1874884346;
assign addr[5043]= 1707199606;
assign addr[5044]= 1504918373;
assign addr[5045]= 1272139887;
assign addr[5046]= 1013581418;
assign addr[5047]= 734482665;
assign addr[5048]= 440499581;
assign addr[5049]= 137589750;
assign addr[5050]= -168108346;
assign addr[5051]= -470399716;
assign addr[5052]= -763158411;
assign addr[5053]= -1040451659;
assign addr[5054]= -1296660098;
assign addr[5055]= -1526591649;
assign addr[5056]= -1725586737;
assign addr[5057]= -1889612716;
assign addr[5058]= -2015345591;
assign addr[5059]= -2100237377;
assign addr[5060]= -2142567738;
assign addr[5061]= -2141478848;
assign addr[5062]= -2096992772;
assign addr[5063]= -2010011024;
assign addr[5064]= -1882296293;
assign addr[5065]= -1716436725;
assign addr[5066]= -1515793473;
assign addr[5067]= -1284432584;
assign addr[5068]= -1027042599;
assign addr[5069]= -748839539;
assign addr[5070]= -455461206;
assign addr[5071]= -152852926;
assign addr[5072]= 152852926;
assign addr[5073]= 455461206;
assign addr[5074]= 748839539;
assign addr[5075]= 1027042599;
assign addr[5076]= 1284432584;
assign addr[5077]= 1515793473;
assign addr[5078]= 1716436725;
assign addr[5079]= 1882296293;
assign addr[5080]= 2010011024;
assign addr[5081]= 2096992772;
assign addr[5082]= 2141478848;
assign addr[5083]= 2142567738;
assign addr[5084]= 2100237377;
assign addr[5085]= 2015345591;
assign addr[5086]= 1889612716;
assign addr[5087]= 1725586737;
assign addr[5088]= 1526591649;
assign addr[5089]= 1296660098;
assign addr[5090]= 1040451659;
assign addr[5091]= 763158411;
assign addr[5092]= 470399716;
assign addr[5093]= 168108346;
assign addr[5094]= -137589750;
assign addr[5095]= -440499581;
assign addr[5096]= -734482665;
assign addr[5097]= -1013581418;
assign addr[5098]= -1272139887;
assign addr[5099]= -1504918373;
assign addr[5100]= -1707199606;
assign addr[5101]= -1874884346;
assign addr[5102]= -2004574453;
assign addr[5103]= -2093641749;
assign addr[5104]= -2140281282;
assign addr[5105]= -2143547897;
assign addr[5106]= -2103375398;
assign addr[5107]= -2020577882;
assign addr[5108]= -1896833245;
assign addr[5109]= -1734649179;
assign addr[5110]= -1537312353;
assign addr[5111]= -1308821808;
assign addr[5112]= -1053807919;
assign addr[5113]= -777438554;
assign addr[5114]= -485314355;
assign addr[5115]= -183355234;
assign addr[5116]= 122319591;
assign addr[5117]= 425515602;
assign addr[5118]= 720088517;
assign addr[5119]= 1000068799;
assign addr[5120]= 1259782632;
assign addr[5121]= 1493966902;
assign addr[5122]= 1697875851;
assign addr[5123]= 1867377253;
assign addr[5124]= 1999036154;
assign addr[5125]= 2090184478;
assign addr[5126]= 2138975100;
assign addr[5127]= 2144419275;
assign addr[5128]= 2106406677;
assign addr[5129]= 2025707632;
assign addr[5130]= 1903957513;
assign addr[5131]= 1743623590;
assign addr[5132]= 1547955041;
assign addr[5133]= 1320917099;
assign addr[5134]= 1067110699;
assign addr[5135]= 791679244;
assign addr[5136]= 500204365;
assign addr[5137]= 198592817;
assign addr[5138]= -107043224;
assign addr[5139]= -410510029;
assign addr[5140]= -705657826;
assign addr[5141]= -986505429;
assign addr[5142]= -1247361445;
assign addr[5143]= -1482939614;
assign addr[5144]= -1688465931;
assign addr[5145]= -1859775393;
assign addr[5146]= -1993396407;
assign addr[5147]= -2086621133;
assign addr[5148]= -2137560369;
assign addr[5149]= -2145181827;
assign addr[5150]= -2109331059;
assign addr[5151]= -2030734582;
assign addr[5152]= -1910985158;
assign addr[5153]= -1752509516;
assign addr[5154]= -1558519173;
assign addr[5155]= -1332945355;
assign addr[5156]= -1080359326;
assign addr[5157]= -805879757;
assign addr[5158]= -515068990;
assign addr[5159]= -213820322;
assign addr[5160]= 91761426;
assign addr[5161]= 395483624;
assign addr[5162]= 691191324;
assign addr[5163]= 972891995;
assign addr[5164]= 1234876957;
assign addr[5165]= 1471837070;
assign addr[5166]= 1678970324;
assign addr[5167]= 1852079154;
assign addr[5168]= 1987655498;
assign addr[5169]= 2082951896;
assign addr[5170]= 2136037160;
assign addr[5171]= 2145835515;
assign addr[5172]= 2112148396;
assign addr[5173]= 2035658475;
assign addr[5174]= 1917915825;
assign addr[5175]= 1761306505;
assign addr[5176]= 1569004214;
assign addr[5177]= 1344905966;
assign addr[5178]= 1093553126;
assign addr[5179]= 820039373;
assign addr[5180]= 529907477;
assign addr[5181]= 229036977;
assign addr[5182]= -76474970;
assign addr[5183]= -380437148;
assign addr[5184]= -676689746;
assign addr[5185]= -959229189;
assign addr[5186]= -1222329801;
assign addr[5187]= -1460659832;
assign addr[5188]= -1669389513;
assign addr[5189]= -1844288924;
assign addr[5190]= -1981813720;
assign addr[5191]= -2079176953;
assign addr[5192]= -2134405552;
assign addr[5193]= -2146380306;
assign addr[5194]= -2114858546;
assign addr[5195]= -2040479063;
assign addr[5196]= -1924749160;
assign addr[5197]= -1770014111;
assign addr[5198]= -1579409630;
assign addr[5199]= -1356798326;
assign addr[5200]= -1106691431;
assign addr[5201]= -834157373;
assign addr[5202]= -544719071;
assign addr[5203]= -244242007;
assign addr[5204]= 61184634;
assign addr[5205]= 365371365;
assign addr[5206]= 662153826;
assign addr[5207]= 945517704;
assign addr[5208]= 1209720613;
assign addr[5209]= 1449408469;
assign addr[5210]= 1659723983;
assign addr[5211]= 1836405100;
assign addr[5212]= 1975871368;
assign addr[5213]= 2075296495;
assign addr[5214]= 2132665626;
assign addr[5215]= 2146816171;
assign addr[5216]= 2117461370;
assign addr[5217]= 2045196100;
assign addr[5218]= 1931484818;
assign addr[5219]= 1778631892;
assign addr[5220]= 1589734894;
assign addr[5221]= 1368621831;
assign addr[5222]= 1119773573;
assign addr[5223]= 848233042;
assign addr[5224]= 559503022;
assign addr[5225]= 259434643;
assign addr[5226]= -45891193;
assign addr[5227]= -350287041;
assign addr[5228]= -647584304;
assign addr[5229]= -931758235;
assign addr[5230]= -1197050035;
assign addr[5231]= -1438083551;
assign addr[5232]= -1649974225;
assign addr[5233]= -1828428082;
assign addr[5234]= -1969828744;
assign addr[5235]= -2071310720;
assign addr[5236]= -2130817471;
assign addr[5237]= -2147143090;
assign addr[5238]= -2119956737;
assign addr[5239]= -2049809346;
assign addr[5240]= -1938122457;
assign addr[5241]= -1787159411;
assign addr[5242]= -1599979481;
assign addr[5243]= -1380375881;
assign addr[5244]= -1132798888;
assign addr[5245]= -862265664;
assign addr[5246]= -574258580;
assign addr[5247]= -274614114;
assign addr[5248]= 30595422;
assign addr[5249]= 335184940;
assign addr[5250]= 632981917;
assign addr[5251]= 917951481;
assign addr[5252]= 1184318708;
assign addr[5253]= 1426685652;
assign addr[5254]= 1640140734;
assign addr[5255]= 1820358275;
assign addr[5256]= 1963686155;
assign addr[5257]= 2067219829;
assign addr[5258]= 2128861181;
assign addr[5259]= 2147361045;
assign addr[5260]= 2122344521;
assign addr[5261]= 2054318569;
assign addr[5262]= 1944661739;
assign addr[5263]= 1795596234;
assign addr[5264]= 1610142873;
assign addr[5265]= 1392059879;
assign addr[5266]= 1145766716;
assign addr[5267]= 876254528;
assign addr[5268]= 588984994;
assign addr[5269]= 289779648;
assign addr[5270]= -15298099;
assign addr[5271]= -320065829;
assign addr[5272]= -618347408;
assign addr[5273]= -904098143;
assign addr[5274]= -1171527280;
assign addr[5275]= -1415215352;
assign addr[5276]= -1630224009;
assign addr[5277]= -1812196087;
assign addr[5278]= -1957443913;
assign addr[5279]= -2063024031;
assign addr[5280]= -2126796855;
assign addr[5281]= -2147470025;
assign addr[5282]= -2124624598;
assign addr[5283]= -2058723538;
assign addr[5284]= -1951102334;
assign addr[5285]= -1803941934;
assign addr[5286]= -1620224553;
assign addr[5287]= -1403673233;
assign addr[5288]= -1158676398;
assign addr[5289]= -890198924;
assign addr[5290]= -603681519;
assign addr[5291]= -304930476;
assign addr[5292]= 0;
assign addr[5293]= 304930476;
assign addr[5294]= 603681519;
assign addr[5295]= 890198924;
assign addr[5296]= 1158676398;
assign addr[5297]= 1403673233;
assign addr[5298]= 1620224553;
assign addr[5299]= 1803941934;
assign addr[5300]= 1951102334;
assign addr[5301]= 2058723538;
assign addr[5302]= 2124624598;
assign addr[5303]= 2147470025;
assign addr[5304]= 2126796855;
assign addr[5305]= 2063024031;
assign addr[5306]= 1957443913;
assign addr[5307]= 1812196087;
assign addr[5308]= 1630224009;
assign addr[5309]= 1415215352;
assign addr[5310]= 1171527280;
assign addr[5311]= 904098143;
assign addr[5312]= 618347408;
assign addr[5313]= 320065829;
assign addr[5314]= 15298099;
assign addr[5315]= -289779648;
assign addr[5316]= -588984994;
assign addr[5317]= -876254528;
assign addr[5318]= -1145766716;
assign addr[5319]= -1392059879;
assign addr[5320]= -1610142873;
assign addr[5321]= -1795596234;
assign addr[5322]= -1944661739;
assign addr[5323]= -2054318569;
assign addr[5324]= -2122344521;
assign addr[5325]= -2147361045;
assign addr[5326]= -2128861181;
assign addr[5327]= -2067219829;
assign addr[5328]= -1963686155;
assign addr[5329]= -1820358275;
assign addr[5330]= -1640140734;
assign addr[5331]= -1426685652;
assign addr[5332]= -1184318708;
assign addr[5333]= -917951481;
assign addr[5334]= -632981917;
assign addr[5335]= -335184940;
assign addr[5336]= -30595422;
assign addr[5337]= 274614114;
assign addr[5338]= 574258580;
assign addr[5339]= 862265664;
assign addr[5340]= 1132798888;
assign addr[5341]= 1380375881;
assign addr[5342]= 1599979481;
assign addr[5343]= 1787159411;
assign addr[5344]= 1938122457;
assign addr[5345]= 2049809346;
assign addr[5346]= 2119956737;
assign addr[5347]= 2147143090;
assign addr[5348]= 2130817471;
assign addr[5349]= 2071310720;
assign addr[5350]= 1969828744;
assign addr[5351]= 1828428082;
assign addr[5352]= 1649974225;
assign addr[5353]= 1438083551;
assign addr[5354]= 1197050035;
assign addr[5355]= 931758235;
assign addr[5356]= 647584304;
assign addr[5357]= 350287041;
assign addr[5358]= 45891193;
assign addr[5359]= -259434643;
assign addr[5360]= -559503022;
assign addr[5361]= -848233042;
assign addr[5362]= -1119773573;
assign addr[5363]= -1368621831;
assign addr[5364]= -1589734894;
assign addr[5365]= -1778631892;
assign addr[5366]= -1931484818;
assign addr[5367]= -2045196100;
assign addr[5368]= -2117461370;
assign addr[5369]= -2146816171;
assign addr[5370]= -2132665626;
assign addr[5371]= -2075296495;
assign addr[5372]= -1975871368;
assign addr[5373]= -1836405100;
assign addr[5374]= -1659723983;
assign addr[5375]= -1449408469;
assign addr[5376]= -1209720613;
assign addr[5377]= -945517704;
assign addr[5378]= -662153826;
assign addr[5379]= -365371365;
assign addr[5380]= -61184634;
assign addr[5381]= 244242007;
assign addr[5382]= 544719071;
assign addr[5383]= 834157373;
assign addr[5384]= 1106691431;
assign addr[5385]= 1356798326;
assign addr[5386]= 1579409630;
assign addr[5387]= 1770014111;
assign addr[5388]= 1924749160;
assign addr[5389]= 2040479063;
assign addr[5390]= 2114858546;
assign addr[5391]= 2146380306;
assign addr[5392]= 2134405552;
assign addr[5393]= 2079176953;
assign addr[5394]= 1981813720;
assign addr[5395]= 1844288924;
assign addr[5396]= 1669389513;
assign addr[5397]= 1460659832;
assign addr[5398]= 1222329801;
assign addr[5399]= 959229189;
assign addr[5400]= 676689746;
assign addr[5401]= 380437148;
assign addr[5402]= 76474970;
assign addr[5403]= -229036977;
assign addr[5404]= -529907477;
assign addr[5405]= -820039373;
assign addr[5406]= -1093553126;
assign addr[5407]= -1344905966;
assign addr[5408]= -1569004214;
assign addr[5409]= -1761306505;
assign addr[5410]= -1917915825;
assign addr[5411]= -2035658475;
assign addr[5412]= -2112148396;
assign addr[5413]= -2145835515;
assign addr[5414]= -2136037160;
assign addr[5415]= -2082951896;
assign addr[5416]= -1987655498;
assign addr[5417]= -1852079154;
assign addr[5418]= -1678970324;
assign addr[5419]= -1471837070;
assign addr[5420]= -1234876957;
assign addr[5421]= -972891995;
assign addr[5422]= -691191324;
assign addr[5423]= -395483624;
assign addr[5424]= -91761426;
assign addr[5425]= 213820322;
assign addr[5426]= 515068990;
assign addr[5427]= 805879757;
assign addr[5428]= 1080359326;
assign addr[5429]= 1332945355;
assign addr[5430]= 1558519173;
assign addr[5431]= 1752509516;
assign addr[5432]= 1910985158;
assign addr[5433]= 2030734582;
assign addr[5434]= 2109331059;
assign addr[5435]= 2145181827;
assign addr[5436]= 2137560369;
assign addr[5437]= 2086621133;
assign addr[5438]= 1993396407;
assign addr[5439]= 1859775393;
assign addr[5440]= 1688465931;
assign addr[5441]= 1482939614;
assign addr[5442]= 1247361445;
assign addr[5443]= 986505429;
assign addr[5444]= 705657826;
assign addr[5445]= 410510029;
assign addr[5446]= 107043224;
assign addr[5447]= -198592817;
assign addr[5448]= -500204365;
assign addr[5449]= -791679244;
assign addr[5450]= -1067110699;
assign addr[5451]= -1320917099;
assign addr[5452]= -1547955041;
assign addr[5453]= -1743623590;
assign addr[5454]= -1903957513;
assign addr[5455]= -2025707632;
assign addr[5456]= -2106406677;
assign addr[5457]= -2144419275;
assign addr[5458]= -2138975100;
assign addr[5459]= -2090184478;
assign addr[5460]= -1999036154;
assign addr[5461]= -1867377253;
assign addr[5462]= -1697875851;
assign addr[5463]= -1493966902;
assign addr[5464]= -1259782632;
assign addr[5465]= -1000068799;
assign addr[5466]= -720088517;
assign addr[5467]= -425515602;
assign addr[5468]= -122319591;
assign addr[5469]= 183355234;
assign addr[5470]= 485314355;
assign addr[5471]= 777438554;
assign addr[5472]= 1053807919;
assign addr[5473]= 1308821808;
assign addr[5474]= 1537312353;
assign addr[5475]= 1734649179;
assign addr[5476]= 1896833245;
assign addr[5477]= 2020577882;
assign addr[5478]= 2103375398;
assign addr[5479]= 2143547897;
assign addr[5480]= 2140281282;
assign addr[5481]= 2093641749;
assign addr[5482]= 2004574453;
assign addr[5483]= 1874884346;
assign addr[5484]= 1707199606;
assign addr[5485]= 1504918373;
assign addr[5486]= 1272139887;
assign addr[5487]= 1013581418;
assign addr[5488]= 734482665;
assign addr[5489]= 440499581;
assign addr[5490]= 137589750;
assign addr[5491]= -168108346;
assign addr[5492]= -470399716;
assign addr[5493]= -763158411;
assign addr[5494]= -1040451659;
assign addr[5495]= -1296660098;
assign addr[5496]= -1526591649;
assign addr[5497]= -1725586737;
assign addr[5498]= -1889612716;
assign addr[5499]= -2015345591;
assign addr[5500]= -2100237377;
assign addr[5501]= -2142567738;
assign addr[5502]= -2141478848;
assign addr[5503]= -2096992772;
assign addr[5504]= -2010011024;
assign addr[5505]= -1882296293;
assign addr[5506]= -1716436725;
assign addr[5507]= -1515793473;
assign addr[5508]= -1284432584;
assign addr[5509]= -1027042599;
assign addr[5510]= -748839539;
assign addr[5511]= -455461206;
assign addr[5512]= -152852926;
assign addr[5513]= 152852926;
assign addr[5514]= 455461206;
assign addr[5515]= 748839539;
assign addr[5516]= 1027042599;
assign addr[5517]= 1284432584;
assign addr[5518]= 1515793473;
assign addr[5519]= 1716436725;
assign addr[5520]= 1882296293;
assign addr[5521]= 2010011024;
assign addr[5522]= 2096992772;
assign addr[5523]= 2141478848;
assign addr[5524]= 2142567738;
assign addr[5525]= 2100237377;
assign addr[5526]= 2015345591;
assign addr[5527]= 1889612716;
assign addr[5528]= 1725586737;
assign addr[5529]= 1526591649;
assign addr[5530]= 1296660098;
assign addr[5531]= 1040451659;
assign addr[5532]= 763158411;
assign addr[5533]= 470399716;
assign addr[5534]= 168108346;
assign addr[5535]= -137589750;
assign addr[5536]= -440499581;
assign addr[5537]= -734482665;
assign addr[5538]= -1013581418;
assign addr[5539]= -1272139887;
assign addr[5540]= -1504918373;
assign addr[5541]= -1707199606;
assign addr[5542]= -1874884346;
assign addr[5543]= -2004574453;
assign addr[5544]= -2093641749;
assign addr[5545]= -2140281282;
assign addr[5546]= -2143547897;
assign addr[5547]= -2103375398;
assign addr[5548]= -2020577882;
assign addr[5549]= -1896833245;
assign addr[5550]= -1734649179;
assign addr[5551]= -1537312353;
assign addr[5552]= -1308821808;
assign addr[5553]= -1053807919;
assign addr[5554]= -777438554;
assign addr[5555]= -485314355;
assign addr[5556]= -183355234;
assign addr[5557]= 122319591;
assign addr[5558]= 425515602;
assign addr[5559]= 720088517;
assign addr[5560]= 1000068799;
assign addr[5561]= 1259782632;
assign addr[5562]= 1493966902;
assign addr[5563]= 1697875851;
assign addr[5564]= 1867377253;
assign addr[5565]= 1999036154;
assign addr[5566]= 2090184478;
assign addr[5567]= 2138975100;
assign addr[5568]= 2144419275;
assign addr[5569]= 2106406677;
assign addr[5570]= 2025707632;
assign addr[5571]= 1903957513;
assign addr[5572]= 1743623590;
assign addr[5573]= 1547955041;
assign addr[5574]= 1320917099;
assign addr[5575]= 1067110699;
assign addr[5576]= 791679244;
assign addr[5577]= 500204365;
assign addr[5578]= 198592817;
assign addr[5579]= -107043224;
assign addr[5580]= -410510029;
assign addr[5581]= -705657826;
assign addr[5582]= -986505429;
assign addr[5583]= -1247361445;
assign addr[5584]= -1482939614;
assign addr[5585]= -1688465931;
assign addr[5586]= -1859775393;
assign addr[5587]= -1993396407;
assign addr[5588]= -2086621133;
assign addr[5589]= -2137560369;
assign addr[5590]= -2145181827;
assign addr[5591]= -2109331059;
assign addr[5592]= -2030734582;
assign addr[5593]= -1910985158;
assign addr[5594]= -1752509516;
assign addr[5595]= -1558519173;
assign addr[5596]= -1332945355;
assign addr[5597]= -1080359326;
assign addr[5598]= -805879757;
assign addr[5599]= -515068990;
assign addr[5600]= -213820322;
assign addr[5601]= 91761426;
assign addr[5602]= 395483624;
assign addr[5603]= 691191324;
assign addr[5604]= 972891995;
assign addr[5605]= 1234876957;
assign addr[5606]= 1471837070;
assign addr[5607]= 1678970324;
assign addr[5608]= 1852079154;
assign addr[5609]= 1987655498;
assign addr[5610]= 2082951896;
assign addr[5611]= 2136037160;
assign addr[5612]= 2145835515;
assign addr[5613]= 2112148396;
assign addr[5614]= 2035658475;
assign addr[5615]= 1917915825;
assign addr[5616]= 1761306505;
assign addr[5617]= 1569004214;
assign addr[5618]= 1344905966;
assign addr[5619]= 1093553126;
assign addr[5620]= 820039373;
assign addr[5621]= 529907477;
assign addr[5622]= 229036977;
assign addr[5623]= -76474970;
assign addr[5624]= -380437148;
assign addr[5625]= -676689746;
assign addr[5626]= -959229189;
assign addr[5627]= -1222329801;
assign addr[5628]= -1460659832;
assign addr[5629]= -1669389513;
assign addr[5630]= -1844288924;
assign addr[5631]= -1981813720;
assign addr[5632]= -2079176953;
assign addr[5633]= -2134405552;
assign addr[5634]= -2146380306;
assign addr[5635]= -2114858546;
assign addr[5636]= -2040479063;
assign addr[5637]= -1924749160;
assign addr[5638]= -1770014111;
assign addr[5639]= -1579409630;
assign addr[5640]= -1356798326;
assign addr[5641]= -1106691431;
assign addr[5642]= -834157373;
assign addr[5643]= -544719071;
assign addr[5644]= -244242007;
assign addr[5645]= 61184634;
assign addr[5646]= 365371365;
assign addr[5647]= 662153826;
assign addr[5648]= 945517704;
assign addr[5649]= 1209720613;
assign addr[5650]= 1449408469;
assign addr[5651]= 1659723983;
assign addr[5652]= 1836405100;
assign addr[5653]= 1975871368;
assign addr[5654]= 2075296495;
assign addr[5655]= 2132665626;
assign addr[5656]= 2146816171;
assign addr[5657]= 2117461370;
assign addr[5658]= 2045196100;
assign addr[5659]= 1931484818;
assign addr[5660]= 1778631892;
assign addr[5661]= 1589734894;
assign addr[5662]= 1368621831;
assign addr[5663]= 1119773573;
assign addr[5664]= 848233042;
assign addr[5665]= 559503022;
assign addr[5666]= 259434643;
assign addr[5667]= -45891193;
assign addr[5668]= -350287041;
assign addr[5669]= -647584304;
assign addr[5670]= -931758235;
assign addr[5671]= -1197050035;
assign addr[5672]= -1438083551;
assign addr[5673]= -1649974225;
assign addr[5674]= -1828428082;
assign addr[5675]= -1969828744;
assign addr[5676]= -2071310720;
assign addr[5677]= -2130817471;
assign addr[5678]= -2147143090;
assign addr[5679]= -2119956737;
assign addr[5680]= -2049809346;
assign addr[5681]= -1938122457;
assign addr[5682]= -1787159411;
assign addr[5683]= -1599979481;
assign addr[5684]= -1380375881;
assign addr[5685]= -1132798888;
assign addr[5686]= -862265664;
assign addr[5687]= -574258580;
assign addr[5688]= -274614114;
assign addr[5689]= 30595422;
assign addr[5690]= 335184940;
assign addr[5691]= 632981917;
assign addr[5692]= 917951481;
assign addr[5693]= 1184318708;
assign addr[5694]= 1426685652;
assign addr[5695]= 1640140734;
assign addr[5696]= 1820358275;
assign addr[5697]= 1963686155;
assign addr[5698]= 2067219829;
assign addr[5699]= 2128861181;
assign addr[5700]= 2147361045;
assign addr[5701]= 2122344521;
assign addr[5702]= 2054318569;
assign addr[5703]= 1944661739;
assign addr[5704]= 1795596234;
assign addr[5705]= 1610142873;
assign addr[5706]= 1392059879;
assign addr[5707]= 1145766716;
assign addr[5708]= 876254528;
assign addr[5709]= 588984994;
assign addr[5710]= 289779648;
assign addr[5711]= -15298099;
assign addr[5712]= -320065829;
assign addr[5713]= -618347408;
assign addr[5714]= -904098143;
assign addr[5715]= -1171527280;
assign addr[5716]= -1415215352;
assign addr[5717]= -1630224009;
assign addr[5718]= -1812196087;
assign addr[5719]= -1957443913;
assign addr[5720]= -2063024031;
assign addr[5721]= -2126796855;
assign addr[5722]= -2147470025;
assign addr[5723]= -2124624598;
assign addr[5724]= -2058723538;
assign addr[5725]= -1951102334;
assign addr[5726]= -1803941934;
assign addr[5727]= -1620224553;
assign addr[5728]= -1403673233;
assign addr[5729]= -1158676398;
assign addr[5730]= -890198924;
assign addr[5731]= -603681519;
assign addr[5732]= -304930476;
assign addr[5733]= 0;
assign addr[5734]= 304930476;
assign addr[5735]= 603681519;
assign addr[5736]= 890198924;
assign addr[5737]= 1158676398;
assign addr[5738]= 1403673233;
assign addr[5739]= 1620224553;
assign addr[5740]= 1803941934;
assign addr[5741]= 1951102334;
assign addr[5742]= 2058723538;
assign addr[5743]= 2124624598;
assign addr[5744]= 2147470025;
assign addr[5745]= 2126796855;
assign addr[5746]= 2063024031;
assign addr[5747]= 1957443913;
assign addr[5748]= 1812196087;
assign addr[5749]= 1630224009;
assign addr[5750]= 1415215352;
assign addr[5751]= 1171527280;
assign addr[5752]= 904098143;
assign addr[5753]= 618347408;
assign addr[5754]= 320065829;
assign addr[5755]= 15298099;
assign addr[5756]= -289779648;
assign addr[5757]= -588984994;
assign addr[5758]= -876254528;
assign addr[5759]= -1145766716;
assign addr[5760]= -1392059879;
assign addr[5761]= -1610142873;
assign addr[5762]= -1795596234;
assign addr[5763]= -1944661739;
assign addr[5764]= -2054318569;
assign addr[5765]= -2122344521;
assign addr[5766]= -2147361045;
assign addr[5767]= -2128861181;
assign addr[5768]= -2067219829;
assign addr[5769]= -1963686155;
assign addr[5770]= -1820358275;
assign addr[5771]= -1640140734;
assign addr[5772]= -1426685652;
assign addr[5773]= -1184318708;
assign addr[5774]= -917951481;
assign addr[5775]= -632981917;
assign addr[5776]= -335184940;
assign addr[5777]= -30595422;
assign addr[5778]= 274614114;
assign addr[5779]= 574258580;
assign addr[5780]= 862265664;
assign addr[5781]= 1132798888;
assign addr[5782]= 1380375881;
assign addr[5783]= 1599979481;
assign addr[5784]= 1787159411;
assign addr[5785]= 1938122457;
assign addr[5786]= 2049809346;
assign addr[5787]= 2119956737;
assign addr[5788]= 2147143090;
assign addr[5789]= 2130817471;
assign addr[5790]= 2071310720;
assign addr[5791]= 1969828744;
assign addr[5792]= 1828428082;
assign addr[5793]= 1649974225;
assign addr[5794]= 1438083551;
assign addr[5795]= 1197050035;
assign addr[5796]= 931758235;
assign addr[5797]= 647584304;
assign addr[5798]= 350287041;
assign addr[5799]= 45891193;
assign addr[5800]= -259434643;
assign addr[5801]= -559503022;
assign addr[5802]= -848233042;
assign addr[5803]= -1119773573;
assign addr[5804]= -1368621831;
assign addr[5805]= -1589734894;
assign addr[5806]= -1778631892;
assign addr[5807]= -1931484818;
assign addr[5808]= -2045196100;
assign addr[5809]= -2117461370;
assign addr[5810]= -2146816171;
assign addr[5811]= -2132665626;
assign addr[5812]= -2075296495;
assign addr[5813]= -1975871368;
assign addr[5814]= -1836405100;
assign addr[5815]= -1659723983;
assign addr[5816]= -1449408469;
assign addr[5817]= -1209720613;
assign addr[5818]= -945517704;
assign addr[5819]= -662153826;
assign addr[5820]= -365371365;
assign addr[5821]= -61184634;
assign addr[5822]= 244242007;
assign addr[5823]= 544719071;
assign addr[5824]= 834157373;
assign addr[5825]= 1106691431;
assign addr[5826]= 1356798326;
assign addr[5827]= 1579409630;
assign addr[5828]= 1770014111;
assign addr[5829]= 1924749160;
assign addr[5830]= 2040479063;
assign addr[5831]= 2114858546;
assign addr[5832]= 2146380306;
assign addr[5833]= 2134405552;
assign addr[5834]= 2079176953;
assign addr[5835]= 1981813720;
assign addr[5836]= 1844288924;
assign addr[5837]= 1669389513;
assign addr[5838]= 1460659832;
assign addr[5839]= 1222329801;
assign addr[5840]= 959229189;
assign addr[5841]= 676689746;
assign addr[5842]= 380437148;
assign addr[5843]= 76474970;
assign addr[5844]= -229036977;
assign addr[5845]= -529907477;
assign addr[5846]= -820039373;
assign addr[5847]= -1093553126;
assign addr[5848]= -1344905966;
assign addr[5849]= -1569004214;
assign addr[5850]= -1761306505;
assign addr[5851]= -1917915825;
assign addr[5852]= -2035658475;
assign addr[5853]= -2112148396;
assign addr[5854]= -2145835515;
assign addr[5855]= -2136037160;
assign addr[5856]= -2082951896;
assign addr[5857]= -1987655498;
assign addr[5858]= -1852079154;
assign addr[5859]= -1678970324;
assign addr[5860]= -1471837070;
assign addr[5861]= -1234876957;
assign addr[5862]= -972891995;
assign addr[5863]= -691191324;
assign addr[5864]= -395483624;
assign addr[5865]= -91761426;
assign addr[5866]= 213820322;
assign addr[5867]= 515068990;
assign addr[5868]= 805879757;
assign addr[5869]= 1080359326;
assign addr[5870]= 1332945355;
assign addr[5871]= 1558519173;
assign addr[5872]= 1752509516;
assign addr[5873]= 1910985158;
assign addr[5874]= 2030734582;
assign addr[5875]= 2109331059;
assign addr[5876]= 2145181827;
assign addr[5877]= 2137560369;
assign addr[5878]= 2086621133;
assign addr[5879]= 1993396407;
assign addr[5880]= 1859775393;
assign addr[5881]= 1688465931;
assign addr[5882]= 1482939614;
assign addr[5883]= 1247361445;
assign addr[5884]= 986505429;
assign addr[5885]= 705657826;
assign addr[5886]= 410510029;
assign addr[5887]= 107043224;
assign addr[5888]= -198592817;
assign addr[5889]= -500204365;
assign addr[5890]= -791679244;
assign addr[5891]= -1067110699;
assign addr[5892]= -1320917099;
assign addr[5893]= -1547955041;
assign addr[5894]= -1743623590;
assign addr[5895]= -1903957513;
assign addr[5896]= -2025707632;
assign addr[5897]= -2106406677;
assign addr[5898]= -2144419275;
assign addr[5899]= -2138975100;
assign addr[5900]= -2090184478;
assign addr[5901]= -1999036154;
assign addr[5902]= -1867377253;
assign addr[5903]= -1697875851;
assign addr[5904]= -1493966902;
assign addr[5905]= -1259782632;
assign addr[5906]= -1000068799;
assign addr[5907]= -720088517;
assign addr[5908]= -425515602;
assign addr[5909]= -122319591;
assign addr[5910]= 183355234;
assign addr[5911]= 485314355;
assign addr[5912]= 777438554;
assign addr[5913]= 1053807919;
assign addr[5914]= 1308821808;
assign addr[5915]= 1537312353;
assign addr[5916]= 1734649179;
assign addr[5917]= 1896833245;
assign addr[5918]= 2020577882;
assign addr[5919]= 2103375398;
assign addr[5920]= 2143547897;
assign addr[5921]= 2140281282;
assign addr[5922]= 2093641749;
assign addr[5923]= 2004574453;
assign addr[5924]= 1874884346;
assign addr[5925]= 1707199606;
assign addr[5926]= 1504918373;
assign addr[5927]= 1272139887;
assign addr[5928]= 1013581418;
assign addr[5929]= 734482665;
assign addr[5930]= 440499581;
assign addr[5931]= 137589750;
assign addr[5932]= -168108346;
assign addr[5933]= -470399716;
assign addr[5934]= -763158411;
assign addr[5935]= -1040451659;
assign addr[5936]= -1296660098;
assign addr[5937]= -1526591649;
assign addr[5938]= -1725586737;
assign addr[5939]= -1889612716;
assign addr[5940]= -2015345591;
assign addr[5941]= -2100237377;
assign addr[5942]= -2142567738;
assign addr[5943]= -2141478848;
assign addr[5944]= -2096992772;
assign addr[5945]= -2010011024;
assign addr[5946]= -1882296293;
assign addr[5947]= -1716436725;
assign addr[5948]= -1515793473;
assign addr[5949]= -1284432584;
assign addr[5950]= -1027042599;
assign addr[5951]= -748839539;
assign addr[5952]= -455461206;
assign addr[5953]= -152852926;
assign addr[5954]= 152852926;
assign addr[5955]= 455461206;
assign addr[5956]= 748839539;
assign addr[5957]= 1027042599;
assign addr[5958]= 1284432584;
assign addr[5959]= 1515793473;
assign addr[5960]= 1716436725;
assign addr[5961]= 1882296293;
assign addr[5962]= 2010011024;
assign addr[5963]= 2096992772;
assign addr[5964]= 2141478848;
assign addr[5965]= 2142567738;
assign addr[5966]= 2100237377;
assign addr[5967]= 2015345591;
assign addr[5968]= 1889612716;
assign addr[5969]= 1725586737;
assign addr[5970]= 1526591649;
assign addr[5971]= 1296660098;
assign addr[5972]= 1040451659;
assign addr[5973]= 763158411;
assign addr[5974]= 470399716;
assign addr[5975]= 168108346;
assign addr[5976]= -137589750;
assign addr[5977]= -440499581;
assign addr[5978]= -734482665;
assign addr[5979]= -1013581418;
assign addr[5980]= -1272139887;
assign addr[5981]= -1504918373;
assign addr[5982]= -1707199606;
assign addr[5983]= -1874884346;
assign addr[5984]= -2004574453;
assign addr[5985]= -2093641749;
assign addr[5986]= -2140281282;
assign addr[5987]= -2143547897;
assign addr[5988]= -2103375398;
assign addr[5989]= -2020577882;
assign addr[5990]= -1896833245;
assign addr[5991]= -1734649179;
assign addr[5992]= -1537312353;
assign addr[5993]= -1308821808;
assign addr[5994]= -1053807919;
assign addr[5995]= -777438554;
assign addr[5996]= -485314355;
assign addr[5997]= -183355234;
assign addr[5998]= 122319591;
assign addr[5999]= 425515602;
assign addr[6000]= 720088517;
assign addr[6001]= 1000068799;
assign addr[6002]= 1259782632;
assign addr[6003]= 1493966902;
assign addr[6004]= 1697875851;
assign addr[6005]= 1867377253;
assign addr[6006]= 1999036154;
assign addr[6007]= 2090184478;
assign addr[6008]= 2138975100;
assign addr[6009]= 2144419275;
assign addr[6010]= 2106406677;
assign addr[6011]= 2025707632;
assign addr[6012]= 1903957513;
assign addr[6013]= 1743623590;
assign addr[6014]= 1547955041;
assign addr[6015]= 1320917099;
assign addr[6016]= 1067110699;
assign addr[6017]= 791679244;
assign addr[6018]= 500204365;
assign addr[6019]= 198592817;
assign addr[6020]= -107043224;
assign addr[6021]= -410510029;
assign addr[6022]= -705657826;
assign addr[6023]= -986505429;
assign addr[6024]= -1247361445;
assign addr[6025]= -1482939614;
assign addr[6026]= -1688465931;
assign addr[6027]= -1859775393;
assign addr[6028]= -1993396407;
assign addr[6029]= -2086621133;
assign addr[6030]= -2137560369;
assign addr[6031]= -2145181827;
assign addr[6032]= -2109331059;
assign addr[6033]= -2030734582;
assign addr[6034]= -1910985158;
assign addr[6035]= -1752509516;
assign addr[6036]= -1558519173;
assign addr[6037]= -1332945355;
assign addr[6038]= -1080359326;
assign addr[6039]= -805879757;
assign addr[6040]= -515068990;
assign addr[6041]= -213820322;
assign addr[6042]= 91761426;
assign addr[6043]= 395483624;
assign addr[6044]= 691191324;
assign addr[6045]= 972891995;
assign addr[6046]= 1234876957;
assign addr[6047]= 1471837070;
assign addr[6048]= 1678970324;
assign addr[6049]= 1852079154;
assign addr[6050]= 1987655498;
assign addr[6051]= 2082951896;
assign addr[6052]= 2136037160;
assign addr[6053]= 2145835515;
assign addr[6054]= 2112148396;
assign addr[6055]= 2035658475;
assign addr[6056]= 1917915825;
assign addr[6057]= 1761306505;
assign addr[6058]= 1569004214;
assign addr[6059]= 1344905966;
assign addr[6060]= 1093553126;
assign addr[6061]= 820039373;
assign addr[6062]= 529907477;
assign addr[6063]= 229036977;
assign addr[6064]= -76474970;
assign addr[6065]= -380437148;
assign addr[6066]= -676689746;
assign addr[6067]= -959229189;
assign addr[6068]= -1222329801;
assign addr[6069]= -1460659832;
assign addr[6070]= -1669389513;
assign addr[6071]= -1844288924;
assign addr[6072]= -1981813720;
assign addr[6073]= -2079176953;
assign addr[6074]= -2134405552;
assign addr[6075]= -2146380306;
assign addr[6076]= -2114858546;
assign addr[6077]= -2040479063;
assign addr[6078]= -1924749160;
assign addr[6079]= -1770014111;
assign addr[6080]= -1579409630;
assign addr[6081]= -1356798326;
assign addr[6082]= -1106691431;
assign addr[6083]= -834157373;
assign addr[6084]= -544719071;
assign addr[6085]= -244242007;
assign addr[6086]= 61184634;
assign addr[6087]= 365371365;
assign addr[6088]= 662153826;
assign addr[6089]= 945517704;
assign addr[6090]= 1209720613;
assign addr[6091]= 1449408469;
assign addr[6092]= 1659723983;
assign addr[6093]= 1836405100;
assign addr[6094]= 1975871368;
assign addr[6095]= 2075296495;
assign addr[6096]= 2132665626;
assign addr[6097]= 2146816171;
assign addr[6098]= 2117461370;
assign addr[6099]= 2045196100;
assign addr[6100]= 1931484818;
assign addr[6101]= 1778631892;
assign addr[6102]= 1589734894;
assign addr[6103]= 1368621831;
assign addr[6104]= 1119773573;
assign addr[6105]= 848233042;
assign addr[6106]= 559503022;
assign addr[6107]= 259434643;
assign addr[6108]= -45891193;
assign addr[6109]= -350287041;
assign addr[6110]= -647584304;
assign addr[6111]= -931758235;
assign addr[6112]= -1197050035;
assign addr[6113]= -1438083551;
assign addr[6114]= -1649974225;
assign addr[6115]= -1828428082;
assign addr[6116]= -1969828744;
assign addr[6117]= -2071310720;
assign addr[6118]= -2130817471;
assign addr[6119]= -2147143090;
assign addr[6120]= -2119956737;
assign addr[6121]= -2049809346;
assign addr[6122]= -1938122457;
assign addr[6123]= -1787159411;
assign addr[6124]= -1599979481;
assign addr[6125]= -1380375881;
assign addr[6126]= -1132798888;
assign addr[6127]= -862265664;
assign addr[6128]= -574258580;
assign addr[6129]= -274614114;
assign addr[6130]= 30595422;
assign addr[6131]= 335184940;
assign addr[6132]= 632981917;
assign addr[6133]= 917951481;
assign addr[6134]= 1184318708;
assign addr[6135]= 1426685652;
assign addr[6136]= 1640140734;
assign addr[6137]= 1820358275;
assign addr[6138]= 1963686155;
assign addr[6139]= 2067219829;
assign addr[6140]= 2128861181;
assign addr[6141]= 2147361045;
assign addr[6142]= 2122344521;
assign addr[6143]= 2054318569;
assign addr[6144]= 1944661739;
assign addr[6145]= 1795596234;
assign addr[6146]= 1610142873;
assign addr[6147]= 1392059879;
assign addr[6148]= 1145766716;
assign addr[6149]= 876254528;
assign addr[6150]= 588984994;
assign addr[6151]= 289779648;
assign addr[6152]= -15298099;
assign addr[6153]= -320065829;
assign addr[6154]= -618347408;
assign addr[6155]= -904098143;
assign addr[6156]= -1171527280;
assign addr[6157]= -1415215352;
assign addr[6158]= -1630224009;
assign addr[6159]= -1812196087;
assign addr[6160]= -1957443913;
assign addr[6161]= -2063024031;
assign addr[6162]= -2126796855;
assign addr[6163]= -2147470025;
assign addr[6164]= -2124624598;
assign addr[6165]= -2058723538;
assign addr[6166]= -1951102334;
assign addr[6167]= -1803941934;
assign addr[6168]= -1620224553;
assign addr[6169]= -1403673233;
assign addr[6170]= -1158676398;
assign addr[6171]= -890198924;
assign addr[6172]= -603681519;
assign addr[6173]= -304930476;
assign addr[6174]= 0;
assign addr[6175]= 304930476;
assign addr[6176]= 603681519;
assign addr[6177]= 890198924;
assign addr[6178]= 1158676398;
assign addr[6179]= 1403673233;
assign addr[6180]= 1620224553;
assign addr[6181]= 1803941934;
assign addr[6182]= 1951102334;
assign addr[6183]= 2058723538;
assign addr[6184]= 2124624598;
assign addr[6185]= 2147470025;
assign addr[6186]= 2126796855;
assign addr[6187]= 2063024031;
assign addr[6188]= 1957443913;
assign addr[6189]= 1812196087;
assign addr[6190]= 1630224009;
assign addr[6191]= 1415215352;
assign addr[6192]= 1171527280;
assign addr[6193]= 904098143;
assign addr[6194]= 618347408;
assign addr[6195]= 320065829;
assign addr[6196]= 15298099;
assign addr[6197]= -289779648;
assign addr[6198]= -588984994;
assign addr[6199]= -876254528;
assign addr[6200]= -1145766716;
assign addr[6201]= -1392059879;
assign addr[6202]= -1610142873;
assign addr[6203]= -1795596234;
assign addr[6204]= -1944661739;
assign addr[6205]= -2054318569;
assign addr[6206]= -2122344521;
assign addr[6207]= -2147361045;
assign addr[6208]= -2128861181;
assign addr[6209]= -2067219829;
assign addr[6210]= -1963686155;
assign addr[6211]= -1820358275;
assign addr[6212]= -1640140734;
assign addr[6213]= -1426685652;
assign addr[6214]= -1184318708;
assign addr[6215]= -917951481;
assign addr[6216]= -632981917;
assign addr[6217]= -335184940;
assign addr[6218]= -30595422;
assign addr[6219]= 274614114;
assign addr[6220]= 574258580;
assign addr[6221]= 862265664;
assign addr[6222]= 1132798888;
assign addr[6223]= 1380375881;
assign addr[6224]= 1599979481;
assign addr[6225]= 1787159411;
assign addr[6226]= 1938122457;
assign addr[6227]= 2049809346;
assign addr[6228]= 2119956737;
assign addr[6229]= 2147143090;
assign addr[6230]= 2130817471;
assign addr[6231]= 2071310720;
assign addr[6232]= 1969828744;
assign addr[6233]= 1828428082;
assign addr[6234]= 1649974225;
assign addr[6235]= 1438083551;
assign addr[6236]= 1197050035;
assign addr[6237]= 931758235;
assign addr[6238]= 647584304;
assign addr[6239]= 350287041;
assign addr[6240]= 45891193;
assign addr[6241]= -259434643;
assign addr[6242]= -559503022;
assign addr[6243]= -848233042;
assign addr[6244]= -1119773573;
assign addr[6245]= -1368621831;
assign addr[6246]= -1589734894;
assign addr[6247]= -1778631892;
assign addr[6248]= -1931484818;
assign addr[6249]= -2045196100;
assign addr[6250]= -2117461370;
assign addr[6251]= -2146816171;
assign addr[6252]= -2132665626;
assign addr[6253]= -2075296495;
assign addr[6254]= -1975871368;
assign addr[6255]= -1836405100;
assign addr[6256]= -1659723983;
assign addr[6257]= -1449408469;
assign addr[6258]= -1209720613;
assign addr[6259]= -945517704;
assign addr[6260]= -662153826;
assign addr[6261]= -365371365;
assign addr[6262]= -61184634;
assign addr[6263]= 244242007;
assign addr[6264]= 544719071;
assign addr[6265]= 834157373;
assign addr[6266]= 1106691431;
assign addr[6267]= 1356798326;
assign addr[6268]= 1579409630;
assign addr[6269]= 1770014111;
assign addr[6270]= 1924749160;
assign addr[6271]= 2040479063;
assign addr[6272]= 2114858546;
assign addr[6273]= 2146380306;
assign addr[6274]= 2134405552;
assign addr[6275]= 2079176953;
assign addr[6276]= 1981813720;
assign addr[6277]= 1844288924;
assign addr[6278]= 1669389513;
assign addr[6279]= 1460659832;
assign addr[6280]= 1222329801;
assign addr[6281]= 959229189;
assign addr[6282]= 676689746;
assign addr[6283]= 380437148;
assign addr[6284]= 76474970;
assign addr[6285]= -229036977;
assign addr[6286]= -529907477;
assign addr[6287]= -820039373;
assign addr[6288]= -1093553126;
assign addr[6289]= -1344905966;
assign addr[6290]= -1569004214;
assign addr[6291]= -1761306505;
assign addr[6292]= -1917915825;
assign addr[6293]= -2035658475;
assign addr[6294]= -2112148396;
assign addr[6295]= -2145835515;
assign addr[6296]= -2136037160;
assign addr[6297]= -2082951896;
assign addr[6298]= -1987655498;
assign addr[6299]= -1852079154;
assign addr[6300]= -1678970324;
assign addr[6301]= -1471837070;
assign addr[6302]= -1234876957;
assign addr[6303]= -972891995;
assign addr[6304]= -691191324;
assign addr[6305]= -395483624;
assign addr[6306]= -91761426;
assign addr[6307]= 213820322;
assign addr[6308]= 515068990;
assign addr[6309]= 805879757;
assign addr[6310]= 1080359326;
assign addr[6311]= 1332945355;
assign addr[6312]= 1558519173;
assign addr[6313]= 1752509516;
assign addr[6314]= 1910985158;
assign addr[6315]= 2030734582;
assign addr[6316]= 2109331059;
assign addr[6317]= 2145181827;
assign addr[6318]= 2137560369;
assign addr[6319]= 2086621133;
assign addr[6320]= 1993396407;
assign addr[6321]= 1859775393;
assign addr[6322]= 1688465931;
assign addr[6323]= 1482939614;
assign addr[6324]= 1247361445;
assign addr[6325]= 986505429;
assign addr[6326]= 705657826;
assign addr[6327]= 410510029;
assign addr[6328]= 107043224;
assign addr[6329]= -198592817;
assign addr[6330]= -500204365;
assign addr[6331]= -791679244;
assign addr[6332]= -1067110699;
assign addr[6333]= -1320917099;
assign addr[6334]= -1547955041;
assign addr[6335]= -1743623590;
assign addr[6336]= -1903957513;
assign addr[6337]= -2025707632;
assign addr[6338]= -2106406677;
assign addr[6339]= -2144419275;
assign addr[6340]= -2138975100;
assign addr[6341]= -2090184478;
assign addr[6342]= -1999036154;
assign addr[6343]= -1867377253;
assign addr[6344]= -1697875851;
assign addr[6345]= -1493966902;
assign addr[6346]= -1259782632;
assign addr[6347]= -1000068799;
assign addr[6348]= -720088517;
assign addr[6349]= -425515602;
assign addr[6350]= -122319591;
assign addr[6351]= 183355234;
assign addr[6352]= 485314355;
assign addr[6353]= 777438554;
assign addr[6354]= 1053807919;
assign addr[6355]= 1308821808;
assign addr[6356]= 1537312353;
assign addr[6357]= 1734649179;
assign addr[6358]= 1896833245;
assign addr[6359]= 2020577882;
assign addr[6360]= 2103375398;
assign addr[6361]= 2143547897;
assign addr[6362]= 2140281282;
assign addr[6363]= 2093641749;
assign addr[6364]= 2004574453;
assign addr[6365]= 1874884346;
assign addr[6366]= 1707199606;
assign addr[6367]= 1504918373;
assign addr[6368]= 1272139887;
assign addr[6369]= 1013581418;
assign addr[6370]= 734482665;
assign addr[6371]= 440499581;
assign addr[6372]= 137589750;
assign addr[6373]= -168108346;
assign addr[6374]= -470399716;
assign addr[6375]= -763158411;
assign addr[6376]= -1040451659;
assign addr[6377]= -1296660098;
assign addr[6378]= -1526591649;
assign addr[6379]= -1725586737;
assign addr[6380]= -1889612716;
assign addr[6381]= -2015345591;
assign addr[6382]= -2100237377;
assign addr[6383]= -2142567738;
assign addr[6384]= -2141478848;
assign addr[6385]= -2096992772;
assign addr[6386]= -2010011024;
assign addr[6387]= -1882296293;
assign addr[6388]= -1716436725;
assign addr[6389]= -1515793473;
assign addr[6390]= -1284432584;
assign addr[6391]= -1027042599;
assign addr[6392]= -748839539;
assign addr[6393]= -455461206;
assign addr[6394]= -152852926;
assign addr[6395]= 152852926;
assign addr[6396]= 455461206;
assign addr[6397]= 748839539;
assign addr[6398]= 1027042599;
assign addr[6399]= 1284432584;
assign addr[6400]= 1515793473;
assign addr[6401]= 1716436725;
assign addr[6402]= 1882296293;
assign addr[6403]= 2010011024;
assign addr[6404]= 2096992772;
assign addr[6405]= 2141478848;
assign addr[6406]= 2142567738;
assign addr[6407]= 2100237377;
assign addr[6408]= 2015345591;
assign addr[6409]= 1889612716;
assign addr[6410]= 1725586737;
assign addr[6411]= 1526591649;
assign addr[6412]= 1296660098;
assign addr[6413]= 1040451659;
assign addr[6414]= 763158411;
assign addr[6415]= 470399716;
assign addr[6416]= 168108346;
assign addr[6417]= -137589750;
assign addr[6418]= -440499581;
assign addr[6419]= -734482665;
assign addr[6420]= -1013581418;
assign addr[6421]= -1272139887;
assign addr[6422]= -1504918373;
assign addr[6423]= -1707199606;
assign addr[6424]= -1874884346;
assign addr[6425]= -2004574453;
assign addr[6426]= -2093641749;
assign addr[6427]= -2140281282;
assign addr[6428]= -2143547897;
assign addr[6429]= -2103375398;
assign addr[6430]= -2020577882;
assign addr[6431]= -1896833245;
assign addr[6432]= -1734649179;
assign addr[6433]= -1537312353;
assign addr[6434]= -1308821808;
assign addr[6435]= -1053807919;
assign addr[6436]= -777438554;
assign addr[6437]= -485314355;
assign addr[6438]= -183355234;
assign addr[6439]= 122319591;
assign addr[6440]= 425515602;
assign addr[6441]= 720088517;
assign addr[6442]= 1000068799;
assign addr[6443]= 1259782632;
assign addr[6444]= 1493966902;
assign addr[6445]= 1697875851;
assign addr[6446]= 1867377253;
assign addr[6447]= 1999036154;
assign addr[6448]= 2090184478;
assign addr[6449]= 2138975100;
assign addr[6450]= 2144419275;
assign addr[6451]= 2106406677;
assign addr[6452]= 2025707632;
assign addr[6453]= 1903957513;
assign addr[6454]= 1743623590;
assign addr[6455]= 1547955041;
assign addr[6456]= 1320917099;
assign addr[6457]= 1067110699;
assign addr[6458]= 791679244;
assign addr[6459]= 500204365;
assign addr[6460]= 198592817;
assign addr[6461]= -107043224;
assign addr[6462]= -410510029;
assign addr[6463]= -705657826;
assign addr[6464]= -986505429;
assign addr[6465]= -1247361445;
assign addr[6466]= -1482939614;
assign addr[6467]= -1688465931;
assign addr[6468]= -1859775393;
assign addr[6469]= -1993396407;
assign addr[6470]= -2086621133;
assign addr[6471]= -2137560369;
assign addr[6472]= -2145181827;
assign addr[6473]= -2109331059;
assign addr[6474]= -2030734582;
assign addr[6475]= -1910985158;
assign addr[6476]= -1752509516;
assign addr[6477]= -1558519173;
assign addr[6478]= -1332945355;
assign addr[6479]= -1080359326;
assign addr[6480]= -805879757;
assign addr[6481]= -515068990;
assign addr[6482]= -213820322;
assign addr[6483]= 91761426;
assign addr[6484]= 395483624;
assign addr[6485]= 691191324;
assign addr[6486]= 972891995;
assign addr[6487]= 1234876957;
assign addr[6488]= 1471837070;
assign addr[6489]= 1678970324;
assign addr[6490]= 1852079154;
assign addr[6491]= 1987655498;
assign addr[6492]= 2082951896;
assign addr[6493]= 2136037160;
assign addr[6494]= 2145835515;
assign addr[6495]= 2112148396;
assign addr[6496]= 2035658475;
assign addr[6497]= 1917915825;
assign addr[6498]= 1761306505;
assign addr[6499]= 1569004214;
assign addr[6500]= 1344905966;
assign addr[6501]= 1093553126;
assign addr[6502]= 820039373;
assign addr[6503]= 529907477;
assign addr[6504]= 229036977;
assign addr[6505]= -76474970;
assign addr[6506]= -380437148;
assign addr[6507]= -676689746;
assign addr[6508]= -959229189;
assign addr[6509]= -1222329801;
assign addr[6510]= -1460659832;
assign addr[6511]= -1669389513;
assign addr[6512]= -1844288924;
assign addr[6513]= -1981813720;
assign addr[6514]= -2079176953;
assign addr[6515]= -2134405552;
assign addr[6516]= -2146380306;
assign addr[6517]= -2114858546;
assign addr[6518]= -2040479063;
assign addr[6519]= -1924749160;
assign addr[6520]= -1770014111;
assign addr[6521]= -1579409630;
assign addr[6522]= -1356798326;
assign addr[6523]= -1106691431;
assign addr[6524]= -834157373;
assign addr[6525]= -544719071;
assign addr[6526]= -244242007;
assign addr[6527]= 61184634;
assign addr[6528]= 365371365;
assign addr[6529]= 662153826;
assign addr[6530]= 945517704;
assign addr[6531]= 1209720613;
assign addr[6532]= 1449408469;
assign addr[6533]= 1659723983;
assign addr[6534]= 1836405100;
assign addr[6535]= 1975871368;
assign addr[6536]= 2075296495;
assign addr[6537]= 2132665626;
assign addr[6538]= 2146816171;
assign addr[6539]= 2117461370;
assign addr[6540]= 2045196100;
assign addr[6541]= 1931484818;
assign addr[6542]= 1778631892;
assign addr[6543]= 1589734894;
assign addr[6544]= 1368621831;
assign addr[6545]= 1119773573;
assign addr[6546]= 848233042;
assign addr[6547]= 559503022;
assign addr[6548]= 259434643;
assign addr[6549]= -45891193;
assign addr[6550]= -350287041;
assign addr[6551]= -647584304;
assign addr[6552]= -931758235;
assign addr[6553]= -1197050035;
assign addr[6554]= -1438083551;
assign addr[6555]= -1649974225;
assign addr[6556]= -1828428082;
assign addr[6557]= -1969828744;
assign addr[6558]= -2071310720;
assign addr[6559]= -2130817471;
assign addr[6560]= -2147143090;
assign addr[6561]= -2119956737;
assign addr[6562]= -2049809346;
assign addr[6563]= -1938122457;
assign addr[6564]= -1787159411;
assign addr[6565]= -1599979481;
assign addr[6566]= -1380375881;
assign addr[6567]= -1132798888;
assign addr[6568]= -862265664;
assign addr[6569]= -574258580;
assign addr[6570]= -274614114;
assign addr[6571]= 30595422;
assign addr[6572]= 335184940;
assign addr[6573]= 632981917;
assign addr[6574]= 917951481;
assign addr[6575]= 1184318708;
assign addr[6576]= 1426685652;
assign addr[6577]= 1640140734;
assign addr[6578]= 1820358275;
assign addr[6579]= 1963686155;
assign addr[6580]= 2067219829;
assign addr[6581]= 2128861181;
assign addr[6582]= 2147361045;
assign addr[6583]= 2122344521;
assign addr[6584]= 2054318569;
assign addr[6585]= 1944661739;
assign addr[6586]= 1795596234;
assign addr[6587]= 1610142873;
assign addr[6588]= 1392059879;
assign addr[6589]= 1145766716;
assign addr[6590]= 876254528;
assign addr[6591]= 588984994;
assign addr[6592]= 289779648;
assign addr[6593]= -15298099;
assign addr[6594]= -320065829;
assign addr[6595]= -618347408;
assign addr[6596]= -904098143;
assign addr[6597]= -1171527280;
assign addr[6598]= -1415215352;
assign addr[6599]= -1630224009;
assign addr[6600]= -1812196087;
assign addr[6601]= -1957443913;
assign addr[6602]= -2063024031;
assign addr[6603]= -2126796855;
assign addr[6604]= -2147470025;
assign addr[6605]= -2124624598;
assign addr[6606]= -2058723538;
assign addr[6607]= -1951102334;
assign addr[6608]= -1803941934;
assign addr[6609]= -1620224553;
assign addr[6610]= -1403673233;
assign addr[6611]= -1158676398;
assign addr[6612]= -890198924;
assign addr[6613]= -603681519;
assign addr[6614]= -304930476;
assign addr[6615]= 0;
assign addr[6616]= 304930476;
assign addr[6617]= 603681519;
assign addr[6618]= 890198924;
assign addr[6619]= 1158676398;
assign addr[6620]= 1403673233;
assign addr[6621]= 1620224553;
assign addr[6622]= 1803941934;
assign addr[6623]= 1951102334;
assign addr[6624]= 2058723538;
assign addr[6625]= 2124624598;
assign addr[6626]= 2147470025;
assign addr[6627]= 2126796855;
assign addr[6628]= 2063024031;
assign addr[6629]= 1957443913;
assign addr[6630]= 1812196087;
assign addr[6631]= 1630224009;
assign addr[6632]= 1415215352;
assign addr[6633]= 1171527280;
assign addr[6634]= 904098143;
assign addr[6635]= 618347408;
assign addr[6636]= 320065829;
assign addr[6637]= 15298099;
assign addr[6638]= -289779648;
assign addr[6639]= -588984994;
assign addr[6640]= -876254528;
assign addr[6641]= -1145766716;
assign addr[6642]= -1392059879;
assign addr[6643]= -1610142873;
assign addr[6644]= -1795596234;
assign addr[6645]= -1944661739;
assign addr[6646]= -2054318569;
assign addr[6647]= -2122344521;
assign addr[6648]= -2147361045;
assign addr[6649]= -2128861181;
assign addr[6650]= -2067219829;
assign addr[6651]= -1963686155;
assign addr[6652]= -1820358275;
assign addr[6653]= -1640140734;
assign addr[6654]= -1426685652;
assign addr[6655]= -1184318708;
assign addr[6656]= -917951481;
assign addr[6657]= -632981917;
assign addr[6658]= -335184940;
assign addr[6659]= -30595422;
assign addr[6660]= 274614114;
assign addr[6661]= 574258580;
assign addr[6662]= 862265664;
assign addr[6663]= 1132798888;
assign addr[6664]= 1380375881;
assign addr[6665]= 1599979481;
assign addr[6666]= 1787159411;
assign addr[6667]= 1938122457;
assign addr[6668]= 2049809346;
assign addr[6669]= 2119956737;
assign addr[6670]= 2147143090;
assign addr[6671]= 2130817471;
assign addr[6672]= 2071310720;
assign addr[6673]= 1969828744;
assign addr[6674]= 1828428082;
assign addr[6675]= 1649974225;
assign addr[6676]= 1438083551;
assign addr[6677]= 1197050035;
assign addr[6678]= 931758235;
assign addr[6679]= 647584304;
assign addr[6680]= 350287041;
assign addr[6681]= 45891193;
assign addr[6682]= -259434643;
assign addr[6683]= -559503022;
assign addr[6684]= -848233042;
assign addr[6685]= -1119773573;
assign addr[6686]= -1368621831;
assign addr[6687]= -1589734894;
assign addr[6688]= -1778631892;
assign addr[6689]= -1931484818;
assign addr[6690]= -2045196100;
assign addr[6691]= -2117461370;
assign addr[6692]= -2146816171;
assign addr[6693]= -2132665626;
assign addr[6694]= -2075296495;
assign addr[6695]= -1975871368;
assign addr[6696]= -1836405100;
assign addr[6697]= -1659723983;
assign addr[6698]= -1449408469;
assign addr[6699]= -1209720613;
assign addr[6700]= -945517704;
assign addr[6701]= -662153826;
assign addr[6702]= -365371365;
assign addr[6703]= -61184634;
assign addr[6704]= 244242007;
assign addr[6705]= 544719071;
assign addr[6706]= 834157373;
assign addr[6707]= 1106691431;
assign addr[6708]= 1356798326;
assign addr[6709]= 1579409630;
assign addr[6710]= 1770014111;
assign addr[6711]= 1924749160;
assign addr[6712]= 2040479063;
assign addr[6713]= 2114858546;
assign addr[6714]= 2146380306;
assign addr[6715]= 2134405552;
assign addr[6716]= 2079176953;
assign addr[6717]= 1981813720;
assign addr[6718]= 1844288924;
assign addr[6719]= 1669389513;
assign addr[6720]= 1460659832;
assign addr[6721]= 1222329801;
assign addr[6722]= 959229189;
assign addr[6723]= 676689746;
assign addr[6724]= 380437148;
assign addr[6725]= 76474970;
assign addr[6726]= -229036977;
assign addr[6727]= -529907477;
assign addr[6728]= -820039373;
assign addr[6729]= -1093553126;
assign addr[6730]= -1344905966;
assign addr[6731]= -1569004214;
assign addr[6732]= -1761306505;
assign addr[6733]= -1917915825;
assign addr[6734]= -2035658475;
assign addr[6735]= -2112148396;
assign addr[6736]= -2145835515;
assign addr[6737]= -2136037160;
assign addr[6738]= -2082951896;
assign addr[6739]= -1987655498;
assign addr[6740]= -1852079154;
assign addr[6741]= -1678970324;
assign addr[6742]= -1471837070;
assign addr[6743]= -1234876957;
assign addr[6744]= -972891995;
assign addr[6745]= -691191324;
assign addr[6746]= -395483624;
assign addr[6747]= -91761426;
assign addr[6748]= 213820322;
assign addr[6749]= 515068990;
assign addr[6750]= 805879757;
assign addr[6751]= 1080359326;
assign addr[6752]= 1332945355;
assign addr[6753]= 1558519173;
assign addr[6754]= 1752509516;
assign addr[6755]= 1910985158;
assign addr[6756]= 2030734582;
assign addr[6757]= 2109331059;
assign addr[6758]= 2145181827;
assign addr[6759]= 2137560369;
assign addr[6760]= 2086621133;
assign addr[6761]= 1993396407;
assign addr[6762]= 1859775393;
assign addr[6763]= 1688465931;
assign addr[6764]= 1482939614;
assign addr[6765]= 1247361445;
assign addr[6766]= 986505429;
assign addr[6767]= 705657826;
assign addr[6768]= 410510029;
assign addr[6769]= 107043224;
assign addr[6770]= -198592817;
assign addr[6771]= -500204365;
assign addr[6772]= -791679244;
assign addr[6773]= -1067110699;
assign addr[6774]= -1320917099;
assign addr[6775]= -1547955041;
assign addr[6776]= -1743623590;
assign addr[6777]= -1903957513;
assign addr[6778]= -2025707632;
assign addr[6779]= -2106406677;
assign addr[6780]= -2144419275;
assign addr[6781]= -2138975100;
assign addr[6782]= -2090184478;
assign addr[6783]= -1999036154;
assign addr[6784]= -1867377253;
assign addr[6785]= -1697875851;
assign addr[6786]= -1493966902;
assign addr[6787]= -1259782632;
assign addr[6788]= -1000068799;
assign addr[6789]= -720088517;
assign addr[6790]= -425515602;
assign addr[6791]= -122319591;
assign addr[6792]= 183355234;
assign addr[6793]= 485314355;
assign addr[6794]= 777438554;
assign addr[6795]= 1053807919;
assign addr[6796]= 1308821808;
assign addr[6797]= 1537312353;
assign addr[6798]= 1734649179;
assign addr[6799]= 1896833245;
assign addr[6800]= 2020577882;
assign addr[6801]= 2103375398;
assign addr[6802]= 2143547897;
assign addr[6803]= 2140281282;
assign addr[6804]= 2093641749;
assign addr[6805]= 2004574453;
assign addr[6806]= 1874884346;
assign addr[6807]= 1707199606;
assign addr[6808]= 1504918373;
assign addr[6809]= 1272139887;
assign addr[6810]= 1013581418;
assign addr[6811]= 734482665;
assign addr[6812]= 440499581;
assign addr[6813]= 137589750;
assign addr[6814]= -168108346;
assign addr[6815]= -470399716;
assign addr[6816]= -763158411;
assign addr[6817]= -1040451659;
assign addr[6818]= -1296660098;
assign addr[6819]= -1526591649;
assign addr[6820]= -1725586737;
assign addr[6821]= -1889612716;
assign addr[6822]= -2015345591;
assign addr[6823]= -2100237377;
assign addr[6824]= -2142567738;
assign addr[6825]= -2141478848;
assign addr[6826]= -2096992772;
assign addr[6827]= -2010011024;
assign addr[6828]= -1882296293;
assign addr[6829]= -1716436725;
assign addr[6830]= -1515793473;
assign addr[6831]= -1284432584;
assign addr[6832]= -1027042599;
assign addr[6833]= -748839539;
assign addr[6834]= -455461206;
assign addr[6835]= -152852926;
assign addr[6836]= 152852926;
assign addr[6837]= 455461206;
assign addr[6838]= 748839539;
assign addr[6839]= 1027042599;
assign addr[6840]= 1284432584;
assign addr[6841]= 1515793473;
assign addr[6842]= 1716436725;
assign addr[6843]= 1882296293;
assign addr[6844]= 2010011024;
assign addr[6845]= 2096992772;
assign addr[6846]= 2141478848;
assign addr[6847]= 2142567738;
assign addr[6848]= 2100237377;
assign addr[6849]= 2015345591;
assign addr[6850]= 1889612716;
assign addr[6851]= 1725586737;
assign addr[6852]= 1526591649;
assign addr[6853]= 1296660098;
assign addr[6854]= 1040451659;
assign addr[6855]= 763158411;
assign addr[6856]= 470399716;
assign addr[6857]= 168108346;
assign addr[6858]= -137589750;
assign addr[6859]= -440499581;
assign addr[6860]= -734482665;
assign addr[6861]= -1013581418;
assign addr[6862]= -1272139887;
assign addr[6863]= -1504918373;
assign addr[6864]= -1707199606;
assign addr[6865]= -1874884346;
assign addr[6866]= -2004574453;
assign addr[6867]= -2093641749;
assign addr[6868]= -2140281282;
assign addr[6869]= -2143547897;
assign addr[6870]= -2103375398;
assign addr[6871]= -2020577882;
assign addr[6872]= -1896833245;
assign addr[6873]= -1734649179;
assign addr[6874]= -1537312353;
assign addr[6875]= -1308821808;
assign addr[6876]= -1053807919;
assign addr[6877]= -777438554;
assign addr[6878]= -485314355;
assign addr[6879]= -183355234;
assign addr[6880]= 122319591;
assign addr[6881]= 425515602;
assign addr[6882]= 720088517;
assign addr[6883]= 1000068799;
assign addr[6884]= 1259782632;
assign addr[6885]= 1493966902;
assign addr[6886]= 1697875851;
assign addr[6887]= 1867377253;
assign addr[6888]= 1999036154;
assign addr[6889]= 2090184478;
assign addr[6890]= 2138975100;
assign addr[6891]= 2144419275;
assign addr[6892]= 2106406677;
assign addr[6893]= 2025707632;
assign addr[6894]= 1903957513;
assign addr[6895]= 1743623590;
assign addr[6896]= 1547955041;
assign addr[6897]= 1320917099;
assign addr[6898]= 1067110699;
assign addr[6899]= 791679244;
assign addr[6900]= 500204365;
assign addr[6901]= 198592817;
assign addr[6902]= -107043224;
assign addr[6903]= -410510029;
assign addr[6904]= -705657826;
assign addr[6905]= -986505429;
assign addr[6906]= -1247361445;
assign addr[6907]= -1482939614;
assign addr[6908]= -1688465931;
assign addr[6909]= -1859775393;
assign addr[6910]= -1993396407;
assign addr[6911]= -2086621133;
assign addr[6912]= -2137560369;
assign addr[6913]= -2145181827;
assign addr[6914]= -2109331059;
assign addr[6915]= -2030734582;
assign addr[6916]= -1910985158;
assign addr[6917]= -1752509516;
assign addr[6918]= -1558519173;
assign addr[6919]= -1332945355;
assign addr[6920]= -1080359326;
assign addr[6921]= -805879757;
assign addr[6922]= -515068990;
assign addr[6923]= -213820322;
assign addr[6924]= 91761426;
assign addr[6925]= 395483624;
assign addr[6926]= 691191324;
assign addr[6927]= 972891995;
assign addr[6928]= 1234876957;
assign addr[6929]= 1471837070;
assign addr[6930]= 1678970324;
assign addr[6931]= 1852079154;
assign addr[6932]= 1987655498;
assign addr[6933]= 2082951896;
assign addr[6934]= 2136037160;
assign addr[6935]= 2145835515;
assign addr[6936]= 2112148396;
assign addr[6937]= 2035658475;
assign addr[6938]= 1917915825;
assign addr[6939]= 1761306505;
assign addr[6940]= 1569004214;
assign addr[6941]= 1344905966;
assign addr[6942]= 1093553126;
assign addr[6943]= 820039373;
assign addr[6944]= 529907477;
assign addr[6945]= 229036977;
assign addr[6946]= -76474970;
assign addr[6947]= -380437148;
assign addr[6948]= -676689746;
assign addr[6949]= -959229189;
assign addr[6950]= -1222329801;
assign addr[6951]= -1460659832;
assign addr[6952]= -1669389513;
assign addr[6953]= -1844288924;
assign addr[6954]= -1981813720;
assign addr[6955]= -2079176953;
assign addr[6956]= -2134405552;
assign addr[6957]= -2146380306;
assign addr[6958]= -2114858546;
assign addr[6959]= -2040479063;
assign addr[6960]= -1924749160;
assign addr[6961]= -1770014111;
assign addr[6962]= -1579409630;
assign addr[6963]= -1356798326;
assign addr[6964]= -1106691431;
assign addr[6965]= -834157373;
assign addr[6966]= -544719071;
assign addr[6967]= -244242007;
assign addr[6968]= 61184634;
assign addr[6969]= 365371365;
assign addr[6970]= 662153826;
assign addr[6971]= 945517704;
assign addr[6972]= 1209720613;
assign addr[6973]= 1449408469;
assign addr[6974]= 1659723983;
assign addr[6975]= 1836405100;
assign addr[6976]= 1975871368;
assign addr[6977]= 2075296495;
assign addr[6978]= 2132665626;
assign addr[6979]= 2146816171;
assign addr[6980]= 2117461370;
assign addr[6981]= 2045196100;
assign addr[6982]= 1931484818;
assign addr[6983]= 1778631892;
assign addr[6984]= 1589734894;
assign addr[6985]= 1368621831;
assign addr[6986]= 1119773573;
assign addr[6987]= 848233042;
assign addr[6988]= 559503022;
assign addr[6989]= 259434643;
assign addr[6990]= -45891193;
assign addr[6991]= -350287041;
assign addr[6992]= -647584304;
assign addr[6993]= -931758235;
assign addr[6994]= -1197050035;
assign addr[6995]= -1438083551;
assign addr[6996]= -1649974225;
assign addr[6997]= -1828428082;
assign addr[6998]= -1969828744;
assign addr[6999]= -2071310720;
assign addr[7000]= -2130817471;
assign addr[7001]= -2147143090;
assign addr[7002]= -2119956737;
assign addr[7003]= -2049809346;
assign addr[7004]= -1938122457;
assign addr[7005]= -1787159411;
assign addr[7006]= -1599979481;
assign addr[7007]= -1380375881;
assign addr[7008]= -1132798888;
assign addr[7009]= -862265664;
assign addr[7010]= -574258580;
assign addr[7011]= -274614114;
assign addr[7012]= 30595422;
assign addr[7013]= 335184940;
assign addr[7014]= 632981917;
assign addr[7015]= 917951481;
assign addr[7016]= 1184318708;
assign addr[7017]= 1426685652;
assign addr[7018]= 1640140734;
assign addr[7019]= 1820358275;
assign addr[7020]= 1963686155;
assign addr[7021]= 2067219829;
assign addr[7022]= 2128861181;
assign addr[7023]= 2147361045;
assign addr[7024]= 2122344521;
assign addr[7025]= 2054318569;
assign addr[7026]= 1944661739;
assign addr[7027]= 1795596234;
assign addr[7028]= 1610142873;
assign addr[7029]= 1392059879;
assign addr[7030]= 1145766716;
assign addr[7031]= 876254528;
assign addr[7032]= 588984994;
assign addr[7033]= 289779648;
assign addr[7034]= -15298099;
assign addr[7035]= -320065829;
assign addr[7036]= -618347408;
assign addr[7037]= -904098143;
assign addr[7038]= -1171527280;
assign addr[7039]= -1415215352;
assign addr[7040]= -1630224009;
assign addr[7041]= -1812196087;
assign addr[7042]= -1957443913;
assign addr[7043]= -2063024031;
assign addr[7044]= -2126796855;
assign addr[7045]= -2147470025;
assign addr[7046]= -2124624598;
assign addr[7047]= -2058723538;
assign addr[7048]= -1951102334;
assign addr[7049]= -1803941934;
assign addr[7050]= -1620224553;
assign addr[7051]= -1403673233;
assign addr[7052]= -1158676398;
assign addr[7053]= -890198924;
assign addr[7054]= -603681519;
assign addr[7055]= -304930476;
assign addr[7056]= 0;
assign addr[7057]= 304930476;
assign addr[7058]= 603681519;
assign addr[7059]= 890198924;
assign addr[7060]= 1158676398;
assign addr[7061]= 1403673233;
assign addr[7062]= 1620224553;
assign addr[7063]= 1803941934;
assign addr[7064]= 1951102334;
assign addr[7065]= 2058723538;
assign addr[7066]= 2124624598;
assign addr[7067]= 2147470025;
assign addr[7068]= 2126796855;
assign addr[7069]= 2063024031;
assign addr[7070]= 1957443913;
assign addr[7071]= 1812196087;
assign addr[7072]= 1630224009;
assign addr[7073]= 1415215352;
assign addr[7074]= 1171527280;
assign addr[7075]= 904098143;
assign addr[7076]= 618347408;
assign addr[7077]= 320065829;
assign addr[7078]= 15298099;
assign addr[7079]= -289779648;
assign addr[7080]= -588984994;
assign addr[7081]= -876254528;
assign addr[7082]= -1145766716;
assign addr[7083]= -1392059879;
assign addr[7084]= -1610142873;
assign addr[7085]= -1795596234;
assign addr[7086]= -1944661739;
assign addr[7087]= -2054318569;
assign addr[7088]= -2122344521;
assign addr[7089]= -2147361045;
assign addr[7090]= -2128861181;
assign addr[7091]= -2067219829;
assign addr[7092]= -1963686155;
assign addr[7093]= -1820358275;
assign addr[7094]= -1640140734;
assign addr[7095]= -1426685652;
assign addr[7096]= -1184318708;
assign addr[7097]= -917951481;
assign addr[7098]= -632981917;
assign addr[7099]= -335184940;
assign addr[7100]= -30595422;
assign addr[7101]= 274614114;
assign addr[7102]= 574258580;
assign addr[7103]= 862265664;
assign addr[7104]= 1132798888;
assign addr[7105]= 1380375881;
assign addr[7106]= 1599979481;
assign addr[7107]= 1787159411;
assign addr[7108]= 1938122457;
assign addr[7109]= 2049809346;
assign addr[7110]= 2119956737;
assign addr[7111]= 2147143090;
assign addr[7112]= 2130817471;
assign addr[7113]= 2071310720;
assign addr[7114]= 1969828744;
assign addr[7115]= 1828428082;
assign addr[7116]= 1649974225;
assign addr[7117]= 1438083551;
assign addr[7118]= 1197050035;
assign addr[7119]= 931758235;
assign addr[7120]= 647584304;
assign addr[7121]= 350287041;
assign addr[7122]= 45891193;
assign addr[7123]= -259434643;
assign addr[7124]= -559503022;
assign addr[7125]= -848233042;
assign addr[7126]= -1119773573;
assign addr[7127]= -1368621831;
assign addr[7128]= -1589734894;
assign addr[7129]= -1778631892;
assign addr[7130]= -1931484818;
assign addr[7131]= -2045196100;
assign addr[7132]= -2117461370;
assign addr[7133]= -2146816171;
assign addr[7134]= -2132665626;
assign addr[7135]= -2075296495;
assign addr[7136]= -1975871368;
assign addr[7137]= -1836405100;
assign addr[7138]= -1659723983;
assign addr[7139]= -1449408469;
assign addr[7140]= -1209720613;
assign addr[7141]= -945517704;
assign addr[7142]= -662153826;
assign addr[7143]= -365371365;
assign addr[7144]= -61184634;
assign addr[7145]= 244242007;
assign addr[7146]= 544719071;
assign addr[7147]= 834157373;
assign addr[7148]= 1106691431;
assign addr[7149]= 1356798326;
assign addr[7150]= 1579409630;
assign addr[7151]= 1770014111;
assign addr[7152]= 1924749160;
assign addr[7153]= 2040479063;
assign addr[7154]= 2114858546;
assign addr[7155]= 2146380306;
assign addr[7156]= 2134405552;
assign addr[7157]= 2079176953;
assign addr[7158]= 1981813720;
assign addr[7159]= 1844288924;
assign addr[7160]= 1669389513;
assign addr[7161]= 1460659832;
assign addr[7162]= 1222329801;
assign addr[7163]= 959229189;
assign addr[7164]= 676689746;
assign addr[7165]= 380437148;
assign addr[7166]= 76474970;
assign addr[7167]= -229036977;
assign addr[7168]= -529907477;
assign addr[7169]= -820039373;
assign addr[7170]= -1093553126;
assign addr[7171]= -1344905966;
assign addr[7172]= -1569004214;
assign addr[7173]= -1761306505;
assign addr[7174]= -1917915825;
assign addr[7175]= -2035658475;
assign addr[7176]= -2112148396;
assign addr[7177]= -2145835515;
assign addr[7178]= -2136037160;
assign addr[7179]= -2082951896;
assign addr[7180]= -1987655498;
assign addr[7181]= -1852079154;
assign addr[7182]= -1678970324;
assign addr[7183]= -1471837070;
assign addr[7184]= -1234876957;
assign addr[7185]= -972891995;
assign addr[7186]= -691191324;
assign addr[7187]= -395483624;
assign addr[7188]= -91761426;
assign addr[7189]= 213820322;
assign addr[7190]= 515068990;
assign addr[7191]= 805879757;
assign addr[7192]= 1080359326;
assign addr[7193]= 1332945355;
assign addr[7194]= 1558519173;
assign addr[7195]= 1752509516;
assign addr[7196]= 1910985158;
assign addr[7197]= 2030734582;
assign addr[7198]= 2109331059;
assign addr[7199]= 2145181827;
assign addr[7200]= 2137560369;
assign addr[7201]= 2086621133;
assign addr[7202]= 1993396407;
assign addr[7203]= 1859775393;
assign addr[7204]= 1688465931;
assign addr[7205]= 1482939614;
assign addr[7206]= 1247361445;
assign addr[7207]= 986505429;
assign addr[7208]= 705657826;
assign addr[7209]= 410510029;
assign addr[7210]= 107043224;
assign addr[7211]= -198592817;
assign addr[7212]= -500204365;
assign addr[7213]= -791679244;
assign addr[7214]= -1067110699;
assign addr[7215]= -1320917099;
assign addr[7216]= -1547955041;
assign addr[7217]= -1743623590;
assign addr[7218]= -1903957513;
assign addr[7219]= -2025707632;
assign addr[7220]= -2106406677;
assign addr[7221]= -2144419275;
assign addr[7222]= -2138975100;
assign addr[7223]= -2090184478;
assign addr[7224]= -1999036154;
assign addr[7225]= -1867377253;
assign addr[7226]= -1697875851;
assign addr[7227]= -1493966902;
assign addr[7228]= -1259782632;
assign addr[7229]= -1000068799;
assign addr[7230]= -720088517;
assign addr[7231]= -425515602;
assign addr[7232]= -122319591;
assign addr[7233]= 183355234;
assign addr[7234]= 485314355;
assign addr[7235]= 777438554;
assign addr[7236]= 1053807919;
assign addr[7237]= 1308821808;
assign addr[7238]= 1537312353;
assign addr[7239]= 1734649179;
assign addr[7240]= 1896833245;
assign addr[7241]= 2020577882;
assign addr[7242]= 2103375398;
assign addr[7243]= 2143547897;
assign addr[7244]= 2140281282;
assign addr[7245]= 2093641749;
assign addr[7246]= 2004574453;
assign addr[7247]= 1874884346;
assign addr[7248]= 1707199606;
assign addr[7249]= 1504918373;
assign addr[7250]= 1272139887;
assign addr[7251]= 1013581418;
assign addr[7252]= 734482665;
assign addr[7253]= 440499581;
assign addr[7254]= 137589750;
assign addr[7255]= -168108346;
assign addr[7256]= -470399716;
assign addr[7257]= -763158411;
assign addr[7258]= -1040451659;
assign addr[7259]= -1296660098;
assign addr[7260]= -1526591649;
assign addr[7261]= -1725586737;
assign addr[7262]= -1889612716;
assign addr[7263]= -2015345591;
assign addr[7264]= -2100237377;
assign addr[7265]= -2142567738;
assign addr[7266]= -2141478848;
assign addr[7267]= -2096992772;
assign addr[7268]= -2010011024;
assign addr[7269]= -1882296293;
assign addr[7270]= -1716436725;
assign addr[7271]= -1515793473;
assign addr[7272]= -1284432584;
assign addr[7273]= -1027042599;
assign addr[7274]= -748839539;
assign addr[7275]= -455461206;
assign addr[7276]= -152852926;
assign addr[7277]= 152852926;
assign addr[7278]= 455461206;
assign addr[7279]= 748839539;
assign addr[7280]= 1027042599;
assign addr[7281]= 1284432584;
assign addr[7282]= 1515793473;
assign addr[7283]= 1716436725;
assign addr[7284]= 1882296293;
assign addr[7285]= 2010011024;
assign addr[7286]= 2096992772;
assign addr[7287]= 2141478848;
assign addr[7288]= 2142567738;
assign addr[7289]= 2100237377;
assign addr[7290]= 2015345591;
assign addr[7291]= 1889612716;
assign addr[7292]= 1725586737;
assign addr[7293]= 1526591649;
assign addr[7294]= 1296660098;
assign addr[7295]= 1040451659;
assign addr[7296]= 763158411;
assign addr[7297]= 470399716;
assign addr[7298]= 168108346;
assign addr[7299]= -137589750;
assign addr[7300]= -440499581;
assign addr[7301]= -734482665;
assign addr[7302]= -1013581418;
assign addr[7303]= -1272139887;
assign addr[7304]= -1504918373;
assign addr[7305]= -1707199606;
assign addr[7306]= -1874884346;
assign addr[7307]= -2004574453;
assign addr[7308]= -2093641749;
assign addr[7309]= -2140281282;
assign addr[7310]= -2143547897;
assign addr[7311]= -2103375398;
assign addr[7312]= -2020577882;
assign addr[7313]= -1896833245;
assign addr[7314]= -1734649179;
assign addr[7315]= -1537312353;
assign addr[7316]= -1308821808;
assign addr[7317]= -1053807919;
assign addr[7318]= -777438554;
assign addr[7319]= -485314355;
assign addr[7320]= -183355234;
assign addr[7321]= 122319591;
assign addr[7322]= 425515602;
assign addr[7323]= 720088517;
assign addr[7324]= 1000068799;
assign addr[7325]= 1259782632;
assign addr[7326]= 1493966902;
assign addr[7327]= 1697875851;
assign addr[7328]= 1867377253;
assign addr[7329]= 1999036154;
assign addr[7330]= 2090184478;
assign addr[7331]= 2138975100;
assign addr[7332]= 2144419275;
assign addr[7333]= 2106406677;
assign addr[7334]= 2025707632;
assign addr[7335]= 1903957513;
assign addr[7336]= 1743623590;
assign addr[7337]= 1547955041;
assign addr[7338]= 1320917099;
assign addr[7339]= 1067110699;
assign addr[7340]= 791679244;
assign addr[7341]= 500204365;
assign addr[7342]= 198592817;
assign addr[7343]= -107043224;
assign addr[7344]= -410510029;
assign addr[7345]= -705657826;
assign addr[7346]= -986505429;
assign addr[7347]= -1247361445;
assign addr[7348]= -1482939614;
assign addr[7349]= -1688465931;
assign addr[7350]= -1859775393;
assign addr[7351]= -1993396407;
assign addr[7352]= -2086621133;
assign addr[7353]= -2137560369;
assign addr[7354]= -2145181827;
assign addr[7355]= -2109331059;
assign addr[7356]= -2030734582;
assign addr[7357]= -1910985158;
assign addr[7358]= -1752509516;
assign addr[7359]= -1558519173;
assign addr[7360]= -1332945355;
assign addr[7361]= -1080359326;
assign addr[7362]= -805879757;
assign addr[7363]= -515068990;
assign addr[7364]= -213820322;
assign addr[7365]= 91761426;
assign addr[7366]= 395483624;
assign addr[7367]= 691191324;
assign addr[7368]= 972891995;
assign addr[7369]= 1234876957;
assign addr[7370]= 1471837070;
assign addr[7371]= 1678970324;
assign addr[7372]= 1852079154;
assign addr[7373]= 1987655498;
assign addr[7374]= 2082951896;
assign addr[7375]= 2136037160;
assign addr[7376]= 2145835515;
assign addr[7377]= 2112148396;
assign addr[7378]= 2035658475;
assign addr[7379]= 1917915825;
assign addr[7380]= 1761306505;
assign addr[7381]= 1569004214;
assign addr[7382]= 1344905966;
assign addr[7383]= 1093553126;
assign addr[7384]= 820039373;
assign addr[7385]= 529907477;
assign addr[7386]= 229036977;
assign addr[7387]= -76474970;
assign addr[7388]= -380437148;
assign addr[7389]= -676689746;
assign addr[7390]= -959229189;
assign addr[7391]= -1222329801;
assign addr[7392]= -1460659832;
assign addr[7393]= -1669389513;
assign addr[7394]= -1844288924;
assign addr[7395]= -1981813720;
assign addr[7396]= -2079176953;
assign addr[7397]= -2134405552;
assign addr[7398]= -2146380306;
assign addr[7399]= -2114858546;
assign addr[7400]= -2040479063;
assign addr[7401]= -1924749160;
assign addr[7402]= -1770014111;
assign addr[7403]= -1579409630;
assign addr[7404]= -1356798326;
assign addr[7405]= -1106691431;
assign addr[7406]= -834157373;
assign addr[7407]= -544719071;
assign addr[7408]= -244242007;
assign addr[7409]= 61184634;
assign addr[7410]= 365371365;
assign addr[7411]= 662153826;
assign addr[7412]= 945517704;
assign addr[7413]= 1209720613;
assign addr[7414]= 1449408469;
assign addr[7415]= 1659723983;
assign addr[7416]= 1836405100;
assign addr[7417]= 1975871368;
assign addr[7418]= 2075296495;
assign addr[7419]= 2132665626;
assign addr[7420]= 2146816171;
assign addr[7421]= 2117461370;
assign addr[7422]= 2045196100;
assign addr[7423]= 1931484818;
assign addr[7424]= 1778631892;
assign addr[7425]= 1589734894;
assign addr[7426]= 1368621831;
assign addr[7427]= 1119773573;
assign addr[7428]= 848233042;
assign addr[7429]= 559503022;
assign addr[7430]= 259434643;
assign addr[7431]= -45891193;
assign addr[7432]= -350287041;
assign addr[7433]= -647584304;
assign addr[7434]= -931758235;
assign addr[7435]= -1197050035;
assign addr[7436]= -1438083551;
assign addr[7437]= -1649974225;
assign addr[7438]= -1828428082;
assign addr[7439]= -1969828744;
assign addr[7440]= -2071310720;
assign addr[7441]= -2130817471;
assign addr[7442]= -2147143090;
assign addr[7443]= -2119956737;
assign addr[7444]= -2049809346;
assign addr[7445]= -1938122457;
assign addr[7446]= -1787159411;
assign addr[7447]= -1599979481;
assign addr[7448]= -1380375881;
assign addr[7449]= -1132798888;
assign addr[7450]= -862265664;
assign addr[7451]= -574258580;
assign addr[7452]= -274614114;
assign addr[7453]= 30595422;
assign addr[7454]= 335184940;
assign addr[7455]= 632981917;
assign addr[7456]= 917951481;
assign addr[7457]= 1184318708;
assign addr[7458]= 1426685652;
assign addr[7459]= 1640140734;
assign addr[7460]= 1820358275;
assign addr[7461]= 1963686155;
assign addr[7462]= 2067219829;
assign addr[7463]= 2128861181;
assign addr[7464]= 2147361045;
assign addr[7465]= 2122344521;
assign addr[7466]= 2054318569;
assign addr[7467]= 1944661739;
assign addr[7468]= 1795596234;
assign addr[7469]= 1610142873;
assign addr[7470]= 1392059879;
assign addr[7471]= 1145766716;
assign addr[7472]= 876254528;
assign addr[7473]= 588984994;
assign addr[7474]= 289779648;
assign addr[7475]= -15298099;
assign addr[7476]= -320065829;
assign addr[7477]= -618347408;
assign addr[7478]= -904098143;
assign addr[7479]= -1171527280;
assign addr[7480]= -1415215352;
assign addr[7481]= -1630224009;
assign addr[7482]= -1812196087;
assign addr[7483]= -1957443913;
assign addr[7484]= -2063024031;
assign addr[7485]= -2126796855;
assign addr[7486]= -2147470025;
assign addr[7487]= -2124624598;
assign addr[7488]= -2058723538;
assign addr[7489]= -1951102334;
assign addr[7490]= -1803941934;
assign addr[7491]= -1620224553;
assign addr[7492]= -1403673233;
assign addr[7493]= -1158676398;
assign addr[7494]= -890198924;
assign addr[7495]= -603681519;
assign addr[7496]= -304930476;
assign addr[7497]= 0;
assign addr[7498]= 304930476;
assign addr[7499]= 603681519;
assign addr[7500]= 890198924;
assign addr[7501]= 1158676398;
assign addr[7502]= 1403673233;
assign addr[7503]= 1620224553;
assign addr[7504]= 1803941934;
assign addr[7505]= 1951102334;
assign addr[7506]= 2058723538;
assign addr[7507]= 2124624598;
assign addr[7508]= 2147470025;
assign addr[7509]= 2126796855;
assign addr[7510]= 2063024031;
assign addr[7511]= 1957443913;
assign addr[7512]= 1812196087;
assign addr[7513]= 1630224009;
assign addr[7514]= 1415215352;
assign addr[7515]= 1171527280;
assign addr[7516]= 904098143;
assign addr[7517]= 618347408;
assign addr[7518]= 320065829;
assign addr[7519]= 15298099;
assign addr[7520]= -289779648;
assign addr[7521]= -588984994;
assign addr[7522]= -876254528;
assign addr[7523]= -1145766716;
assign addr[7524]= -1392059879;
assign addr[7525]= -1610142873;
assign addr[7526]= -1795596234;
assign addr[7527]= -1944661739;
assign addr[7528]= -2054318569;
assign addr[7529]= -2122344521;
assign addr[7530]= -2147361045;
assign addr[7531]= -2128861181;
assign addr[7532]= -2067219829;
assign addr[7533]= -1963686155;
assign addr[7534]= -1820358275;
assign addr[7535]= -1640140734;
assign addr[7536]= -1426685652;
assign addr[7537]= -1184318708;
assign addr[7538]= -917951481;
assign addr[7539]= -632981917;
assign addr[7540]= -335184940;
assign addr[7541]= -30595422;
assign addr[7542]= 274614114;
assign addr[7543]= 574258580;
assign addr[7544]= 862265664;
assign addr[7545]= 1132798888;
assign addr[7546]= 1380375881;
assign addr[7547]= 1599979481;
assign addr[7548]= 1787159411;
assign addr[7549]= 1938122457;
assign addr[7550]= 2049809346;
assign addr[7551]= 2119956737;
assign addr[7552]= 2147143090;
assign addr[7553]= 2130817471;
assign addr[7554]= 2071310720;
assign addr[7555]= 1969828744;
assign addr[7556]= 1828428082;
assign addr[7557]= 1649974225;
assign addr[7558]= 1438083551;
assign addr[7559]= 1197050035;
assign addr[7560]= 931758235;
assign addr[7561]= 647584304;
assign addr[7562]= 350287041;
assign addr[7563]= 45891193;
assign addr[7564]= -259434643;
assign addr[7565]= -559503022;
assign addr[7566]= -848233042;
assign addr[7567]= -1119773573;
assign addr[7568]= -1368621831;
assign addr[7569]= -1589734894;
assign addr[7570]= -1778631892;
assign addr[7571]= -1931484818;
assign addr[7572]= -2045196100;
assign addr[7573]= -2117461370;
assign addr[7574]= -2146816171;
assign addr[7575]= -2132665626;
assign addr[7576]= -2075296495;
assign addr[7577]= -1975871368;
assign addr[7578]= -1836405100;
assign addr[7579]= -1659723983;
assign addr[7580]= -1449408469;
assign addr[7581]= -1209720613;
assign addr[7582]= -945517704;
assign addr[7583]= -662153826;
assign addr[7584]= -365371365;
assign addr[7585]= -61184634;
assign addr[7586]= 244242007;
assign addr[7587]= 544719071;
assign addr[7588]= 834157373;
assign addr[7589]= 1106691431;
assign addr[7590]= 1356798326;
assign addr[7591]= 1579409630;
assign addr[7592]= 1770014111;
assign addr[7593]= 1924749160;
assign addr[7594]= 2040479063;
assign addr[7595]= 2114858546;
assign addr[7596]= 2146380306;
assign addr[7597]= 2134405552;
assign addr[7598]= 2079176953;
assign addr[7599]= 1981813720;
assign addr[7600]= 1844288924;
assign addr[7601]= 1669389513;
assign addr[7602]= 1460659832;
assign addr[7603]= 1222329801;
assign addr[7604]= 959229189;
assign addr[7605]= 676689746;
assign addr[7606]= 380437148;
assign addr[7607]= 76474970;
assign addr[7608]= -229036977;
assign addr[7609]= -529907477;
assign addr[7610]= -820039373;
assign addr[7611]= -1093553126;
assign addr[7612]= -1344905966;
assign addr[7613]= -1569004214;
assign addr[7614]= -1761306505;
assign addr[7615]= -1917915825;
assign addr[7616]= -2035658475;
assign addr[7617]= -2112148396;
assign addr[7618]= -2145835515;
assign addr[7619]= -2136037160;
assign addr[7620]= -2082951896;
assign addr[7621]= -1987655498;
assign addr[7622]= -1852079154;
assign addr[7623]= -1678970324;
assign addr[7624]= -1471837070;
assign addr[7625]= -1234876957;
assign addr[7626]= -972891995;
assign addr[7627]= -691191324;
assign addr[7628]= -395483624;
assign addr[7629]= -91761426;
assign addr[7630]= 213820322;
assign addr[7631]= 515068990;
assign addr[7632]= 805879757;
assign addr[7633]= 1080359326;
assign addr[7634]= 1332945355;
assign addr[7635]= 1558519173;
assign addr[7636]= 1752509516;
assign addr[7637]= 1910985158;
assign addr[7638]= 2030734582;
assign addr[7639]= 2109331059;
assign addr[7640]= 2145181827;
assign addr[7641]= 2137560369;
assign addr[7642]= 2086621133;
assign addr[7643]= 1993396407;
assign addr[7644]= 1859775393;
assign addr[7645]= 1688465931;
assign addr[7646]= 1482939614;
assign addr[7647]= 1247361445;
assign addr[7648]= 986505429;
assign addr[7649]= 705657826;
assign addr[7650]= 410510029;
assign addr[7651]= 107043224;
assign addr[7652]= -198592817;
assign addr[7653]= -500204365;
assign addr[7654]= -791679244;
assign addr[7655]= -1067110699;
assign addr[7656]= -1320917099;
assign addr[7657]= -1547955041;
assign addr[7658]= -1743623590;
assign addr[7659]= -1903957513;
assign addr[7660]= -2025707632;
assign addr[7661]= -2106406677;
assign addr[7662]= -2144419275;
assign addr[7663]= -2138975100;
assign addr[7664]= -2090184478;
assign addr[7665]= -1999036154;
assign addr[7666]= -1867377253;
assign addr[7667]= -1697875851;
assign addr[7668]= -1493966902;
assign addr[7669]= -1259782632;
assign addr[7670]= -1000068799;
assign addr[7671]= -720088517;
assign addr[7672]= -425515602;
assign addr[7673]= -122319591;
assign addr[7674]= 183355234;
assign addr[7675]= 485314355;
assign addr[7676]= 777438554;
assign addr[7677]= 1053807919;
assign addr[7678]= 1308821808;
assign addr[7679]= 1537312353;
assign addr[7680]= 1734649179;
assign addr[7681]= 1896833245;
assign addr[7682]= 2020577882;
assign addr[7683]= 2103375398;
assign addr[7684]= 2143547897;
assign addr[7685]= 2140281282;
assign addr[7686]= 2093641749;
assign addr[7687]= 2004574453;
assign addr[7688]= 1874884346;
assign addr[7689]= 1707199606;
assign addr[7690]= 1504918373;
assign addr[7691]= 1272139887;
assign addr[7692]= 1013581418;
assign addr[7693]= 734482665;
assign addr[7694]= 440499581;
assign addr[7695]= 137589750;
assign addr[7696]= -168108346;
assign addr[7697]= -470399716;
assign addr[7698]= -763158411;
assign addr[7699]= -1040451659;
assign addr[7700]= -1296660098;
assign addr[7701]= -1526591649;
assign addr[7702]= -1725586737;
assign addr[7703]= -1889612716;
assign addr[7704]= -2015345591;
assign addr[7705]= -2100237377;
assign addr[7706]= -2142567738;
assign addr[7707]= -2141478848;
assign addr[7708]= -2096992772;
assign addr[7709]= -2010011024;
assign addr[7710]= -1882296293;
assign addr[7711]= -1716436725;
assign addr[7712]= -1515793473;
assign addr[7713]= -1284432584;
assign addr[7714]= -1027042599;
assign addr[7715]= -748839539;
assign addr[7716]= -455461206;
assign addr[7717]= -152852926;
assign addr[7718]= 152852926;
assign addr[7719]= 455461206;
assign addr[7720]= 748839539;
assign addr[7721]= 1027042599;
assign addr[7722]= 1284432584;
assign addr[7723]= 1515793473;
assign addr[7724]= 1716436725;
assign addr[7725]= 1882296293;
assign addr[7726]= 2010011024;
assign addr[7727]= 2096992772;
assign addr[7728]= 2141478848;
assign addr[7729]= 2142567738;
assign addr[7730]= 2100237377;
assign addr[7731]= 2015345591;
assign addr[7732]= 1889612716;
assign addr[7733]= 1725586737;
assign addr[7734]= 1526591649;
assign addr[7735]= 1296660098;
assign addr[7736]= 1040451659;
assign addr[7737]= 763158411;
assign addr[7738]= 470399716;
assign addr[7739]= 168108346;
assign addr[7740]= -137589750;
assign addr[7741]= -440499581;
assign addr[7742]= -734482665;
assign addr[7743]= -1013581418;
assign addr[7744]= -1272139887;
assign addr[7745]= -1504918373;
assign addr[7746]= -1707199606;
assign addr[7747]= -1874884346;
assign addr[7748]= -2004574453;
assign addr[7749]= -2093641749;
assign addr[7750]= -2140281282;
assign addr[7751]= -2143547897;
assign addr[7752]= -2103375398;
assign addr[7753]= -2020577882;
assign addr[7754]= -1896833245;
assign addr[7755]= -1734649179;
assign addr[7756]= -1537312353;
assign addr[7757]= -1308821808;
assign addr[7758]= -1053807919;
assign addr[7759]= -777438554;
assign addr[7760]= -485314355;
assign addr[7761]= -183355234;
assign addr[7762]= 122319591;
assign addr[7763]= 425515602;
assign addr[7764]= 720088517;
assign addr[7765]= 1000068799;
assign addr[7766]= 1259782632;
assign addr[7767]= 1493966902;
assign addr[7768]= 1697875851;
assign addr[7769]= 1867377253;
assign addr[7770]= 1999036154;
assign addr[7771]= 2090184478;
assign addr[7772]= 2138975100;
assign addr[7773]= 2144419275;
assign addr[7774]= 2106406677;
assign addr[7775]= 2025707632;
assign addr[7776]= 1903957513;
assign addr[7777]= 1743623590;
assign addr[7778]= 1547955041;
assign addr[7779]= 1320917099;
assign addr[7780]= 1067110699;
assign addr[7781]= 791679244;
assign addr[7782]= 500204365;
assign addr[7783]= 198592817;
assign addr[7784]= -107043224;
assign addr[7785]= -410510029;
assign addr[7786]= -705657826;
assign addr[7787]= -986505429;
assign addr[7788]= -1247361445;
assign addr[7789]= -1482939614;
assign addr[7790]= -1688465931;
assign addr[7791]= -1859775393;
assign addr[7792]= -1993396407;
assign addr[7793]= -2086621133;
assign addr[7794]= -2137560369;
assign addr[7795]= -2145181827;
assign addr[7796]= -2109331059;
assign addr[7797]= -2030734582;
assign addr[7798]= -1910985158;
assign addr[7799]= -1752509516;
assign addr[7800]= -1558519173;
assign addr[7801]= -1332945355;
assign addr[7802]= -1080359326;
assign addr[7803]= -805879757;
assign addr[7804]= -515068990;
assign addr[7805]= -213820322;
assign addr[7806]= 91761426;
assign addr[7807]= 395483624;
assign addr[7808]= 691191324;
assign addr[7809]= 972891995;
assign addr[7810]= 1234876957;
assign addr[7811]= 1471837070;
assign addr[7812]= 1678970324;
assign addr[7813]= 1852079154;
assign addr[7814]= 1987655498;
assign addr[7815]= 2082951896;
assign addr[7816]= 2136037160;
assign addr[7817]= 2145835515;
assign addr[7818]= 2112148396;
assign addr[7819]= 2035658475;
assign addr[7820]= 1917915825;
assign addr[7821]= 1761306505;
assign addr[7822]= 1569004214;
assign addr[7823]= 1344905966;
assign addr[7824]= 1093553126;
assign addr[7825]= 820039373;
assign addr[7826]= 529907477;
assign addr[7827]= 229036977;
assign addr[7828]= -76474970;
assign addr[7829]= -380437148;
assign addr[7830]= -676689746;
assign addr[7831]= -959229189;
assign addr[7832]= -1222329801;
assign addr[7833]= -1460659832;
assign addr[7834]= -1669389513;
assign addr[7835]= -1844288924;
assign addr[7836]= -1981813720;
assign addr[7837]= -2079176953;
assign addr[7838]= -2134405552;
assign addr[7839]= -2146380306;
assign addr[7840]= -2114858546;
assign addr[7841]= -2040479063;
assign addr[7842]= -1924749160;
assign addr[7843]= -1770014111;
assign addr[7844]= -1579409630;
assign addr[7845]= -1356798326;
assign addr[7846]= -1106691431;
assign addr[7847]= -834157373;
assign addr[7848]= -544719071;
assign addr[7849]= -244242007;
assign addr[7850]= 61184634;
assign addr[7851]= 365371365;
assign addr[7852]= 662153826;
assign addr[7853]= 945517704;
assign addr[7854]= 1209720613;
assign addr[7855]= 1449408469;
assign addr[7856]= 1659723983;
assign addr[7857]= 1836405100;
assign addr[7858]= 1975871368;
assign addr[7859]= 2075296495;
assign addr[7860]= 2132665626;
assign addr[7861]= 2146816171;
assign addr[7862]= 2117461370;
assign addr[7863]= 2045196100;
assign addr[7864]= 1931484818;
assign addr[7865]= 1778631892;
assign addr[7866]= 1589734894;
assign addr[7867]= 1368621831;
assign addr[7868]= 1119773573;
assign addr[7869]= 848233042;
assign addr[7870]= 559503022;
assign addr[7871]= 259434643;
assign addr[7872]= -45891193;
assign addr[7873]= -350287041;
assign addr[7874]= -647584304;
assign addr[7875]= -931758235;
assign addr[7876]= -1197050035;
assign addr[7877]= -1438083551;
assign addr[7878]= -1649974225;
assign addr[7879]= -1828428082;
assign addr[7880]= -1969828744;
assign addr[7881]= -2071310720;
assign addr[7882]= -2130817471;
assign addr[7883]= -2147143090;
assign addr[7884]= -2119956737;
assign addr[7885]= -2049809346;
assign addr[7886]= -1938122457;
assign addr[7887]= -1787159411;
assign addr[7888]= -1599979481;
assign addr[7889]= -1380375881;
assign addr[7890]= -1132798888;
assign addr[7891]= -862265664;
assign addr[7892]= -574258580;
assign addr[7893]= -274614114;
assign addr[7894]= 30595422;
assign addr[7895]= 335184940;
assign addr[7896]= 632981917;
assign addr[7897]= 917951481;
assign addr[7898]= 1184318708;
assign addr[7899]= 1426685652;
assign addr[7900]= 1640140734;
assign addr[7901]= 1820358275;
assign addr[7902]= 1963686155;
assign addr[7903]= 2067219829;
assign addr[7904]= 2128861181;
assign addr[7905]= 2147361045;
assign addr[7906]= 2122344521;
assign addr[7907]= 2054318569;
assign addr[7908]= 1944661739;
assign addr[7909]= 1795596234;
assign addr[7910]= 1610142873;
assign addr[7911]= 1392059879;
assign addr[7912]= 1145766716;
assign addr[7913]= 876254528;
assign addr[7914]= 588984994;
assign addr[7915]= 289779648;
assign addr[7916]= -15298099;
assign addr[7917]= -320065829;
assign addr[7918]= -618347408;
assign addr[7919]= -904098143;
assign addr[7920]= -1171527280;
assign addr[7921]= -1415215352;
assign addr[7922]= -1630224009;
assign addr[7923]= -1812196087;
assign addr[7924]= -1957443913;
assign addr[7925]= -2063024031;
assign addr[7926]= -2126796855;
assign addr[7927]= -2147470025;
assign addr[7928]= -2124624598;
assign addr[7929]= -2058723538;
assign addr[7930]= -1951102334;
assign addr[7931]= -1803941934;
assign addr[7932]= -1620224553;
assign addr[7933]= -1403673233;
assign addr[7934]= -1158676398;
assign addr[7935]= -890198924;
assign addr[7936]= -603681519;
assign addr[7937]= -304930476;
assign addr[7938]= 0;
assign addr[7939]= 304930476;
assign addr[7940]= 603681519;
assign addr[7941]= 890198924;
assign addr[7942]= 1158676398;
assign addr[7943]= 1403673233;
assign addr[7944]= 1620224553;
assign addr[7945]= 1803941934;
assign addr[7946]= 1951102334;
assign addr[7947]= 2058723538;
assign addr[7948]= 2124624598;
assign addr[7949]= 2147470025;
assign addr[7950]= 2126796855;
assign addr[7951]= 2063024031;
assign addr[7952]= 1957443913;
assign addr[7953]= 1812196087;
assign addr[7954]= 1630224009;
assign addr[7955]= 1415215352;
assign addr[7956]= 1171527280;
assign addr[7957]= 904098143;
assign addr[7958]= 618347408;
assign addr[7959]= 320065829;
assign addr[7960]= 15298099;
assign addr[7961]= -289779648;
assign addr[7962]= -588984994;
assign addr[7963]= -876254528;
assign addr[7964]= -1145766716;
assign addr[7965]= -1392059879;
assign addr[7966]= -1610142873;
assign addr[7967]= -1795596234;
assign addr[7968]= -1944661739;
assign addr[7969]= -2054318569;
assign addr[7970]= -2122344521;
assign addr[7971]= -2147361045;
assign addr[7972]= -2128861181;
assign addr[7973]= -2067219829;
assign addr[7974]= -1963686155;
assign addr[7975]= -1820358275;
assign addr[7976]= -1640140734;
assign addr[7977]= -1426685652;
assign addr[7978]= -1184318708;
assign addr[7979]= -917951481;
assign addr[7980]= -632981917;
assign addr[7981]= -335184940;
assign addr[7982]= -30595422;
assign addr[7983]= 274614114;
assign addr[7984]= 574258580;
assign addr[7985]= 862265664;
assign addr[7986]= 1132798888;
assign addr[7987]= 1380375881;
assign addr[7988]= 1599979481;
assign addr[7989]= 1787159411;
assign addr[7990]= 1938122457;
assign addr[7991]= 2049809346;
assign addr[7992]= 2119956737;
assign addr[7993]= 2147143090;
assign addr[7994]= 2130817471;
assign addr[7995]= 2071310720;
assign addr[7996]= 1969828744;
assign addr[7997]= 1828428082;
assign addr[7998]= 1649974225;
assign addr[7999]= 1438083551;
assign addr[8000]= 1197050035;
assign addr[8001]= 931758235;
assign addr[8002]= 647584304;
assign addr[8003]= 350287041;
assign addr[8004]= 45891193;
assign addr[8005]= -259434643;
assign addr[8006]= -559503022;
assign addr[8007]= -848233042;
assign addr[8008]= -1119773573;
assign addr[8009]= -1368621831;
assign addr[8010]= -1589734894;
assign addr[8011]= -1778631892;
assign addr[8012]= -1931484818;
assign addr[8013]= -2045196100;
assign addr[8014]= -2117461370;
assign addr[8015]= -2146816171;
assign addr[8016]= -2132665626;
assign addr[8017]= -2075296495;
assign addr[8018]= -1975871368;
assign addr[8019]= -1836405100;
assign addr[8020]= -1659723983;
assign addr[8021]= -1449408469;
assign addr[8022]= -1209720613;
assign addr[8023]= -945517704;
assign addr[8024]= -662153826;
assign addr[8025]= -365371365;
assign addr[8026]= -61184634;
assign addr[8027]= 244242007;
assign addr[8028]= 544719071;
assign addr[8029]= 834157373;
assign addr[8030]= 1106691431;
assign addr[8031]= 1356798326;
assign addr[8032]= 1579409630;
assign addr[8033]= 1770014111;
assign addr[8034]= 1924749160;
assign addr[8035]= 2040479063;
assign addr[8036]= 2114858546;
assign addr[8037]= 2146380306;
assign addr[8038]= 2134405552;
assign addr[8039]= 2079176953;
assign addr[8040]= 1981813720;
assign addr[8041]= 1844288924;
assign addr[8042]= 1669389513;
assign addr[8043]= 1460659832;
assign addr[8044]= 1222329801;
assign addr[8045]= 959229189;
assign addr[8046]= 676689746;
assign addr[8047]= 380437148;
assign addr[8048]= 76474970;
assign addr[8049]= -229036977;
assign addr[8050]= -529907477;
assign addr[8051]= -820039373;
assign addr[8052]= -1093553126;
assign addr[8053]= -1344905966;
assign addr[8054]= -1569004214;
assign addr[8055]= -1761306505;
assign addr[8056]= -1917915825;
assign addr[8057]= -2035658475;
assign addr[8058]= -2112148396;
assign addr[8059]= -2145835515;
assign addr[8060]= -2136037160;
assign addr[8061]= -2082951896;
assign addr[8062]= -1987655498;
assign addr[8063]= -1852079154;
assign addr[8064]= -1678970324;
assign addr[8065]= -1471837070;
assign addr[8066]= -1234876957;
assign addr[8067]= -972891995;
assign addr[8068]= -691191324;
assign addr[8069]= -395483624;
assign addr[8070]= -91761426;
assign addr[8071]= 213820322;
assign addr[8072]= 515068990;
assign addr[8073]= 805879757;
assign addr[8074]= 1080359326;
assign addr[8075]= 1332945355;
assign addr[8076]= 1558519173;
assign addr[8077]= 1752509516;
assign addr[8078]= 1910985158;
assign addr[8079]= 2030734582;
assign addr[8080]= 2109331059;
assign addr[8081]= 2145181827;
assign addr[8082]= 2137560369;
assign addr[8083]= 2086621133;
assign addr[8084]= 1993396407;
assign addr[8085]= 1859775393;
assign addr[8086]= 1688465931;
assign addr[8087]= 1482939614;
assign addr[8088]= 1247361445;
assign addr[8089]= 986505429;
assign addr[8090]= 705657826;
assign addr[8091]= 410510029;
assign addr[8092]= 107043224;
assign addr[8093]= -198592817;
assign addr[8094]= -500204365;
assign addr[8095]= -791679244;
assign addr[8096]= -1067110699;
assign addr[8097]= -1320917099;
assign addr[8098]= -1547955041;
assign addr[8099]= -1743623590;
assign addr[8100]= -1903957513;
assign addr[8101]= -2025707632;
assign addr[8102]= -2106406677;
assign addr[8103]= -2144419275;
assign addr[8104]= -2138975100;
assign addr[8105]= -2090184478;
assign addr[8106]= -1999036154;
assign addr[8107]= -1867377253;
assign addr[8108]= -1697875851;
assign addr[8109]= -1493966902;
assign addr[8110]= -1259782632;
assign addr[8111]= -1000068799;
assign addr[8112]= -720088517;
assign addr[8113]= -425515602;
assign addr[8114]= -122319591;
assign addr[8115]= 183355234;
assign addr[8116]= 485314355;
assign addr[8117]= 777438554;
assign addr[8118]= 1053807919;
assign addr[8119]= 1308821808;
assign addr[8120]= 1537312353;
assign addr[8121]= 1734649179;
assign addr[8122]= 1896833245;
assign addr[8123]= 2020577882;
assign addr[8124]= 2103375398;
assign addr[8125]= 2143547897;
assign addr[8126]= 2140281282;
assign addr[8127]= 2093641749;
assign addr[8128]= 2004574453;
assign addr[8129]= 1874884346;
assign addr[8130]= 1707199606;
assign addr[8131]= 1504918373;
assign addr[8132]= 1272139887;
assign addr[8133]= 1013581418;
assign addr[8134]= 734482665;
assign addr[8135]= 440499581;
assign addr[8136]= 137589750;
assign addr[8137]= -168108346;
assign addr[8138]= -470399716;
assign addr[8139]= -763158411;
assign addr[8140]= -1040451659;
assign addr[8141]= -1296660098;
assign addr[8142]= -1526591649;
assign addr[8143]= -1725586737;
assign addr[8144]= -1889612716;
assign addr[8145]= -2015345591;
assign addr[8146]= -2100237377;
assign addr[8147]= -2142567738;
assign addr[8148]= -2141478848;
assign addr[8149]= -2096992772;
assign addr[8150]= -2010011024;
assign addr[8151]= -1882296293;
assign addr[8152]= -1716436725;
assign addr[8153]= -1515793473;
assign addr[8154]= -1284432584;
assign addr[8155]= -1027042599;
assign addr[8156]= -748839539;
assign addr[8157]= -455461206;
assign addr[8158]= -152852926;
assign addr[8159]= 152852926;
assign addr[8160]= 455461206;
assign addr[8161]= 748839539;
assign addr[8162]= 1027042599;
assign addr[8163]= 1284432584;
assign addr[8164]= 1515793473;
assign addr[8165]= 1716436725;
assign addr[8166]= 1882296293;
assign addr[8167]= 2010011024;
assign addr[8168]= 2096992772;
assign addr[8169]= 2141478848;
assign addr[8170]= 2142567738;
assign addr[8171]= 2100237377;
assign addr[8172]= 2015345591;
assign addr[8173]= 1889612716;
assign addr[8174]= 1725586737;
assign addr[8175]= 1526591649;
assign addr[8176]= 1296660098;
assign addr[8177]= 1040451659;
assign addr[8178]= 763158411;
assign addr[8179]= 470399716;
assign addr[8180]= 168108346;
assign addr[8181]= -137589750;
assign addr[8182]= -440499581;
assign addr[8183]= -734482665;
assign addr[8184]= -1013581418;
assign addr[8185]= -1272139887;
assign addr[8186]= -1504918373;
assign addr[8187]= -1707199606;
assign addr[8188]= -1874884346;
assign addr[8189]= -2004574453;
assign addr[8190]= -2093641749;
assign addr[8191]= -2140281282;
assign addr[8192]= -2143547897;
assign addr[8193]= -2103375398;
assign addr[8194]= -2020577882;
assign addr[8195]= -1896833245;
assign addr[8196]= -1734649179;
assign addr[8197]= -1537312353;
assign addr[8198]= -1308821808;
assign addr[8199]= -1053807919;
assign addr[8200]= -777438554;
assign addr[8201]= -485314355;
assign addr[8202]= -183355234;
assign addr[8203]= 122319591;
assign addr[8204]= 425515602;
assign addr[8205]= 720088517;
assign addr[8206]= 1000068799;
assign addr[8207]= 1259782632;
assign addr[8208]= 1493966902;
assign addr[8209]= 1697875851;
assign addr[8210]= 1867377253;
assign addr[8211]= 1999036154;
assign addr[8212]= 2090184478;
assign addr[8213]= 2138975100;
assign addr[8214]= 2144419275;
assign addr[8215]= 2106406677;
assign addr[8216]= 2025707632;
assign addr[8217]= 1903957513;
assign addr[8218]= 1743623590;
assign addr[8219]= 1547955041;
assign addr[8220]= 1320917099;
assign addr[8221]= 1067110699;
assign addr[8222]= 791679244;
assign addr[8223]= 500204365;
assign addr[8224]= 198592817;
assign addr[8225]= -107043224;
assign addr[8226]= -410510029;
assign addr[8227]= -705657826;
assign addr[8228]= -986505429;
assign addr[8229]= -1247361445;
assign addr[8230]= -1482939614;
assign addr[8231]= -1688465931;
assign addr[8232]= -1859775393;
assign addr[8233]= -1993396407;
assign addr[8234]= -2086621133;
assign addr[8235]= -2137560369;
assign addr[8236]= -2145181827;
assign addr[8237]= -2109331059;
assign addr[8238]= -2030734582;
assign addr[8239]= -1910985158;
assign addr[8240]= -1752509516;
assign addr[8241]= -1558519173;
assign addr[8242]= -1332945355;
assign addr[8243]= -1080359326;
assign addr[8244]= -805879757;
assign addr[8245]= -515068990;
assign addr[8246]= -213820322;
assign addr[8247]= 91761426;
assign addr[8248]= 395483624;
assign addr[8249]= 691191324;
assign addr[8250]= 972891995;
assign addr[8251]= 1234876957;
assign addr[8252]= 1471837070;
assign addr[8253]= 1678970324;
assign addr[8254]= 1852079154;
assign addr[8255]= 1987655498;
assign addr[8256]= 2082951896;
assign addr[8257]= 2136037160;
assign addr[8258]= 2145835515;
assign addr[8259]= 2112148396;
assign addr[8260]= 2035658475;
assign addr[8261]= 1917915825;
assign addr[8262]= 1761306505;
assign addr[8263]= 1569004214;
assign addr[8264]= 1344905966;
assign addr[8265]= 1093553126;
assign addr[8266]= 820039373;
assign addr[8267]= 529907477;
assign addr[8268]= 229036977;
assign addr[8269]= -76474970;
assign addr[8270]= -380437148;
assign addr[8271]= -676689746;
assign addr[8272]= -959229189;
assign addr[8273]= -1222329801;
assign addr[8274]= -1460659832;
assign addr[8275]= -1669389513;
assign addr[8276]= -1844288924;
assign addr[8277]= -1981813720;
assign addr[8278]= -2079176953;
assign addr[8279]= -2134405552;
assign addr[8280]= -2146380306;
assign addr[8281]= -2114858546;
assign addr[8282]= -2040479063;
assign addr[8283]= -1924749160;
assign addr[8284]= -1770014111;
assign addr[8285]= -1579409630;
assign addr[8286]= -1356798326;
assign addr[8287]= -1106691431;
assign addr[8288]= -834157373;
assign addr[8289]= -544719071;
assign addr[8290]= -244242007;
assign addr[8291]= 61184634;
assign addr[8292]= 365371365;
assign addr[8293]= 662153826;
assign addr[8294]= 945517704;
assign addr[8295]= 1209720613;
assign addr[8296]= 1449408469;
assign addr[8297]= 1659723983;
assign addr[8298]= 1836405100;
assign addr[8299]= 1975871368;
assign addr[8300]= 2075296495;
assign addr[8301]= 2132665626;
assign addr[8302]= 2146816171;
assign addr[8303]= 2117461370;
assign addr[8304]= 2045196100;
assign addr[8305]= 1931484818;
assign addr[8306]= 1778631892;
assign addr[8307]= 1589734894;
assign addr[8308]= 1368621831;
assign addr[8309]= 1119773573;
assign addr[8310]= 848233042;
assign addr[8311]= 559503022;
assign addr[8312]= 259434643;
assign addr[8313]= -45891193;
assign addr[8314]= -350287041;
assign addr[8315]= -647584304;
assign addr[8316]= -931758235;
assign addr[8317]= -1197050035;
assign addr[8318]= -1438083551;
assign addr[8319]= -1649974225;
assign addr[8320]= -1828428082;
assign addr[8321]= -1969828744;
assign addr[8322]= -2071310720;
assign addr[8323]= -2130817471;
assign addr[8324]= -2147143090;
assign addr[8325]= -2119956737;
assign addr[8326]= -2049809346;
assign addr[8327]= -1938122457;
assign addr[8328]= -1787159411;
assign addr[8329]= -1599979481;
assign addr[8330]= -1380375881;
assign addr[8331]= -1132798888;
assign addr[8332]= -862265664;
assign addr[8333]= -574258580;
assign addr[8334]= -274614114;
assign addr[8335]= 30595422;
assign addr[8336]= 335184940;
assign addr[8337]= 632981917;
assign addr[8338]= 917951481;
assign addr[8339]= 1184318708;
assign addr[8340]= 1426685652;
assign addr[8341]= 1640140734;
assign addr[8342]= 1820358275;
assign addr[8343]= 1963686155;
assign addr[8344]= 2067219829;
assign addr[8345]= 2128861181;
assign addr[8346]= 2147361045;
assign addr[8347]= 2122344521;
assign addr[8348]= 2054318569;
assign addr[8349]= 1944661739;
assign addr[8350]= 1795596234;
assign addr[8351]= 1610142873;
assign addr[8352]= 1392059879;
assign addr[8353]= 1145766716;
assign addr[8354]= 876254528;
assign addr[8355]= 588984994;
assign addr[8356]= 289779648;
assign addr[8357]= -15298099;
assign addr[8358]= -320065829;
assign addr[8359]= -618347408;
assign addr[8360]= -904098143;
assign addr[8361]= -1171527280;
assign addr[8362]= -1415215352;
assign addr[8363]= -1630224009;
assign addr[8364]= -1812196087;
assign addr[8365]= -1957443913;
assign addr[8366]= -2063024031;
assign addr[8367]= -2126796855;
assign addr[8368]= -2147470025;
assign addr[8369]= -2124624598;
assign addr[8370]= -2058723538;
assign addr[8371]= -1951102334;
assign addr[8372]= -1803941934;
assign addr[8373]= -1620224553;
assign addr[8374]= -1403673233;
assign addr[8375]= -1158676398;
assign addr[8376]= -890198924;
assign addr[8377]= -603681519;
assign addr[8378]= -304930476;
assign addr[8379]= 0;
assign addr[8380]= 304930476;
assign addr[8381]= 603681519;
assign addr[8382]= 890198924;
assign addr[8383]= 1158676398;
assign addr[8384]= 1403673233;
assign addr[8385]= 1620224553;
assign addr[8386]= 1803941934;
assign addr[8387]= 1951102334;
assign addr[8388]= 2058723538;
assign addr[8389]= 2124624598;
assign addr[8390]= 2147470025;
assign addr[8391]= 2126796855;
assign addr[8392]= 2063024031;
assign addr[8393]= 1957443913;
assign addr[8394]= 1812196087;
assign addr[8395]= 1630224009;
assign addr[8396]= 1415215352;
assign addr[8397]= 1171527280;
assign addr[8398]= 904098143;
assign addr[8399]= 618347408;
assign addr[8400]= 320065829;
assign addr[8401]= 15298099;
assign addr[8402]= -289779648;
assign addr[8403]= -588984994;
assign addr[8404]= -876254528;
assign addr[8405]= -1145766716;
assign addr[8406]= -1392059879;
assign addr[8407]= -1610142873;
assign addr[8408]= -1795596234;
assign addr[8409]= -1944661739;
assign addr[8410]= -2054318569;
assign addr[8411]= -2122344521;
assign addr[8412]= -2147361045;
assign addr[8413]= -2128861181;
assign addr[8414]= -2067219829;
assign addr[8415]= -1963686155;
assign addr[8416]= -1820358275;
assign addr[8417]= -1640140734;
assign addr[8418]= -1426685652;
assign addr[8419]= -1184318708;
assign addr[8420]= -917951481;
assign addr[8421]= -632981917;
assign addr[8422]= -335184940;
assign addr[8423]= -30595422;
assign addr[8424]= 274614114;
assign addr[8425]= 574258580;
assign addr[8426]= 862265664;
assign addr[8427]= 1132798888;
assign addr[8428]= 1380375881;
assign addr[8429]= 1599979481;
assign addr[8430]= 1787159411;
assign addr[8431]= 1938122457;
assign addr[8432]= 2049809346;
assign addr[8433]= 2119956737;
assign addr[8434]= 2147143090;
assign addr[8435]= 2130817471;
assign addr[8436]= 2071310720;
assign addr[8437]= 1969828744;
assign addr[8438]= 1828428082;
assign addr[8439]= 1649974225;
assign addr[8440]= 1438083551;
assign addr[8441]= 1197050035;
assign addr[8442]= 931758235;
assign addr[8443]= 647584304;
assign addr[8444]= 350287041;
assign addr[8445]= 45891193;
assign addr[8446]= -259434643;
assign addr[8447]= -559503022;
assign addr[8448]= -848233042;
assign addr[8449]= -1119773573;
assign addr[8450]= -1368621831;
assign addr[8451]= -1589734894;
assign addr[8452]= -1778631892;
assign addr[8453]= -1931484818;
assign addr[8454]= -2045196100;
assign addr[8455]= -2117461370;
assign addr[8456]= -2146816171;
assign addr[8457]= -2132665626;
assign addr[8458]= -2075296495;
assign addr[8459]= -1975871368;
assign addr[8460]= -1836405100;
assign addr[8461]= -1659723983;
assign addr[8462]= -1449408469;
assign addr[8463]= -1209720613;
assign addr[8464]= -945517704;
assign addr[8465]= -662153826;
assign addr[8466]= -365371365;
assign addr[8467]= -61184634;
assign addr[8468]= 244242007;
assign addr[8469]= 544719071;
assign addr[8470]= 834157373;
assign addr[8471]= 1106691431;
assign addr[8472]= 1356798326;
assign addr[8473]= 1579409630;
assign addr[8474]= 1770014111;
assign addr[8475]= 1924749160;
assign addr[8476]= 2040479063;
assign addr[8477]= 2114858546;
assign addr[8478]= 2146380306;
assign addr[8479]= 2134405552;
assign addr[8480]= 2079176953;
assign addr[8481]= 1981813720;
assign addr[8482]= 1844288924;
assign addr[8483]= 1669389513;
assign addr[8484]= 1460659832;
assign addr[8485]= 1222329801;
assign addr[8486]= 959229189;
assign addr[8487]= 676689746;
assign addr[8488]= 380437148;
assign addr[8489]= 76474970;
assign addr[8490]= -229036977;
assign addr[8491]= -529907477;
assign addr[8492]= -820039373;
assign addr[8493]= -1093553126;
assign addr[8494]= -1344905966;
assign addr[8495]= -1569004214;
assign addr[8496]= -1761306505;
assign addr[8497]= -1917915825;
assign addr[8498]= -2035658475;
assign addr[8499]= -2112148396;
assign addr[8500]= -2145835515;
assign addr[8501]= -2136037160;
assign addr[8502]= -2082951896;
assign addr[8503]= -1987655498;
assign addr[8504]= -1852079154;
assign addr[8505]= -1678970324;
assign addr[8506]= -1471837070;
assign addr[8507]= -1234876957;
assign addr[8508]= -972891995;
assign addr[8509]= -691191324;
assign addr[8510]= -395483624;
assign addr[8511]= -91761426;
assign addr[8512]= 213820322;
assign addr[8513]= 515068990;
assign addr[8514]= 805879757;
assign addr[8515]= 1080359326;
assign addr[8516]= 1332945355;
assign addr[8517]= 1558519173;
assign addr[8518]= 1752509516;
assign addr[8519]= 1910985158;
assign addr[8520]= 2030734582;
assign addr[8521]= 2109331059;
assign addr[8522]= 2145181827;
assign addr[8523]= 2137560369;
assign addr[8524]= 2086621133;
assign addr[8525]= 1993396407;
assign addr[8526]= 1859775393;
assign addr[8527]= 1688465931;
assign addr[8528]= 1482939614;
assign addr[8529]= 1247361445;
assign addr[8530]= 986505429;
assign addr[8531]= 705657826;
assign addr[8532]= 410510029;
assign addr[8533]= 107043224;
assign addr[8534]= -198592817;
assign addr[8535]= -500204365;
assign addr[8536]= -791679244;
assign addr[8537]= -1067110699;
assign addr[8538]= -1320917099;
assign addr[8539]= -1547955041;
assign addr[8540]= -1743623590;
assign addr[8541]= -1903957513;
assign addr[8542]= -2025707632;
assign addr[8543]= -2106406677;
assign addr[8544]= -2144419275;
assign addr[8545]= -2138975100;
assign addr[8546]= -2090184478;
assign addr[8547]= -1999036154;
assign addr[8548]= -1867377253;
assign addr[8549]= -1697875851;
assign addr[8550]= -1493966902;
assign addr[8551]= -1259782632;
assign addr[8552]= -1000068799;
assign addr[8553]= -720088517;
assign addr[8554]= -425515602;
assign addr[8555]= -122319591;
assign addr[8556]= 183355234;
assign addr[8557]= 485314355;
assign addr[8558]= 777438554;
assign addr[8559]= 1053807919;
assign addr[8560]= 1308821808;
assign addr[8561]= 1537312353;
assign addr[8562]= 1734649179;
assign addr[8563]= 1896833245;
assign addr[8564]= 2020577882;
assign addr[8565]= 2103375398;
assign addr[8566]= 2143547897;
assign addr[8567]= 2140281282;
assign addr[8568]= 2093641749;
assign addr[8569]= 2004574453;
assign addr[8570]= 1874884346;
assign addr[8571]= 1707199606;
assign addr[8572]= 1504918373;
assign addr[8573]= 1272139887;
assign addr[8574]= 1013581418;
assign addr[8575]= 734482665;
assign addr[8576]= 440499581;
assign addr[8577]= 137589750;
assign addr[8578]= -168108346;
assign addr[8579]= -470399716;
assign addr[8580]= -763158411;
assign addr[8581]= -1040451659;
assign addr[8582]= -1296660098;
assign addr[8583]= -1526591649;
assign addr[8584]= -1725586737;
assign addr[8585]= -1889612716;
assign addr[8586]= -2015345591;
assign addr[8587]= -2100237377;
assign addr[8588]= -2142567738;
assign addr[8589]= -2141478848;
assign addr[8590]= -2096992772;
assign addr[8591]= -2010011024;
assign addr[8592]= -1882296293;
assign addr[8593]= -1716436725;
assign addr[8594]= -1515793473;
assign addr[8595]= -1284432584;
assign addr[8596]= -1027042599;
assign addr[8597]= -748839539;
assign addr[8598]= -455461206;
assign addr[8599]= -152852926;
assign addr[8600]= 152852926;
assign addr[8601]= 455461206;
assign addr[8602]= 748839539;
assign addr[8603]= 1027042599;
assign addr[8604]= 1284432584;
assign addr[8605]= 1515793473;
assign addr[8606]= 1716436725;
assign addr[8607]= 1882296293;
assign addr[8608]= 2010011024;
assign addr[8609]= 2096992772;
assign addr[8610]= 2141478848;
assign addr[8611]= 2142567738;
assign addr[8612]= 2100237377;
assign addr[8613]= 2015345591;
assign addr[8614]= 1889612716;
assign addr[8615]= 1725586737;
assign addr[8616]= 1526591649;
assign addr[8617]= 1296660098;
assign addr[8618]= 1040451659;
assign addr[8619]= 763158411;
assign addr[8620]= 470399716;
assign addr[8621]= 168108346;
assign addr[8622]= -137589750;
assign addr[8623]= -440499581;
assign addr[8624]= -734482665;
assign addr[8625]= -1013581418;
assign addr[8626]= -1272139887;
assign addr[8627]= -1504918373;
assign addr[8628]= -1707199606;
assign addr[8629]= -1874884346;
assign addr[8630]= -2004574453;
assign addr[8631]= -2093641749;
assign addr[8632]= -2140281282;
assign addr[8633]= -2143547897;
assign addr[8634]= -2103375398;
assign addr[8635]= -2020577882;
assign addr[8636]= -1896833245;
assign addr[8637]= -1734649179;
assign addr[8638]= -1537312353;
assign addr[8639]= -1308821808;
assign addr[8640]= -1053807919;
assign addr[8641]= -777438554;
assign addr[8642]= -485314355;
assign addr[8643]= -183355234;
assign addr[8644]= 122319591;
assign addr[8645]= 425515602;
assign addr[8646]= 720088517;
assign addr[8647]= 1000068799;
assign addr[8648]= 1259782632;
assign addr[8649]= 1493966902;
assign addr[8650]= 1697875851;
assign addr[8651]= 1867377253;
assign addr[8652]= 1999036154;
assign addr[8653]= 2090184478;
assign addr[8654]= 2138975100;
assign addr[8655]= 2144419275;
assign addr[8656]= 2106406677;
assign addr[8657]= 2025707632;
assign addr[8658]= 1903957513;
assign addr[8659]= 1743623590;
assign addr[8660]= 1547955041;
assign addr[8661]= 1320917099;
assign addr[8662]= 1067110699;
assign addr[8663]= 791679244;
assign addr[8664]= 500204365;
assign addr[8665]= 198592817;
assign addr[8666]= -107043224;
assign addr[8667]= -410510029;
assign addr[8668]= -705657826;
assign addr[8669]= -986505429;
assign addr[8670]= -1247361445;
assign addr[8671]= -1482939614;
assign addr[8672]= -1688465931;
assign addr[8673]= -1859775393;
assign addr[8674]= -1993396407;
assign addr[8675]= -2086621133;
assign addr[8676]= -2137560369;
assign addr[8677]= -2145181827;
assign addr[8678]= -2109331059;
assign addr[8679]= -2030734582;
assign addr[8680]= -1910985158;
assign addr[8681]= -1752509516;
assign addr[8682]= -1558519173;
assign addr[8683]= -1332945355;
assign addr[8684]= -1080359326;
assign addr[8685]= -805879757;
assign addr[8686]= -515068990;
assign addr[8687]= -213820322;
assign addr[8688]= 91761426;
assign addr[8689]= 395483624;
assign addr[8690]= 691191324;
assign addr[8691]= 972891995;
assign addr[8692]= 1234876957;
assign addr[8693]= 1471837070;
assign addr[8694]= 1678970324;
assign addr[8695]= 1852079154;
assign addr[8696]= 1987655498;
assign addr[8697]= 2082951896;
assign addr[8698]= 2136037160;
assign addr[8699]= 2145835515;
assign addr[8700]= 2112148396;
assign addr[8701]= 2035658475;
assign addr[8702]= 1917915825;
assign addr[8703]= 1761306505;
assign addr[8704]= 1569004214;
assign addr[8705]= 1344905966;
assign addr[8706]= 1093553126;
assign addr[8707]= 820039373;
assign addr[8708]= 529907477;
assign addr[8709]= 229036977;
assign addr[8710]= -76474970;
assign addr[8711]= -380437148;
assign addr[8712]= -676689746;
assign addr[8713]= -959229189;
assign addr[8714]= -1222329801;
assign addr[8715]= -1460659832;
assign addr[8716]= -1669389513;
assign addr[8717]= -1844288924;
assign addr[8718]= -1981813720;
assign addr[8719]= -2079176953;
assign addr[8720]= -2134405552;
assign addr[8721]= -2146380306;
assign addr[8722]= -2114858546;
assign addr[8723]= -2040479063;
assign addr[8724]= -1924749160;
assign addr[8725]= -1770014111;
assign addr[8726]= -1579409630;
assign addr[8727]= -1356798326;
assign addr[8728]= -1106691431;
assign addr[8729]= -834157373;
assign addr[8730]= -544719071;
assign addr[8731]= -244242007;
assign addr[8732]= 61184634;
assign addr[8733]= 365371365;
assign addr[8734]= 662153826;
assign addr[8735]= 945517704;
assign addr[8736]= 1209720613;
assign addr[8737]= 1449408469;
assign addr[8738]= 1659723983;
assign addr[8739]= 1836405100;
assign addr[8740]= 1975871368;
assign addr[8741]= 2075296495;
assign addr[8742]= 2132665626;
assign addr[8743]= 2146816171;
assign addr[8744]= 2117461370;
assign addr[8745]= 2045196100;
assign addr[8746]= 1931484818;
assign addr[8747]= 1778631892;
assign addr[8748]= 1589734894;
assign addr[8749]= 1368621831;
assign addr[8750]= 1119773573;
assign addr[8751]= 848233042;
assign addr[8752]= 559503022;
assign addr[8753]= 259434643;
assign addr[8754]= -45891193;
assign addr[8755]= -350287041;
assign addr[8756]= -647584304;
assign addr[8757]= -931758235;
assign addr[8758]= -1197050035;
assign addr[8759]= -1438083551;
assign addr[8760]= -1649974225;
assign addr[8761]= -1828428082;
assign addr[8762]= -1969828744;
assign addr[8763]= -2071310720;
assign addr[8764]= -2130817471;
assign addr[8765]= -2147143090;
assign addr[8766]= -2119956737;
assign addr[8767]= -2049809346;
assign addr[8768]= -1938122457;
assign addr[8769]= -1787159411;
assign addr[8770]= -1599979481;
assign addr[8771]= -1380375881;
assign addr[8772]= -1132798888;
assign addr[8773]= -862265664;
assign addr[8774]= -574258580;
assign addr[8775]= -274614114;
assign addr[8776]= 30595422;
assign addr[8777]= 335184940;
assign addr[8778]= 632981917;
assign addr[8779]= 917951481;
assign addr[8780]= 1184318708;
assign addr[8781]= 1426685652;
assign addr[8782]= 1640140734;
assign addr[8783]= 1820358275;
assign addr[8784]= 1963686155;
assign addr[8785]= 2067219829;
assign addr[8786]= 2128861181;
assign addr[8787]= 2147361045;
assign addr[8788]= 2122344521;
assign addr[8789]= 2054318569;
assign addr[8790]= 1944661739;
assign addr[8791]= 1795596234;
assign addr[8792]= 1610142873;
assign addr[8793]= 1392059879;
assign addr[8794]= 1145766716;
assign addr[8795]= 876254528;
assign addr[8796]= 588984994;
assign addr[8797]= 289779648;
assign addr[8798]= -15298099;
assign addr[8799]= -320065829;
assign addr[8800]= -618347408;
assign addr[8801]= -904098143;
assign addr[8802]= -1171527280;
assign addr[8803]= -1415215352;
assign addr[8804]= -1630224009;
assign addr[8805]= -1812196087;
assign addr[8806]= -1957443913;
assign addr[8807]= -2063024031;
assign addr[8808]= -2126796855;
assign addr[8809]= -2147470025;
assign addr[8810]= -2124624598;
assign addr[8811]= -2058723538;
assign addr[8812]= -1951102334;
assign addr[8813]= -1803941934;
assign addr[8814]= -1620224553;
assign addr[8815]= -1403673233;
assign addr[8816]= -1158676398;
assign addr[8817]= -890198924;
assign addr[8818]= -603681519;
assign addr[8819]= -304930476;
assign addr[8820]= 0;
assign addr[8821]= 304930476;
assign addr[8822]= 603681519;
assign addr[8823]= 890198924;
assign addr[8824]= 1158676398;
assign addr[8825]= 1403673233;
assign addr[8826]= 1620224553;
assign addr[8827]= 1803941934;
assign addr[8828]= 1951102334;
assign addr[8829]= 2058723538;
assign addr[8830]= 2124624598;
assign addr[8831]= 2147470025;
assign addr[8832]= 2126796855;
assign addr[8833]= 2063024031;
assign addr[8834]= 1957443913;
assign addr[8835]= 1812196087;
assign addr[8836]= 1630224009;
assign addr[8837]= 1415215352;
assign addr[8838]= 1171527280;
assign addr[8839]= 904098143;
assign addr[8840]= 618347408;
assign addr[8841]= 320065829;
assign addr[8842]= 15298099;
assign addr[8843]= -289779648;
assign addr[8844]= -588984994;
assign addr[8845]= -876254528;
assign addr[8846]= -1145766716;
assign addr[8847]= -1392059879;
assign addr[8848]= -1610142873;
assign addr[8849]= -1795596234;
assign addr[8850]= -1944661739;
assign addr[8851]= -2054318569;
assign addr[8852]= -2122344521;
assign addr[8853]= -2147361045;
assign addr[8854]= -2128861181;
assign addr[8855]= -2067219829;
assign addr[8856]= -1963686155;
assign addr[8857]= -1820358275;
assign addr[8858]= -1640140734;
assign addr[8859]= -1426685652;
assign addr[8860]= -1184318708;
assign addr[8861]= -917951481;
assign addr[8862]= -632981917;
assign addr[8863]= -335184940;
assign addr[8864]= -30595422;
assign addr[8865]= 274614114;
assign addr[8866]= 574258580;
assign addr[8867]= 862265664;
assign addr[8868]= 1132798888;
assign addr[8869]= 1380375881;
assign addr[8870]= 1599979481;
assign addr[8871]= 1787159411;
assign addr[8872]= 1938122457;
assign addr[8873]= 2049809346;
assign addr[8874]= 2119956737;
assign addr[8875]= 2147143090;
assign addr[8876]= 2130817471;
assign addr[8877]= 2071310720;
assign addr[8878]= 1969828744;
assign addr[8879]= 1828428082;
assign addr[8880]= 1649974225;
assign addr[8881]= 1438083551;
assign addr[8882]= 1197050035;
assign addr[8883]= 931758235;
assign addr[8884]= 647584304;
assign addr[8885]= 350287041;
assign addr[8886]= 45891193;
assign addr[8887]= -259434643;
assign addr[8888]= -559503022;
assign addr[8889]= -848233042;
assign addr[8890]= -1119773573;
assign addr[8891]= -1368621831;
assign addr[8892]= -1589734894;
assign addr[8893]= -1778631892;
assign addr[8894]= -1931484818;
assign addr[8895]= -2045196100;
assign addr[8896]= -2117461370;
assign addr[8897]= -2146816171;
assign addr[8898]= -2132665626;
assign addr[8899]= -2075296495;
assign addr[8900]= -1975871368;
assign addr[8901]= -1836405100;
assign addr[8902]= -1659723983;
assign addr[8903]= -1449408469;
assign addr[8904]= -1209720613;
assign addr[8905]= -945517704;
assign addr[8906]= -662153826;
assign addr[8907]= -365371365;
assign addr[8908]= -61184634;
assign addr[8909]= 244242007;
assign addr[8910]= 544719071;
assign addr[8911]= 834157373;
assign addr[8912]= 1106691431;
assign addr[8913]= 1356798326;
assign addr[8914]= 1579409630;
assign addr[8915]= 1770014111;
assign addr[8916]= 1924749160;
assign addr[8917]= 2040479063;
assign addr[8918]= 2114858546;
assign addr[8919]= 2146380306;
assign addr[8920]= 2134405552;
assign addr[8921]= 2079176953;
assign addr[8922]= 1981813720;
assign addr[8923]= 1844288924;
assign addr[8924]= 1669389513;
assign addr[8925]= 1460659832;
assign addr[8926]= 1222329801;
assign addr[8927]= 959229189;
assign addr[8928]= 676689746;
assign addr[8929]= 380437148;
assign addr[8930]= 76474970;
assign addr[8931]= -229036977;
assign addr[8932]= -529907477;
assign addr[8933]= -820039373;
assign addr[8934]= -1093553126;
assign addr[8935]= -1344905966;
assign addr[8936]= -1569004214;
assign addr[8937]= -1761306505;
assign addr[8938]= -1917915825;
assign addr[8939]= -2035658475;
assign addr[8940]= -2112148396;
assign addr[8941]= -2145835515;
assign addr[8942]= -2136037160;
assign addr[8943]= -2082951896;
assign addr[8944]= -1987655498;
assign addr[8945]= -1852079154;
assign addr[8946]= -1678970324;
assign addr[8947]= -1471837070;
assign addr[8948]= -1234876957;
assign addr[8949]= -972891995;
assign addr[8950]= -691191324;
assign addr[8951]= -395483624;
assign addr[8952]= -91761426;
assign addr[8953]= 213820322;
assign addr[8954]= 515068990;
assign addr[8955]= 805879757;
assign addr[8956]= 1080359326;
assign addr[8957]= 1332945355;
assign addr[8958]= 1558519173;
assign addr[8959]= 1752509516;
assign addr[8960]= 1910985158;
assign addr[8961]= 2030734582;
assign addr[8962]= 2109331059;
assign addr[8963]= 2145181827;
assign addr[8964]= 2137560369;
assign addr[8965]= 2086621133;
assign addr[8966]= 1993396407;
assign addr[8967]= 1859775393;
assign addr[8968]= 1688465931;
assign addr[8969]= 1482939614;
assign addr[8970]= 1247361445;
assign addr[8971]= 986505429;
assign addr[8972]= 705657826;
assign addr[8973]= 410510029;
assign addr[8974]= 107043224;
assign addr[8975]= -198592817;
assign addr[8976]= -500204365;
assign addr[8977]= -791679244;
assign addr[8978]= -1067110699;
assign addr[8979]= -1320917099;
assign addr[8980]= -1547955041;
assign addr[8981]= -1743623590;
assign addr[8982]= -1903957513;
assign addr[8983]= -2025707632;
assign addr[8984]= -2106406677;
assign addr[8985]= -2144419275;
assign addr[8986]= -2138975100;
assign addr[8987]= -2090184478;
assign addr[8988]= -1999036154;
assign addr[8989]= -1867377253;
assign addr[8990]= -1697875851;
assign addr[8991]= -1493966902;
assign addr[8992]= -1259782632;
assign addr[8993]= -1000068799;
assign addr[8994]= -720088517;
assign addr[8995]= -425515602;
assign addr[8996]= -122319591;
assign addr[8997]= 183355234;
assign addr[8998]= 485314355;
assign addr[8999]= 777438554;
assign addr[9000]= 1053807919;
assign addr[9001]= 1308821808;
assign addr[9002]= 1537312353;
assign addr[9003]= 1734649179;
assign addr[9004]= 1896833245;
assign addr[9005]= 2020577882;
assign addr[9006]= 2103375398;
assign addr[9007]= 2143547897;
assign addr[9008]= 2140281282;
assign addr[9009]= 2093641749;
assign addr[9010]= 2004574453;
assign addr[9011]= 1874884346;
assign addr[9012]= 1707199606;
assign addr[9013]= 1504918373;
assign addr[9014]= 1272139887;
assign addr[9015]= 1013581418;
assign addr[9016]= 734482665;
assign addr[9017]= 440499581;
assign addr[9018]= 137589750;
assign addr[9019]= -168108346;
assign addr[9020]= -470399716;
assign addr[9021]= -763158411;
assign addr[9022]= -1040451659;
assign addr[9023]= -1296660098;
assign addr[9024]= -1526591649;
assign addr[9025]= -1725586737;
assign addr[9026]= -1889612716;
assign addr[9027]= -2015345591;
assign addr[9028]= -2100237377;
assign addr[9029]= -2142567738;
assign addr[9030]= -2141478848;
assign addr[9031]= -2096992772;
assign addr[9032]= -2010011024;
assign addr[9033]= -1882296293;
assign addr[9034]= -1716436725;
assign addr[9035]= -1515793473;
assign addr[9036]= -1284432584;
assign addr[9037]= -1027042599;
assign addr[9038]= -748839539;
assign addr[9039]= -455461206;
assign addr[9040]= -152852926;
assign addr[9041]= 152852926;
assign addr[9042]= 455461206;
assign addr[9043]= 748839539;
assign addr[9044]= 1027042599;
assign addr[9045]= 1284432584;
assign addr[9046]= 1515793473;
assign addr[9047]= 1716436725;
assign addr[9048]= 1882296293;
assign addr[9049]= 2010011024;
assign addr[9050]= 2096992772;
assign addr[9051]= 2141478848;
assign addr[9052]= 2142567738;
assign addr[9053]= 2100237377;
assign addr[9054]= 2015345591;
assign addr[9055]= 1889612716;
assign addr[9056]= 1725586737;
assign addr[9057]= 1526591649;
assign addr[9058]= 1296660098;
assign addr[9059]= 1040451659;
assign addr[9060]= 763158411;
assign addr[9061]= 470399716;
assign addr[9062]= 168108346;
assign addr[9063]= -137589750;
assign addr[9064]= -440499581;
assign addr[9065]= -734482665;
assign addr[9066]= -1013581418;
assign addr[9067]= -1272139887;
assign addr[9068]= -1504918373;
assign addr[9069]= -1707199606;
assign addr[9070]= -1874884346;
assign addr[9071]= -2004574453;
assign addr[9072]= -2093641749;
assign addr[9073]= -2140281282;
assign addr[9074]= -2143547897;
assign addr[9075]= -2103375398;
assign addr[9076]= -2020577882;
assign addr[9077]= -1896833245;
assign addr[9078]= -1734649179;
assign addr[9079]= -1537312353;
assign addr[9080]= -1308821808;
assign addr[9081]= -1053807919;
assign addr[9082]= -777438554;
assign addr[9083]= -485314355;
assign addr[9084]= -183355234;
assign addr[9085]= 122319591;
assign addr[9086]= 425515602;
assign addr[9087]= 720088517;
assign addr[9088]= 1000068799;
assign addr[9089]= 1259782632;
assign addr[9090]= 1493966902;
assign addr[9091]= 1697875851;
assign addr[9092]= 1867377253;
assign addr[9093]= 1999036154;
assign addr[9094]= 2090184478;
assign addr[9095]= 2138975100;
assign addr[9096]= 2144419275;
assign addr[9097]= 2106406677;
assign addr[9098]= 2025707632;
assign addr[9099]= 1903957513;
assign addr[9100]= 1743623590;
assign addr[9101]= 1547955041;
assign addr[9102]= 1320917099;
assign addr[9103]= 1067110699;
assign addr[9104]= 791679244;
assign addr[9105]= 500204365;
assign addr[9106]= 198592817;
assign addr[9107]= -107043224;
assign addr[9108]= -410510029;
assign addr[9109]= -705657826;
assign addr[9110]= -986505429;
assign addr[9111]= -1247361445;
assign addr[9112]= -1482939614;
assign addr[9113]= -1688465931;
assign addr[9114]= -1859775393;
assign addr[9115]= -1993396407;
assign addr[9116]= -2086621133;
assign addr[9117]= -2137560369;
assign addr[9118]= -2145181827;
assign addr[9119]= -2109331059;
assign addr[9120]= -2030734582;
assign addr[9121]= -1910985158;
assign addr[9122]= -1752509516;
assign addr[9123]= -1558519173;
assign addr[9124]= -1332945355;
assign addr[9125]= -1080359326;
assign addr[9126]= -805879757;
assign addr[9127]= -515068990;
assign addr[9128]= -213820322;
assign addr[9129]= 91761426;
assign addr[9130]= 395483624;
assign addr[9131]= 691191324;
assign addr[9132]= 972891995;
assign addr[9133]= 1234876957;
assign addr[9134]= 1471837070;
assign addr[9135]= 1678970324;
assign addr[9136]= 1852079154;
assign addr[9137]= 1987655498;
assign addr[9138]= 2082951896;
assign addr[9139]= 2136037160;
assign addr[9140]= 2145835515;
assign addr[9141]= 2112148396;
assign addr[9142]= 2035658475;
assign addr[9143]= 1917915825;
assign addr[9144]= 1761306505;
assign addr[9145]= 1569004214;
assign addr[9146]= 1344905966;
assign addr[9147]= 1093553126;
assign addr[9148]= 820039373;
assign addr[9149]= 529907477;
assign addr[9150]= 229036977;
assign addr[9151]= -76474970;
assign addr[9152]= -380437148;
assign addr[9153]= -676689746;
assign addr[9154]= -959229189;
assign addr[9155]= -1222329801;
assign addr[9156]= -1460659832;
assign addr[9157]= -1669389513;
assign addr[9158]= -1844288924;
assign addr[9159]= -1981813720;
assign addr[9160]= -2079176953;
assign addr[9161]= -2134405552;
assign addr[9162]= -2146380306;
assign addr[9163]= -2114858546;
assign addr[9164]= -2040479063;
assign addr[9165]= -1924749160;
assign addr[9166]= -1770014111;
assign addr[9167]= -1579409630;
assign addr[9168]= -1356798326;
assign addr[9169]= -1106691431;
assign addr[9170]= -834157373;
assign addr[9171]= -544719071;
assign addr[9172]= -244242007;
assign addr[9173]= 61184634;
assign addr[9174]= 365371365;
assign addr[9175]= 662153826;
assign addr[9176]= 945517704;
assign addr[9177]= 1209720613;
assign addr[9178]= 1449408469;
assign addr[9179]= 1659723983;
assign addr[9180]= 1836405100;
assign addr[9181]= 1975871368;
assign addr[9182]= 2075296495;
assign addr[9183]= 2132665626;
assign addr[9184]= 2146816171;
assign addr[9185]= 2117461370;
assign addr[9186]= 2045196100;
assign addr[9187]= 1931484818;
assign addr[9188]= 1778631892;
assign addr[9189]= 1589734894;
assign addr[9190]= 1368621831;
assign addr[9191]= 1119773573;
assign addr[9192]= 848233042;
assign addr[9193]= 559503022;
assign addr[9194]= 259434643;
assign addr[9195]= -45891193;
assign addr[9196]= -350287041;
assign addr[9197]= -647584304;
assign addr[9198]= -931758235;
assign addr[9199]= -1197050035;
assign addr[9200]= -1438083551;
assign addr[9201]= -1649974225;
assign addr[9202]= -1828428082;
assign addr[9203]= -1969828744;
assign addr[9204]= -2071310720;
assign addr[9205]= -2130817471;
assign addr[9206]= -2147143090;
assign addr[9207]= -2119956737;
assign addr[9208]= -2049809346;
assign addr[9209]= -1938122457;
assign addr[9210]= -1787159411;
assign addr[9211]= -1599979481;
assign addr[9212]= -1380375881;
assign addr[9213]= -1132798888;
assign addr[9214]= -862265664;
assign addr[9215]= -574258580;
assign addr[9216]= -274614114;
assign addr[9217]= 30595422;
assign addr[9218]= 335184940;
assign addr[9219]= 632981917;
assign addr[9220]= 917951481;
assign addr[9221]= 1184318708;
assign addr[9222]= 1426685652;
assign addr[9223]= 1640140734;
assign addr[9224]= 1820358275;
assign addr[9225]= 1963686155;
assign addr[9226]= 2067219829;
assign addr[9227]= 2128861181;
assign addr[9228]= 2147361045;
assign addr[9229]= 2122344521;
assign addr[9230]= 2054318569;
assign addr[9231]= 1944661739;
assign addr[9232]= 1795596234;
assign addr[9233]= 1610142873;
assign addr[9234]= 1392059879;
assign addr[9235]= 1145766716;
assign addr[9236]= 876254528;
assign addr[9237]= 588984994;
assign addr[9238]= 289779648;
assign addr[9239]= -15298099;
assign addr[9240]= -320065829;
assign addr[9241]= -618347408;
assign addr[9242]= -904098143;
assign addr[9243]= -1171527280;
assign addr[9244]= -1415215352;
assign addr[9245]= -1630224009;
assign addr[9246]= -1812196087;
assign addr[9247]= -1957443913;
assign addr[9248]= -2063024031;
assign addr[9249]= -2126796855;
assign addr[9250]= -2147470025;
assign addr[9251]= -2124624598;
assign addr[9252]= -2058723538;
assign addr[9253]= -1951102334;
assign addr[9254]= -1803941934;
assign addr[9255]= -1620224553;
assign addr[9256]= -1403673233;
assign addr[9257]= -1158676398;
assign addr[9258]= -890198924;
assign addr[9259]= -603681519;
assign addr[9260]= -304930476;
assign addr[9261]= 0;
assign addr[9262]= 304930476;
assign addr[9263]= 603681519;
assign addr[9264]= 890198924;
assign addr[9265]= 1158676398;
assign addr[9266]= 1403673233;
assign addr[9267]= 1620224553;
assign addr[9268]= 1803941934;
assign addr[9269]= 1951102334;
assign addr[9270]= 2058723538;
assign addr[9271]= 2124624598;
assign addr[9272]= 2147470025;
assign addr[9273]= 2126796855;
assign addr[9274]= 2063024031;
assign addr[9275]= 1957443913;
assign addr[9276]= 1812196087;
assign addr[9277]= 1630224009;
assign addr[9278]= 1415215352;
assign addr[9279]= 1171527280;
assign addr[9280]= 904098143;
assign addr[9281]= 618347408;
assign addr[9282]= 320065829;
assign addr[9283]= 15298099;
assign addr[9284]= -289779648;
assign addr[9285]= -588984994;
assign addr[9286]= -876254528;
assign addr[9287]= -1145766716;
assign addr[9288]= -1392059879;
assign addr[9289]= -1610142873;
assign addr[9290]= -1795596234;
assign addr[9291]= -1944661739;
assign addr[9292]= -2054318569;
assign addr[9293]= -2122344521;
assign addr[9294]= -2147361045;
assign addr[9295]= -2128861181;
assign addr[9296]= -2067219829;
assign addr[9297]= -1963686155;
assign addr[9298]= -1820358275;
assign addr[9299]= -1640140734;
assign addr[9300]= -1426685652;
assign addr[9301]= -1184318708;
assign addr[9302]= -917951481;
assign addr[9303]= -632981917;
assign addr[9304]= -335184940;
assign addr[9305]= -30595422;
assign addr[9306]= 274614114;
assign addr[9307]= 574258580;
assign addr[9308]= 862265664;
assign addr[9309]= 1132798888;
assign addr[9310]= 1380375881;
assign addr[9311]= 1599979481;
assign addr[9312]= 1787159411;
assign addr[9313]= 1938122457;
assign addr[9314]= 2049809346;
assign addr[9315]= 2119956737;
assign addr[9316]= 2147143090;
assign addr[9317]= 2130817471;
assign addr[9318]= 2071310720;
assign addr[9319]= 1969828744;
assign addr[9320]= 1828428082;
assign addr[9321]= 1649974225;
assign addr[9322]= 1438083551;
assign addr[9323]= 1197050035;
assign addr[9324]= 931758235;
assign addr[9325]= 647584304;
assign addr[9326]= 350287041;
assign addr[9327]= 45891193;
assign addr[9328]= -259434643;
assign addr[9329]= -559503022;
assign addr[9330]= -848233042;
assign addr[9331]= -1119773573;
assign addr[9332]= -1368621831;
assign addr[9333]= -1589734894;
assign addr[9334]= -1778631892;
assign addr[9335]= -1931484818;
assign addr[9336]= -2045196100;
assign addr[9337]= -2117461370;
assign addr[9338]= -2146816171;
assign addr[9339]= -2132665626;
assign addr[9340]= -2075296495;
assign addr[9341]= -1975871368;
assign addr[9342]= -1836405100;
assign addr[9343]= -1659723983;
assign addr[9344]= -1449408469;
assign addr[9345]= -1209720613;
assign addr[9346]= -945517704;
assign addr[9347]= -662153826;
assign addr[9348]= -365371365;
assign addr[9349]= -61184634;
assign addr[9350]= 244242007;
assign addr[9351]= 544719071;
assign addr[9352]= 834157373;
assign addr[9353]= 1106691431;
assign addr[9354]= 1356798326;
assign addr[9355]= 1579409630;
assign addr[9356]= 1770014111;
assign addr[9357]= 1924749160;
assign addr[9358]= 2040479063;
assign addr[9359]= 2114858546;
assign addr[9360]= 2146380306;
assign addr[9361]= 2134405552;
assign addr[9362]= 2079176953;
assign addr[9363]= 1981813720;
assign addr[9364]= 1844288924;
assign addr[9365]= 1669389513;
assign addr[9366]= 1460659832;
assign addr[9367]= 1222329801;
assign addr[9368]= 959229189;
assign addr[9369]= 676689746;
assign addr[9370]= 380437148;
assign addr[9371]= 76474970;
assign addr[9372]= -229036977;
assign addr[9373]= -529907477;
assign addr[9374]= -820039373;
assign addr[9375]= -1093553126;
assign addr[9376]= -1344905966;
assign addr[9377]= -1569004214;
assign addr[9378]= -1761306505;
assign addr[9379]= -1917915825;
assign addr[9380]= -2035658475;
assign addr[9381]= -2112148396;
assign addr[9382]= -2145835515;
assign addr[9383]= -2136037160;
assign addr[9384]= -2082951896;
assign addr[9385]= -1987655498;
assign addr[9386]= -1852079154;
assign addr[9387]= -1678970324;
assign addr[9388]= -1471837070;
assign addr[9389]= -1234876957;
assign addr[9390]= -972891995;
assign addr[9391]= -691191324;
assign addr[9392]= -395483624;
assign addr[9393]= -91761426;
assign addr[9394]= 213820322;
assign addr[9395]= 515068990;
assign addr[9396]= 805879757;
assign addr[9397]= 1080359326;
assign addr[9398]= 1332945355;
assign addr[9399]= 1558519173;
assign addr[9400]= 1752509516;
assign addr[9401]= 1910985158;
assign addr[9402]= 2030734582;
assign addr[9403]= 2109331059;
assign addr[9404]= 2145181827;
assign addr[9405]= 2137560369;
assign addr[9406]= 2086621133;
assign addr[9407]= 1993396407;
assign addr[9408]= 1859775393;
assign addr[9409]= 1688465931;
assign addr[9410]= 1482939614;
assign addr[9411]= 1247361445;
assign addr[9412]= 986505429;
assign addr[9413]= 705657826;
assign addr[9414]= 410510029;
assign addr[9415]= 107043224;
assign addr[9416]= -198592817;
assign addr[9417]= -500204365;
assign addr[9418]= -791679244;
assign addr[9419]= -1067110699;
assign addr[9420]= -1320917099;
assign addr[9421]= -1547955041;
assign addr[9422]= -1743623590;
assign addr[9423]= -1903957513;
assign addr[9424]= -2025707632;
assign addr[9425]= -2106406677;
assign addr[9426]= -2144419275;
assign addr[9427]= -2138975100;
assign addr[9428]= -2090184478;
assign addr[9429]= -1999036154;
assign addr[9430]= -1867377253;
assign addr[9431]= -1697875851;
assign addr[9432]= -1493966902;
assign addr[9433]= -1259782632;
assign addr[9434]= -1000068799;
assign addr[9435]= -720088517;
assign addr[9436]= -425515602;
assign addr[9437]= -122319591;
assign addr[9438]= 183355234;
assign addr[9439]= 485314355;
assign addr[9440]= 777438554;
assign addr[9441]= 1053807919;
assign addr[9442]= 1308821808;
assign addr[9443]= 1537312353;
assign addr[9444]= 1734649179;
assign addr[9445]= 1896833245;
assign addr[9446]= 2020577882;
assign addr[9447]= 2103375398;
assign addr[9448]= 2143547897;
assign addr[9449]= 2140281282;
assign addr[9450]= 2093641749;
assign addr[9451]= 2004574453;
assign addr[9452]= 1874884346;
assign addr[9453]= 1707199606;
assign addr[9454]= 1504918373;
assign addr[9455]= 1272139887;
assign addr[9456]= 1013581418;
assign addr[9457]= 734482665;
assign addr[9458]= 440499581;
assign addr[9459]= 137589750;
assign addr[9460]= -168108346;
assign addr[9461]= -470399716;
assign addr[9462]= -763158411;
assign addr[9463]= -1040451659;
assign addr[9464]= -1296660098;
assign addr[9465]= -1526591649;
assign addr[9466]= -1725586737;
assign addr[9467]= -1889612716;
assign addr[9468]= -2015345591;
assign addr[9469]= -2100237377;
assign addr[9470]= -2142567738;
assign addr[9471]= -2141478848;
assign addr[9472]= -2096992772;
assign addr[9473]= -2010011024;
assign addr[9474]= -1882296293;
assign addr[9475]= -1716436725;
assign addr[9476]= -1515793473;
assign addr[9477]= -1284432584;
assign addr[9478]= -1027042599;
assign addr[9479]= -748839539;
assign addr[9480]= -455461206;
assign addr[9481]= -152852926;
assign addr[9482]= 152852926;
assign addr[9483]= 455461206;
assign addr[9484]= 748839539;
assign addr[9485]= 1027042599;
assign addr[9486]= 1284432584;
assign addr[9487]= 1515793473;
assign addr[9488]= 1716436725;
assign addr[9489]= 1882296293;
assign addr[9490]= 2010011024;
assign addr[9491]= 2096992772;
assign addr[9492]= 2141478848;
assign addr[9493]= 2142567738;
assign addr[9494]= 2100237377;
assign addr[9495]= 2015345591;
assign addr[9496]= 1889612716;
assign addr[9497]= 1725586737;
assign addr[9498]= 1526591649;
assign addr[9499]= 1296660098;
assign addr[9500]= 1040451659;
assign addr[9501]= 763158411;
assign addr[9502]= 470399716;
assign addr[9503]= 168108346;
assign addr[9504]= -137589750;
assign addr[9505]= -440499581;
assign addr[9506]= -734482665;
assign addr[9507]= -1013581418;
assign addr[9508]= -1272139887;
assign addr[9509]= -1504918373;
assign addr[9510]= -1707199606;
assign addr[9511]= -1874884346;
assign addr[9512]= -2004574453;
assign addr[9513]= -2093641749;
assign addr[9514]= -2140281282;
assign addr[9515]= -2143547897;
assign addr[9516]= -2103375398;
assign addr[9517]= -2020577882;
assign addr[9518]= -1896833245;
assign addr[9519]= -1734649179;
assign addr[9520]= -1537312353;
assign addr[9521]= -1308821808;
assign addr[9522]= -1053807919;
assign addr[9523]= -777438554;
assign addr[9524]= -485314355;
assign addr[9525]= -183355234;
assign addr[9526]= 122319591;
assign addr[9527]= 425515602;
assign addr[9528]= 720088517;
assign addr[9529]= 1000068799;
assign addr[9530]= 1259782632;
assign addr[9531]= 1493966902;
assign addr[9532]= 1697875851;
assign addr[9533]= 1867377253;
assign addr[9534]= 1999036154;
assign addr[9535]= 2090184478;
assign addr[9536]= 2138975100;
assign addr[9537]= 2144419275;
assign addr[9538]= 2106406677;
assign addr[9539]= 2025707632;
assign addr[9540]= 1903957513;
assign addr[9541]= 1743623590;
assign addr[9542]= 1547955041;
assign addr[9543]= 1320917099;
assign addr[9544]= 1067110699;
assign addr[9545]= 791679244;
assign addr[9546]= 500204365;
assign addr[9547]= 198592817;
assign addr[9548]= -107043224;
assign addr[9549]= -410510029;
assign addr[9550]= -705657826;
assign addr[9551]= -986505429;
assign addr[9552]= -1247361445;
assign addr[9553]= -1482939614;
assign addr[9554]= -1688465931;
assign addr[9555]= -1859775393;
assign addr[9556]= -1993396407;
assign addr[9557]= -2086621133;
assign addr[9558]= -2137560369;
assign addr[9559]= -2145181827;
assign addr[9560]= -2109331059;
assign addr[9561]= -2030734582;
assign addr[9562]= -1910985158;
assign addr[9563]= -1752509516;
assign addr[9564]= -1558519173;
assign addr[9565]= -1332945355;
assign addr[9566]= -1080359326;
assign addr[9567]= -805879757;
assign addr[9568]= -515068990;
assign addr[9569]= -213820322;
assign addr[9570]= 91761426;
assign addr[9571]= 395483624;
assign addr[9572]= 691191324;
assign addr[9573]= 972891995;
assign addr[9574]= 1234876957;
assign addr[9575]= 1471837070;
assign addr[9576]= 1678970324;
assign addr[9577]= 1852079154;
assign addr[9578]= 1987655498;
assign addr[9579]= 2082951896;
assign addr[9580]= 2136037160;
assign addr[9581]= 2145835515;
assign addr[9582]= 2112148396;
assign addr[9583]= 2035658475;
assign addr[9584]= 1917915825;
assign addr[9585]= 1761306505;
assign addr[9586]= 1569004214;
assign addr[9587]= 1344905966;
assign addr[9588]= 1093553126;
assign addr[9589]= 820039373;
assign addr[9590]= 529907477;
assign addr[9591]= 229036977;
assign addr[9592]= -76474970;
assign addr[9593]= -380437148;
assign addr[9594]= -676689746;
assign addr[9595]= -959229189;
assign addr[9596]= -1222329801;
assign addr[9597]= -1460659832;
assign addr[9598]= -1669389513;
assign addr[9599]= -1844288924;
assign addr[9600]= -1981813720;
assign addr[9601]= -2079176953;
assign addr[9602]= -2134405552;
assign addr[9603]= -2146380306;
assign addr[9604]= -2114858546;
assign addr[9605]= -2040479063;
assign addr[9606]= -1924749160;
assign addr[9607]= -1770014111;
assign addr[9608]= -1579409630;
assign addr[9609]= -1356798326;
assign addr[9610]= -1106691431;
assign addr[9611]= -834157373;
assign addr[9612]= -544719071;
assign addr[9613]= -244242007;
assign addr[9614]= 61184634;
assign addr[9615]= 365371365;
assign addr[9616]= 662153826;
assign addr[9617]= 945517704;
assign addr[9618]= 1209720613;
assign addr[9619]= 1449408469;
assign addr[9620]= 1659723983;
assign addr[9621]= 1836405100;
assign addr[9622]= 1975871368;
assign addr[9623]= 2075296495;
assign addr[9624]= 2132665626;
assign addr[9625]= 2146816171;
assign addr[9626]= 2117461370;
assign addr[9627]= 2045196100;
assign addr[9628]= 1931484818;
assign addr[9629]= 1778631892;
assign addr[9630]= 1589734894;
assign addr[9631]= 1368621831;
assign addr[9632]= 1119773573;
assign addr[9633]= 848233042;
assign addr[9634]= 559503022;
assign addr[9635]= 259434643;
assign addr[9636]= -45891193;
assign addr[9637]= -350287041;
assign addr[9638]= -647584304;
assign addr[9639]= -931758235;
assign addr[9640]= -1197050035;
assign addr[9641]= -1438083551;
assign addr[9642]= -1649974225;
assign addr[9643]= -1828428082;
assign addr[9644]= -1969828744;
assign addr[9645]= -2071310720;
assign addr[9646]= -2130817471;
assign addr[9647]= -2147143090;
assign addr[9648]= -2119956737;
assign addr[9649]= -2049809346;
assign addr[9650]= -1938122457;
assign addr[9651]= -1787159411;
assign addr[9652]= -1599979481;
assign addr[9653]= -1380375881;
assign addr[9654]= -1132798888;
assign addr[9655]= -862265664;
assign addr[9656]= -574258580;
assign addr[9657]= -274614114;
assign addr[9658]= 30595422;
assign addr[9659]= 335184940;
assign addr[9660]= 632981917;
assign addr[9661]= 917951481;
assign addr[9662]= 1184318708;
assign addr[9663]= 1426685652;
assign addr[9664]= 1640140734;
assign addr[9665]= 1820358275;
assign addr[9666]= 1963686155;
assign addr[9667]= 2067219829;
assign addr[9668]= 2128861181;
assign addr[9669]= 2147361045;
assign addr[9670]= 2122344521;
assign addr[9671]= 2054318569;
assign addr[9672]= 1944661739;
assign addr[9673]= 1795596234;
assign addr[9674]= 1610142873;
assign addr[9675]= 1392059879;
assign addr[9676]= 1145766716;
assign addr[9677]= 876254528;
assign addr[9678]= 588984994;
assign addr[9679]= 289779648;
assign addr[9680]= -15298099;
assign addr[9681]= -320065829;
assign addr[9682]= -618347408;
assign addr[9683]= -904098143;
assign addr[9684]= -1171527280;
assign addr[9685]= -1415215352;
assign addr[9686]= -1630224009;
assign addr[9687]= -1812196087;
assign addr[9688]= -1957443913;
assign addr[9689]= -2063024031;
assign addr[9690]= -2126796855;
assign addr[9691]= -2147470025;
assign addr[9692]= -2124624598;
assign addr[9693]= -2058723538;
assign addr[9694]= -1951102334;
assign addr[9695]= -1803941934;
assign addr[9696]= -1620224553;
assign addr[9697]= -1403673233;
assign addr[9698]= -1158676398;
assign addr[9699]= -890198924;
assign addr[9700]= -603681519;
assign addr[9701]= -304930476;
assign addr[9702]= 0;
assign addr[9703]= 304930476;
assign addr[9704]= 603681519;
assign addr[9705]= 890198924;
assign addr[9706]= 1158676398;
assign addr[9707]= 1403673233;
assign addr[9708]= 1620224553;
assign addr[9709]= 1803941934;
assign addr[9710]= 1951102334;
assign addr[9711]= 2058723538;
assign addr[9712]= 2124624598;
assign addr[9713]= 2147470025;
assign addr[9714]= 2126796855;
assign addr[9715]= 2063024031;
assign addr[9716]= 1957443913;
assign addr[9717]= 1812196087;
assign addr[9718]= 1630224009;
assign addr[9719]= 1415215352;
assign addr[9720]= 1171527280;
assign addr[9721]= 904098143;
assign addr[9722]= 618347408;
assign addr[9723]= 320065829;
assign addr[9724]= 15298099;
assign addr[9725]= -289779648;
assign addr[9726]= -588984994;
assign addr[9727]= -876254528;
assign addr[9728]= -1145766716;
assign addr[9729]= -1392059879;
assign addr[9730]= -1610142873;
assign addr[9731]= -1795596234;
assign addr[9732]= -1944661739;
assign addr[9733]= -2054318569;
assign addr[9734]= -2122344521;
assign addr[9735]= -2147361045;
assign addr[9736]= -2128861181;
assign addr[9737]= -2067219829;
assign addr[9738]= -1963686155;
assign addr[9739]= -1820358275;
assign addr[9740]= -1640140734;
assign addr[9741]= -1426685652;
assign addr[9742]= -1184318708;
assign addr[9743]= -917951481;
assign addr[9744]= -632981917;
assign addr[9745]= -335184940;
assign addr[9746]= -30595422;
assign addr[9747]= 274614114;
assign addr[9748]= 574258580;
assign addr[9749]= 862265664;
assign addr[9750]= 1132798888;
assign addr[9751]= 1380375881;
assign addr[9752]= 1599979481;
assign addr[9753]= 1787159411;
assign addr[9754]= 1938122457;
assign addr[9755]= 2049809346;
assign addr[9756]= 2119956737;
assign addr[9757]= 2147143090;
assign addr[9758]= 2130817471;
assign addr[9759]= 2071310720;
assign addr[9760]= 1969828744;
assign addr[9761]= 1828428082;
assign addr[9762]= 1649974225;
assign addr[9763]= 1438083551;
assign addr[9764]= 1197050035;
assign addr[9765]= 931758235;
assign addr[9766]= 647584304;
assign addr[9767]= 350287041;
assign addr[9768]= 45891193;
assign addr[9769]= -259434643;
assign addr[9770]= -559503022;
assign addr[9771]= -848233042;
assign addr[9772]= -1119773573;
assign addr[9773]= -1368621831;
assign addr[9774]= -1589734894;
assign addr[9775]= -1778631892;
assign addr[9776]= -1931484818;
assign addr[9777]= -2045196100;
assign addr[9778]= -2117461370;
assign addr[9779]= -2146816171;
assign addr[9780]= -2132665626;
assign addr[9781]= -2075296495;
assign addr[9782]= -1975871368;
assign addr[9783]= -1836405100;
assign addr[9784]= -1659723983;
assign addr[9785]= -1449408469;
assign addr[9786]= -1209720613;
assign addr[9787]= -945517704;
assign addr[9788]= -662153826;
assign addr[9789]= -365371365;
assign addr[9790]= -61184634;
assign addr[9791]= 244242007;
assign addr[9792]= 544719071;
assign addr[9793]= 834157373;
assign addr[9794]= 1106691431;
assign addr[9795]= 1356798326;
assign addr[9796]= 1579409630;
assign addr[9797]= 1770014111;
assign addr[9798]= 1924749160;
assign addr[9799]= 2040479063;
assign addr[9800]= 2114858546;
assign addr[9801]= 2146380306;
assign addr[9802]= 2134405552;
assign addr[9803]= 2079176953;
assign addr[9804]= 1981813720;
assign addr[9805]= 1844288924;
assign addr[9806]= 1669389513;
assign addr[9807]= 1460659832;
assign addr[9808]= 1222329801;
assign addr[9809]= 959229189;
assign addr[9810]= 676689746;
assign addr[9811]= 380437148;
assign addr[9812]= 76474970;
assign addr[9813]= -229036977;
assign addr[9814]= -529907477;
assign addr[9815]= -820039373;
assign addr[9816]= -1093553126;
assign addr[9817]= -1344905966;
assign addr[9818]= -1569004214;
assign addr[9819]= -1761306505;
assign addr[9820]= -1917915825;
assign addr[9821]= -2035658475;
assign addr[9822]= -2112148396;
assign addr[9823]= -2145835515;
assign addr[9824]= -2136037160;
assign addr[9825]= -2082951896;
assign addr[9826]= -1987655498;
assign addr[9827]= -1852079154;
assign addr[9828]= -1678970324;
assign addr[9829]= -1471837070;
assign addr[9830]= -1234876957;
assign addr[9831]= -972891995;
assign addr[9832]= -691191324;
assign addr[9833]= -395483624;
assign addr[9834]= -91761426;
assign addr[9835]= 213820322;
assign addr[9836]= 515068990;
assign addr[9837]= 805879757;
assign addr[9838]= 1080359326;
assign addr[9839]= 1332945355;
assign addr[9840]= 1558519173;
assign addr[9841]= 1752509516;
assign addr[9842]= 1910985158;
assign addr[9843]= 2030734582;
assign addr[9844]= 2109331059;
assign addr[9845]= 2145181827;
assign addr[9846]= 2137560369;
assign addr[9847]= 2086621133;
assign addr[9848]= 1993396407;
assign addr[9849]= 1859775393;
assign addr[9850]= 1688465931;
assign addr[9851]= 1482939614;
assign addr[9852]= 1247361445;
assign addr[9853]= 986505429;
assign addr[9854]= 705657826;
assign addr[9855]= 410510029;
assign addr[9856]= 107043224;
assign addr[9857]= -198592817;
assign addr[9858]= -500204365;
assign addr[9859]= -791679244;
assign addr[9860]= -1067110699;
assign addr[9861]= -1320917099;
assign addr[9862]= -1547955041;
assign addr[9863]= -1743623590;
assign addr[9864]= -1903957513;
assign addr[9865]= -2025707632;
assign addr[9866]= -2106406677;
assign addr[9867]= -2144419275;
assign addr[9868]= -2138975100;
assign addr[9869]= -2090184478;
assign addr[9870]= -1999036154;
assign addr[9871]= -1867377253;
assign addr[9872]= -1697875851;
assign addr[9873]= -1493966902;
assign addr[9874]= -1259782632;
assign addr[9875]= -1000068799;
assign addr[9876]= -720088517;
assign addr[9877]= -425515602;
assign addr[9878]= -122319591;
assign addr[9879]= 183355234;
assign addr[9880]= 485314355;
assign addr[9881]= 777438554;
assign addr[9882]= 1053807919;
assign addr[9883]= 1308821808;
assign addr[9884]= 1537312353;
assign addr[9885]= 1734649179;
assign addr[9886]= 1896833245;
assign addr[9887]= 2020577882;
assign addr[9888]= 2103375398;
assign addr[9889]= 2143547897;
assign addr[9890]= 2140281282;
assign addr[9891]= 2093641749;
assign addr[9892]= 2004574453;
assign addr[9893]= 1874884346;
assign addr[9894]= 1707199606;
assign addr[9895]= 1504918373;
assign addr[9896]= 1272139887;
assign addr[9897]= 1013581418;
assign addr[9898]= 734482665;
assign addr[9899]= 440499581;
assign addr[9900]= 137589750;
assign addr[9901]= -168108346;
assign addr[9902]= -470399716;
assign addr[9903]= -763158411;
assign addr[9904]= -1040451659;
assign addr[9905]= -1296660098;
assign addr[9906]= -1526591649;
assign addr[9907]= -1725586737;
assign addr[9908]= -1889612716;
assign addr[9909]= -2015345591;
assign addr[9910]= -2100237377;
assign addr[9911]= -2142567738;
assign addr[9912]= -2141478848;
assign addr[9913]= -2096992772;
assign addr[9914]= -2010011024;
assign addr[9915]= -1882296293;
assign addr[9916]= -1716436725;
assign addr[9917]= -1515793473;
assign addr[9918]= -1284432584;
assign addr[9919]= -1027042599;
assign addr[9920]= -748839539;
assign addr[9921]= -455461206;
assign addr[9922]= -152852926;
assign addr[9923]= 152852926;
assign addr[9924]= 455461206;
assign addr[9925]= 748839539;
assign addr[9926]= 1027042599;
assign addr[9927]= 1284432584;
assign addr[9928]= 1515793473;
assign addr[9929]= 1716436725;
assign addr[9930]= 1882296293;
assign addr[9931]= 2010011024;
assign addr[9932]= 2096992772;
assign addr[9933]= 2141478848;
assign addr[9934]= 2142567738;
assign addr[9935]= 2100237377;
assign addr[9936]= 2015345591;
assign addr[9937]= 1889612716;
assign addr[9938]= 1725586737;
assign addr[9939]= 1526591649;
assign addr[9940]= 1296660098;
assign addr[9941]= 1040451659;
assign addr[9942]= 763158411;
assign addr[9943]= 470399716;
assign addr[9944]= 168108346;
assign addr[9945]= -137589750;
assign addr[9946]= -440499581;
assign addr[9947]= -734482665;
assign addr[9948]= -1013581418;
assign addr[9949]= -1272139887;
assign addr[9950]= -1504918373;
assign addr[9951]= -1707199606;
assign addr[9952]= -1874884346;
assign addr[9953]= -2004574453;
assign addr[9954]= -2093641749;
assign addr[9955]= -2140281282;
assign addr[9956]= -2143547897;
assign addr[9957]= -2103375398;
assign addr[9958]= -2020577882;
assign addr[9959]= -1896833245;
assign addr[9960]= -1734649179;
assign addr[9961]= -1537312353;
assign addr[9962]= -1308821808;
assign addr[9963]= -1053807919;
assign addr[9964]= -777438554;
assign addr[9965]= -485314355;
assign addr[9966]= -183355234;
assign addr[9967]= 122319591;
assign addr[9968]= 425515602;
assign addr[9969]= 720088517;
assign addr[9970]= 1000068799;
assign addr[9971]= 1259782632;
assign addr[9972]= 1493966902;
assign addr[9973]= 1697875851;
assign addr[9974]= 1867377253;
assign addr[9975]= 1999036154;
assign addr[9976]= 2090184478;
assign addr[9977]= 2138975100;
assign addr[9978]= 2144419275;
assign addr[9979]= 2106406677;
assign addr[9980]= 2025707632;
assign addr[9981]= 1903957513;
assign addr[9982]= 1743623590;
assign addr[9983]= 1547955041;
assign addr[9984]= 1320917099;
assign addr[9985]= 1067110699;
assign addr[9986]= 791679244;
assign addr[9987]= 500204365;
assign addr[9988]= 198592817;
assign addr[9989]= -107043224;
assign addr[9990]= -410510029;
assign addr[9991]= -705657826;
assign addr[9992]= -986505429;
assign addr[9993]= -1247361445;
assign addr[9994]= -1482939614;
assign addr[9995]= -1688465931;
assign addr[9996]= -1859775393;
assign addr[9997]= -1993396407;
assign addr[9998]= -2086621133;
assign addr[9999]= -2137560369;
assign addr[10000]= -2145181827;
assign addr[10001]= -2109331059;
assign addr[10002]= -2030734582;
assign addr[10003]= -1910985158;
assign addr[10004]= -1752509516;
assign addr[10005]= -1558519173;
assign addr[10006]= -1332945355;
assign addr[10007]= -1080359326;
assign addr[10008]= -805879757;
assign addr[10009]= -515068990;
assign addr[10010]= -213820322;
assign addr[10011]= 91761426;
assign addr[10012]= 395483624;
assign addr[10013]= 691191324;
assign addr[10014]= 972891995;
assign addr[10015]= 1234876957;
assign addr[10016]= 1471837070;
assign addr[10017]= 1678970324;
assign addr[10018]= 1852079154;
assign addr[10019]= 1987655498;
assign addr[10020]= 2082951896;
assign addr[10021]= 2136037160;
assign addr[10022]= 2145835515;
assign addr[10023]= 2112148396;
assign addr[10024]= 2035658475;
assign addr[10025]= 1917915825;
assign addr[10026]= 1761306505;
assign addr[10027]= 1569004214;
assign addr[10028]= 1344905966;
assign addr[10029]= 1093553126;
assign addr[10030]= 820039373;
assign addr[10031]= 529907477;
assign addr[10032]= 229036977;
assign addr[10033]= -76474970;
assign addr[10034]= -380437148;
assign addr[10035]= -676689746;
assign addr[10036]= -959229189;
assign addr[10037]= -1222329801;
assign addr[10038]= -1460659832;
assign addr[10039]= -1669389513;
assign addr[10040]= -1844288924;
assign addr[10041]= -1981813720;
assign addr[10042]= -2079176953;
assign addr[10043]= -2134405552;
assign addr[10044]= -2146380306;
assign addr[10045]= -2114858546;
assign addr[10046]= -2040479063;
assign addr[10047]= -1924749160;
assign addr[10048]= -1770014111;
assign addr[10049]= -1579409630;
assign addr[10050]= -1356798326;
assign addr[10051]= -1106691431;
assign addr[10052]= -834157373;
assign addr[10053]= -544719071;
assign addr[10054]= -244242007;
assign addr[10055]= 61184634;
assign addr[10056]= 365371365;
assign addr[10057]= 662153826;
assign addr[10058]= 945517704;
assign addr[10059]= 1209720613;
assign addr[10060]= 1449408469;
assign addr[10061]= 1659723983;
assign addr[10062]= 1836405100;
assign addr[10063]= 1975871368;
assign addr[10064]= 2075296495;
assign addr[10065]= 2132665626;
assign addr[10066]= 2146816171;
assign addr[10067]= 2117461370;
assign addr[10068]= 2045196100;
assign addr[10069]= 1931484818;
assign addr[10070]= 1778631892;
assign addr[10071]= 1589734894;
assign addr[10072]= 1368621831;
assign addr[10073]= 1119773573;
assign addr[10074]= 848233042;
assign addr[10075]= 559503022;
assign addr[10076]= 259434643;
assign addr[10077]= -45891193;
assign addr[10078]= -350287041;
assign addr[10079]= -647584304;
assign addr[10080]= -931758235;
assign addr[10081]= -1197050035;
assign addr[10082]= -1438083551;
assign addr[10083]= -1649974225;
assign addr[10084]= -1828428082;
assign addr[10085]= -1969828744;
assign addr[10086]= -2071310720;
assign addr[10087]= -2130817471;
assign addr[10088]= -2147143090;
assign addr[10089]= -2119956737;
assign addr[10090]= -2049809346;
assign addr[10091]= -1938122457;
assign addr[10092]= -1787159411;
assign addr[10093]= -1599979481;
assign addr[10094]= -1380375881;
assign addr[10095]= -1132798888;
assign addr[10096]= -862265664;
assign addr[10097]= -574258580;
assign addr[10098]= -274614114;
assign addr[10099]= 30595422;
assign addr[10100]= 335184940;
assign addr[10101]= 632981917;
assign addr[10102]= 917951481;
assign addr[10103]= 1184318708;
assign addr[10104]= 1426685652;
assign addr[10105]= 1640140734;
assign addr[10106]= 1820358275;
assign addr[10107]= 1963686155;
assign addr[10108]= 2067219829;
assign addr[10109]= 2128861181;
assign addr[10110]= 2147361045;
assign addr[10111]= 2122344521;
assign addr[10112]= 2054318569;
assign addr[10113]= 1944661739;
assign addr[10114]= 1795596234;
assign addr[10115]= 1610142873;
assign addr[10116]= 1392059879;
assign addr[10117]= 1145766716;
assign addr[10118]= 876254528;
assign addr[10119]= 588984994;
assign addr[10120]= 289779648;
assign addr[10121]= -15298099;
assign addr[10122]= -320065829;
assign addr[10123]= -618347408;
assign addr[10124]= -904098143;
assign addr[10125]= -1171527280;
assign addr[10126]= -1415215352;
assign addr[10127]= -1630224009;
assign addr[10128]= -1812196087;
assign addr[10129]= -1957443913;
assign addr[10130]= -2063024031;
assign addr[10131]= -2126796855;
assign addr[10132]= -2147470025;
assign addr[10133]= -2124624598;
assign addr[10134]= -2058723538;
assign addr[10135]= -1951102334;
assign addr[10136]= -1803941934;
assign addr[10137]= -1620224553;
assign addr[10138]= -1403673233;
assign addr[10139]= -1158676398;
assign addr[10140]= -890198924;
assign addr[10141]= -603681519;
assign addr[10142]= -304930476;
assign addr[10143]= 0;
assign addr[10144]= 304930476;
assign addr[10145]= 603681519;
assign addr[10146]= 890198924;
assign addr[10147]= 1158676398;
assign addr[10148]= 1403673233;
assign addr[10149]= 1620224553;
assign addr[10150]= 1803941934;
assign addr[10151]= 1951102334;
assign addr[10152]= 2058723538;
assign addr[10153]= 2124624598;
assign addr[10154]= 2147470025;
assign addr[10155]= 2126796855;
assign addr[10156]= 2063024031;
assign addr[10157]= 1957443913;
assign addr[10158]= 1812196087;
assign addr[10159]= 1630224009;
assign addr[10160]= 1415215352;
assign addr[10161]= 1171527280;
assign addr[10162]= 904098143;
assign addr[10163]= 618347408;
assign addr[10164]= 320065829;
assign addr[10165]= 15298099;
assign addr[10166]= -289779648;
assign addr[10167]= -588984994;
assign addr[10168]= -876254528;
assign addr[10169]= -1145766716;
assign addr[10170]= -1392059879;
assign addr[10171]= -1610142873;
assign addr[10172]= -1795596234;
assign addr[10173]= -1944661739;
assign addr[10174]= -2054318569;
assign addr[10175]= -2122344521;
assign addr[10176]= -2147361045;
assign addr[10177]= -2128861181;
assign addr[10178]= -2067219829;
assign addr[10179]= -1963686155;
assign addr[10180]= -1820358275;
assign addr[10181]= -1640140734;
assign addr[10182]= -1426685652;
assign addr[10183]= -1184318708;
assign addr[10184]= -917951481;
assign addr[10185]= -632981917;
assign addr[10186]= -335184940;
assign addr[10187]= -30595422;
assign addr[10188]= 274614114;
assign addr[10189]= 574258580;
assign addr[10190]= 862265664;
assign addr[10191]= 1132798888;
assign addr[10192]= 1380375881;
assign addr[10193]= 1599979481;
assign addr[10194]= 1787159411;
assign addr[10195]= 1938122457;
assign addr[10196]= 2049809346;
assign addr[10197]= 2119956737;
assign addr[10198]= 2147143090;
assign addr[10199]= 2130817471;
assign addr[10200]= 2071310720;
assign addr[10201]= 1969828744;
assign addr[10202]= 1828428082;
assign addr[10203]= 1649974225;
assign addr[10204]= 1438083551;
assign addr[10205]= 1197050035;
assign addr[10206]= 931758235;
assign addr[10207]= 647584304;
assign addr[10208]= 350287041;
assign addr[10209]= 45891193;
assign addr[10210]= -259434643;
assign addr[10211]= -559503022;
assign addr[10212]= -848233042;
assign addr[10213]= -1119773573;
assign addr[10214]= -1368621831;
assign addr[10215]= -1589734894;
assign addr[10216]= -1778631892;
assign addr[10217]= -1931484818;
assign addr[10218]= -2045196100;
assign addr[10219]= -2117461370;
assign addr[10220]= -2146816171;
assign addr[10221]= -2132665626;
assign addr[10222]= -2075296495;
assign addr[10223]= -1975871368;
assign addr[10224]= -1836405100;
assign addr[10225]= -1659723983;
assign addr[10226]= -1449408469;
assign addr[10227]= -1209720613;
assign addr[10228]= -945517704;
assign addr[10229]= -662153826;
assign addr[10230]= -365371365;
assign addr[10231]= -61184634;
assign addr[10232]= 244242007;
assign addr[10233]= 544719071;
assign addr[10234]= 834157373;
assign addr[10235]= 1106691431;
assign addr[10236]= 1356798326;
assign addr[10237]= 1579409630;
assign addr[10238]= 1770014111;
assign addr[10239]= 1924749160;
assign addr[10240]= 2040479063;
assign addr[10241]= 2114858546;
assign addr[10242]= 2146380306;
assign addr[10243]= 2134405552;
assign addr[10244]= 2079176953;
assign addr[10245]= 1981813720;
assign addr[10246]= 1844288924;
assign addr[10247]= 1669389513;
assign addr[10248]= 1460659832;
assign addr[10249]= 1222329801;
assign addr[10250]= 959229189;
assign addr[10251]= 676689746;
assign addr[10252]= 380437148;
assign addr[10253]= 76474970;
assign addr[10254]= -229036977;
assign addr[10255]= -529907477;
assign addr[10256]= -820039373;
assign addr[10257]= -1093553126;
assign addr[10258]= -1344905966;
assign addr[10259]= -1569004214;
assign addr[10260]= -1761306505;
assign addr[10261]= -1917915825;
assign addr[10262]= -2035658475;
assign addr[10263]= -2112148396;
assign addr[10264]= -2145835515;
assign addr[10265]= -2136037160;
assign addr[10266]= -2082951896;
assign addr[10267]= -1987655498;
assign addr[10268]= -1852079154;
assign addr[10269]= -1678970324;
assign addr[10270]= -1471837070;
assign addr[10271]= -1234876957;
assign addr[10272]= -972891995;
assign addr[10273]= -691191324;
assign addr[10274]= -395483624;
assign addr[10275]= -91761426;
assign addr[10276]= 213820322;
assign addr[10277]= 515068990;
assign addr[10278]= 805879757;
assign addr[10279]= 1080359326;
assign addr[10280]= 1332945355;
assign addr[10281]= 1558519173;
assign addr[10282]= 1752509516;
assign addr[10283]= 1910985158;
assign addr[10284]= 2030734582;
assign addr[10285]= 2109331059;
assign addr[10286]= 2145181827;
assign addr[10287]= 2137560369;
assign addr[10288]= 2086621133;
assign addr[10289]= 1993396407;
assign addr[10290]= 1859775393;
assign addr[10291]= 1688465931;
assign addr[10292]= 1482939614;
assign addr[10293]= 1247361445;
assign addr[10294]= 986505429;
assign addr[10295]= 705657826;
assign addr[10296]= 410510029;
assign addr[10297]= 107043224;
assign addr[10298]= -198592817;
assign addr[10299]= -500204365;
assign addr[10300]= -791679244;
assign addr[10301]= -1067110699;
assign addr[10302]= -1320917099;
assign addr[10303]= -1547955041;
assign addr[10304]= -1743623590;
assign addr[10305]= -1903957513;
assign addr[10306]= -2025707632;
assign addr[10307]= -2106406677;
assign addr[10308]= -2144419275;
assign addr[10309]= -2138975100;
assign addr[10310]= -2090184478;
assign addr[10311]= -1999036154;
assign addr[10312]= -1867377253;
assign addr[10313]= -1697875851;
assign addr[10314]= -1493966902;
assign addr[10315]= -1259782632;
assign addr[10316]= -1000068799;
assign addr[10317]= -720088517;
assign addr[10318]= -425515602;
assign addr[10319]= -122319591;
assign addr[10320]= 183355234;
assign addr[10321]= 485314355;
assign addr[10322]= 777438554;
assign addr[10323]= 1053807919;
assign addr[10324]= 1308821808;
assign addr[10325]= 1537312353;
assign addr[10326]= 1734649179;
assign addr[10327]= 1896833245;
assign addr[10328]= 2020577882;
assign addr[10329]= 2103375398;
assign addr[10330]= 2143547897;
assign addr[10331]= 2140281282;
assign addr[10332]= 2093641749;
assign addr[10333]= 2004574453;
assign addr[10334]= 1874884346;
assign addr[10335]= 1707199606;
assign addr[10336]= 1504918373;
assign addr[10337]= 1272139887;
assign addr[10338]= 1013581418;
assign addr[10339]= 734482665;
assign addr[10340]= 440499581;
assign addr[10341]= 137589750;
assign addr[10342]= -168108346;
assign addr[10343]= -470399716;
assign addr[10344]= -763158411;
assign addr[10345]= -1040451659;
assign addr[10346]= -1296660098;
assign addr[10347]= -1526591649;
assign addr[10348]= -1725586737;
assign addr[10349]= -1889612716;
assign addr[10350]= -2015345591;
assign addr[10351]= -2100237377;
assign addr[10352]= -2142567738;
assign addr[10353]= -2141478848;
assign addr[10354]= -2096992772;
assign addr[10355]= -2010011024;
assign addr[10356]= -1882296293;
assign addr[10357]= -1716436725;
assign addr[10358]= -1515793473;
assign addr[10359]= -1284432584;
assign addr[10360]= -1027042599;
assign addr[10361]= -748839539;
assign addr[10362]= -455461206;
assign addr[10363]= -152852926;
assign addr[10364]= 152852926;
assign addr[10365]= 455461206;
assign addr[10366]= 748839539;
assign addr[10367]= 1027042599;
assign addr[10368]= 1284432584;
assign addr[10369]= 1515793473;
assign addr[10370]= 1716436725;
assign addr[10371]= 1882296293;
assign addr[10372]= 2010011024;
assign addr[10373]= 2096992772;
assign addr[10374]= 2141478848;
assign addr[10375]= 2142567738;
assign addr[10376]= 2100237377;
assign addr[10377]= 2015345591;
assign addr[10378]= 1889612716;
assign addr[10379]= 1725586737;
assign addr[10380]= 1526591649;
assign addr[10381]= 1296660098;
assign addr[10382]= 1040451659;
assign addr[10383]= 763158411;
assign addr[10384]= 470399716;
assign addr[10385]= 168108346;
assign addr[10386]= -137589750;
assign addr[10387]= -440499581;
assign addr[10388]= -734482665;
assign addr[10389]= -1013581418;
assign addr[10390]= -1272139887;
assign addr[10391]= -1504918373;
assign addr[10392]= -1707199606;
assign addr[10393]= -1874884346;
assign addr[10394]= -2004574453;
assign addr[10395]= -2093641749;
assign addr[10396]= -2140281282;
assign addr[10397]= -2143547897;
assign addr[10398]= -2103375398;
assign addr[10399]= -2020577882;
assign addr[10400]= -1896833245;
assign addr[10401]= -1734649179;
assign addr[10402]= -1537312353;
assign addr[10403]= -1308821808;
assign addr[10404]= -1053807919;
assign addr[10405]= -777438554;
assign addr[10406]= -485314355;
assign addr[10407]= -183355234;
assign addr[10408]= 122319591;
assign addr[10409]= 425515602;
assign addr[10410]= 720088517;
assign addr[10411]= 1000068799;
assign addr[10412]= 1259782632;
assign addr[10413]= 1493966902;
assign addr[10414]= 1697875851;
assign addr[10415]= 1867377253;
assign addr[10416]= 1999036154;
assign addr[10417]= 2090184478;
assign addr[10418]= 2138975100;
assign addr[10419]= 2144419275;
assign addr[10420]= 2106406677;
assign addr[10421]= 2025707632;
assign addr[10422]= 1903957513;
assign addr[10423]= 1743623590;
assign addr[10424]= 1547955041;
assign addr[10425]= 1320917099;
assign addr[10426]= 1067110699;
assign addr[10427]= 791679244;
assign addr[10428]= 500204365;
assign addr[10429]= 198592817;
assign addr[10430]= -107043224;
assign addr[10431]= -410510029;
assign addr[10432]= -705657826;
assign addr[10433]= -986505429;
assign addr[10434]= -1247361445;
assign addr[10435]= -1482939614;
assign addr[10436]= -1688465931;
assign addr[10437]= -1859775393;
assign addr[10438]= -1993396407;
assign addr[10439]= -2086621133;
assign addr[10440]= -2137560369;
assign addr[10441]= -2145181827;
assign addr[10442]= -2109331059;
assign addr[10443]= -2030734582;
assign addr[10444]= -1910985158;
assign addr[10445]= -1752509516;
assign addr[10446]= -1558519173;
assign addr[10447]= -1332945355;
assign addr[10448]= -1080359326;
assign addr[10449]= -805879757;
assign addr[10450]= -515068990;
assign addr[10451]= -213820322;
assign addr[10452]= 91761426;
assign addr[10453]= 395483624;
assign addr[10454]= 691191324;
assign addr[10455]= 972891995;
assign addr[10456]= 1234876957;
assign addr[10457]= 1471837070;
assign addr[10458]= 1678970324;
assign addr[10459]= 1852079154;
assign addr[10460]= 1987655498;
assign addr[10461]= 2082951896;
assign addr[10462]= 2136037160;
assign addr[10463]= 2145835515;
assign addr[10464]= 2112148396;
assign addr[10465]= 2035658475;
assign addr[10466]= 1917915825;
assign addr[10467]= 1761306505;
assign addr[10468]= 1569004214;
assign addr[10469]= 1344905966;
assign addr[10470]= 1093553126;
assign addr[10471]= 820039373;
assign addr[10472]= 529907477;
assign addr[10473]= 229036977;
assign addr[10474]= -76474970;
assign addr[10475]= -380437148;
assign addr[10476]= -676689746;
assign addr[10477]= -959229189;
assign addr[10478]= -1222329801;
assign addr[10479]= -1460659832;
assign addr[10480]= -1669389513;
assign addr[10481]= -1844288924;
assign addr[10482]= -1981813720;
assign addr[10483]= -2079176953;
assign addr[10484]= -2134405552;
assign addr[10485]= -2146380306;
assign addr[10486]= -2114858546;
assign addr[10487]= -2040479063;
assign addr[10488]= -1924749160;
assign addr[10489]= -1770014111;
assign addr[10490]= -1579409630;
assign addr[10491]= -1356798326;
assign addr[10492]= -1106691431;
assign addr[10493]= -834157373;
assign addr[10494]= -544719071;
assign addr[10495]= -244242007;
assign addr[10496]= 61184634;
assign addr[10497]= 365371365;
assign addr[10498]= 662153826;
assign addr[10499]= 945517704;
assign addr[10500]= 1209720613;
assign addr[10501]= 1449408469;
assign addr[10502]= 1659723983;
assign addr[10503]= 1836405100;
assign addr[10504]= 1975871368;
assign addr[10505]= 2075296495;
assign addr[10506]= 2132665626;
assign addr[10507]= 2146816171;
assign addr[10508]= 2117461370;
assign addr[10509]= 2045196100;
assign addr[10510]= 1931484818;
assign addr[10511]= 1778631892;
assign addr[10512]= 1589734894;
assign addr[10513]= 1368621831;
assign addr[10514]= 1119773573;
assign addr[10515]= 848233042;
assign addr[10516]= 559503022;
assign addr[10517]= 259434643;
assign addr[10518]= -45891193;
assign addr[10519]= -350287041;
assign addr[10520]= -647584304;
assign addr[10521]= -931758235;
assign addr[10522]= -1197050035;
assign addr[10523]= -1438083551;
assign addr[10524]= -1649974225;
assign addr[10525]= -1828428082;
assign addr[10526]= -1969828744;
assign addr[10527]= -2071310720;
assign addr[10528]= -2130817471;
assign addr[10529]= -2147143090;
assign addr[10530]= -2119956737;
assign addr[10531]= -2049809346;
assign addr[10532]= -1938122457;
assign addr[10533]= -1787159411;
assign addr[10534]= -1599979481;
assign addr[10535]= -1380375881;
assign addr[10536]= -1132798888;
assign addr[10537]= -862265664;
assign addr[10538]= -574258580;
assign addr[10539]= -274614114;
assign addr[10540]= 30595422;
assign addr[10541]= 335184940;
assign addr[10542]= 632981917;
assign addr[10543]= 917951481;
assign addr[10544]= 1184318708;
assign addr[10545]= 1426685652;
assign addr[10546]= 1640140734;
assign addr[10547]= 1820358275;
assign addr[10548]= 1963686155;
assign addr[10549]= 2067219829;
assign addr[10550]= 2128861181;
assign addr[10551]= 2147361045;
assign addr[10552]= 2122344521;
assign addr[10553]= 2054318569;
assign addr[10554]= 1944661739;
assign addr[10555]= 1795596234;
assign addr[10556]= 1610142873;
assign addr[10557]= 1392059879;
assign addr[10558]= 1145766716;
assign addr[10559]= 876254528;
assign addr[10560]= 588984994;
assign addr[10561]= 289779648;
assign addr[10562]= -15298099;
assign addr[10563]= -320065829;
assign addr[10564]= -618347408;
assign addr[10565]= -904098143;
assign addr[10566]= -1171527280;
assign addr[10567]= -1415215352;
assign addr[10568]= -1630224009;
assign addr[10569]= -1812196087;
assign addr[10570]= -1957443913;
assign addr[10571]= -2063024031;
assign addr[10572]= -2126796855;
assign addr[10573]= -2147470025;
assign addr[10574]= -2124624598;
assign addr[10575]= -2058723538;
assign addr[10576]= -1951102334;
assign addr[10577]= -1803941934;
assign addr[10578]= -1620224553;
assign addr[10579]= -1403673233;
assign addr[10580]= -1158676398;
assign addr[10581]= -890198924;
assign addr[10582]= -603681519;
assign addr[10583]= -304930476;
assign addr[10584]= 0;
assign addr[10585]= 304930476;
assign addr[10586]= 603681519;
assign addr[10587]= 890198924;
assign addr[10588]= 1158676398;
assign addr[10589]= 1403673233;
assign addr[10590]= 1620224553;
assign addr[10591]= 1803941934;
assign addr[10592]= 1951102334;
assign addr[10593]= 2058723538;
assign addr[10594]= 2124624598;
assign addr[10595]= 2147470025;
assign addr[10596]= 2126796855;
assign addr[10597]= 2063024031;
assign addr[10598]= 1957443913;
assign addr[10599]= 1812196087;
assign addr[10600]= 1630224009;
assign addr[10601]= 1415215352;
assign addr[10602]= 1171527280;
assign addr[10603]= 904098143;
assign addr[10604]= 618347408;
assign addr[10605]= 320065829;
assign addr[10606]= 15298099;
assign addr[10607]= -289779648;
assign addr[10608]= -588984994;
assign addr[10609]= -876254528;
assign addr[10610]= -1145766716;
assign addr[10611]= -1392059879;
assign addr[10612]= -1610142873;
assign addr[10613]= -1795596234;
assign addr[10614]= -1944661739;
assign addr[10615]= -2054318569;
assign addr[10616]= -2122344521;
assign addr[10617]= -2147361045;
assign addr[10618]= -2128861181;
assign addr[10619]= -2067219829;
assign addr[10620]= -1963686155;
assign addr[10621]= -1820358275;
assign addr[10622]= -1640140734;
assign addr[10623]= -1426685652;
assign addr[10624]= -1184318708;
assign addr[10625]= -917951481;
assign addr[10626]= -632981917;
assign addr[10627]= -335184940;
assign addr[10628]= -30595422;
assign addr[10629]= 274614114;
assign addr[10630]= 574258580;
assign addr[10631]= 862265664;
assign addr[10632]= 1132798888;
assign addr[10633]= 1380375881;
assign addr[10634]= 1599979481;
assign addr[10635]= 1787159411;
assign addr[10636]= 1938122457;
assign addr[10637]= 2049809346;
assign addr[10638]= 2119956737;
assign addr[10639]= 2147143090;
assign addr[10640]= 2130817471;
assign addr[10641]= 2071310720;
assign addr[10642]= 1969828744;
assign addr[10643]= 1828428082;
assign addr[10644]= 1649974225;
assign addr[10645]= 1438083551;
assign addr[10646]= 1197050035;
assign addr[10647]= 931758235;
assign addr[10648]= 647584304;
assign addr[10649]= 350287041;
assign addr[10650]= 45891193;
assign addr[10651]= -259434643;
assign addr[10652]= -559503022;
assign addr[10653]= -848233042;
assign addr[10654]= -1119773573;
assign addr[10655]= -1368621831;
assign addr[10656]= -1589734894;
assign addr[10657]= -1778631892;
assign addr[10658]= -1931484818;
assign addr[10659]= -2045196100;
assign addr[10660]= -2117461370;
assign addr[10661]= -2146816171;
assign addr[10662]= -2132665626;
assign addr[10663]= -2075296495;
assign addr[10664]= -1975871368;
assign addr[10665]= -1836405100;
assign addr[10666]= -1659723983;
assign addr[10667]= -1449408469;
assign addr[10668]= -1209720613;
assign addr[10669]= -945517704;
assign addr[10670]= -662153826;
assign addr[10671]= -365371365;
assign addr[10672]= -61184634;
assign addr[10673]= 244242007;
assign addr[10674]= 544719071;
assign addr[10675]= 834157373;
assign addr[10676]= 1106691431;
assign addr[10677]= 1356798326;
assign addr[10678]= 1579409630;
assign addr[10679]= 1770014111;
assign addr[10680]= 1924749160;
assign addr[10681]= 2040479063;
assign addr[10682]= 2114858546;
assign addr[10683]= 2146380306;
assign addr[10684]= 2134405552;
assign addr[10685]= 2079176953;
assign addr[10686]= 1981813720;
assign addr[10687]= 1844288924;
assign addr[10688]= 1669389513;
assign addr[10689]= 1460659832;
assign addr[10690]= 1222329801;
assign addr[10691]= 959229189;
assign addr[10692]= 676689746;
assign addr[10693]= 380437148;
assign addr[10694]= 76474970;
assign addr[10695]= -229036977;
assign addr[10696]= -529907477;
assign addr[10697]= -820039373;
assign addr[10698]= -1093553126;
assign addr[10699]= -1344905966;
assign addr[10700]= -1569004214;
assign addr[10701]= -1761306505;
assign addr[10702]= -1917915825;
assign addr[10703]= -2035658475;
assign addr[10704]= -2112148396;
assign addr[10705]= -2145835515;
assign addr[10706]= -2136037160;
assign addr[10707]= -2082951896;
assign addr[10708]= -1987655498;
assign addr[10709]= -1852079154;
assign addr[10710]= -1678970324;
assign addr[10711]= -1471837070;
assign addr[10712]= -1234876957;
assign addr[10713]= -972891995;
assign addr[10714]= -691191324;
assign addr[10715]= -395483624;
assign addr[10716]= -91761426;
assign addr[10717]= 213820322;
assign addr[10718]= 515068990;
assign addr[10719]= 805879757;
assign addr[10720]= 1080359326;
assign addr[10721]= 1332945355;
assign addr[10722]= 1558519173;
assign addr[10723]= 1752509516;
assign addr[10724]= 1910985158;
assign addr[10725]= 2030734582;
assign addr[10726]= 2109331059;
assign addr[10727]= 2145181827;
assign addr[10728]= 2137560369;
assign addr[10729]= 2086621133;
assign addr[10730]= 1993396407;
assign addr[10731]= 1859775393;
assign addr[10732]= 1688465931;
assign addr[10733]= 1482939614;
assign addr[10734]= 1247361445;
assign addr[10735]= 986505429;
assign addr[10736]= 705657826;
assign addr[10737]= 410510029;
assign addr[10738]= 107043224;
assign addr[10739]= -198592817;
assign addr[10740]= -500204365;
assign addr[10741]= -791679244;
assign addr[10742]= -1067110699;
assign addr[10743]= -1320917099;
assign addr[10744]= -1547955041;
assign addr[10745]= -1743623590;
assign addr[10746]= -1903957513;
assign addr[10747]= -2025707632;
assign addr[10748]= -2106406677;
assign addr[10749]= -2144419275;
assign addr[10750]= -2138975100;
assign addr[10751]= -2090184478;
assign addr[10752]= -1999036154;
assign addr[10753]= -1867377253;
assign addr[10754]= -1697875851;
assign addr[10755]= -1493966902;
assign addr[10756]= -1259782632;
assign addr[10757]= -1000068799;
assign addr[10758]= -720088517;
assign addr[10759]= -425515602;
assign addr[10760]= -122319591;
assign addr[10761]= 183355234;
assign addr[10762]= 485314355;
assign addr[10763]= 777438554;
assign addr[10764]= 1053807919;
assign addr[10765]= 1308821808;
assign addr[10766]= 1537312353;
assign addr[10767]= 1734649179;
assign addr[10768]= 1896833245;
assign addr[10769]= 2020577882;
assign addr[10770]= 2103375398;
assign addr[10771]= 2143547897;
assign addr[10772]= 2140281282;
assign addr[10773]= 2093641749;
assign addr[10774]= 2004574453;
assign addr[10775]= 1874884346;
assign addr[10776]= 1707199606;
assign addr[10777]= 1504918373;
assign addr[10778]= 1272139887;
assign addr[10779]= 1013581418;
assign addr[10780]= 734482665;
assign addr[10781]= 440499581;
assign addr[10782]= 137589750;
assign addr[10783]= -168108346;
assign addr[10784]= -470399716;
assign addr[10785]= -763158411;
assign addr[10786]= -1040451659;
assign addr[10787]= -1296660098;
assign addr[10788]= -1526591649;
assign addr[10789]= -1725586737;
assign addr[10790]= -1889612716;
assign addr[10791]= -2015345591;
assign addr[10792]= -2100237377;
assign addr[10793]= -2142567738;
assign addr[10794]= -2141478848;
assign addr[10795]= -2096992772;
assign addr[10796]= -2010011024;
assign addr[10797]= -1882296293;
assign addr[10798]= -1716436725;
assign addr[10799]= -1515793473;
assign addr[10800]= -1284432584;
assign addr[10801]= -1027042599;
assign addr[10802]= -748839539;
assign addr[10803]= -455461206;
assign addr[10804]= -152852926;
assign addr[10805]= 152852926;
assign addr[10806]= 455461206;
assign addr[10807]= 748839539;
assign addr[10808]= 1027042599;
assign addr[10809]= 1284432584;
assign addr[10810]= 1515793473;
assign addr[10811]= 1716436725;
assign addr[10812]= 1882296293;
assign addr[10813]= 2010011024;
assign addr[10814]= 2096992772;
assign addr[10815]= 2141478848;
assign addr[10816]= 2142567738;
assign addr[10817]= 2100237377;
assign addr[10818]= 2015345591;
assign addr[10819]= 1889612716;
assign addr[10820]= 1725586737;
assign addr[10821]= 1526591649;
assign addr[10822]= 1296660098;
assign addr[10823]= 1040451659;
assign addr[10824]= 763158411;
assign addr[10825]= 470399716;
assign addr[10826]= 168108346;
assign addr[10827]= -137589750;
assign addr[10828]= -440499581;
assign addr[10829]= -734482665;
assign addr[10830]= -1013581418;
assign addr[10831]= -1272139887;
assign addr[10832]= -1504918373;
assign addr[10833]= -1707199606;
assign addr[10834]= -1874884346;
assign addr[10835]= -2004574453;
assign addr[10836]= -2093641749;
assign addr[10837]= -2140281282;
assign addr[10838]= -2143547897;
assign addr[10839]= -2103375398;
assign addr[10840]= -2020577882;
assign addr[10841]= -1896833245;
assign addr[10842]= -1734649179;
assign addr[10843]= -1537312353;
assign addr[10844]= -1308821808;
assign addr[10845]= -1053807919;
assign addr[10846]= -777438554;
assign addr[10847]= -485314355;
assign addr[10848]= -183355234;
assign addr[10849]= 122319591;
assign addr[10850]= 425515602;
assign addr[10851]= 720088517;
assign addr[10852]= 1000068799;
assign addr[10853]= 1259782632;
assign addr[10854]= 1493966902;
assign addr[10855]= 1697875851;
assign addr[10856]= 1867377253;
assign addr[10857]= 1999036154;
assign addr[10858]= 2090184478;
assign addr[10859]= 2138975100;
assign addr[10860]= 2144419275;
assign addr[10861]= 2106406677;
assign addr[10862]= 2025707632;
assign addr[10863]= 1903957513;
assign addr[10864]= 1743623590;
assign addr[10865]= 1547955041;
assign addr[10866]= 1320917099;
assign addr[10867]= 1067110699;
assign addr[10868]= 791679244;
assign addr[10869]= 500204365;
assign addr[10870]= 198592817;
assign addr[10871]= -107043224;
assign addr[10872]= -410510029;
assign addr[10873]= -705657826;
assign addr[10874]= -986505429;
assign addr[10875]= -1247361445;
assign addr[10876]= -1482939614;
assign addr[10877]= -1688465931;
assign addr[10878]= -1859775393;
assign addr[10879]= -1993396407;
assign addr[10880]= -2086621133;
assign addr[10881]= -2137560369;
assign addr[10882]= -2145181827;
assign addr[10883]= -2109331059;
assign addr[10884]= -2030734582;
assign addr[10885]= -1910985158;
assign addr[10886]= -1752509516;
assign addr[10887]= -1558519173;
assign addr[10888]= -1332945355;
assign addr[10889]= -1080359326;
assign addr[10890]= -805879757;
assign addr[10891]= -515068990;
assign addr[10892]= -213820322;
assign addr[10893]= 91761426;
assign addr[10894]= 395483624;
assign addr[10895]= 691191324;
assign addr[10896]= 972891995;
assign addr[10897]= 1234876957;
assign addr[10898]= 1471837070;
assign addr[10899]= 1678970324;
assign addr[10900]= 1852079154;
assign addr[10901]= 1987655498;
assign addr[10902]= 2082951896;
assign addr[10903]= 2136037160;
assign addr[10904]= 2145835515;
assign addr[10905]= 2112148396;
assign addr[10906]= 2035658475;
assign addr[10907]= 1917915825;
assign addr[10908]= 1761306505;
assign addr[10909]= 1569004214;
assign addr[10910]= 1344905966;
assign addr[10911]= 1093553126;
assign addr[10912]= 820039373;
assign addr[10913]= 529907477;
assign addr[10914]= 229036977;
assign addr[10915]= -76474970;
assign addr[10916]= -380437148;
assign addr[10917]= -676689746;
assign addr[10918]= -959229189;
assign addr[10919]= -1222329801;
assign addr[10920]= -1460659832;
assign addr[10921]= -1669389513;
assign addr[10922]= -1844288924;
assign addr[10923]= -1981813720;
assign addr[10924]= -2079176953;
assign addr[10925]= -2134405552;
assign addr[10926]= -2146380306;
assign addr[10927]= -2114858546;
assign addr[10928]= -2040479063;
assign addr[10929]= -1924749160;
assign addr[10930]= -1770014111;
assign addr[10931]= -1579409630;
assign addr[10932]= -1356798326;
assign addr[10933]= -1106691431;
assign addr[10934]= -834157373;
assign addr[10935]= -544719071;
assign addr[10936]= -244242007;
assign addr[10937]= 61184634;
assign addr[10938]= 365371365;
assign addr[10939]= 662153826;
assign addr[10940]= 945517704;
assign addr[10941]= 1209720613;
assign addr[10942]= 1449408469;
assign addr[10943]= 1659723983;
assign addr[10944]= 1836405100;
assign addr[10945]= 1975871368;
assign addr[10946]= 2075296495;
assign addr[10947]= 2132665626;
assign addr[10948]= 2146816171;
assign addr[10949]= 2117461370;
assign addr[10950]= 2045196100;
assign addr[10951]= 1931484818;
assign addr[10952]= 1778631892;
assign addr[10953]= 1589734894;
assign addr[10954]= 1368621831;
assign addr[10955]= 1119773573;
assign addr[10956]= 848233042;
assign addr[10957]= 559503022;
assign addr[10958]= 259434643;
assign addr[10959]= -45891193;
assign addr[10960]= -350287041;
assign addr[10961]= -647584304;
assign addr[10962]= -931758235;
assign addr[10963]= -1197050035;
assign addr[10964]= -1438083551;
assign addr[10965]= -1649974225;
assign addr[10966]= -1828428082;
assign addr[10967]= -1969828744;
assign addr[10968]= -2071310720;
assign addr[10969]= -2130817471;
assign addr[10970]= -2147143090;
assign addr[10971]= -2119956737;
assign addr[10972]= -2049809346;
assign addr[10973]= -1938122457;
assign addr[10974]= -1787159411;
assign addr[10975]= -1599979481;
assign addr[10976]= -1380375881;
assign addr[10977]= -1132798888;
assign addr[10978]= -862265664;
assign addr[10979]= -574258580;
assign addr[10980]= -274614114;
assign addr[10981]= 30595422;
assign addr[10982]= 335184940;
assign addr[10983]= 632981917;
assign addr[10984]= 917951481;
assign addr[10985]= 1184318708;
assign addr[10986]= 1426685652;
assign addr[10987]= 1640140734;
assign addr[10988]= 1820358275;
assign addr[10989]= 1963686155;
assign addr[10990]= 2067219829;
assign addr[10991]= 2128861181;
assign addr[10992]= 2147361045;
assign addr[10993]= 2122344521;
assign addr[10994]= 2054318569;
assign addr[10995]= 1944661739;
assign addr[10996]= 1795596234;
assign addr[10997]= 1610142873;
assign addr[10998]= 1392059879;
assign addr[10999]= 1145766716;
assign addr[11000]= 876254528;
assign addr[11001]= 588984994;
assign addr[11002]= 289779648;
assign addr[11003]= -15298099;
assign addr[11004]= -320065829;
assign addr[11005]= -618347408;
assign addr[11006]= -904098143;
assign addr[11007]= -1171527280;
assign addr[11008]= -1415215352;
assign addr[11009]= -1630224009;
assign addr[11010]= -1812196087;
assign addr[11011]= -1957443913;
assign addr[11012]= -2063024031;
assign addr[11013]= -2126796855;
assign addr[11014]= -2147470025;
assign addr[11015]= -2124624598;
assign addr[11016]= -2058723538;
assign addr[11017]= -1951102334;
assign addr[11018]= -1803941934;
assign addr[11019]= -1620224553;
assign addr[11020]= -1403673233;
assign addr[11021]= -1158676398;
assign addr[11022]= -890198924;
assign addr[11023]= -603681519;
assign addr[11024]= -304930476;
assign addr[11025]= 0;
assign addr[11026]= 304930476;
assign addr[11027]= 603681519;
assign addr[11028]= 890198924;
assign addr[11029]= 1158676398;
assign addr[11030]= 1403673233;
assign addr[11031]= 1620224553;
assign addr[11032]= 1803941934;
assign addr[11033]= 1951102334;
assign addr[11034]= 2058723538;
assign addr[11035]= 2124624598;
assign addr[11036]= 2147470025;
assign addr[11037]= 2126796855;
assign addr[11038]= 2063024031;
assign addr[11039]= 1957443913;
assign addr[11040]= 1812196087;
assign addr[11041]= 1630224009;
assign addr[11042]= 1415215352;
assign addr[11043]= 1171527280;
assign addr[11044]= 904098143;
assign addr[11045]= 618347408;
assign addr[11046]= 320065829;
assign addr[11047]= 15298099;
assign addr[11048]= -289779648;
assign addr[11049]= -588984994;
assign addr[11050]= -876254528;
assign addr[11051]= -1145766716;
assign addr[11052]= -1392059879;
assign addr[11053]= -1610142873;
assign addr[11054]= -1795596234;
assign addr[11055]= -1944661739;
assign addr[11056]= -2054318569;
assign addr[11057]= -2122344521;
assign addr[11058]= -2147361045;
assign addr[11059]= -2128861181;
assign addr[11060]= -2067219829;
assign addr[11061]= -1963686155;
assign addr[11062]= -1820358275;
assign addr[11063]= -1640140734;
assign addr[11064]= -1426685652;
assign addr[11065]= -1184318708;
assign addr[11066]= -917951481;
assign addr[11067]= -632981917;
assign addr[11068]= -335184940;
assign addr[11069]= -30595422;
assign addr[11070]= 274614114;
assign addr[11071]= 574258580;
assign addr[11072]= 862265664;
assign addr[11073]= 1132798888;
assign addr[11074]= 1380375881;
assign addr[11075]= 1599979481;
assign addr[11076]= 1787159411;
assign addr[11077]= 1938122457;
assign addr[11078]= 2049809346;
assign addr[11079]= 2119956737;
assign addr[11080]= 2147143090;
assign addr[11081]= 2130817471;
assign addr[11082]= 2071310720;
assign addr[11083]= 1969828744;
assign addr[11084]= 1828428082;
assign addr[11085]= 1649974225;
assign addr[11086]= 1438083551;
assign addr[11087]= 1197050035;
assign addr[11088]= 931758235;
assign addr[11089]= 647584304;
assign addr[11090]= 350287041;
assign addr[11091]= 45891193;
assign addr[11092]= -259434643;
assign addr[11093]= -559503022;
assign addr[11094]= -848233042;
assign addr[11095]= -1119773573;
assign addr[11096]= -1368621831;
assign addr[11097]= -1589734894;
assign addr[11098]= -1778631892;
assign addr[11099]= -1931484818;
assign addr[11100]= -2045196100;
assign addr[11101]= -2117461370;
assign addr[11102]= -2146816171;
assign addr[11103]= -2132665626;
assign addr[11104]= -2075296495;
assign addr[11105]= -1975871368;
assign addr[11106]= -1836405100;
assign addr[11107]= -1659723983;
assign addr[11108]= -1449408469;
assign addr[11109]= -1209720613;
assign addr[11110]= -945517704;
assign addr[11111]= -662153826;
assign addr[11112]= -365371365;
assign addr[11113]= -61184634;
assign addr[11114]= 244242007;
assign addr[11115]= 544719071;
assign addr[11116]= 834157373;
assign addr[11117]= 1106691431;
assign addr[11118]= 1356798326;
assign addr[11119]= 1579409630;
assign addr[11120]= 1770014111;
assign addr[11121]= 1924749160;
assign addr[11122]= 2040479063;
assign addr[11123]= 2114858546;
assign addr[11124]= 2146380306;
assign addr[11125]= 2134405552;
assign addr[11126]= 2079176953;
assign addr[11127]= 1981813720;
assign addr[11128]= 1844288924;
assign addr[11129]= 1669389513;
assign addr[11130]= 1460659832;
assign addr[11131]= 1222329801;
assign addr[11132]= 959229189;
assign addr[11133]= 676689746;
assign addr[11134]= 380437148;
assign addr[11135]= 76474970;
assign addr[11136]= -229036977;
assign addr[11137]= -529907477;
assign addr[11138]= -820039373;
assign addr[11139]= -1093553126;
assign addr[11140]= -1344905966;
assign addr[11141]= -1569004214;
assign addr[11142]= -1761306505;
assign addr[11143]= -1917915825;
assign addr[11144]= -2035658475;
assign addr[11145]= -2112148396;
assign addr[11146]= -2145835515;
assign addr[11147]= -2136037160;
assign addr[11148]= -2082951896;
assign addr[11149]= -1987655498;
assign addr[11150]= -1852079154;
assign addr[11151]= -1678970324;
assign addr[11152]= -1471837070;
assign addr[11153]= -1234876957;
assign addr[11154]= -972891995;
assign addr[11155]= -691191324;
assign addr[11156]= -395483624;
assign addr[11157]= -91761426;
assign addr[11158]= 213820322;
assign addr[11159]= 515068990;
assign addr[11160]= 805879757;
assign addr[11161]= 1080359326;
assign addr[11162]= 1332945355;
assign addr[11163]= 1558519173;
assign addr[11164]= 1752509516;
assign addr[11165]= 1910985158;
assign addr[11166]= 2030734582;
assign addr[11167]= 2109331059;
assign addr[11168]= 2145181827;
assign addr[11169]= 2137560369;
assign addr[11170]= 2086621133;
assign addr[11171]= 1993396407;
assign addr[11172]= 1859775393;
assign addr[11173]= 1688465931;
assign addr[11174]= 1482939614;
assign addr[11175]= 1247361445;
assign addr[11176]= 986505429;
assign addr[11177]= 705657826;
assign addr[11178]= 410510029;
assign addr[11179]= 107043224;
assign addr[11180]= -198592817;
assign addr[11181]= -500204365;
assign addr[11182]= -791679244;
assign addr[11183]= -1067110699;
assign addr[11184]= -1320917099;
assign addr[11185]= -1547955041;
assign addr[11186]= -1743623590;
assign addr[11187]= -1903957513;
assign addr[11188]= -2025707632;
assign addr[11189]= -2106406677;
assign addr[11190]= -2144419275;
assign addr[11191]= -2138975100;
assign addr[11192]= -2090184478;
assign addr[11193]= -1999036154;
assign addr[11194]= -1867377253;
assign addr[11195]= -1697875851;
assign addr[11196]= -1493966902;
assign addr[11197]= -1259782632;
assign addr[11198]= -1000068799;
assign addr[11199]= -720088517;
assign addr[11200]= -425515602;
assign addr[11201]= -122319591;
assign addr[11202]= 183355234;
assign addr[11203]= 485314355;
assign addr[11204]= 777438554;
assign addr[11205]= 1053807919;
assign addr[11206]= 1308821808;
assign addr[11207]= 1537312353;
assign addr[11208]= 1734649179;
assign addr[11209]= 1896833245;
assign addr[11210]= 2020577882;
assign addr[11211]= 2103375398;
assign addr[11212]= 2143547897;
assign addr[11213]= 2140281282;
assign addr[11214]= 2093641749;
assign addr[11215]= 2004574453;
assign addr[11216]= 1874884346;
assign addr[11217]= 1707199606;
assign addr[11218]= 1504918373;
assign addr[11219]= 1272139887;
assign addr[11220]= 1013581418;
assign addr[11221]= 734482665;
assign addr[11222]= 440499581;
assign addr[11223]= 137589750;
assign addr[11224]= -168108346;
assign addr[11225]= -470399716;
assign addr[11226]= -763158411;
assign addr[11227]= -1040451659;
assign addr[11228]= -1296660098;
assign addr[11229]= -1526591649;
assign addr[11230]= -1725586737;
assign addr[11231]= -1889612716;
assign addr[11232]= -2015345591;
assign addr[11233]= -2100237377;
assign addr[11234]= -2142567738;
assign addr[11235]= -2141478848;
assign addr[11236]= -2096992772;
assign addr[11237]= -2010011024;
assign addr[11238]= -1882296293;
assign addr[11239]= -1716436725;
assign addr[11240]= -1515793473;
assign addr[11241]= -1284432584;
assign addr[11242]= -1027042599;
assign addr[11243]= -748839539;
assign addr[11244]= -455461206;
assign addr[11245]= -152852926;
assign addr[11246]= 152852926;
assign addr[11247]= 455461206;
assign addr[11248]= 748839539;
assign addr[11249]= 1027042599;
assign addr[11250]= 1284432584;
assign addr[11251]= 1515793473;
assign addr[11252]= 1716436725;
assign addr[11253]= 1882296293;
assign addr[11254]= 2010011024;
assign addr[11255]= 2096992772;
assign addr[11256]= 2141478848;
assign addr[11257]= 2142567738;
assign addr[11258]= 2100237377;
assign addr[11259]= 2015345591;
assign addr[11260]= 1889612716;
assign addr[11261]= 1725586737;
assign addr[11262]= 1526591649;
assign addr[11263]= 1296660098;
assign addr[11264]= 1040451659;
assign addr[11265]= 763158411;
assign addr[11266]= 470399716;
assign addr[11267]= 168108346;
assign addr[11268]= -137589750;
assign addr[11269]= -440499581;
assign addr[11270]= -734482665;
assign addr[11271]= -1013581418;
assign addr[11272]= -1272139887;
assign addr[11273]= -1504918373;
assign addr[11274]= -1707199606;
assign addr[11275]= -1874884346;
assign addr[11276]= -2004574453;
assign addr[11277]= -2093641749;
assign addr[11278]= -2140281282;
assign addr[11279]= -2143547897;
assign addr[11280]= -2103375398;
assign addr[11281]= -2020577882;
assign addr[11282]= -1896833245;
assign addr[11283]= -1734649179;
assign addr[11284]= -1537312353;
assign addr[11285]= -1308821808;
assign addr[11286]= -1053807919;
assign addr[11287]= -777438554;
assign addr[11288]= -485314355;
assign addr[11289]= -183355234;
assign addr[11290]= 122319591;
assign addr[11291]= 425515602;
assign addr[11292]= 720088517;
assign addr[11293]= 1000068799;
assign addr[11294]= 1259782632;
assign addr[11295]= 1493966902;
assign addr[11296]= 1697875851;
assign addr[11297]= 1867377253;
assign addr[11298]= 1999036154;
assign addr[11299]= 2090184478;
assign addr[11300]= 2138975100;
assign addr[11301]= 2144419275;
assign addr[11302]= 2106406677;
assign addr[11303]= 2025707632;
assign addr[11304]= 1903957513;
assign addr[11305]= 1743623590;
assign addr[11306]= 1547955041;
assign addr[11307]= 1320917099;
assign addr[11308]= 1067110699;
assign addr[11309]= 791679244;
assign addr[11310]= 500204365;
assign addr[11311]= 198592817;
assign addr[11312]= -107043224;
assign addr[11313]= -410510029;
assign addr[11314]= -705657826;
assign addr[11315]= -986505429;
assign addr[11316]= -1247361445;
assign addr[11317]= -1482939614;
assign addr[11318]= -1688465931;
assign addr[11319]= -1859775393;
assign addr[11320]= -1993396407;
assign addr[11321]= -2086621133;
assign addr[11322]= -2137560369;
assign addr[11323]= -2145181827;
assign addr[11324]= -2109331059;
assign addr[11325]= -2030734582;
assign addr[11326]= -1910985158;
assign addr[11327]= -1752509516;
assign addr[11328]= -1558519173;
assign addr[11329]= -1332945355;
assign addr[11330]= -1080359326;
assign addr[11331]= -805879757;
assign addr[11332]= -515068990;
assign addr[11333]= -213820322;
assign addr[11334]= 91761426;
assign addr[11335]= 395483624;
assign addr[11336]= 691191324;
assign addr[11337]= 972891995;
assign addr[11338]= 1234876957;
assign addr[11339]= 1471837070;
assign addr[11340]= 1678970324;
assign addr[11341]= 1852079154;
assign addr[11342]= 1987655498;
assign addr[11343]= 2082951896;
assign addr[11344]= 2136037160;
assign addr[11345]= 2145835515;
assign addr[11346]= 2112148396;
assign addr[11347]= 2035658475;
assign addr[11348]= 1917915825;
assign addr[11349]= 1761306505;
assign addr[11350]= 1569004214;
assign addr[11351]= 1344905966;
assign addr[11352]= 1093553126;
assign addr[11353]= 820039373;
assign addr[11354]= 529907477;
assign addr[11355]= 229036977;
assign addr[11356]= -76474970;
assign addr[11357]= -380437148;
assign addr[11358]= -676689746;
assign addr[11359]= -959229189;
assign addr[11360]= -1222329801;
assign addr[11361]= -1460659832;
assign addr[11362]= -1669389513;
assign addr[11363]= -1844288924;
assign addr[11364]= -1981813720;
assign addr[11365]= -2079176953;
assign addr[11366]= -2134405552;
assign addr[11367]= -2146380306;
assign addr[11368]= -2114858546;
assign addr[11369]= -2040479063;
assign addr[11370]= -1924749160;
assign addr[11371]= -1770014111;
assign addr[11372]= -1579409630;
assign addr[11373]= -1356798326;
assign addr[11374]= -1106691431;
assign addr[11375]= -834157373;
assign addr[11376]= -544719071;
assign addr[11377]= -244242007;
assign addr[11378]= 61184634;
assign addr[11379]= 365371365;
assign addr[11380]= 662153826;
assign addr[11381]= 945517704;
assign addr[11382]= 1209720613;
assign addr[11383]= 1449408469;
assign addr[11384]= 1659723983;
assign addr[11385]= 1836405100;
assign addr[11386]= 1975871368;
assign addr[11387]= 2075296495;
assign addr[11388]= 2132665626;
assign addr[11389]= 2146816171;
assign addr[11390]= 2117461370;
assign addr[11391]= 2045196100;
assign addr[11392]= 1931484818;
assign addr[11393]= 1778631892;
assign addr[11394]= 1589734894;
assign addr[11395]= 1368621831;
assign addr[11396]= 1119773573;
assign addr[11397]= 848233042;
assign addr[11398]= 559503022;
assign addr[11399]= 259434643;
assign addr[11400]= -45891193;
assign addr[11401]= -350287041;
assign addr[11402]= -647584304;
assign addr[11403]= -931758235;
assign addr[11404]= -1197050035;
assign addr[11405]= -1438083551;
assign addr[11406]= -1649974225;
assign addr[11407]= -1828428082;
assign addr[11408]= -1969828744;
assign addr[11409]= -2071310720;
assign addr[11410]= -2130817471;
assign addr[11411]= -2147143090;
assign addr[11412]= -2119956737;
assign addr[11413]= -2049809346;
assign addr[11414]= -1938122457;
assign addr[11415]= -1787159411;
assign addr[11416]= -1599979481;
assign addr[11417]= -1380375881;
assign addr[11418]= -1132798888;
assign addr[11419]= -862265664;
assign addr[11420]= -574258580;
assign addr[11421]= -274614114;
assign addr[11422]= 30595422;
assign addr[11423]= 335184940;
assign addr[11424]= 632981917;
assign addr[11425]= 917951481;
assign addr[11426]= 1184318708;
assign addr[11427]= 1426685652;
assign addr[11428]= 1640140734;
assign addr[11429]= 1820358275;
assign addr[11430]= 1963686155;
assign addr[11431]= 2067219829;
assign addr[11432]= 2128861181;
assign addr[11433]= 2147361045;
assign addr[11434]= 2122344521;
assign addr[11435]= 2054318569;
assign addr[11436]= 1944661739;
assign addr[11437]= 1795596234;
assign addr[11438]= 1610142873;
assign addr[11439]= 1392059879;
assign addr[11440]= 1145766716;
assign addr[11441]= 876254528;
assign addr[11442]= 588984994;
assign addr[11443]= 289779648;
assign addr[11444]= -15298099;
assign addr[11445]= -320065829;
assign addr[11446]= -618347408;
assign addr[11447]= -904098143;
assign addr[11448]= -1171527280;
assign addr[11449]= -1415215352;
assign addr[11450]= -1630224009;
assign addr[11451]= -1812196087;
assign addr[11452]= -1957443913;
assign addr[11453]= -2063024031;
assign addr[11454]= -2126796855;
assign addr[11455]= -2147470025;
assign addr[11456]= -2124624598;
assign addr[11457]= -2058723538;
assign addr[11458]= -1951102334;
assign addr[11459]= -1803941934;
assign addr[11460]= -1620224553;
assign addr[11461]= -1403673233;
assign addr[11462]= -1158676398;
assign addr[11463]= -890198924;
assign addr[11464]= -603681519;
assign addr[11465]= -304930476;
assign addr[11466]= 0;
assign addr[11467]= 304930476;
assign addr[11468]= 603681519;
assign addr[11469]= 890198924;
assign addr[11470]= 1158676398;
assign addr[11471]= 1403673233;
assign addr[11472]= 1620224553;
assign addr[11473]= 1803941934;
assign addr[11474]= 1951102334;
assign addr[11475]= 2058723538;
assign addr[11476]= 2124624598;
assign addr[11477]= 2147470025;
assign addr[11478]= 2126796855;
assign addr[11479]= 2063024031;
assign addr[11480]= 1957443913;
assign addr[11481]= 1812196087;
assign addr[11482]= 1630224009;
assign addr[11483]= 1415215352;
assign addr[11484]= 1171527280;
assign addr[11485]= 904098143;
assign addr[11486]= 618347408;
assign addr[11487]= 320065829;
assign addr[11488]= 15298099;
assign addr[11489]= -289779648;
assign addr[11490]= -588984994;
assign addr[11491]= -876254528;
assign addr[11492]= -1145766716;
assign addr[11493]= -1392059879;
assign addr[11494]= -1610142873;
assign addr[11495]= -1795596234;
assign addr[11496]= -1944661739;
assign addr[11497]= -2054318569;
assign addr[11498]= -2122344521;
assign addr[11499]= -2147361045;
assign addr[11500]= -2128861181;
assign addr[11501]= -2067219829;
assign addr[11502]= -1963686155;
assign addr[11503]= -1820358275;
assign addr[11504]= -1640140734;
assign addr[11505]= -1426685652;
assign addr[11506]= -1184318708;
assign addr[11507]= -917951481;
assign addr[11508]= -632981917;
assign addr[11509]= -335184940;
assign addr[11510]= -30595422;
assign addr[11511]= 274614114;
assign addr[11512]= 574258580;
assign addr[11513]= 862265664;
assign addr[11514]= 1132798888;
assign addr[11515]= 1380375881;
assign addr[11516]= 1599979481;
assign addr[11517]= 1787159411;
assign addr[11518]= 1938122457;
assign addr[11519]= 2049809346;
assign addr[11520]= 2119956737;
assign addr[11521]= 2147143090;
assign addr[11522]= 2130817471;
assign addr[11523]= 2071310720;
assign addr[11524]= 1969828744;
assign addr[11525]= 1828428082;
assign addr[11526]= 1649974225;
assign addr[11527]= 1438083551;
assign addr[11528]= 1197050035;
assign addr[11529]= 931758235;
assign addr[11530]= 647584304;
assign addr[11531]= 350287041;
assign addr[11532]= 45891193;
assign addr[11533]= -259434643;
assign addr[11534]= -559503022;
assign addr[11535]= -848233042;
assign addr[11536]= -1119773573;
assign addr[11537]= -1368621831;
assign addr[11538]= -1589734894;
assign addr[11539]= -1778631892;
assign addr[11540]= -1931484818;
assign addr[11541]= -2045196100;
assign addr[11542]= -2117461370;
assign addr[11543]= -2146816171;
assign addr[11544]= -2132665626;
assign addr[11545]= -2075296495;
assign addr[11546]= -1975871368;
assign addr[11547]= -1836405100;
assign addr[11548]= -1659723983;
assign addr[11549]= -1449408469;
assign addr[11550]= -1209720613;
assign addr[11551]= -945517704;
assign addr[11552]= -662153826;
assign addr[11553]= -365371365;
assign addr[11554]= -61184634;
assign addr[11555]= 244242007;
assign addr[11556]= 544719071;
assign addr[11557]= 834157373;
assign addr[11558]= 1106691431;
assign addr[11559]= 1356798326;
assign addr[11560]= 1579409630;
assign addr[11561]= 1770014111;
assign addr[11562]= 1924749160;
assign addr[11563]= 2040479063;
assign addr[11564]= 2114858546;
assign addr[11565]= 2146380306;
assign addr[11566]= 2134405552;
assign addr[11567]= 2079176953;
assign addr[11568]= 1981813720;
assign addr[11569]= 1844288924;
assign addr[11570]= 1669389513;
assign addr[11571]= 1460659832;
assign addr[11572]= 1222329801;
assign addr[11573]= 959229189;
assign addr[11574]= 676689746;
assign addr[11575]= 380437148;
assign addr[11576]= 76474970;
assign addr[11577]= -229036977;
assign addr[11578]= -529907477;
assign addr[11579]= -820039373;
assign addr[11580]= -1093553126;
assign addr[11581]= -1344905966;
assign addr[11582]= -1569004214;
assign addr[11583]= -1761306505;
assign addr[11584]= -1917915825;
assign addr[11585]= -2035658475;
assign addr[11586]= -2112148396;
assign addr[11587]= -2145835515;
assign addr[11588]= -2136037160;
assign addr[11589]= -2082951896;
assign addr[11590]= -1987655498;
assign addr[11591]= -1852079154;
assign addr[11592]= -1678970324;
assign addr[11593]= -1471837070;
assign addr[11594]= -1234876957;
assign addr[11595]= -972891995;
assign addr[11596]= -691191324;
assign addr[11597]= -395483624;
assign addr[11598]= -91761426;
assign addr[11599]= 213820322;
assign addr[11600]= 515068990;
assign addr[11601]= 805879757;
assign addr[11602]= 1080359326;
assign addr[11603]= 1332945355;
assign addr[11604]= 1558519173;
assign addr[11605]= 1752509516;
assign addr[11606]= 1910985158;
assign addr[11607]= 2030734582;
assign addr[11608]= 2109331059;
assign addr[11609]= 2145181827;
assign addr[11610]= 2137560369;
assign addr[11611]= 2086621133;
assign addr[11612]= 1993396407;
assign addr[11613]= 1859775393;
assign addr[11614]= 1688465931;
assign addr[11615]= 1482939614;
assign addr[11616]= 1247361445;
assign addr[11617]= 986505429;
assign addr[11618]= 705657826;
assign addr[11619]= 410510029;
assign addr[11620]= 107043224;
assign addr[11621]= -198592817;
assign addr[11622]= -500204365;
assign addr[11623]= -791679244;
assign addr[11624]= -1067110699;
assign addr[11625]= -1320917099;
assign addr[11626]= -1547955041;
assign addr[11627]= -1743623590;
assign addr[11628]= -1903957513;
assign addr[11629]= -2025707632;
assign addr[11630]= -2106406677;
assign addr[11631]= -2144419275;
assign addr[11632]= -2138975100;
assign addr[11633]= -2090184478;
assign addr[11634]= -1999036154;
assign addr[11635]= -1867377253;
assign addr[11636]= -1697875851;
assign addr[11637]= -1493966902;
assign addr[11638]= -1259782632;
assign addr[11639]= -1000068799;
assign addr[11640]= -720088517;
assign addr[11641]= -425515602;
assign addr[11642]= -122319591;
assign addr[11643]= 183355234;
assign addr[11644]= 485314355;
assign addr[11645]= 777438554;
assign addr[11646]= 1053807919;
assign addr[11647]= 1308821808;
assign addr[11648]= 1537312353;
assign addr[11649]= 1734649179;
assign addr[11650]= 1896833245;
assign addr[11651]= 2020577882;
assign addr[11652]= 2103375398;
assign addr[11653]= 2143547897;
assign addr[11654]= 2140281282;
assign addr[11655]= 2093641749;
assign addr[11656]= 2004574453;
assign addr[11657]= 1874884346;
assign addr[11658]= 1707199606;
assign addr[11659]= 1504918373;
assign addr[11660]= 1272139887;
assign addr[11661]= 1013581418;
assign addr[11662]= 734482665;
assign addr[11663]= 440499581;
assign addr[11664]= 137589750;
assign addr[11665]= -168108346;
assign addr[11666]= -470399716;
assign addr[11667]= -763158411;
assign addr[11668]= -1040451659;
assign addr[11669]= -1296660098;
assign addr[11670]= -1526591649;
assign addr[11671]= -1725586737;
assign addr[11672]= -1889612716;
assign addr[11673]= -2015345591;
assign addr[11674]= -2100237377;
assign addr[11675]= -2142567738;
assign addr[11676]= -2141478848;
assign addr[11677]= -2096992772;
assign addr[11678]= -2010011024;
assign addr[11679]= -1882296293;
assign addr[11680]= -1716436725;
assign addr[11681]= -1515793473;
assign addr[11682]= -1284432584;
assign addr[11683]= -1027042599;
assign addr[11684]= -748839539;
assign addr[11685]= -455461206;
assign addr[11686]= -152852926;
assign addr[11687]= 152852926;
assign addr[11688]= 455461206;
assign addr[11689]= 748839539;
assign addr[11690]= 1027042599;
assign addr[11691]= 1284432584;
assign addr[11692]= 1515793473;
assign addr[11693]= 1716436725;
assign addr[11694]= 1882296293;
assign addr[11695]= 2010011024;
assign addr[11696]= 2096992772;
assign addr[11697]= 2141478848;
assign addr[11698]= 2142567738;
assign addr[11699]= 2100237377;
assign addr[11700]= 2015345591;
assign addr[11701]= 1889612716;
assign addr[11702]= 1725586737;
assign addr[11703]= 1526591649;
assign addr[11704]= 1296660098;
assign addr[11705]= 1040451659;
assign addr[11706]= 763158411;
assign addr[11707]= 470399716;
assign addr[11708]= 168108346;
assign addr[11709]= -137589750;
assign addr[11710]= -440499581;
assign addr[11711]= -734482665;
assign addr[11712]= -1013581418;
assign addr[11713]= -1272139887;
assign addr[11714]= -1504918373;
assign addr[11715]= -1707199606;
assign addr[11716]= -1874884346;
assign addr[11717]= -2004574453;
assign addr[11718]= -2093641749;
assign addr[11719]= -2140281282;
assign addr[11720]= -2143547897;
assign addr[11721]= -2103375398;
assign addr[11722]= -2020577882;
assign addr[11723]= -1896833245;
assign addr[11724]= -1734649179;
assign addr[11725]= -1537312353;
assign addr[11726]= -1308821808;
assign addr[11727]= -1053807919;
assign addr[11728]= -777438554;
assign addr[11729]= -485314355;
assign addr[11730]= -183355234;
assign addr[11731]= 122319591;
assign addr[11732]= 425515602;
assign addr[11733]= 720088517;
assign addr[11734]= 1000068799;
assign addr[11735]= 1259782632;
assign addr[11736]= 1493966902;
assign addr[11737]= 1697875851;
assign addr[11738]= 1867377253;
assign addr[11739]= 1999036154;
assign addr[11740]= 2090184478;
assign addr[11741]= 2138975100;
assign addr[11742]= 2144419275;
assign addr[11743]= 2106406677;
assign addr[11744]= 2025707632;
assign addr[11745]= 1903957513;
assign addr[11746]= 1743623590;
assign addr[11747]= 1547955041;
assign addr[11748]= 1320917099;
assign addr[11749]= 1067110699;
assign addr[11750]= 791679244;
assign addr[11751]= 500204365;
assign addr[11752]= 198592817;
assign addr[11753]= -107043224;
assign addr[11754]= -410510029;
assign addr[11755]= -705657826;
assign addr[11756]= -986505429;
assign addr[11757]= -1247361445;
assign addr[11758]= -1482939614;
assign addr[11759]= -1688465931;
assign addr[11760]= -1859775393;
assign addr[11761]= -1993396407;
assign addr[11762]= -2086621133;
assign addr[11763]= -2137560369;
assign addr[11764]= -2145181827;
assign addr[11765]= -2109331059;
assign addr[11766]= -2030734582;
assign addr[11767]= -1910985158;
assign addr[11768]= -1752509516;
assign addr[11769]= -1558519173;
assign addr[11770]= -1332945355;
assign addr[11771]= -1080359326;
assign addr[11772]= -805879757;
assign addr[11773]= -515068990;
assign addr[11774]= -213820322;
assign addr[11775]= 91761426;
assign addr[11776]= 395483624;
assign addr[11777]= 691191324;
assign addr[11778]= 972891995;
assign addr[11779]= 1234876957;
assign addr[11780]= 1471837070;
assign addr[11781]= 1678970324;
assign addr[11782]= 1852079154;
assign addr[11783]= 1987655498;
assign addr[11784]= 2082951896;
assign addr[11785]= 2136037160;
assign addr[11786]= 2145835515;
assign addr[11787]= 2112148396;
assign addr[11788]= 2035658475;
assign addr[11789]= 1917915825;
assign addr[11790]= 1761306505;
assign addr[11791]= 1569004214;
assign addr[11792]= 1344905966;
assign addr[11793]= 1093553126;
assign addr[11794]= 820039373;
assign addr[11795]= 529907477;
assign addr[11796]= 229036977;
assign addr[11797]= -76474970;
assign addr[11798]= -380437148;
assign addr[11799]= -676689746;
assign addr[11800]= -959229189;
assign addr[11801]= -1222329801;
assign addr[11802]= -1460659832;
assign addr[11803]= -1669389513;
assign addr[11804]= -1844288924;
assign addr[11805]= -1981813720;
assign addr[11806]= -2079176953;
assign addr[11807]= -2134405552;
assign addr[11808]= -2146380306;
assign addr[11809]= -2114858546;
assign addr[11810]= -2040479063;
assign addr[11811]= -1924749160;
assign addr[11812]= -1770014111;
assign addr[11813]= -1579409630;
assign addr[11814]= -1356798326;
assign addr[11815]= -1106691431;
assign addr[11816]= -834157373;
assign addr[11817]= -544719071;
assign addr[11818]= -244242007;
assign addr[11819]= 61184634;
assign addr[11820]= 365371365;
assign addr[11821]= 662153826;
assign addr[11822]= 945517704;
assign addr[11823]= 1209720613;
assign addr[11824]= 1449408469;
assign addr[11825]= 1659723983;
assign addr[11826]= 1836405100;
assign addr[11827]= 1975871368;
assign addr[11828]= 2075296495;
assign addr[11829]= 2132665626;
assign addr[11830]= 2146816171;
assign addr[11831]= 2117461370;
assign addr[11832]= 2045196100;
assign addr[11833]= 1931484818;
assign addr[11834]= 1778631892;
assign addr[11835]= 1589734894;
assign addr[11836]= 1368621831;
assign addr[11837]= 1119773573;
assign addr[11838]= 848233042;
assign addr[11839]= 559503022;
assign addr[11840]= 259434643;
assign addr[11841]= -45891193;
assign addr[11842]= -350287041;
assign addr[11843]= -647584304;
assign addr[11844]= -931758235;
assign addr[11845]= -1197050035;
assign addr[11846]= -1438083551;
assign addr[11847]= -1649974225;
assign addr[11848]= -1828428082;
assign addr[11849]= -1969828744;
assign addr[11850]= -2071310720;
assign addr[11851]= -2130817471;
assign addr[11852]= -2147143090;
assign addr[11853]= -2119956737;
assign addr[11854]= -2049809346;
assign addr[11855]= -1938122457;
assign addr[11856]= -1787159411;
assign addr[11857]= -1599979481;
assign addr[11858]= -1380375881;
assign addr[11859]= -1132798888;
assign addr[11860]= -862265664;
assign addr[11861]= -574258580;
assign addr[11862]= -274614114;
assign addr[11863]= 30595422;
assign addr[11864]= 335184940;
assign addr[11865]= 632981917;
assign addr[11866]= 917951481;
assign addr[11867]= 1184318708;
assign addr[11868]= 1426685652;
assign addr[11869]= 1640140734;
assign addr[11870]= 1820358275;
assign addr[11871]= 1963686155;
assign addr[11872]= 2067219829;
assign addr[11873]= 2128861181;
assign addr[11874]= 2147361045;
assign addr[11875]= 2122344521;
assign addr[11876]= 2054318569;
assign addr[11877]= 1944661739;
assign addr[11878]= 1795596234;
assign addr[11879]= 1610142873;
assign addr[11880]= 1392059879;
assign addr[11881]= 1145766716;
assign addr[11882]= 876254528;
assign addr[11883]= 588984994;
assign addr[11884]= 289779648;
assign addr[11885]= -15298099;
assign addr[11886]= -320065829;
assign addr[11887]= -618347408;
assign addr[11888]= -904098143;
assign addr[11889]= -1171527280;
assign addr[11890]= -1415215352;
assign addr[11891]= -1630224009;
assign addr[11892]= -1812196087;
assign addr[11893]= -1957443913;
assign addr[11894]= -2063024031;
assign addr[11895]= -2126796855;
assign addr[11896]= -2147470025;
assign addr[11897]= -2124624598;
assign addr[11898]= -2058723538;
assign addr[11899]= -1951102334;
assign addr[11900]= -1803941934;
assign addr[11901]= -1620224553;
assign addr[11902]= -1403673233;
assign addr[11903]= -1158676398;
assign addr[11904]= -890198924;
assign addr[11905]= -603681519;
assign addr[11906]= -304930476;
assign addr[11907]= 0;
assign addr[11908]= 304930476;
assign addr[11909]= 603681519;
assign addr[11910]= 890198924;
assign addr[11911]= 1158676398;
assign addr[11912]= 1403673233;
assign addr[11913]= 1620224553;
assign addr[11914]= 1803941934;
assign addr[11915]= 1951102334;
assign addr[11916]= 2058723538;
assign addr[11917]= 2124624598;
assign addr[11918]= 2147470025;
assign addr[11919]= 2126796855;
assign addr[11920]= 2063024031;
assign addr[11921]= 1957443913;
assign addr[11922]= 1812196087;
assign addr[11923]= 1630224009;
assign addr[11924]= 1415215352;
assign addr[11925]= 1171527280;
assign addr[11926]= 904098143;
assign addr[11927]= 618347408;
assign addr[11928]= 320065829;
assign addr[11929]= 15298099;
assign addr[11930]= -289779648;
assign addr[11931]= -588984994;
assign addr[11932]= -876254528;
assign addr[11933]= -1145766716;
assign addr[11934]= -1392059879;
assign addr[11935]= -1610142873;
assign addr[11936]= -1795596234;
assign addr[11937]= -1944661739;
assign addr[11938]= -2054318569;
assign addr[11939]= -2122344521;
assign addr[11940]= -2147361045;
assign addr[11941]= -2128861181;
assign addr[11942]= -2067219829;
assign addr[11943]= -1963686155;
assign addr[11944]= -1820358275;
assign addr[11945]= -1640140734;
assign addr[11946]= -1426685652;
assign addr[11947]= -1184318708;
assign addr[11948]= -917951481;
assign addr[11949]= -632981917;
assign addr[11950]= -335184940;
assign addr[11951]= -30595422;
assign addr[11952]= 274614114;
assign addr[11953]= 574258580;
assign addr[11954]= 862265664;
assign addr[11955]= 1132798888;
assign addr[11956]= 1380375881;
assign addr[11957]= 1599979481;
assign addr[11958]= 1787159411;
assign addr[11959]= 1938122457;
assign addr[11960]= 2049809346;
assign addr[11961]= 2119956737;
assign addr[11962]= 2147143090;
assign addr[11963]= 2130817471;
assign addr[11964]= 2071310720;
assign addr[11965]= 1969828744;
assign addr[11966]= 1828428082;
assign addr[11967]= 1649974225;
assign addr[11968]= 1438083551;
assign addr[11969]= 1197050035;
assign addr[11970]= 931758235;
assign addr[11971]= 647584304;
assign addr[11972]= 350287041;
assign addr[11973]= 45891193;
assign addr[11974]= -259434643;
assign addr[11975]= -559503022;
assign addr[11976]= -848233042;
assign addr[11977]= -1119773573;
assign addr[11978]= -1368621831;
assign addr[11979]= -1589734894;
assign addr[11980]= -1778631892;
assign addr[11981]= -1931484818;
assign addr[11982]= -2045196100;
assign addr[11983]= -2117461370;
assign addr[11984]= -2146816171;
assign addr[11985]= -2132665626;
assign addr[11986]= -2075296495;
assign addr[11987]= -1975871368;
assign addr[11988]= -1836405100;
assign addr[11989]= -1659723983;
assign addr[11990]= -1449408469;
assign addr[11991]= -1209720613;
assign addr[11992]= -945517704;
assign addr[11993]= -662153826;
assign addr[11994]= -365371365;
assign addr[11995]= -61184634;
assign addr[11996]= 244242007;
assign addr[11997]= 544719071;
assign addr[11998]= 834157373;
assign addr[11999]= 1106691431;
assign addr[12000]= 1356798326;
assign addr[12001]= 1579409630;
assign addr[12002]= 1770014111;
assign addr[12003]= 1924749160;
assign addr[12004]= 2040479063;
assign addr[12005]= 2114858546;
assign addr[12006]= 2146380306;
assign addr[12007]= 2134405552;
assign addr[12008]= 2079176953;
assign addr[12009]= 1981813720;
assign addr[12010]= 1844288924;
assign addr[12011]= 1669389513;
assign addr[12012]= 1460659832;
assign addr[12013]= 1222329801;
assign addr[12014]= 959229189;
assign addr[12015]= 676689746;
assign addr[12016]= 380437148;
assign addr[12017]= 76474970;
assign addr[12018]= -229036977;
assign addr[12019]= -529907477;
assign addr[12020]= -820039373;
assign addr[12021]= -1093553126;
assign addr[12022]= -1344905966;
assign addr[12023]= -1569004214;
assign addr[12024]= -1761306505;
assign addr[12025]= -1917915825;
assign addr[12026]= -2035658475;
assign addr[12027]= -2112148396;
assign addr[12028]= -2145835515;
assign addr[12029]= -2136037160;
assign addr[12030]= -2082951896;
assign addr[12031]= -1987655498;
assign addr[12032]= -1852079154;
assign addr[12033]= -1678970324;
assign addr[12034]= -1471837070;
assign addr[12035]= -1234876957;
assign addr[12036]= -972891995;
assign addr[12037]= -691191324;
assign addr[12038]= -395483624;
assign addr[12039]= -91761426;
assign addr[12040]= 213820322;
assign addr[12041]= 515068990;
assign addr[12042]= 805879757;
assign addr[12043]= 1080359326;
assign addr[12044]= 1332945355;
assign addr[12045]= 1558519173;
assign addr[12046]= 1752509516;
assign addr[12047]= 1910985158;
assign addr[12048]= 2030734582;
assign addr[12049]= 2109331059;
assign addr[12050]= 2145181827;
assign addr[12051]= 2137560369;
assign addr[12052]= 2086621133;
assign addr[12053]= 1993396407;
assign addr[12054]= 1859775393;
assign addr[12055]= 1688465931;
assign addr[12056]= 1482939614;
assign addr[12057]= 1247361445;
assign addr[12058]= 986505429;
assign addr[12059]= 705657826;
assign addr[12060]= 410510029;
assign addr[12061]= 107043224;
assign addr[12062]= -198592817;
assign addr[12063]= -500204365;
assign addr[12064]= -791679244;
assign addr[12065]= -1067110699;
assign addr[12066]= -1320917099;
assign addr[12067]= -1547955041;
assign addr[12068]= -1743623590;
assign addr[12069]= -1903957513;
assign addr[12070]= -2025707632;
assign addr[12071]= -2106406677;
assign addr[12072]= -2144419275;
assign addr[12073]= -2138975100;
assign addr[12074]= -2090184478;
assign addr[12075]= -1999036154;
assign addr[12076]= -1867377253;
assign addr[12077]= -1697875851;
assign addr[12078]= -1493966902;
assign addr[12079]= -1259782632;
assign addr[12080]= -1000068799;
assign addr[12081]= -720088517;
assign addr[12082]= -425515602;
assign addr[12083]= -122319591;
assign addr[12084]= 183355234;
assign addr[12085]= 485314355;
assign addr[12086]= 777438554;
assign addr[12087]= 1053807919;
assign addr[12088]= 1308821808;
assign addr[12089]= 1537312353;
assign addr[12090]= 1734649179;
assign addr[12091]= 1896833245;
assign addr[12092]= 2020577882;
assign addr[12093]= 2103375398;
assign addr[12094]= 2143547897;
assign addr[12095]= 2140281282;
assign addr[12096]= 2093641749;
assign addr[12097]= 2004574453;
assign addr[12098]= 1874884346;
assign addr[12099]= 1707199606;
assign addr[12100]= 1504918373;
assign addr[12101]= 1272139887;
assign addr[12102]= 1013581418;
assign addr[12103]= 734482665;
assign addr[12104]= 440499581;
assign addr[12105]= 137589750;
assign addr[12106]= -168108346;
assign addr[12107]= -470399716;
assign addr[12108]= -763158411;
assign addr[12109]= -1040451659;
assign addr[12110]= -1296660098;
assign addr[12111]= -1526591649;
assign addr[12112]= -1725586737;
assign addr[12113]= -1889612716;
assign addr[12114]= -2015345591;
assign addr[12115]= -2100237377;
assign addr[12116]= -2142567738;
assign addr[12117]= -2141478848;
assign addr[12118]= -2096992772;
assign addr[12119]= -2010011024;
assign addr[12120]= -1882296293;
assign addr[12121]= -1716436725;
assign addr[12122]= -1515793473;
assign addr[12123]= -1284432584;
assign addr[12124]= -1027042599;
assign addr[12125]= -748839539;
assign addr[12126]= -455461206;
assign addr[12127]= -152852926;
assign addr[12128]= 152852926;
assign addr[12129]= 455461206;
assign addr[12130]= 748839539;
assign addr[12131]= 1027042599;
assign addr[12132]= 1284432584;
assign addr[12133]= 1515793473;
assign addr[12134]= 1716436725;
assign addr[12135]= 1882296293;
assign addr[12136]= 2010011024;
assign addr[12137]= 2096992772;
assign addr[12138]= 2141478848;
assign addr[12139]= 2142567738;
assign addr[12140]= 2100237377;
assign addr[12141]= 2015345591;
assign addr[12142]= 1889612716;
assign addr[12143]= 1725586737;
assign addr[12144]= 1526591649;
assign addr[12145]= 1296660098;
assign addr[12146]= 1040451659;
assign addr[12147]= 763158411;
assign addr[12148]= 470399716;
assign addr[12149]= 168108346;
assign addr[12150]= -137589750;
assign addr[12151]= -440499581;
assign addr[12152]= -734482665;
assign addr[12153]= -1013581418;
assign addr[12154]= -1272139887;
assign addr[12155]= -1504918373;
assign addr[12156]= -1707199606;
assign addr[12157]= -1874884346;
assign addr[12158]= -2004574453;
assign addr[12159]= -2093641749;
assign addr[12160]= -2140281282;
assign addr[12161]= -2143547897;
assign addr[12162]= -2103375398;
assign addr[12163]= -2020577882;
assign addr[12164]= -1896833245;
assign addr[12165]= -1734649179;
assign addr[12166]= -1537312353;
assign addr[12167]= -1308821808;
assign addr[12168]= -1053807919;
assign addr[12169]= -777438554;
assign addr[12170]= -485314355;
assign addr[12171]= -183355234;
assign addr[12172]= 122319591;
assign addr[12173]= 425515602;
assign addr[12174]= 720088517;
assign addr[12175]= 1000068799;
assign addr[12176]= 1259782632;
assign addr[12177]= 1493966902;
assign addr[12178]= 1697875851;
assign addr[12179]= 1867377253;
assign addr[12180]= 1999036154;
assign addr[12181]= 2090184478;
assign addr[12182]= 2138975100;
assign addr[12183]= 2144419275;
assign addr[12184]= 2106406677;
assign addr[12185]= 2025707632;
assign addr[12186]= 1903957513;
assign addr[12187]= 1743623590;
assign addr[12188]= 1547955041;
assign addr[12189]= 1320917099;
assign addr[12190]= 1067110699;
assign addr[12191]= 791679244;
assign addr[12192]= 500204365;
assign addr[12193]= 198592817;
assign addr[12194]= -107043224;
assign addr[12195]= -410510029;
assign addr[12196]= -705657826;
assign addr[12197]= -986505429;
assign addr[12198]= -1247361445;
assign addr[12199]= -1482939614;
assign addr[12200]= -1688465931;
assign addr[12201]= -1859775393;
assign addr[12202]= -1993396407;
assign addr[12203]= -2086621133;
assign addr[12204]= -2137560369;
assign addr[12205]= -2145181827;
assign addr[12206]= -2109331059;
assign addr[12207]= -2030734582;
assign addr[12208]= -1910985158;
assign addr[12209]= -1752509516;
assign addr[12210]= -1558519173;
assign addr[12211]= -1332945355;
assign addr[12212]= -1080359326;
assign addr[12213]= -805879757;
assign addr[12214]= -515068990;
assign addr[12215]= -213820322;
assign addr[12216]= 91761426;
assign addr[12217]= 395483624;
assign addr[12218]= 691191324;
assign addr[12219]= 972891995;
assign addr[12220]= 1234876957;
assign addr[12221]= 1471837070;
assign addr[12222]= 1678970324;
assign addr[12223]= 1852079154;
assign addr[12224]= 1987655498;
assign addr[12225]= 2082951896;
assign addr[12226]= 2136037160;
assign addr[12227]= 2145835515;
assign addr[12228]= 2112148396;
assign addr[12229]= 2035658475;
assign addr[12230]= 1917915825;
assign addr[12231]= 1761306505;
assign addr[12232]= 1569004214;
assign addr[12233]= 1344905966;
assign addr[12234]= 1093553126;
assign addr[12235]= 820039373;
assign addr[12236]= 529907477;
assign addr[12237]= 229036977;
assign addr[12238]= -76474970;
assign addr[12239]= -380437148;
assign addr[12240]= -676689746;
assign addr[12241]= -959229189;
assign addr[12242]= -1222329801;
assign addr[12243]= -1460659832;
assign addr[12244]= -1669389513;
assign addr[12245]= -1844288924;
assign addr[12246]= -1981813720;
assign addr[12247]= -2079176953;
assign addr[12248]= -2134405552;
assign addr[12249]= -2146380306;
assign addr[12250]= -2114858546;
assign addr[12251]= -2040479063;
assign addr[12252]= -1924749160;
assign addr[12253]= -1770014111;
assign addr[12254]= -1579409630;
assign addr[12255]= -1356798326;
assign addr[12256]= -1106691431;
assign addr[12257]= -834157373;
assign addr[12258]= -544719071;
assign addr[12259]= -244242007;
assign addr[12260]= 61184634;
assign addr[12261]= 365371365;
assign addr[12262]= 662153826;
assign addr[12263]= 945517704;
assign addr[12264]= 1209720613;
assign addr[12265]= 1449408469;
assign addr[12266]= 1659723983;
assign addr[12267]= 1836405100;
assign addr[12268]= 1975871368;
assign addr[12269]= 2075296495;
assign addr[12270]= 2132665626;
assign addr[12271]= 2146816171;
assign addr[12272]= 2117461370;
assign addr[12273]= 2045196100;
assign addr[12274]= 1931484818;
assign addr[12275]= 1778631892;
assign addr[12276]= 1589734894;
assign addr[12277]= 1368621831;
assign addr[12278]= 1119773573;
assign addr[12279]= 848233042;
assign addr[12280]= 559503022;
assign addr[12281]= 259434643;
assign addr[12282]= -45891193;
assign addr[12283]= -350287041;
assign addr[12284]= -647584304;
assign addr[12285]= -931758235;
assign addr[12286]= -1197050035;
assign addr[12287]= -1438083551;
assign addr[12288]= -1649974225;
assign addr[12289]= -1828428082;
assign addr[12290]= -1969828744;
assign addr[12291]= -2071310720;
assign addr[12292]= -2130817471;
assign addr[12293]= -2147143090;
assign addr[12294]= -2119956737;
assign addr[12295]= -2049809346;
assign addr[12296]= -1938122457;
assign addr[12297]= -1787159411;
assign addr[12298]= -1599979481;
assign addr[12299]= -1380375881;
assign addr[12300]= -1132798888;
assign addr[12301]= -862265664;
assign addr[12302]= -574258580;
assign addr[12303]= -274614114;
assign addr[12304]= 30595422;
assign addr[12305]= 335184940;
assign addr[12306]= 632981917;
assign addr[12307]= 917951481;
assign addr[12308]= 1184318708;
assign addr[12309]= 1426685652;
assign addr[12310]= 1640140734;
assign addr[12311]= 1820358275;
assign addr[12312]= 1963686155;
assign addr[12313]= 2067219829;
assign addr[12314]= 2128861181;
assign addr[12315]= 2147361045;
assign addr[12316]= 2122344521;
assign addr[12317]= 2054318569;
assign addr[12318]= 1944661739;
assign addr[12319]= 1795596234;
assign addr[12320]= 1610142873;
assign addr[12321]= 1392059879;
assign addr[12322]= 1145766716;
assign addr[12323]= 876254528;
assign addr[12324]= 588984994;
assign addr[12325]= 289779648;
assign addr[12326]= -15298099;
assign addr[12327]= -320065829;
assign addr[12328]= -618347408;
assign addr[12329]= -904098143;
assign addr[12330]= -1171527280;
assign addr[12331]= -1415215352;
assign addr[12332]= -1630224009;
assign addr[12333]= -1812196087;
assign addr[12334]= -1957443913;
assign addr[12335]= -2063024031;
assign addr[12336]= -2126796855;
assign addr[12337]= -2147470025;
assign addr[12338]= -2124624598;
assign addr[12339]= -2058723538;
assign addr[12340]= -1951102334;
assign addr[12341]= -1803941934;
assign addr[12342]= -1620224553;
assign addr[12343]= -1403673233;
assign addr[12344]= -1158676398;
assign addr[12345]= -890198924;
assign addr[12346]= -603681519;
assign addr[12347]= -304930476;
assign addr[12348]= 0;
assign addr[12349]= 304930476;
assign addr[12350]= 603681519;
assign addr[12351]= 890198924;
assign addr[12352]= 1158676398;
assign addr[12353]= 1403673233;
assign addr[12354]= 1620224553;
assign addr[12355]= 1803941934;
assign addr[12356]= 1951102334;
assign addr[12357]= 2058723538;
assign addr[12358]= 2124624598;
assign addr[12359]= 2147470025;
assign addr[12360]= 2126796855;
assign addr[12361]= 2063024031;
assign addr[12362]= 1957443913;
assign addr[12363]= 1812196087;
assign addr[12364]= 1630224009;
assign addr[12365]= 1415215352;
assign addr[12366]= 1171527280;
assign addr[12367]= 904098143;
assign addr[12368]= 618347408;
assign addr[12369]= 320065829;
assign addr[12370]= 15298099;
assign addr[12371]= -289779648;
assign addr[12372]= -588984994;
assign addr[12373]= -876254528;
assign addr[12374]= -1145766716;
assign addr[12375]= -1392059879;
assign addr[12376]= -1610142873;
assign addr[12377]= -1795596234;
assign addr[12378]= -1944661739;
assign addr[12379]= -2054318569;
assign addr[12380]= -2122344521;
assign addr[12381]= -2147361045;
assign addr[12382]= -2128861181;
assign addr[12383]= -2067219829;
assign addr[12384]= -1963686155;
assign addr[12385]= -1820358275;
assign addr[12386]= -1640140734;
assign addr[12387]= -1426685652;
assign addr[12388]= -1184318708;
assign addr[12389]= -917951481;
assign addr[12390]= -632981917;
assign addr[12391]= -335184940;
assign addr[12392]= -30595422;
assign addr[12393]= 274614114;
assign addr[12394]= 574258580;
assign addr[12395]= 862265664;
assign addr[12396]= 1132798888;
assign addr[12397]= 1380375881;
assign addr[12398]= 1599979481;
assign addr[12399]= 1787159411;
assign addr[12400]= 1938122457;
assign addr[12401]= 2049809346;
assign addr[12402]= 2119956737;
assign addr[12403]= 2147143090;
assign addr[12404]= 2130817471;
assign addr[12405]= 2071310720;
assign addr[12406]= 1969828744;
assign addr[12407]= 1828428082;
assign addr[12408]= 1649974225;
assign addr[12409]= 1438083551;
assign addr[12410]= 1197050035;
assign addr[12411]= 931758235;
assign addr[12412]= 647584304;
assign addr[12413]= 350287041;
assign addr[12414]= 45891193;
assign addr[12415]= -259434643;
assign addr[12416]= -559503022;
assign addr[12417]= -848233042;
assign addr[12418]= -1119773573;
assign addr[12419]= -1368621831;
assign addr[12420]= -1589734894;
assign addr[12421]= -1778631892;
assign addr[12422]= -1931484818;
assign addr[12423]= -2045196100;
assign addr[12424]= -2117461370;
assign addr[12425]= -2146816171;
assign addr[12426]= -2132665626;
assign addr[12427]= -2075296495;
assign addr[12428]= -1975871368;
assign addr[12429]= -1836405100;
assign addr[12430]= -1659723983;
assign addr[12431]= -1449408469;
assign addr[12432]= -1209720613;
assign addr[12433]= -945517704;
assign addr[12434]= -662153826;
assign addr[12435]= -365371365;
assign addr[12436]= -61184634;
assign addr[12437]= 244242007;
assign addr[12438]= 544719071;
assign addr[12439]= 834157373;
assign addr[12440]= 1106691431;
assign addr[12441]= 1356798326;
assign addr[12442]= 1579409630;
assign addr[12443]= 1770014111;
assign addr[12444]= 1924749160;
assign addr[12445]= 2040479063;
assign addr[12446]= 2114858546;
assign addr[12447]= 2146380306;
assign addr[12448]= 2134405552;
assign addr[12449]= 2079176953;
assign addr[12450]= 1981813720;
assign addr[12451]= 1844288924;
assign addr[12452]= 1669389513;
assign addr[12453]= 1460659832;
assign addr[12454]= 1222329801;
assign addr[12455]= 959229189;
assign addr[12456]= 676689746;
assign addr[12457]= 380437148;
assign addr[12458]= 76474970;
assign addr[12459]= -229036977;
assign addr[12460]= -529907477;
assign addr[12461]= -820039373;
assign addr[12462]= -1093553126;
assign addr[12463]= -1344905966;
assign addr[12464]= -1569004214;
assign addr[12465]= -1761306505;
assign addr[12466]= -1917915825;
assign addr[12467]= -2035658475;
assign addr[12468]= -2112148396;
assign addr[12469]= -2145835515;
assign addr[12470]= -2136037160;
assign addr[12471]= -2082951896;
assign addr[12472]= -1987655498;
assign addr[12473]= -1852079154;
assign addr[12474]= -1678970324;
assign addr[12475]= -1471837070;
assign addr[12476]= -1234876957;
assign addr[12477]= -972891995;
assign addr[12478]= -691191324;
assign addr[12479]= -395483624;
assign addr[12480]= -91761426;
assign addr[12481]= 213820322;
assign addr[12482]= 515068990;
assign addr[12483]= 805879757;
assign addr[12484]= 1080359326;
assign addr[12485]= 1332945355;
assign addr[12486]= 1558519173;
assign addr[12487]= 1752509516;
assign addr[12488]= 1910985158;
assign addr[12489]= 2030734582;
assign addr[12490]= 2109331059;
assign addr[12491]= 2145181827;
assign addr[12492]= 2137560369;
assign addr[12493]= 2086621133;
assign addr[12494]= 1993396407;
assign addr[12495]= 1859775393;
assign addr[12496]= 1688465931;
assign addr[12497]= 1482939614;
assign addr[12498]= 1247361445;
assign addr[12499]= 986505429;
assign addr[12500]= 705657826;
assign addr[12501]= 410510029;
assign addr[12502]= 107043224;
assign addr[12503]= -198592817;
assign addr[12504]= -500204365;
assign addr[12505]= -791679244;
assign addr[12506]= -1067110699;
assign addr[12507]= -1320917099;
assign addr[12508]= -1547955041;
assign addr[12509]= -1743623590;
assign addr[12510]= -1903957513;
assign addr[12511]= -2025707632;
assign addr[12512]= -2106406677;
assign addr[12513]= -2144419275;
assign addr[12514]= -2138975100;
assign addr[12515]= -2090184478;
assign addr[12516]= -1999036154;
assign addr[12517]= -1867377253;
assign addr[12518]= -1697875851;
assign addr[12519]= -1493966902;
assign addr[12520]= -1259782632;
assign addr[12521]= -1000068799;
assign addr[12522]= -720088517;
assign addr[12523]= -425515602;
assign addr[12524]= -122319591;
assign addr[12525]= 183355234;
assign addr[12526]= 485314355;
assign addr[12527]= 777438554;
assign addr[12528]= 1053807919;
assign addr[12529]= 1308821808;
assign addr[12530]= 1537312353;
assign addr[12531]= 1734649179;
assign addr[12532]= 1896833245;
assign addr[12533]= 2020577882;
assign addr[12534]= 2103375398;
assign addr[12535]= 2143547897;
assign addr[12536]= 2140281282;
assign addr[12537]= 2093641749;
assign addr[12538]= 2004574453;
assign addr[12539]= 1874884346;
assign addr[12540]= 1707199606;
assign addr[12541]= 1504918373;
assign addr[12542]= 1272139887;
assign addr[12543]= 1013581418;
assign addr[12544]= 734482665;
assign addr[12545]= 440499581;
assign addr[12546]= 137589750;
assign addr[12547]= -168108346;
assign addr[12548]= -470399716;
assign addr[12549]= -763158411;
assign addr[12550]= -1040451659;
assign addr[12551]= -1296660098;
assign addr[12552]= -1526591649;
assign addr[12553]= -1725586737;
assign addr[12554]= -1889612716;
assign addr[12555]= -2015345591;
assign addr[12556]= -2100237377;
assign addr[12557]= -2142567738;
assign addr[12558]= -2141478848;
assign addr[12559]= -2096992772;
assign addr[12560]= -2010011024;
assign addr[12561]= -1882296293;
assign addr[12562]= -1716436725;
assign addr[12563]= -1515793473;
assign addr[12564]= -1284432584;
assign addr[12565]= -1027042599;
assign addr[12566]= -748839539;
assign addr[12567]= -455461206;
assign addr[12568]= -152852926;
assign addr[12569]= 152852926;
assign addr[12570]= 455461206;
assign addr[12571]= 748839539;
assign addr[12572]= 1027042599;
assign addr[12573]= 1284432584;
assign addr[12574]= 1515793473;
assign addr[12575]= 1716436725;
assign addr[12576]= 1882296293;
assign addr[12577]= 2010011024;
assign addr[12578]= 2096992772;
assign addr[12579]= 2141478848;
assign addr[12580]= 2142567738;
assign addr[12581]= 2100237377;
assign addr[12582]= 2015345591;
assign addr[12583]= 1889612716;
assign addr[12584]= 1725586737;
assign addr[12585]= 1526591649;
assign addr[12586]= 1296660098;
assign addr[12587]= 1040451659;
assign addr[12588]= 763158411;
assign addr[12589]= 470399716;
assign addr[12590]= 168108346;
assign addr[12591]= -137589750;
assign addr[12592]= -440499581;
assign addr[12593]= -734482665;
assign addr[12594]= -1013581418;
assign addr[12595]= -1272139887;
assign addr[12596]= -1504918373;
assign addr[12597]= -1707199606;
assign addr[12598]= -1874884346;
assign addr[12599]= -2004574453;
assign addr[12600]= -2093641749;
assign addr[12601]= -2140281282;
assign addr[12602]= -2143547897;
assign addr[12603]= -2103375398;
assign addr[12604]= -2020577882;
assign addr[12605]= -1896833245;
assign addr[12606]= -1734649179;
assign addr[12607]= -1537312353;
assign addr[12608]= -1308821808;
assign addr[12609]= -1053807919;
assign addr[12610]= -777438554;
assign addr[12611]= -485314355;
assign addr[12612]= -183355234;
assign addr[12613]= 122319591;
assign addr[12614]= 425515602;
assign addr[12615]= 720088517;
assign addr[12616]= 1000068799;
assign addr[12617]= 1259782632;
assign addr[12618]= 1493966902;
assign addr[12619]= 1697875851;
assign addr[12620]= 1867377253;
assign addr[12621]= 1999036154;
assign addr[12622]= 2090184478;
assign addr[12623]= 2138975100;
assign addr[12624]= 2144419275;
assign addr[12625]= 2106406677;
assign addr[12626]= 2025707632;
assign addr[12627]= 1903957513;
assign addr[12628]= 1743623590;
assign addr[12629]= 1547955041;
assign addr[12630]= 1320917099;
assign addr[12631]= 1067110699;
assign addr[12632]= 791679244;
assign addr[12633]= 500204365;
assign addr[12634]= 198592817;
assign addr[12635]= -107043224;
assign addr[12636]= -410510029;
assign addr[12637]= -705657826;
assign addr[12638]= -986505429;
assign addr[12639]= -1247361445;
assign addr[12640]= -1482939614;
assign addr[12641]= -1688465931;
assign addr[12642]= -1859775393;
assign addr[12643]= -1993396407;
assign addr[12644]= -2086621133;
assign addr[12645]= -2137560369;
assign addr[12646]= -2145181827;
assign addr[12647]= -2109331059;
assign addr[12648]= -2030734582;
assign addr[12649]= -1910985158;
assign addr[12650]= -1752509516;
assign addr[12651]= -1558519173;
assign addr[12652]= -1332945355;
assign addr[12653]= -1080359326;
assign addr[12654]= -805879757;
assign addr[12655]= -515068990;
assign addr[12656]= -213820322;
assign addr[12657]= 91761426;
assign addr[12658]= 395483624;
assign addr[12659]= 691191324;
assign addr[12660]= 972891995;
assign addr[12661]= 1234876957;
assign addr[12662]= 1471837070;
assign addr[12663]= 1678970324;
assign addr[12664]= 1852079154;
assign addr[12665]= 1987655498;
assign addr[12666]= 2082951896;
assign addr[12667]= 2136037160;
assign addr[12668]= 2145835515;
assign addr[12669]= 2112148396;
assign addr[12670]= 2035658475;
assign addr[12671]= 1917915825;
assign addr[12672]= 1761306505;
assign addr[12673]= 1569004214;
assign addr[12674]= 1344905966;
assign addr[12675]= 1093553126;
assign addr[12676]= 820039373;
assign addr[12677]= 529907477;
assign addr[12678]= 229036977;
assign addr[12679]= -76474970;
assign addr[12680]= -380437148;
assign addr[12681]= -676689746;
assign addr[12682]= -959229189;
assign addr[12683]= -1222329801;
assign addr[12684]= -1460659832;
assign addr[12685]= -1669389513;
assign addr[12686]= -1844288924;
assign addr[12687]= -1981813720;
assign addr[12688]= -2079176953;
assign addr[12689]= -2134405552;
assign addr[12690]= -2146380306;
assign addr[12691]= -2114858546;
assign addr[12692]= -2040479063;
assign addr[12693]= -1924749160;
assign addr[12694]= -1770014111;
assign addr[12695]= -1579409630;
assign addr[12696]= -1356798326;
assign addr[12697]= -1106691431;
assign addr[12698]= -834157373;
assign addr[12699]= -544719071;
assign addr[12700]= -244242007;
assign addr[12701]= 61184634;
assign addr[12702]= 365371365;
assign addr[12703]= 662153826;
assign addr[12704]= 945517704;
assign addr[12705]= 1209720613;
assign addr[12706]= 1449408469;
assign addr[12707]= 1659723983;
assign addr[12708]= 1836405100;
assign addr[12709]= 1975871368;
assign addr[12710]= 2075296495;
assign addr[12711]= 2132665626;
assign addr[12712]= 2146816171;
assign addr[12713]= 2117461370;
assign addr[12714]= 2045196100;
assign addr[12715]= 1931484818;
assign addr[12716]= 1778631892;
assign addr[12717]= 1589734894;
assign addr[12718]= 1368621831;
assign addr[12719]= 1119773573;
assign addr[12720]= 848233042;
assign addr[12721]= 559503022;
assign addr[12722]= 259434643;
assign addr[12723]= -45891193;
assign addr[12724]= -350287041;
assign addr[12725]= -647584304;
assign addr[12726]= -931758235;
assign addr[12727]= -1197050035;
assign addr[12728]= -1438083551;
assign addr[12729]= -1649974225;
assign addr[12730]= -1828428082;
assign addr[12731]= -1969828744;
assign addr[12732]= -2071310720;
assign addr[12733]= -2130817471;
assign addr[12734]= -2147143090;
assign addr[12735]= -2119956737;
assign addr[12736]= -2049809346;
assign addr[12737]= -1938122457;
assign addr[12738]= -1787159411;
assign addr[12739]= -1599979481;
assign addr[12740]= -1380375881;
assign addr[12741]= -1132798888;
assign addr[12742]= -862265664;
assign addr[12743]= -574258580;
assign addr[12744]= -274614114;
assign addr[12745]= 30595422;
assign addr[12746]= 335184940;
assign addr[12747]= 632981917;
assign addr[12748]= 917951481;
assign addr[12749]= 1184318708;
assign addr[12750]= 1426685652;
assign addr[12751]= 1640140734;
assign addr[12752]= 1820358275;
assign addr[12753]= 1963686155;
assign addr[12754]= 2067219829;
assign addr[12755]= 2128861181;
assign addr[12756]= 2147361045;
assign addr[12757]= 2122344521;
assign addr[12758]= 2054318569;
assign addr[12759]= 1944661739;
assign addr[12760]= 1795596234;
assign addr[12761]= 1610142873;
assign addr[12762]= 1392059879;
assign addr[12763]= 1145766716;
assign addr[12764]= 876254528;
assign addr[12765]= 588984994;
assign addr[12766]= 289779648;
assign addr[12767]= -15298099;
assign addr[12768]= -320065829;
assign addr[12769]= -618347408;
assign addr[12770]= -904098143;
assign addr[12771]= -1171527280;
assign addr[12772]= -1415215352;
assign addr[12773]= -1630224009;
assign addr[12774]= -1812196087;
assign addr[12775]= -1957443913;
assign addr[12776]= -2063024031;
assign addr[12777]= -2126796855;
assign addr[12778]= -2147470025;
assign addr[12779]= -2124624598;
assign addr[12780]= -2058723538;
assign addr[12781]= -1951102334;
assign addr[12782]= -1803941934;
assign addr[12783]= -1620224553;
assign addr[12784]= -1403673233;
assign addr[12785]= -1158676398;
assign addr[12786]= -890198924;
assign addr[12787]= -603681519;
assign addr[12788]= -304930476;
assign addr[12789]= 0;
assign addr[12790]= 304930476;
assign addr[12791]= 603681519;
assign addr[12792]= 890198924;
assign addr[12793]= 1158676398;
assign addr[12794]= 1403673233;
assign addr[12795]= 1620224553;
assign addr[12796]= 1803941934;
assign addr[12797]= 1951102334;
assign addr[12798]= 2058723538;
assign addr[12799]= 2124624598;
assign addr[12800]= 2147470025;
assign addr[12801]= 2126796855;
assign addr[12802]= 2063024031;
assign addr[12803]= 1957443913;
assign addr[12804]= 1812196087;
assign addr[12805]= 1630224009;
assign addr[12806]= 1415215352;
assign addr[12807]= 1171527280;
assign addr[12808]= 904098143;
assign addr[12809]= 618347408;
assign addr[12810]= 320065829;
assign addr[12811]= 15298099;
assign addr[12812]= -289779648;
assign addr[12813]= -588984994;
assign addr[12814]= -876254528;
assign addr[12815]= -1145766716;
assign addr[12816]= -1392059879;
assign addr[12817]= -1610142873;
assign addr[12818]= -1795596234;
assign addr[12819]= -1944661739;
assign addr[12820]= -2054318569;
assign addr[12821]= -2122344521;
assign addr[12822]= -2147361045;
assign addr[12823]= -2128861181;
assign addr[12824]= -2067219829;
assign addr[12825]= -1963686155;
assign addr[12826]= -1820358275;
assign addr[12827]= -1640140734;
assign addr[12828]= -1426685652;
assign addr[12829]= -1184318708;
assign addr[12830]= -917951481;
assign addr[12831]= -632981917;
assign addr[12832]= -335184940;
assign addr[12833]= -30595422;
assign addr[12834]= 274614114;
assign addr[12835]= 574258580;
assign addr[12836]= 862265664;
assign addr[12837]= 1132798888;
assign addr[12838]= 1380375881;
assign addr[12839]= 1599979481;
assign addr[12840]= 1787159411;
assign addr[12841]= 1938122457;
assign addr[12842]= 2049809346;
assign addr[12843]= 2119956737;
assign addr[12844]= 2147143090;
assign addr[12845]= 2130817471;
assign addr[12846]= 2071310720;
assign addr[12847]= 1969828744;
assign addr[12848]= 1828428082;
assign addr[12849]= 1649974225;
assign addr[12850]= 1438083551;
assign addr[12851]= 1197050035;
assign addr[12852]= 931758235;
assign addr[12853]= 647584304;
assign addr[12854]= 350287041;
assign addr[12855]= 45891193;
assign addr[12856]= -259434643;
assign addr[12857]= -559503022;
assign addr[12858]= -848233042;
assign addr[12859]= -1119773573;
assign addr[12860]= -1368621831;
assign addr[12861]= -1589734894;
assign addr[12862]= -1778631892;
assign addr[12863]= -1931484818;
assign addr[12864]= -2045196100;
assign addr[12865]= -2117461370;
assign addr[12866]= -2146816171;
assign addr[12867]= -2132665626;
assign addr[12868]= -2075296495;
assign addr[12869]= -1975871368;
assign addr[12870]= -1836405100;
assign addr[12871]= -1659723983;
assign addr[12872]= -1449408469;
assign addr[12873]= -1209720613;
assign addr[12874]= -945517704;
assign addr[12875]= -662153826;
assign addr[12876]= -365371365;
assign addr[12877]= -61184634;
assign addr[12878]= 244242007;
assign addr[12879]= 544719071;
assign addr[12880]= 834157373;
assign addr[12881]= 1106691431;
assign addr[12882]= 1356798326;
assign addr[12883]= 1579409630;
assign addr[12884]= 1770014111;
assign addr[12885]= 1924749160;
assign addr[12886]= 2040479063;
assign addr[12887]= 2114858546;
assign addr[12888]= 2146380306;
assign addr[12889]= 2134405552;
assign addr[12890]= 2079176953;
assign addr[12891]= 1981813720;
assign addr[12892]= 1844288924;
assign addr[12893]= 1669389513;
assign addr[12894]= 1460659832;
assign addr[12895]= 1222329801;
assign addr[12896]= 959229189;
assign addr[12897]= 676689746;
assign addr[12898]= 380437148;
assign addr[12899]= 76474970;
assign addr[12900]= -229036977;
assign addr[12901]= -529907477;
assign addr[12902]= -820039373;
assign addr[12903]= -1093553126;
assign addr[12904]= -1344905966;
assign addr[12905]= -1569004214;
assign addr[12906]= -1761306505;
assign addr[12907]= -1917915825;
assign addr[12908]= -2035658475;
assign addr[12909]= -2112148396;
assign addr[12910]= -2145835515;
assign addr[12911]= -2136037160;
assign addr[12912]= -2082951896;
assign addr[12913]= -1987655498;
assign addr[12914]= -1852079154;
assign addr[12915]= -1678970324;
assign addr[12916]= -1471837070;
assign addr[12917]= -1234876957;
assign addr[12918]= -972891995;
assign addr[12919]= -691191324;
assign addr[12920]= -395483624;
assign addr[12921]= -91761426;
assign addr[12922]= 213820322;
assign addr[12923]= 515068990;
assign addr[12924]= 805879757;
assign addr[12925]= 1080359326;
assign addr[12926]= 1332945355;
assign addr[12927]= 1558519173;
assign addr[12928]= 1752509516;
assign addr[12929]= 1910985158;
assign addr[12930]= 2030734582;
assign addr[12931]= 2109331059;
assign addr[12932]= 2145181827;
assign addr[12933]= 2137560369;
assign addr[12934]= 2086621133;
assign addr[12935]= 1993396407;
assign addr[12936]= 1859775393;
assign addr[12937]= 1688465931;
assign addr[12938]= 1482939614;
assign addr[12939]= 1247361445;
assign addr[12940]= 986505429;
assign addr[12941]= 705657826;
assign addr[12942]= 410510029;
assign addr[12943]= 107043224;
assign addr[12944]= -198592817;
assign addr[12945]= -500204365;
assign addr[12946]= -791679244;
assign addr[12947]= -1067110699;
assign addr[12948]= -1320917099;
assign addr[12949]= -1547955041;
assign addr[12950]= -1743623590;
assign addr[12951]= -1903957513;
assign addr[12952]= -2025707632;
assign addr[12953]= -2106406677;
assign addr[12954]= -2144419275;
assign addr[12955]= -2138975100;
assign addr[12956]= -2090184478;
assign addr[12957]= -1999036154;
assign addr[12958]= -1867377253;
assign addr[12959]= -1697875851;
assign addr[12960]= -1493966902;
assign addr[12961]= -1259782632;
assign addr[12962]= -1000068799;
assign addr[12963]= -720088517;
assign addr[12964]= -425515602;
assign addr[12965]= -122319591;
assign addr[12966]= 183355234;
assign addr[12967]= 485314355;
assign addr[12968]= 777438554;
assign addr[12969]= 1053807919;
assign addr[12970]= 1308821808;
assign addr[12971]= 1537312353;
assign addr[12972]= 1734649179;
assign addr[12973]= 1896833245;
assign addr[12974]= 2020577882;
assign addr[12975]= 2103375398;
assign addr[12976]= 2143547897;
assign addr[12977]= 2140281282;
assign addr[12978]= 2093641749;
assign addr[12979]= 2004574453;
assign addr[12980]= 1874884346;
assign addr[12981]= 1707199606;
assign addr[12982]= 1504918373;
assign addr[12983]= 1272139887;
assign addr[12984]= 1013581418;
assign addr[12985]= 734482665;
assign addr[12986]= 440499581;
assign addr[12987]= 137589750;
assign addr[12988]= -168108346;
assign addr[12989]= -470399716;
assign addr[12990]= -763158411;
assign addr[12991]= -1040451659;
assign addr[12992]= -1296660098;
assign addr[12993]= -1526591649;
assign addr[12994]= -1725586737;
assign addr[12995]= -1889612716;
assign addr[12996]= -2015345591;
assign addr[12997]= -2100237377;
assign addr[12998]= -2142567738;
assign addr[12999]= -2141478848;
assign addr[13000]= -2096992772;
assign addr[13001]= -2010011024;
assign addr[13002]= -1882296293;
assign addr[13003]= -1716436725;
assign addr[13004]= -1515793473;
assign addr[13005]= -1284432584;
assign addr[13006]= -1027042599;
assign addr[13007]= -748839539;
assign addr[13008]= -455461206;
assign addr[13009]= -152852926;
assign addr[13010]= 152852926;
assign addr[13011]= 455461206;
assign addr[13012]= 748839539;
assign addr[13013]= 1027042599;
assign addr[13014]= 1284432584;
assign addr[13015]= 1515793473;
assign addr[13016]= 1716436725;
assign addr[13017]= 1882296293;
assign addr[13018]= 2010011024;
assign addr[13019]= 2096992772;
assign addr[13020]= 2141478848;
assign addr[13021]= 2142567738;
assign addr[13022]= 2100237377;
assign addr[13023]= 2015345591;
assign addr[13024]= 1889612716;
assign addr[13025]= 1725586737;
assign addr[13026]= 1526591649;
assign addr[13027]= 1296660098;
assign addr[13028]= 1040451659;
assign addr[13029]= 763158411;
assign addr[13030]= 470399716;
assign addr[13031]= 168108346;
assign addr[13032]= -137589750;
assign addr[13033]= -440499581;
assign addr[13034]= -734482665;
assign addr[13035]= -1013581418;
assign addr[13036]= -1272139887;
assign addr[13037]= -1504918373;
assign addr[13038]= -1707199606;
assign addr[13039]= -1874884346;
assign addr[13040]= -2004574453;
assign addr[13041]= -2093641749;
assign addr[13042]= -2140281282;
assign addr[13043]= -2143547897;
assign addr[13044]= -2103375398;
assign addr[13045]= -2020577882;
assign addr[13046]= -1896833245;
assign addr[13047]= -1734649179;
assign addr[13048]= -1537312353;
assign addr[13049]= -1308821808;
assign addr[13050]= -1053807919;
assign addr[13051]= -777438554;
assign addr[13052]= -485314355;
assign addr[13053]= -183355234;
assign addr[13054]= 122319591;
assign addr[13055]= 425515602;
assign addr[13056]= 720088517;
assign addr[13057]= 1000068799;
assign addr[13058]= 1259782632;
assign addr[13059]= 1493966902;
assign addr[13060]= 1697875851;
assign addr[13061]= 1867377253;
assign addr[13062]= 1999036154;
assign addr[13063]= 2090184478;
assign addr[13064]= 2138975100;
assign addr[13065]= 2144419275;
assign addr[13066]= 2106406677;
assign addr[13067]= 2025707632;
assign addr[13068]= 1903957513;
assign addr[13069]= 1743623590;
assign addr[13070]= 1547955041;
assign addr[13071]= 1320917099;
assign addr[13072]= 1067110699;
assign addr[13073]= 791679244;
assign addr[13074]= 500204365;
assign addr[13075]= 198592817;
assign addr[13076]= -107043224;
assign addr[13077]= -410510029;
assign addr[13078]= -705657826;
assign addr[13079]= -986505429;
assign addr[13080]= -1247361445;
assign addr[13081]= -1482939614;
assign addr[13082]= -1688465931;
assign addr[13083]= -1859775393;
assign addr[13084]= -1993396407;
assign addr[13085]= -2086621133;
assign addr[13086]= -2137560369;
assign addr[13087]= -2145181827;
assign addr[13088]= -2109331059;
assign addr[13089]= -2030734582;
assign addr[13090]= -1910985158;
assign addr[13091]= -1752509516;
assign addr[13092]= -1558519173;
assign addr[13093]= -1332945355;
assign addr[13094]= -1080359326;
assign addr[13095]= -805879757;
assign addr[13096]= -515068990;
assign addr[13097]= -213820322;
assign addr[13098]= 91761426;
assign addr[13099]= 395483624;
assign addr[13100]= 691191324;
assign addr[13101]= 972891995;
assign addr[13102]= 1234876957;
assign addr[13103]= 1471837070;
assign addr[13104]= 1678970324;
assign addr[13105]= 1852079154;
assign addr[13106]= 1987655498;
assign addr[13107]= 2082951896;
assign addr[13108]= 2136037160;
assign addr[13109]= 2145835515;
assign addr[13110]= 2112148396;
assign addr[13111]= 2035658475;
assign addr[13112]= 1917915825;
assign addr[13113]= 1761306505;
assign addr[13114]= 1569004214;
assign addr[13115]= 1344905966;
assign addr[13116]= 1093553126;
assign addr[13117]= 820039373;
assign addr[13118]= 529907477;
assign addr[13119]= 229036977;
assign addr[13120]= -76474970;
assign addr[13121]= -380437148;
assign addr[13122]= -676689746;
assign addr[13123]= -959229189;
assign addr[13124]= -1222329801;
assign addr[13125]= -1460659832;
assign addr[13126]= -1669389513;
assign addr[13127]= -1844288924;
assign addr[13128]= -1981813720;
assign addr[13129]= -2079176953;
assign addr[13130]= -2134405552;
assign addr[13131]= -2146380306;
assign addr[13132]= -2114858546;
assign addr[13133]= -2040479063;
assign addr[13134]= -1924749160;
assign addr[13135]= -1770014111;
assign addr[13136]= -1579409630;
assign addr[13137]= -1356798326;
assign addr[13138]= -1106691431;
assign addr[13139]= -834157373;
assign addr[13140]= -544719071;
assign addr[13141]= -244242007;
assign addr[13142]= 61184634;
assign addr[13143]= 365371365;
assign addr[13144]= 662153826;
assign addr[13145]= 945517704;
assign addr[13146]= 1209720613;
assign addr[13147]= 1449408469;
assign addr[13148]= 1659723983;
assign addr[13149]= 1836405100;
assign addr[13150]= 1975871368;
assign addr[13151]= 2075296495;
assign addr[13152]= 2132665626;
assign addr[13153]= 2146816171;
assign addr[13154]= 2117461370;
assign addr[13155]= 2045196100;
assign addr[13156]= 1931484818;
assign addr[13157]= 1778631892;
assign addr[13158]= 1589734894;
assign addr[13159]= 1368621831;
assign addr[13160]= 1119773573;
assign addr[13161]= 848233042;
assign addr[13162]= 559503022;
assign addr[13163]= 259434643;
assign addr[13164]= -45891193;
assign addr[13165]= -350287041;
assign addr[13166]= -647584304;
assign addr[13167]= -931758235;
assign addr[13168]= -1197050035;
assign addr[13169]= -1438083551;
assign addr[13170]= -1649974225;
assign addr[13171]= -1828428082;
assign addr[13172]= -1969828744;
assign addr[13173]= -2071310720;
assign addr[13174]= -2130817471;
assign addr[13175]= -2147143090;
assign addr[13176]= -2119956737;
assign addr[13177]= -2049809346;
assign addr[13178]= -1938122457;
assign addr[13179]= -1787159411;
assign addr[13180]= -1599979481;
assign addr[13181]= -1380375881;
assign addr[13182]= -1132798888;
assign addr[13183]= -862265664;
assign addr[13184]= -574258580;
assign addr[13185]= -274614114;
assign addr[13186]= 30595422;
assign addr[13187]= 335184940;
assign addr[13188]= 632981917;
assign addr[13189]= 917951481;
assign addr[13190]= 1184318708;
assign addr[13191]= 1426685652;
assign addr[13192]= 1640140734;
assign addr[13193]= 1820358275;
assign addr[13194]= 1963686155;
assign addr[13195]= 2067219829;
assign addr[13196]= 2128861181;
assign addr[13197]= 2147361045;
assign addr[13198]= 2122344521;
assign addr[13199]= 2054318569;
assign addr[13200]= 1944661739;
assign addr[13201]= 1795596234;
assign addr[13202]= 1610142873;
assign addr[13203]= 1392059879;
assign addr[13204]= 1145766716;
assign addr[13205]= 876254528;
assign addr[13206]= 588984994;
assign addr[13207]= 289779648;
assign addr[13208]= -15298099;
assign addr[13209]= -320065829;
assign addr[13210]= -618347408;
assign addr[13211]= -904098143;
assign addr[13212]= -1171527280;
assign addr[13213]= -1415215352;
assign addr[13214]= -1630224009;
assign addr[13215]= -1812196087;
assign addr[13216]= -1957443913;
assign addr[13217]= -2063024031;
assign addr[13218]= -2126796855;
assign addr[13219]= -2147470025;
assign addr[13220]= -2124624598;
assign addr[13221]= -2058723538;
assign addr[13222]= -1951102334;
assign addr[13223]= -1803941934;
assign addr[13224]= -1620224553;
assign addr[13225]= -1403673233;
assign addr[13226]= -1158676398;
assign addr[13227]= -890198924;
assign addr[13228]= -603681519;
assign addr[13229]= -304930476;
assign addr[13230]= 0;
assign addr[13231]= 304930476;
assign addr[13232]= 603681519;
assign addr[13233]= 890198924;
assign addr[13234]= 1158676398;
assign addr[13235]= 1403673233;
assign addr[13236]= 1620224553;
assign addr[13237]= 1803941934;
assign addr[13238]= 1951102334;
assign addr[13239]= 2058723538;
assign addr[13240]= 2124624598;
assign addr[13241]= 2147470025;
assign addr[13242]= 2126796855;
assign addr[13243]= 2063024031;
assign addr[13244]= 1957443913;
assign addr[13245]= 1812196087;
assign addr[13246]= 1630224009;
assign addr[13247]= 1415215352;
assign addr[13248]= 1171527280;
assign addr[13249]= 904098143;
assign addr[13250]= 618347408;
assign addr[13251]= 320065829;
assign addr[13252]= 15298099;
assign addr[13253]= -289779648;
assign addr[13254]= -588984994;
assign addr[13255]= -876254528;
assign addr[13256]= -1145766716;
assign addr[13257]= -1392059879;
assign addr[13258]= -1610142873;
assign addr[13259]= -1795596234;
assign addr[13260]= -1944661739;
assign addr[13261]= -2054318569;
assign addr[13262]= -2122344521;
assign addr[13263]= -2147361045;
assign addr[13264]= -2128861181;
assign addr[13265]= -2067219829;
assign addr[13266]= -1963686155;
assign addr[13267]= -1820358275;
assign addr[13268]= -1640140734;
assign addr[13269]= -1426685652;
assign addr[13270]= -1184318708;
assign addr[13271]= -917951481;
assign addr[13272]= -632981917;
assign addr[13273]= -335184940;
assign addr[13274]= -30595422;
assign addr[13275]= 274614114;
assign addr[13276]= 574258580;
assign addr[13277]= 862265664;
assign addr[13278]= 1132798888;
assign addr[13279]= 1380375881;
assign addr[13280]= 1599979481;
assign addr[13281]= 1787159411;
assign addr[13282]= 1938122457;
assign addr[13283]= 2049809346;
assign addr[13284]= 2119956737;
assign addr[13285]= 2147143090;
assign addr[13286]= 2130817471;
assign addr[13287]= 2071310720;
assign addr[13288]= 1969828744;
assign addr[13289]= 1828428082;
assign addr[13290]= 1649974225;
assign addr[13291]= 1438083551;
assign addr[13292]= 1197050035;
assign addr[13293]= 931758235;
assign addr[13294]= 647584304;
assign addr[13295]= 350287041;
assign addr[13296]= 45891193;
assign addr[13297]= -259434643;
assign addr[13298]= -559503022;
assign addr[13299]= -848233042;
assign addr[13300]= -1119773573;
assign addr[13301]= -1368621831;
assign addr[13302]= -1589734894;
assign addr[13303]= -1778631892;
assign addr[13304]= -1931484818;
assign addr[13305]= -2045196100;
assign addr[13306]= -2117461370;
assign addr[13307]= -2146816171;
assign addr[13308]= -2132665626;
assign addr[13309]= -2075296495;
assign addr[13310]= -1975871368;
assign addr[13311]= -1836405100;
assign addr[13312]= -1659723983;
assign addr[13313]= -1449408469;
assign addr[13314]= -1209720613;
assign addr[13315]= -945517704;
assign addr[13316]= -662153826;
assign addr[13317]= -365371365;
assign addr[13318]= -61184634;
assign addr[13319]= 244242007;
assign addr[13320]= 544719071;
assign addr[13321]= 834157373;
assign addr[13322]= 1106691431;
assign addr[13323]= 1356798326;
assign addr[13324]= 1579409630;
assign addr[13325]= 1770014111;
assign addr[13326]= 1924749160;
assign addr[13327]= 2040479063;
assign addr[13328]= 2114858546;
assign addr[13329]= 2146380306;
assign addr[13330]= 2134405552;
assign addr[13331]= 2079176953;
assign addr[13332]= 1981813720;
assign addr[13333]= 1844288924;
assign addr[13334]= 1669389513;
assign addr[13335]= 1460659832;
assign addr[13336]= 1222329801;
assign addr[13337]= 959229189;
assign addr[13338]= 676689746;
assign addr[13339]= 380437148;
assign addr[13340]= 76474970;
assign addr[13341]= -229036977;
assign addr[13342]= -529907477;
assign addr[13343]= -820039373;
assign addr[13344]= -1093553126;
assign addr[13345]= -1344905966;
assign addr[13346]= -1569004214;
assign addr[13347]= -1761306505;
assign addr[13348]= -1917915825;
assign addr[13349]= -2035658475;
assign addr[13350]= -2112148396;
assign addr[13351]= -2145835515;
assign addr[13352]= -2136037160;
assign addr[13353]= -2082951896;
assign addr[13354]= -1987655498;
assign addr[13355]= -1852079154;
assign addr[13356]= -1678970324;
assign addr[13357]= -1471837070;
assign addr[13358]= -1234876957;
assign addr[13359]= -972891995;
assign addr[13360]= -691191324;
assign addr[13361]= -395483624;
assign addr[13362]= -91761426;
assign addr[13363]= 213820322;
assign addr[13364]= 515068990;
assign addr[13365]= 805879757;
assign addr[13366]= 1080359326;
assign addr[13367]= 1332945355;
assign addr[13368]= 1558519173;
assign addr[13369]= 1752509516;
assign addr[13370]= 1910985158;
assign addr[13371]= 2030734582;
assign addr[13372]= 2109331059;
assign addr[13373]= 2145181827;
assign addr[13374]= 2137560369;
assign addr[13375]= 2086621133;
assign addr[13376]= 1993396407;
assign addr[13377]= 1859775393;
assign addr[13378]= 1688465931;
assign addr[13379]= 1482939614;
assign addr[13380]= 1247361445;
assign addr[13381]= 986505429;
assign addr[13382]= 705657826;
assign addr[13383]= 410510029;
assign addr[13384]= 107043224;
assign addr[13385]= -198592817;
assign addr[13386]= -500204365;
assign addr[13387]= -791679244;
assign addr[13388]= -1067110699;
assign addr[13389]= -1320917099;
assign addr[13390]= -1547955041;
assign addr[13391]= -1743623590;
assign addr[13392]= -1903957513;
assign addr[13393]= -2025707632;
assign addr[13394]= -2106406677;
assign addr[13395]= -2144419275;
assign addr[13396]= -2138975100;
assign addr[13397]= -2090184478;
assign addr[13398]= -1999036154;
assign addr[13399]= -1867377253;
assign addr[13400]= -1697875851;
assign addr[13401]= -1493966902;
assign addr[13402]= -1259782632;
assign addr[13403]= -1000068799;
assign addr[13404]= -720088517;
assign addr[13405]= -425515602;
assign addr[13406]= -122319591;
assign addr[13407]= 183355234;
assign addr[13408]= 485314355;
assign addr[13409]= 777438554;
assign addr[13410]= 1053807919;
assign addr[13411]= 1308821808;
assign addr[13412]= 1537312353;
assign addr[13413]= 1734649179;
assign addr[13414]= 1896833245;
assign addr[13415]= 2020577882;
assign addr[13416]= 2103375398;
assign addr[13417]= 2143547897;
assign addr[13418]= 2140281282;
assign addr[13419]= 2093641749;
assign addr[13420]= 2004574453;
assign addr[13421]= 1874884346;
assign addr[13422]= 1707199606;
assign addr[13423]= 1504918373;
assign addr[13424]= 1272139887;
assign addr[13425]= 1013581418;
assign addr[13426]= 734482665;
assign addr[13427]= 440499581;
assign addr[13428]= 137589750;
assign addr[13429]= -168108346;
assign addr[13430]= -470399716;
assign addr[13431]= -763158411;
assign addr[13432]= -1040451659;
assign addr[13433]= -1296660098;
assign addr[13434]= -1526591649;
assign addr[13435]= -1725586737;
assign addr[13436]= -1889612716;
assign addr[13437]= -2015345591;
assign addr[13438]= -2100237377;
assign addr[13439]= -2142567738;
assign addr[13440]= -2141478848;
assign addr[13441]= -2096992772;
assign addr[13442]= -2010011024;
assign addr[13443]= -1882296293;
assign addr[13444]= -1716436725;
assign addr[13445]= -1515793473;
assign addr[13446]= -1284432584;
assign addr[13447]= -1027042599;
assign addr[13448]= -748839539;
assign addr[13449]= -455461206;
assign addr[13450]= -152852926;
assign addr[13451]= 152852926;
assign addr[13452]= 455461206;
assign addr[13453]= 748839539;
assign addr[13454]= 1027042599;
assign addr[13455]= 1284432584;
assign addr[13456]= 1515793473;
assign addr[13457]= 1716436725;
assign addr[13458]= 1882296293;
assign addr[13459]= 2010011024;
assign addr[13460]= 2096992772;
assign addr[13461]= 2141478848;
assign addr[13462]= 2142567738;
assign addr[13463]= 2100237377;
assign addr[13464]= 2015345591;
assign addr[13465]= 1889612716;
assign addr[13466]= 1725586737;
assign addr[13467]= 1526591649;
assign addr[13468]= 1296660098;
assign addr[13469]= 1040451659;
assign addr[13470]= 763158411;
assign addr[13471]= 470399716;
assign addr[13472]= 168108346;
assign addr[13473]= -137589750;
assign addr[13474]= -440499581;
assign addr[13475]= -734482665;
assign addr[13476]= -1013581418;
assign addr[13477]= -1272139887;
assign addr[13478]= -1504918373;
assign addr[13479]= -1707199606;
assign addr[13480]= -1874884346;
assign addr[13481]= -2004574453;
assign addr[13482]= -2093641749;
assign addr[13483]= -2140281282;
assign addr[13484]= -2143547897;
assign addr[13485]= -2103375398;
assign addr[13486]= -2020577882;
assign addr[13487]= -1896833245;
assign addr[13488]= -1734649179;
assign addr[13489]= -1537312353;
assign addr[13490]= -1308821808;
assign addr[13491]= -1053807919;
assign addr[13492]= -777438554;
assign addr[13493]= -485314355;
assign addr[13494]= -183355234;
assign addr[13495]= 122319591;
assign addr[13496]= 425515602;
assign addr[13497]= 720088517;
assign addr[13498]= 1000068799;
assign addr[13499]= 1259782632;
assign addr[13500]= 1493966902;
assign addr[13501]= 1697875851;
assign addr[13502]= 1867377253;
assign addr[13503]= 1999036154;
assign addr[13504]= 2090184478;
assign addr[13505]= 2138975100;
assign addr[13506]= 2144419275;
assign addr[13507]= 2106406677;
assign addr[13508]= 2025707632;
assign addr[13509]= 1903957513;
assign addr[13510]= 1743623590;
assign addr[13511]= 1547955041;
assign addr[13512]= 1320917099;
assign addr[13513]= 1067110699;
assign addr[13514]= 791679244;
assign addr[13515]= 500204365;
assign addr[13516]= 198592817;
assign addr[13517]= -107043224;
assign addr[13518]= -410510029;
assign addr[13519]= -705657826;
assign addr[13520]= -986505429;
assign addr[13521]= -1247361445;
assign addr[13522]= -1482939614;
assign addr[13523]= -1688465931;
assign addr[13524]= -1859775393;
assign addr[13525]= -1993396407;
assign addr[13526]= -2086621133;
assign addr[13527]= -2137560369;
assign addr[13528]= -2145181827;
assign addr[13529]= -2109331059;
assign addr[13530]= -2030734582;
assign addr[13531]= -1910985158;
assign addr[13532]= -1752509516;
assign addr[13533]= -1558519173;
assign addr[13534]= -1332945355;
assign addr[13535]= -1080359326;
assign addr[13536]= -805879757;
assign addr[13537]= -515068990;
assign addr[13538]= -213820322;
assign addr[13539]= 91761426;
assign addr[13540]= 395483624;
assign addr[13541]= 691191324;
assign addr[13542]= 972891995;
assign addr[13543]= 1234876957;
assign addr[13544]= 1471837070;
assign addr[13545]= 1678970324;
assign addr[13546]= 1852079154;
assign addr[13547]= 1987655498;
assign addr[13548]= 2082951896;
assign addr[13549]= 2136037160;
assign addr[13550]= 2145835515;
assign addr[13551]= 2112148396;
assign addr[13552]= 2035658475;
assign addr[13553]= 1917915825;
assign addr[13554]= 1761306505;
assign addr[13555]= 1569004214;
assign addr[13556]= 1344905966;
assign addr[13557]= 1093553126;
assign addr[13558]= 820039373;
assign addr[13559]= 529907477;
assign addr[13560]= 229036977;
assign addr[13561]= -76474970;
assign addr[13562]= -380437148;
assign addr[13563]= -676689746;
assign addr[13564]= -959229189;
assign addr[13565]= -1222329801;
assign addr[13566]= -1460659832;
assign addr[13567]= -1669389513;
assign addr[13568]= -1844288924;
assign addr[13569]= -1981813720;
assign addr[13570]= -2079176953;
assign addr[13571]= -2134405552;
assign addr[13572]= -2146380306;
assign addr[13573]= -2114858546;
assign addr[13574]= -2040479063;
assign addr[13575]= -1924749160;
assign addr[13576]= -1770014111;
assign addr[13577]= -1579409630;
assign addr[13578]= -1356798326;
assign addr[13579]= -1106691431;
assign addr[13580]= -834157373;
assign addr[13581]= -544719071;
assign addr[13582]= -244242007;
assign addr[13583]= 61184634;
assign addr[13584]= 365371365;
assign addr[13585]= 662153826;
assign addr[13586]= 945517704;
assign addr[13587]= 1209720613;
assign addr[13588]= 1449408469;
assign addr[13589]= 1659723983;
assign addr[13590]= 1836405100;
assign addr[13591]= 1975871368;
assign addr[13592]= 2075296495;
assign addr[13593]= 2132665626;
assign addr[13594]= 2146816171;
assign addr[13595]= 2117461370;
assign addr[13596]= 2045196100;
assign addr[13597]= 1931484818;
assign addr[13598]= 1778631892;
assign addr[13599]= 1589734894;
assign addr[13600]= 1368621831;
assign addr[13601]= 1119773573;
assign addr[13602]= 848233042;
assign addr[13603]= 559503022;
assign addr[13604]= 259434643;
assign addr[13605]= -45891193;
assign addr[13606]= -350287041;
assign addr[13607]= -647584304;
assign addr[13608]= -931758235;
assign addr[13609]= -1197050035;
assign addr[13610]= -1438083551;
assign addr[13611]= -1649974225;
assign addr[13612]= -1828428082;
assign addr[13613]= -1969828744;
assign addr[13614]= -2071310720;
assign addr[13615]= -2130817471;
assign addr[13616]= -2147143090;
assign addr[13617]= -2119956737;
assign addr[13618]= -2049809346;
assign addr[13619]= -1938122457;
assign addr[13620]= -1787159411;
assign addr[13621]= -1599979481;
assign addr[13622]= -1380375881;
assign addr[13623]= -1132798888;
assign addr[13624]= -862265664;
assign addr[13625]= -574258580;
assign addr[13626]= -274614114;
assign addr[13627]= 30595422;
assign addr[13628]= 335184940;
assign addr[13629]= 632981917;
assign addr[13630]= 917951481;
assign addr[13631]= 1184318708;
assign addr[13632]= 1426685652;
assign addr[13633]= 1640140734;
assign addr[13634]= 1820358275;
assign addr[13635]= 1963686155;
assign addr[13636]= 2067219829;
assign addr[13637]= 2128861181;
assign addr[13638]= 2147361045;
assign addr[13639]= 2122344521;
assign addr[13640]= 2054318569;
assign addr[13641]= 1944661739;
assign addr[13642]= 1795596234;
assign addr[13643]= 1610142873;
assign addr[13644]= 1392059879;
assign addr[13645]= 1145766716;
assign addr[13646]= 876254528;
assign addr[13647]= 588984994;
assign addr[13648]= 289779648;
assign addr[13649]= -15298099;
assign addr[13650]= -320065829;
assign addr[13651]= -618347408;
assign addr[13652]= -904098143;
assign addr[13653]= -1171527280;
assign addr[13654]= -1415215352;
assign addr[13655]= -1630224009;
assign addr[13656]= -1812196087;
assign addr[13657]= -1957443913;
assign addr[13658]= -2063024031;
assign addr[13659]= -2126796855;
assign addr[13660]= -2147470025;
assign addr[13661]= -2124624598;
assign addr[13662]= -2058723538;
assign addr[13663]= -1951102334;
assign addr[13664]= -1803941934;
assign addr[13665]= -1620224553;
assign addr[13666]= -1403673233;
assign addr[13667]= -1158676398;
assign addr[13668]= -890198924;
assign addr[13669]= -603681519;
assign addr[13670]= -304930476;
assign addr[13671]= 0;
assign addr[13672]= 304930476;
assign addr[13673]= 603681519;
assign addr[13674]= 890198924;
assign addr[13675]= 1158676398;
assign addr[13676]= 1403673233;
assign addr[13677]= 1620224553;
assign addr[13678]= 1803941934;
assign addr[13679]= 1951102334;
assign addr[13680]= 2058723538;
assign addr[13681]= 2124624598;
assign addr[13682]= 2147470025;
assign addr[13683]= 2126796855;
assign addr[13684]= 2063024031;
assign addr[13685]= 1957443913;
assign addr[13686]= 1812196087;
assign addr[13687]= 1630224009;
assign addr[13688]= 1415215352;
assign addr[13689]= 1171527280;
assign addr[13690]= 904098143;
assign addr[13691]= 618347408;
assign addr[13692]= 320065829;
assign addr[13693]= 15298099;
assign addr[13694]= -289779648;
assign addr[13695]= -588984994;
assign addr[13696]= -876254528;
assign addr[13697]= -1145766716;
assign addr[13698]= -1392059879;
assign addr[13699]= -1610142873;
assign addr[13700]= -1795596234;
assign addr[13701]= -1944661739;
assign addr[13702]= -2054318569;
assign addr[13703]= -2122344521;
assign addr[13704]= -2147361045;
assign addr[13705]= -2128861181;
assign addr[13706]= -2067219829;
assign addr[13707]= -1963686155;
assign addr[13708]= -1820358275;
assign addr[13709]= -1640140734;
assign addr[13710]= -1426685652;
assign addr[13711]= -1184318708;
assign addr[13712]= -917951481;
assign addr[13713]= -632981917;
assign addr[13714]= -335184940;
assign addr[13715]= -30595422;
assign addr[13716]= 274614114;
assign addr[13717]= 574258580;
assign addr[13718]= 862265664;
assign addr[13719]= 1132798888;
assign addr[13720]= 1380375881;
assign addr[13721]= 1599979481;
assign addr[13722]= 1787159411;
assign addr[13723]= 1938122457;
assign addr[13724]= 2049809346;
assign addr[13725]= 2119956737;
assign addr[13726]= 2147143090;
assign addr[13727]= 2130817471;
assign addr[13728]= 2071310720;
assign addr[13729]= 1969828744;
assign addr[13730]= 1828428082;
assign addr[13731]= 1649974225;
assign addr[13732]= 1438083551;
assign addr[13733]= 1197050035;
assign addr[13734]= 931758235;
assign addr[13735]= 647584304;
assign addr[13736]= 350287041;
assign addr[13737]= 45891193;
assign addr[13738]= -259434643;
assign addr[13739]= -559503022;
assign addr[13740]= -848233042;
assign addr[13741]= -1119773573;
assign addr[13742]= -1368621831;
assign addr[13743]= -1589734894;
assign addr[13744]= -1778631892;
assign addr[13745]= -1931484818;
assign addr[13746]= -2045196100;
assign addr[13747]= -2117461370;
assign addr[13748]= -2146816171;
assign addr[13749]= -2132665626;
assign addr[13750]= -2075296495;
assign addr[13751]= -1975871368;
assign addr[13752]= -1836405100;
assign addr[13753]= -1659723983;
assign addr[13754]= -1449408469;
assign addr[13755]= -1209720613;
assign addr[13756]= -945517704;
assign addr[13757]= -662153826;
assign addr[13758]= -365371365;
assign addr[13759]= -61184634;
assign addr[13760]= 244242007;
assign addr[13761]= 544719071;
assign addr[13762]= 834157373;
assign addr[13763]= 1106691431;
assign addr[13764]= 1356798326;
assign addr[13765]= 1579409630;
assign addr[13766]= 1770014111;
assign addr[13767]= 1924749160;
assign addr[13768]= 2040479063;
assign addr[13769]= 2114858546;
assign addr[13770]= 2146380306;
assign addr[13771]= 2134405552;
assign addr[13772]= 2079176953;
assign addr[13773]= 1981813720;
assign addr[13774]= 1844288924;
assign addr[13775]= 1669389513;
assign addr[13776]= 1460659832;
assign addr[13777]= 1222329801;
assign addr[13778]= 959229189;
assign addr[13779]= 676689746;
assign addr[13780]= 380437148;
assign addr[13781]= 76474970;
assign addr[13782]= -229036977;
assign addr[13783]= -529907477;
assign addr[13784]= -820039373;
assign addr[13785]= -1093553126;
assign addr[13786]= -1344905966;
assign addr[13787]= -1569004214;
assign addr[13788]= -1761306505;
assign addr[13789]= -1917915825;
assign addr[13790]= -2035658475;
assign addr[13791]= -2112148396;
assign addr[13792]= -2145835515;
assign addr[13793]= -2136037160;
assign addr[13794]= -2082951896;
assign addr[13795]= -1987655498;
assign addr[13796]= -1852079154;
assign addr[13797]= -1678970324;
assign addr[13798]= -1471837070;
assign addr[13799]= -1234876957;
assign addr[13800]= -972891995;
assign addr[13801]= -691191324;
assign addr[13802]= -395483624;
assign addr[13803]= -91761426;
assign addr[13804]= 213820322;
assign addr[13805]= 515068990;
assign addr[13806]= 805879757;
assign addr[13807]= 1080359326;
assign addr[13808]= 1332945355;
assign addr[13809]= 1558519173;
assign addr[13810]= 1752509516;
assign addr[13811]= 1910985158;
assign addr[13812]= 2030734582;
assign addr[13813]= 2109331059;
assign addr[13814]= 2145181827;
assign addr[13815]= 2137560369;
assign addr[13816]= 2086621133;
assign addr[13817]= 1993396407;
assign addr[13818]= 1859775393;
assign addr[13819]= 1688465931;
assign addr[13820]= 1482939614;
assign addr[13821]= 1247361445;
assign addr[13822]= 986505429;
assign addr[13823]= 705657826;
assign addr[13824]= 410510029;
assign addr[13825]= 107043224;
assign addr[13826]= -198592817;
assign addr[13827]= -500204365;
assign addr[13828]= -791679244;
assign addr[13829]= -1067110699;
assign addr[13830]= -1320917099;
assign addr[13831]= -1547955041;
assign addr[13832]= -1743623590;
assign addr[13833]= -1903957513;
assign addr[13834]= -2025707632;
assign addr[13835]= -2106406677;
assign addr[13836]= -2144419275;
assign addr[13837]= -2138975100;
assign addr[13838]= -2090184478;
assign addr[13839]= -1999036154;
assign addr[13840]= -1867377253;
assign addr[13841]= -1697875851;
assign addr[13842]= -1493966902;
assign addr[13843]= -1259782632;
assign addr[13844]= -1000068799;
assign addr[13845]= -720088517;
assign addr[13846]= -425515602;
assign addr[13847]= -122319591;
assign addr[13848]= 183355234;
assign addr[13849]= 485314355;
assign addr[13850]= 777438554;
assign addr[13851]= 1053807919;
assign addr[13852]= 1308821808;
assign addr[13853]= 1537312353;
assign addr[13854]= 1734649179;
assign addr[13855]= 1896833245;
assign addr[13856]= 2020577882;
assign addr[13857]= 2103375398;
assign addr[13858]= 2143547897;
assign addr[13859]= 2140281282;
assign addr[13860]= 2093641749;
assign addr[13861]= 2004574453;
assign addr[13862]= 1874884346;
assign addr[13863]= 1707199606;
assign addr[13864]= 1504918373;
assign addr[13865]= 1272139887;
assign addr[13866]= 1013581418;
assign addr[13867]= 734482665;
assign addr[13868]= 440499581;
assign addr[13869]= 137589750;
assign addr[13870]= -168108346;
assign addr[13871]= -470399716;
assign addr[13872]= -763158411;
assign addr[13873]= -1040451659;
assign addr[13874]= -1296660098;
assign addr[13875]= -1526591649;
assign addr[13876]= -1725586737;
assign addr[13877]= -1889612716;
assign addr[13878]= -2015345591;
assign addr[13879]= -2100237377;
assign addr[13880]= -2142567738;
assign addr[13881]= -2141478848;
assign addr[13882]= -2096992772;
assign addr[13883]= -2010011024;
assign addr[13884]= -1882296293;
assign addr[13885]= -1716436725;
assign addr[13886]= -1515793473;
assign addr[13887]= -1284432584;
assign addr[13888]= -1027042599;
assign addr[13889]= -748839539;
assign addr[13890]= -455461206;
assign addr[13891]= -152852926;
assign addr[13892]= 152852926;
assign addr[13893]= 455461206;
assign addr[13894]= 748839539;
assign addr[13895]= 1027042599;
assign addr[13896]= 1284432584;
assign addr[13897]= 1515793473;
assign addr[13898]= 1716436725;
assign addr[13899]= 1882296293;
assign addr[13900]= 2010011024;
assign addr[13901]= 2096992772;
assign addr[13902]= 2141478848;
assign addr[13903]= 2142567738;
assign addr[13904]= 2100237377;
assign addr[13905]= 2015345591;
assign addr[13906]= 1889612716;
assign addr[13907]= 1725586737;
assign addr[13908]= 1526591649;
assign addr[13909]= 1296660098;
assign addr[13910]= 1040451659;
assign addr[13911]= 763158411;
assign addr[13912]= 470399716;
assign addr[13913]= 168108346;
assign addr[13914]= -137589750;
assign addr[13915]= -440499581;
assign addr[13916]= -734482665;
assign addr[13917]= -1013581418;
assign addr[13918]= -1272139887;
assign addr[13919]= -1504918373;
assign addr[13920]= -1707199606;
assign addr[13921]= -1874884346;
assign addr[13922]= -2004574453;
assign addr[13923]= -2093641749;
assign addr[13924]= -2140281282;
assign addr[13925]= -2143547897;
assign addr[13926]= -2103375398;
assign addr[13927]= -2020577882;
assign addr[13928]= -1896833245;
assign addr[13929]= -1734649179;
assign addr[13930]= -1537312353;
assign addr[13931]= -1308821808;
assign addr[13932]= -1053807919;
assign addr[13933]= -777438554;
assign addr[13934]= -485314355;
assign addr[13935]= -183355234;
assign addr[13936]= 122319591;
assign addr[13937]= 425515602;
assign addr[13938]= 720088517;
assign addr[13939]= 1000068799;
assign addr[13940]= 1259782632;
assign addr[13941]= 1493966902;
assign addr[13942]= 1697875851;
assign addr[13943]= 1867377253;
assign addr[13944]= 1999036154;
assign addr[13945]= 2090184478;
assign addr[13946]= 2138975100;
assign addr[13947]= 2144419275;
assign addr[13948]= 2106406677;
assign addr[13949]= 2025707632;
assign addr[13950]= 1903957513;
assign addr[13951]= 1743623590;
assign addr[13952]= 1547955041;
assign addr[13953]= 1320917099;
assign addr[13954]= 1067110699;
assign addr[13955]= 791679244;
assign addr[13956]= 500204365;
assign addr[13957]= 198592817;
assign addr[13958]= -107043224;
assign addr[13959]= -410510029;
assign addr[13960]= -705657826;
assign addr[13961]= -986505429;
assign addr[13962]= -1247361445;
assign addr[13963]= -1482939614;
assign addr[13964]= -1688465931;
assign addr[13965]= -1859775393;
assign addr[13966]= -1993396407;
assign addr[13967]= -2086621133;
assign addr[13968]= -2137560369;
assign addr[13969]= -2145181827;
assign addr[13970]= -2109331059;
assign addr[13971]= -2030734582;
assign addr[13972]= -1910985158;
assign addr[13973]= -1752509516;
assign addr[13974]= -1558519173;
assign addr[13975]= -1332945355;
assign addr[13976]= -1080359326;
assign addr[13977]= -805879757;
assign addr[13978]= -515068990;
assign addr[13979]= -213820322;
assign addr[13980]= 91761426;
assign addr[13981]= 395483624;
assign addr[13982]= 691191324;
assign addr[13983]= 972891995;
assign addr[13984]= 1234876957;
assign addr[13985]= 1471837070;
assign addr[13986]= 1678970324;
assign addr[13987]= 1852079154;
assign addr[13988]= 1987655498;
assign addr[13989]= 2082951896;
assign addr[13990]= 2136037160;
assign addr[13991]= 2145835515;
assign addr[13992]= 2112148396;
assign addr[13993]= 2035658475;
assign addr[13994]= 1917915825;
assign addr[13995]= 1761306505;
assign addr[13996]= 1569004214;
assign addr[13997]= 1344905966;
assign addr[13998]= 1093553126;
assign addr[13999]= 820039373;
assign addr[14000]= 529907477;
assign addr[14001]= 229036977;
assign addr[14002]= -76474970;
assign addr[14003]= -380437148;
assign addr[14004]= -676689746;
assign addr[14005]= -959229189;
assign addr[14006]= -1222329801;
assign addr[14007]= -1460659832;
assign addr[14008]= -1669389513;
assign addr[14009]= -1844288924;
assign addr[14010]= -1981813720;
assign addr[14011]= -2079176953;
assign addr[14012]= -2134405552;
assign addr[14013]= -2146380306;
assign addr[14014]= -2114858546;
assign addr[14015]= -2040479063;
assign addr[14016]= -1924749160;
assign addr[14017]= -1770014111;
assign addr[14018]= -1579409630;
assign addr[14019]= -1356798326;
assign addr[14020]= -1106691431;
assign addr[14021]= -834157373;
assign addr[14022]= -544719071;
assign addr[14023]= -244242007;
assign addr[14024]= 61184634;
assign addr[14025]= 365371365;
assign addr[14026]= 662153826;
assign addr[14027]= 945517704;
assign addr[14028]= 1209720613;
assign addr[14029]= 1449408469;
assign addr[14030]= 1659723983;
assign addr[14031]= 1836405100;
assign addr[14032]= 1975871368;
assign addr[14033]= 2075296495;
assign addr[14034]= 2132665626;
assign addr[14035]= 2146816171;
assign addr[14036]= 2117461370;
assign addr[14037]= 2045196100;
assign addr[14038]= 1931484818;
assign addr[14039]= 1778631892;
assign addr[14040]= 1589734894;
assign addr[14041]= 1368621831;
assign addr[14042]= 1119773573;
assign addr[14043]= 848233042;
assign addr[14044]= 559503022;
assign addr[14045]= 259434643;
assign addr[14046]= -45891193;
assign addr[14047]= -350287041;
assign addr[14048]= -647584304;
assign addr[14049]= -931758235;
assign addr[14050]= -1197050035;
assign addr[14051]= -1438083551;
assign addr[14052]= -1649974225;
assign addr[14053]= -1828428082;
assign addr[14054]= -1969828744;
assign addr[14055]= -2071310720;
assign addr[14056]= -2130817471;
assign addr[14057]= -2147143090;
assign addr[14058]= -2119956737;
assign addr[14059]= -2049809346;
assign addr[14060]= -1938122457;
assign addr[14061]= -1787159411;
assign addr[14062]= -1599979481;
assign addr[14063]= -1380375881;
assign addr[14064]= -1132798888;
assign addr[14065]= -862265664;
assign addr[14066]= -574258580;
assign addr[14067]= -274614114;
assign addr[14068]= 30595422;
assign addr[14069]= 335184940;
assign addr[14070]= 632981917;
assign addr[14071]= 917951481;
assign addr[14072]= 1184318708;
assign addr[14073]= 1426685652;
assign addr[14074]= 1640140734;
assign addr[14075]= 1820358275;
assign addr[14076]= 1963686155;
assign addr[14077]= 2067219829;
assign addr[14078]= 2128861181;
assign addr[14079]= 2147361045;
assign addr[14080]= 2122344521;
assign addr[14081]= 2054318569;
assign addr[14082]= 1944661739;
assign addr[14083]= 1795596234;
assign addr[14084]= 1610142873;
assign addr[14085]= 1392059879;
assign addr[14086]= 1145766716;
assign addr[14087]= 876254528;
assign addr[14088]= 588984994;
assign addr[14089]= 289779648;
assign addr[14090]= -15298099;
assign addr[14091]= -320065829;
assign addr[14092]= -618347408;
assign addr[14093]= -904098143;
assign addr[14094]= -1171527280;
assign addr[14095]= -1415215352;
assign addr[14096]= -1630224009;
assign addr[14097]= -1812196087;
assign addr[14098]= -1957443913;
assign addr[14099]= -2063024031;
assign addr[14100]= -2126796855;
assign addr[14101]= -2147470025;
assign addr[14102]= -2124624598;
assign addr[14103]= -2058723538;
assign addr[14104]= -1951102334;
assign addr[14105]= -1803941934;
assign addr[14106]= -1620224553;
assign addr[14107]= -1403673233;
assign addr[14108]= -1158676398;
assign addr[14109]= -890198924;
assign addr[14110]= -603681519;
assign addr[14111]= -304930476;
assign addr[14112]= 0;
assign addr[14113]= 304930476;
assign addr[14114]= 603681519;
assign addr[14115]= 890198924;
assign addr[14116]= 1158676398;
assign addr[14117]= 1403673233;
assign addr[14118]= 1620224553;
assign addr[14119]= 1803941934;
assign addr[14120]= 1951102334;
assign addr[14121]= 2058723538;
assign addr[14122]= 2124624598;
assign addr[14123]= 2147470025;
assign addr[14124]= 2126796855;
assign addr[14125]= 2063024031;
assign addr[14126]= 1957443913;
assign addr[14127]= 1812196087;
assign addr[14128]= 1630224009;
assign addr[14129]= 1415215352;
assign addr[14130]= 1171527280;
assign addr[14131]= 904098143;
assign addr[14132]= 618347408;
assign addr[14133]= 320065829;
assign addr[14134]= 15298099;
assign addr[14135]= -289779648;
assign addr[14136]= -588984994;
assign addr[14137]= -876254528;
assign addr[14138]= -1145766716;
assign addr[14139]= -1392059879;
assign addr[14140]= -1610142873;
assign addr[14141]= -1795596234;
assign addr[14142]= -1944661739;
assign addr[14143]= -2054318569;
assign addr[14144]= -2122344521;
assign addr[14145]= -2147361045;
assign addr[14146]= -2128861181;
assign addr[14147]= -2067219829;
assign addr[14148]= -1963686155;
assign addr[14149]= -1820358275;
assign addr[14150]= -1640140734;
assign addr[14151]= -1426685652;
assign addr[14152]= -1184318708;
assign addr[14153]= -917951481;
assign addr[14154]= -632981917;
assign addr[14155]= -335184940;
assign addr[14156]= -30595422;
assign addr[14157]= 274614114;
assign addr[14158]= 574258580;
assign addr[14159]= 862265664;
assign addr[14160]= 1132798888;
assign addr[14161]= 1380375881;
assign addr[14162]= 1599979481;
assign addr[14163]= 1787159411;
assign addr[14164]= 1938122457;
assign addr[14165]= 2049809346;
assign addr[14166]= 2119956737;
assign addr[14167]= 2147143090;
assign addr[14168]= 2130817471;
assign addr[14169]= 2071310720;
assign addr[14170]= 1969828744;
assign addr[14171]= 1828428082;
assign addr[14172]= 1649974225;
assign addr[14173]= 1438083551;
assign addr[14174]= 1197050035;
assign addr[14175]= 931758235;
assign addr[14176]= 647584304;
assign addr[14177]= 350287041;
assign addr[14178]= 45891193;
assign addr[14179]= -259434643;
assign addr[14180]= -559503022;
assign addr[14181]= -848233042;
assign addr[14182]= -1119773573;
assign addr[14183]= -1368621831;
assign addr[14184]= -1589734894;
assign addr[14185]= -1778631892;
assign addr[14186]= -1931484818;
assign addr[14187]= -2045196100;
assign addr[14188]= -2117461370;
assign addr[14189]= -2146816171;
assign addr[14190]= -2132665626;
assign addr[14191]= -2075296495;
assign addr[14192]= -1975871368;
assign addr[14193]= -1836405100;
assign addr[14194]= -1659723983;
assign addr[14195]= -1449408469;
assign addr[14196]= -1209720613;
assign addr[14197]= -945517704;
assign addr[14198]= -662153826;
assign addr[14199]= -365371365;
assign addr[14200]= -61184634;
assign addr[14201]= 244242007;
assign addr[14202]= 544719071;
assign addr[14203]= 834157373;
assign addr[14204]= 1106691431;
assign addr[14205]= 1356798326;
assign addr[14206]= 1579409630;
assign addr[14207]= 1770014111;
assign addr[14208]= 1924749160;
assign addr[14209]= 2040479063;
assign addr[14210]= 2114858546;
assign addr[14211]= 2146380306;
assign addr[14212]= 2134405552;
assign addr[14213]= 2079176953;
assign addr[14214]= 1981813720;
assign addr[14215]= 1844288924;
assign addr[14216]= 1669389513;
assign addr[14217]= 1460659832;
assign addr[14218]= 1222329801;
assign addr[14219]= 959229189;
assign addr[14220]= 676689746;
assign addr[14221]= 380437148;
assign addr[14222]= 76474970;
assign addr[14223]= -229036977;
assign addr[14224]= -529907477;
assign addr[14225]= -820039373;
assign addr[14226]= -1093553126;
assign addr[14227]= -1344905966;
assign addr[14228]= -1569004214;
assign addr[14229]= -1761306505;
assign addr[14230]= -1917915825;
assign addr[14231]= -2035658475;
assign addr[14232]= -2112148396;
assign addr[14233]= -2145835515;
assign addr[14234]= -2136037160;
assign addr[14235]= -2082951896;
assign addr[14236]= -1987655498;
assign addr[14237]= -1852079154;
assign addr[14238]= -1678970324;
assign addr[14239]= -1471837070;
assign addr[14240]= -1234876957;
assign addr[14241]= -972891995;
assign addr[14242]= -691191324;
assign addr[14243]= -395483624;
assign addr[14244]= -91761426;
assign addr[14245]= 213820322;
assign addr[14246]= 515068990;
assign addr[14247]= 805879757;
assign addr[14248]= 1080359326;
assign addr[14249]= 1332945355;
assign addr[14250]= 1558519173;
assign addr[14251]= 1752509516;
assign addr[14252]= 1910985158;
assign addr[14253]= 2030734582;
assign addr[14254]= 2109331059;
assign addr[14255]= 2145181827;
assign addr[14256]= 2137560369;
assign addr[14257]= 2086621133;
assign addr[14258]= 1993396407;
assign addr[14259]= 1859775393;
assign addr[14260]= 1688465931;
assign addr[14261]= 1482939614;
assign addr[14262]= 1247361445;
assign addr[14263]= 986505429;
assign addr[14264]= 705657826;
assign addr[14265]= 410510029;
assign addr[14266]= 107043224;
assign addr[14267]= -198592817;
assign addr[14268]= -500204365;
assign addr[14269]= -791679244;
assign addr[14270]= -1067110699;
assign addr[14271]= -1320917099;
assign addr[14272]= -1547955041;
assign addr[14273]= -1743623590;
assign addr[14274]= -1903957513;
assign addr[14275]= -2025707632;
assign addr[14276]= -2106406677;
assign addr[14277]= -2144419275;
assign addr[14278]= -2138975100;
assign addr[14279]= -2090184478;
assign addr[14280]= -1999036154;
assign addr[14281]= -1867377253;
assign addr[14282]= -1697875851;
assign addr[14283]= -1493966902;
assign addr[14284]= -1259782632;
assign addr[14285]= -1000068799;
assign addr[14286]= -720088517;
assign addr[14287]= -425515602;
assign addr[14288]= -122319591;
assign addr[14289]= 183355234;
assign addr[14290]= 485314355;
assign addr[14291]= 777438554;
assign addr[14292]= 1053807919;
assign addr[14293]= 1308821808;
assign addr[14294]= 1537312353;
assign addr[14295]= 1734649179;
assign addr[14296]= 1896833245;
assign addr[14297]= 2020577882;
assign addr[14298]= 2103375398;
assign addr[14299]= 2143547897;
assign addr[14300]= 2140281282;
assign addr[14301]= 2093641749;
assign addr[14302]= 2004574453;
assign addr[14303]= 1874884346;
assign addr[14304]= 1707199606;
assign addr[14305]= 1504918373;
assign addr[14306]= 1272139887;
assign addr[14307]= 1013581418;
assign addr[14308]= 734482665;
assign addr[14309]= 440499581;
assign addr[14310]= 137589750;
assign addr[14311]= -168108346;
assign addr[14312]= -470399716;
assign addr[14313]= -763158411;
assign addr[14314]= -1040451659;
assign addr[14315]= -1296660098;
assign addr[14316]= -1526591649;
assign addr[14317]= -1725586737;
assign addr[14318]= -1889612716;
assign addr[14319]= -2015345591;
assign addr[14320]= -2100237377;
assign addr[14321]= -2142567738;
assign addr[14322]= -2141478848;
assign addr[14323]= -2096992772;
assign addr[14324]= -2010011024;
assign addr[14325]= -1882296293;
assign addr[14326]= -1716436725;
assign addr[14327]= -1515793473;
assign addr[14328]= -1284432584;
assign addr[14329]= -1027042599;
assign addr[14330]= -748839539;
assign addr[14331]= -455461206;
assign addr[14332]= -152852926;
assign addr[14333]= 152852926;
assign addr[14334]= 455461206;
assign addr[14335]= 748839539;
assign addr[14336]= 1027042599;
assign addr[14337]= 1284432584;
assign addr[14338]= 1515793473;
assign addr[14339]= 1716436725;
assign addr[14340]= 1882296293;
assign addr[14341]= 2010011024;
assign addr[14342]= 2096992772;
assign addr[14343]= 2141478848;
assign addr[14344]= 2142567738;
assign addr[14345]= 2100237377;
assign addr[14346]= 2015345591;
assign addr[14347]= 1889612716;
assign addr[14348]= 1725586737;
assign addr[14349]= 1526591649;
assign addr[14350]= 1296660098;
assign addr[14351]= 1040451659;
assign addr[14352]= 763158411;
assign addr[14353]= 470399716;
assign addr[14354]= 168108346;
assign addr[14355]= -137589750;
assign addr[14356]= -440499581;
assign addr[14357]= -734482665;
assign addr[14358]= -1013581418;
assign addr[14359]= -1272139887;
assign addr[14360]= -1504918373;
assign addr[14361]= -1707199606;
assign addr[14362]= -1874884346;
assign addr[14363]= -2004574453;
assign addr[14364]= -2093641749;
assign addr[14365]= -2140281282;
assign addr[14366]= -2143547897;
assign addr[14367]= -2103375398;
assign addr[14368]= -2020577882;
assign addr[14369]= -1896833245;
assign addr[14370]= -1734649179;
assign addr[14371]= -1537312353;
assign addr[14372]= -1308821808;
assign addr[14373]= -1053807919;
assign addr[14374]= -777438554;
assign addr[14375]= -485314355;
assign addr[14376]= -183355234;
assign addr[14377]= 122319591;
assign addr[14378]= 425515602;
assign addr[14379]= 720088517;
assign addr[14380]= 1000068799;
assign addr[14381]= 1259782632;
assign addr[14382]= 1493966902;
assign addr[14383]= 1697875851;
assign addr[14384]= 1867377253;
assign addr[14385]= 1999036154;
assign addr[14386]= 2090184478;
assign addr[14387]= 2138975100;
assign addr[14388]= 2144419275;
assign addr[14389]= 2106406677;
assign addr[14390]= 2025707632;
assign addr[14391]= 1903957513;
assign addr[14392]= 1743623590;
assign addr[14393]= 1547955041;
assign addr[14394]= 1320917099;
assign addr[14395]= 1067110699;
assign addr[14396]= 791679244;
assign addr[14397]= 500204365;
assign addr[14398]= 198592817;
assign addr[14399]= -107043224;
assign addr[14400]= -410510029;
assign addr[14401]= -705657826;
assign addr[14402]= -986505429;
assign addr[14403]= -1247361445;
assign addr[14404]= -1482939614;
assign addr[14405]= -1688465931;
assign addr[14406]= -1859775393;
assign addr[14407]= -1993396407;
assign addr[14408]= -2086621133;
assign addr[14409]= -2137560369;
assign addr[14410]= -2145181827;
assign addr[14411]= -2109331059;
assign addr[14412]= -2030734582;
assign addr[14413]= -1910985158;
assign addr[14414]= -1752509516;
assign addr[14415]= -1558519173;
assign addr[14416]= -1332945355;
assign addr[14417]= -1080359326;
assign addr[14418]= -805879757;
assign addr[14419]= -515068990;
assign addr[14420]= -213820322;
assign addr[14421]= 91761426;
assign addr[14422]= 395483624;
assign addr[14423]= 691191324;
assign addr[14424]= 972891995;
assign addr[14425]= 1234876957;
assign addr[14426]= 1471837070;
assign addr[14427]= 1678970324;
assign addr[14428]= 1852079154;
assign addr[14429]= 1987655498;
assign addr[14430]= 2082951896;
assign addr[14431]= 2136037160;
assign addr[14432]= 2145835515;
assign addr[14433]= 2112148396;
assign addr[14434]= 2035658475;
assign addr[14435]= 1917915825;
assign addr[14436]= 1761306505;
assign addr[14437]= 1569004214;
assign addr[14438]= 1344905966;
assign addr[14439]= 1093553126;
assign addr[14440]= 820039373;
assign addr[14441]= 529907477;
assign addr[14442]= 229036977;
assign addr[14443]= -76474970;
assign addr[14444]= -380437148;
assign addr[14445]= -676689746;
assign addr[14446]= -959229189;
assign addr[14447]= -1222329801;
assign addr[14448]= -1460659832;
assign addr[14449]= -1669389513;
assign addr[14450]= -1844288924;
assign addr[14451]= -1981813720;
assign addr[14452]= -2079176953;
assign addr[14453]= -2134405552;
assign addr[14454]= -2146380306;
assign addr[14455]= -2114858546;
assign addr[14456]= -2040479063;
assign addr[14457]= -1924749160;
assign addr[14458]= -1770014111;
assign addr[14459]= -1579409630;
assign addr[14460]= -1356798326;
assign addr[14461]= -1106691431;
assign addr[14462]= -834157373;
assign addr[14463]= -544719071;
assign addr[14464]= -244242007;
assign addr[14465]= 61184634;
assign addr[14466]= 365371365;
assign addr[14467]= 662153826;
assign addr[14468]= 945517704;
assign addr[14469]= 1209720613;
assign addr[14470]= 1449408469;
assign addr[14471]= 1659723983;
assign addr[14472]= 1836405100;
assign addr[14473]= 1975871368;
assign addr[14474]= 2075296495;
assign addr[14475]= 2132665626;
assign addr[14476]= 2146816171;
assign addr[14477]= 2117461370;
assign addr[14478]= 2045196100;
assign addr[14479]= 1931484818;
assign addr[14480]= 1778631892;
assign addr[14481]= 1589734894;
assign addr[14482]= 1368621831;
assign addr[14483]= 1119773573;
assign addr[14484]= 848233042;
assign addr[14485]= 559503022;
assign addr[14486]= 259434643;
assign addr[14487]= -45891193;
assign addr[14488]= -350287041;
assign addr[14489]= -647584304;
assign addr[14490]= -931758235;
assign addr[14491]= -1197050035;
assign addr[14492]= -1438083551;
assign addr[14493]= -1649974225;
assign addr[14494]= -1828428082;
assign addr[14495]= -1969828744;
assign addr[14496]= -2071310720;
assign addr[14497]= -2130817471;
assign addr[14498]= -2147143090;
assign addr[14499]= -2119956737;
assign addr[14500]= -2049809346;
assign addr[14501]= -1938122457;
assign addr[14502]= -1787159411;
assign addr[14503]= -1599979481;
assign addr[14504]= -1380375881;
assign addr[14505]= -1132798888;
assign addr[14506]= -862265664;
assign addr[14507]= -574258580;
assign addr[14508]= -274614114;
assign addr[14509]= 30595422;
assign addr[14510]= 335184940;
assign addr[14511]= 632981917;
assign addr[14512]= 917951481;
assign addr[14513]= 1184318708;
assign addr[14514]= 1426685652;
assign addr[14515]= 1640140734;
assign addr[14516]= 1820358275;
assign addr[14517]= 1963686155;
assign addr[14518]= 2067219829;
assign addr[14519]= 2128861181;
assign addr[14520]= 2147361045;
assign addr[14521]= 2122344521;
assign addr[14522]= 2054318569;
assign addr[14523]= 1944661739;
assign addr[14524]= 1795596234;
assign addr[14525]= 1610142873;
assign addr[14526]= 1392059879;
assign addr[14527]= 1145766716;
assign addr[14528]= 876254528;
assign addr[14529]= 588984994;
assign addr[14530]= 289779648;
assign addr[14531]= -15298099;
assign addr[14532]= -320065829;
assign addr[14533]= -618347408;
assign addr[14534]= -904098143;
assign addr[14535]= -1171527280;
assign addr[14536]= -1415215352;
assign addr[14537]= -1630224009;
assign addr[14538]= -1812196087;
assign addr[14539]= -1957443913;
assign addr[14540]= -2063024031;
assign addr[14541]= -2126796855;
assign addr[14542]= -2147470025;
assign addr[14543]= -2124624598;
assign addr[14544]= -2058723538;
assign addr[14545]= -1951102334;
assign addr[14546]= -1803941934;
assign addr[14547]= -1620224553;
assign addr[14548]= -1403673233;
assign addr[14549]= -1158676398;
assign addr[14550]= -890198924;
assign addr[14551]= -603681519;
assign addr[14552]= -304930476;
assign addr[14553]= 0;
assign addr[14554]= 304930476;
assign addr[14555]= 603681519;
assign addr[14556]= 890198924;
assign addr[14557]= 1158676398;
assign addr[14558]= 1403673233;
assign addr[14559]= 1620224553;
assign addr[14560]= 1803941934;
assign addr[14561]= 1951102334;
assign addr[14562]= 2058723538;
assign addr[14563]= 2124624598;
assign addr[14564]= 2147470025;
assign addr[14565]= 2126796855;
assign addr[14566]= 2063024031;
assign addr[14567]= 1957443913;
assign addr[14568]= 1812196087;
assign addr[14569]= 1630224009;
assign addr[14570]= 1415215352;
assign addr[14571]= 1171527280;
assign addr[14572]= 904098143;
assign addr[14573]= 618347408;
assign addr[14574]= 320065829;
assign addr[14575]= 15298099;
assign addr[14576]= -289779648;
assign addr[14577]= -588984994;
assign addr[14578]= -876254528;
assign addr[14579]= -1145766716;
assign addr[14580]= -1392059879;
assign addr[14581]= -1610142873;
assign addr[14582]= -1795596234;
assign addr[14583]= -1944661739;
assign addr[14584]= -2054318569;
assign addr[14585]= -2122344521;
assign addr[14586]= -2147361045;
assign addr[14587]= -2128861181;
assign addr[14588]= -2067219829;
assign addr[14589]= -1963686155;
assign addr[14590]= -1820358275;
assign addr[14591]= -1640140734;
assign addr[14592]= -1426685652;
assign addr[14593]= -1184318708;
assign addr[14594]= -917951481;
assign addr[14595]= -632981917;
assign addr[14596]= -335184940;
assign addr[14597]= -30595422;
assign addr[14598]= 274614114;
assign addr[14599]= 574258580;
assign addr[14600]= 862265664;
assign addr[14601]= 1132798888;
assign addr[14602]= 1380375881;
assign addr[14603]= 1599979481;
assign addr[14604]= 1787159411;
assign addr[14605]= 1938122457;
assign addr[14606]= 2049809346;
assign addr[14607]= 2119956737;
assign addr[14608]= 2147143090;
assign addr[14609]= 2130817471;
assign addr[14610]= 2071310720;
assign addr[14611]= 1969828744;
assign addr[14612]= 1828428082;
assign addr[14613]= 1649974225;
assign addr[14614]= 1438083551;
assign addr[14615]= 1197050035;
assign addr[14616]= 931758235;
assign addr[14617]= 647584304;
assign addr[14618]= 350287041;
assign addr[14619]= 45891193;
assign addr[14620]= -259434643;
assign addr[14621]= -559503022;
assign addr[14622]= -848233042;
assign addr[14623]= -1119773573;
assign addr[14624]= -1368621831;
assign addr[14625]= -1589734894;
assign addr[14626]= -1778631892;
assign addr[14627]= -1931484818;
assign addr[14628]= -2045196100;
assign addr[14629]= -2117461370;
assign addr[14630]= -2146816171;
assign addr[14631]= -2132665626;
assign addr[14632]= -2075296495;
assign addr[14633]= -1975871368;
assign addr[14634]= -1836405100;
assign addr[14635]= -1659723983;
assign addr[14636]= -1449408469;
assign addr[14637]= -1209720613;
assign addr[14638]= -945517704;
assign addr[14639]= -662153826;
assign addr[14640]= -365371365;
assign addr[14641]= -61184634;
assign addr[14642]= 244242007;
assign addr[14643]= 544719071;
assign addr[14644]= 834157373;
assign addr[14645]= 1106691431;
assign addr[14646]= 1356798326;
assign addr[14647]= 1579409630;
assign addr[14648]= 1770014111;
assign addr[14649]= 1924749160;
assign addr[14650]= 2040479063;
assign addr[14651]= 2114858546;
assign addr[14652]= 2146380306;
assign addr[14653]= 2134405552;
assign addr[14654]= 2079176953;
assign addr[14655]= 1981813720;
assign addr[14656]= 1844288924;
assign addr[14657]= 1669389513;
assign addr[14658]= 1460659832;
assign addr[14659]= 1222329801;
assign addr[14660]= 959229189;
assign addr[14661]= 676689746;
assign addr[14662]= 380437148;
assign addr[14663]= 76474970;
assign addr[14664]= -229036977;
assign addr[14665]= -529907477;
assign addr[14666]= -820039373;
assign addr[14667]= -1093553126;
assign addr[14668]= -1344905966;
assign addr[14669]= -1569004214;
assign addr[14670]= -1761306505;
assign addr[14671]= -1917915825;
assign addr[14672]= -2035658475;
assign addr[14673]= -2112148396;
assign addr[14674]= -2145835515;
assign addr[14675]= -2136037160;
assign addr[14676]= -2082951896;
assign addr[14677]= -1987655498;
assign addr[14678]= -1852079154;
assign addr[14679]= -1678970324;
assign addr[14680]= -1471837070;
assign addr[14681]= -1234876957;
assign addr[14682]= -972891995;
assign addr[14683]= -691191324;
assign addr[14684]= -395483624;
assign addr[14685]= -91761426;
assign addr[14686]= 213820322;
assign addr[14687]= 515068990;
assign addr[14688]= 805879757;
assign addr[14689]= 1080359326;
assign addr[14690]= 1332945355;
assign addr[14691]= 1558519173;
assign addr[14692]= 1752509516;
assign addr[14693]= 1910985158;
assign addr[14694]= 2030734582;
assign addr[14695]= 2109331059;
assign addr[14696]= 2145181827;
assign addr[14697]= 2137560369;
assign addr[14698]= 2086621133;
assign addr[14699]= 1993396407;
assign addr[14700]= 1859775393;
assign addr[14701]= 1688465931;
assign addr[14702]= 1482939614;
assign addr[14703]= 1247361445;
assign addr[14704]= 986505429;
assign addr[14705]= 705657826;
assign addr[14706]= 410510029;
assign addr[14707]= 107043224;
assign addr[14708]= -198592817;
assign addr[14709]= -500204365;
assign addr[14710]= -791679244;
assign addr[14711]= -1067110699;
assign addr[14712]= -1320917099;
assign addr[14713]= -1547955041;
assign addr[14714]= -1743623590;
assign addr[14715]= -1903957513;
assign addr[14716]= -2025707632;
assign addr[14717]= -2106406677;
assign addr[14718]= -2144419275;
assign addr[14719]= -2138975100;
assign addr[14720]= -2090184478;
assign addr[14721]= -1999036154;
assign addr[14722]= -1867377253;
assign addr[14723]= -1697875851;
assign addr[14724]= -1493966902;
assign addr[14725]= -1259782632;
assign addr[14726]= -1000068799;
assign addr[14727]= -720088517;
assign addr[14728]= -425515602;
assign addr[14729]= -122319591;
assign addr[14730]= 183355234;
assign addr[14731]= 485314355;
assign addr[14732]= 777438554;
assign addr[14733]= 1053807919;
assign addr[14734]= 1308821808;
assign addr[14735]= 1537312353;
assign addr[14736]= 1734649179;
assign addr[14737]= 1896833245;
assign addr[14738]= 2020577882;
assign addr[14739]= 2103375398;
assign addr[14740]= 2143547897;
assign addr[14741]= 2140281282;
assign addr[14742]= 2093641749;
assign addr[14743]= 2004574453;
assign addr[14744]= 1874884346;
assign addr[14745]= 1707199606;
assign addr[14746]= 1504918373;
assign addr[14747]= 1272139887;
assign addr[14748]= 1013581418;
assign addr[14749]= 734482665;
assign addr[14750]= 440499581;
assign addr[14751]= 137589750;
assign addr[14752]= -168108346;
assign addr[14753]= -470399716;
assign addr[14754]= -763158411;
assign addr[14755]= -1040451659;
assign addr[14756]= -1296660098;
assign addr[14757]= -1526591649;
assign addr[14758]= -1725586737;
assign addr[14759]= -1889612716;
assign addr[14760]= -2015345591;
assign addr[14761]= -2100237377;
assign addr[14762]= -2142567738;
assign addr[14763]= -2141478848;
assign addr[14764]= -2096992772;
assign addr[14765]= -2010011024;
assign addr[14766]= -1882296293;
assign addr[14767]= -1716436725;
assign addr[14768]= -1515793473;
assign addr[14769]= -1284432584;
assign addr[14770]= -1027042599;
assign addr[14771]= -748839539;
assign addr[14772]= -455461206;
assign addr[14773]= -152852926;
assign addr[14774]= 152852926;
assign addr[14775]= 455461206;
assign addr[14776]= 748839539;
assign addr[14777]= 1027042599;
assign addr[14778]= 1284432584;
assign addr[14779]= 1515793473;
assign addr[14780]= 1716436725;
assign addr[14781]= 1882296293;
assign addr[14782]= 2010011024;
assign addr[14783]= 2096992772;
assign addr[14784]= 2141478848;
assign addr[14785]= 2142567738;
assign addr[14786]= 2100237377;
assign addr[14787]= 2015345591;
assign addr[14788]= 1889612716;
assign addr[14789]= 1725586737;
assign addr[14790]= 1526591649;
assign addr[14791]= 1296660098;
assign addr[14792]= 1040451659;
assign addr[14793]= 763158411;
assign addr[14794]= 470399716;
assign addr[14795]= 168108346;
assign addr[14796]= -137589750;
assign addr[14797]= -440499581;
assign addr[14798]= -734482665;
assign addr[14799]= -1013581418;
assign addr[14800]= -1272139887;
assign addr[14801]= -1504918373;
assign addr[14802]= -1707199606;
assign addr[14803]= -1874884346;
assign addr[14804]= -2004574453;
assign addr[14805]= -2093641749;
assign addr[14806]= -2140281282;
assign addr[14807]= -2143547897;
assign addr[14808]= -2103375398;
assign addr[14809]= -2020577882;
assign addr[14810]= -1896833245;
assign addr[14811]= -1734649179;
assign addr[14812]= -1537312353;
assign addr[14813]= -1308821808;
assign addr[14814]= -1053807919;
assign addr[14815]= -777438554;
assign addr[14816]= -485314355;
assign addr[14817]= -183355234;
assign addr[14818]= 122319591;
assign addr[14819]= 425515602;
assign addr[14820]= 720088517;
assign addr[14821]= 1000068799;
assign addr[14822]= 1259782632;
assign addr[14823]= 1493966902;
assign addr[14824]= 1697875851;
assign addr[14825]= 1867377253;
assign addr[14826]= 1999036154;
assign addr[14827]= 2090184478;
assign addr[14828]= 2138975100;
assign addr[14829]= 2144419275;
assign addr[14830]= 2106406677;
assign addr[14831]= 2025707632;
assign addr[14832]= 1903957513;
assign addr[14833]= 1743623590;
assign addr[14834]= 1547955041;
assign addr[14835]= 1320917099;
assign addr[14836]= 1067110699;
assign addr[14837]= 791679244;
assign addr[14838]= 500204365;
assign addr[14839]= 198592817;
assign addr[14840]= -107043224;
assign addr[14841]= -410510029;
assign addr[14842]= -705657826;
assign addr[14843]= -986505429;
assign addr[14844]= -1247361445;
assign addr[14845]= -1482939614;
assign addr[14846]= -1688465931;
assign addr[14847]= -1859775393;
assign addr[14848]= -1993396407;
assign addr[14849]= -2086621133;
assign addr[14850]= -2137560369;
assign addr[14851]= -2145181827;
assign addr[14852]= -2109331059;
assign addr[14853]= -2030734582;
assign addr[14854]= -1910985158;
assign addr[14855]= -1752509516;
assign addr[14856]= -1558519173;
assign addr[14857]= -1332945355;
assign addr[14858]= -1080359326;
assign addr[14859]= -805879757;
assign addr[14860]= -515068990;
assign addr[14861]= -213820322;
assign addr[14862]= 91761426;
assign addr[14863]= 395483624;
assign addr[14864]= 691191324;
assign addr[14865]= 972891995;
assign addr[14866]= 1234876957;
assign addr[14867]= 1471837070;
assign addr[14868]= 1678970324;
assign addr[14869]= 1852079154;
assign addr[14870]= 1987655498;
assign addr[14871]= 2082951896;
assign addr[14872]= 2136037160;
assign addr[14873]= 2145835515;
assign addr[14874]= 2112148396;
assign addr[14875]= 2035658475;
assign addr[14876]= 1917915825;
assign addr[14877]= 1761306505;
assign addr[14878]= 1569004214;
assign addr[14879]= 1344905966;
assign addr[14880]= 1093553126;
assign addr[14881]= 820039373;
assign addr[14882]= 529907477;
assign addr[14883]= 229036977;
assign addr[14884]= -76474970;
assign addr[14885]= -380437148;
assign addr[14886]= -676689746;
assign addr[14887]= -959229189;
assign addr[14888]= -1222329801;
assign addr[14889]= -1460659832;
assign addr[14890]= -1669389513;
assign addr[14891]= -1844288924;
assign addr[14892]= -1981813720;
assign addr[14893]= -2079176953;
assign addr[14894]= -2134405552;
assign addr[14895]= -2146380306;
assign addr[14896]= -2114858546;
assign addr[14897]= -2040479063;
assign addr[14898]= -1924749160;
assign addr[14899]= -1770014111;
assign addr[14900]= -1579409630;
assign addr[14901]= -1356798326;
assign addr[14902]= -1106691431;
assign addr[14903]= -834157373;
assign addr[14904]= -544719071;
assign addr[14905]= -244242007;
assign addr[14906]= 61184634;
assign addr[14907]= 365371365;
assign addr[14908]= 662153826;
assign addr[14909]= 945517704;
assign addr[14910]= 1209720613;
assign addr[14911]= 1449408469;
assign addr[14912]= 1659723983;
assign addr[14913]= 1836405100;
assign addr[14914]= 1975871368;
assign addr[14915]= 2075296495;
assign addr[14916]= 2132665626;
assign addr[14917]= 2146816171;
assign addr[14918]= 2117461370;
assign addr[14919]= 2045196100;
assign addr[14920]= 1931484818;
assign addr[14921]= 1778631892;
assign addr[14922]= 1589734894;
assign addr[14923]= 1368621831;
assign addr[14924]= 1119773573;
assign addr[14925]= 848233042;
assign addr[14926]= 559503022;
assign addr[14927]= 259434643;
assign addr[14928]= -45891193;
assign addr[14929]= -350287041;
assign addr[14930]= -647584304;
assign addr[14931]= -931758235;
assign addr[14932]= -1197050035;
assign addr[14933]= -1438083551;
assign addr[14934]= -1649974225;
assign addr[14935]= -1828428082;
assign addr[14936]= -1969828744;
assign addr[14937]= -2071310720;
assign addr[14938]= -2130817471;
assign addr[14939]= -2147143090;
assign addr[14940]= -2119956737;
assign addr[14941]= -2049809346;
assign addr[14942]= -1938122457;
assign addr[14943]= -1787159411;
assign addr[14944]= -1599979481;
assign addr[14945]= -1380375881;
assign addr[14946]= -1132798888;
assign addr[14947]= -862265664;
assign addr[14948]= -574258580;
assign addr[14949]= -274614114;
assign addr[14950]= 30595422;
assign addr[14951]= 335184940;
assign addr[14952]= 632981917;
assign addr[14953]= 917951481;
assign addr[14954]= 1184318708;
assign addr[14955]= 1426685652;
assign addr[14956]= 1640140734;
assign addr[14957]= 1820358275;
assign addr[14958]= 1963686155;
assign addr[14959]= 2067219829;
assign addr[14960]= 2128861181;
assign addr[14961]= 2147361045;
assign addr[14962]= 2122344521;
assign addr[14963]= 2054318569;
assign addr[14964]= 1944661739;
assign addr[14965]= 1795596234;
assign addr[14966]= 1610142873;
assign addr[14967]= 1392059879;
assign addr[14968]= 1145766716;
assign addr[14969]= 876254528;
assign addr[14970]= 588984994;
assign addr[14971]= 289779648;
assign addr[14972]= -15298099;
assign addr[14973]= -320065829;
assign addr[14974]= -618347408;
assign addr[14975]= -904098143;
assign addr[14976]= -1171527280;
assign addr[14977]= -1415215352;
assign addr[14978]= -1630224009;
assign addr[14979]= -1812196087;
assign addr[14980]= -1957443913;
assign addr[14981]= -2063024031;
assign addr[14982]= -2126796855;
assign addr[14983]= -2147470025;
assign addr[14984]= -2124624598;
assign addr[14985]= -2058723538;
assign addr[14986]= -1951102334;
assign addr[14987]= -1803941934;
assign addr[14988]= -1620224553;
assign addr[14989]= -1403673233;
assign addr[14990]= -1158676398;
assign addr[14991]= -890198924;
assign addr[14992]= -603681519;
assign addr[14993]= -304930476;
assign addr[14994]= 0;
assign addr[14995]= 304930476;
assign addr[14996]= 603681519;
assign addr[14997]= 890198924;
assign addr[14998]= 1158676398;
assign addr[14999]= 1403673233;
assign addr[15000]= 1620224553;
assign addr[15001]= 1803941934;
assign addr[15002]= 1951102334;
assign addr[15003]= 2058723538;
assign addr[15004]= 2124624598;
assign addr[15005]= 2147470025;
assign addr[15006]= 2126796855;
assign addr[15007]= 2063024031;
assign addr[15008]= 1957443913;
assign addr[15009]= 1812196087;
assign addr[15010]= 1630224009;
assign addr[15011]= 1415215352;
assign addr[15012]= 1171527280;
assign addr[15013]= 904098143;
assign addr[15014]= 618347408;
assign addr[15015]= 320065829;
assign addr[15016]= 15298099;
assign addr[15017]= -289779648;
assign addr[15018]= -588984994;
assign addr[15019]= -876254528;
assign addr[15020]= -1145766716;
assign addr[15021]= -1392059879;
assign addr[15022]= -1610142873;
assign addr[15023]= -1795596234;
assign addr[15024]= -1944661739;
assign addr[15025]= -2054318569;
assign addr[15026]= -2122344521;
assign addr[15027]= -2147361045;
assign addr[15028]= -2128861181;
assign addr[15029]= -2067219829;
assign addr[15030]= -1963686155;
assign addr[15031]= -1820358275;
assign addr[15032]= -1640140734;
assign addr[15033]= -1426685652;
assign addr[15034]= -1184318708;
assign addr[15035]= -917951481;
assign addr[15036]= -632981917;
assign addr[15037]= -335184940;
assign addr[15038]= -30595422;
assign addr[15039]= 274614114;
assign addr[15040]= 574258580;
assign addr[15041]= 862265664;
assign addr[15042]= 1132798888;
assign addr[15043]= 1380375881;
assign addr[15044]= 1599979481;
assign addr[15045]= 1787159411;
assign addr[15046]= 1938122457;
assign addr[15047]= 2049809346;
assign addr[15048]= 2119956737;
assign addr[15049]= 2147143090;
assign addr[15050]= 2130817471;
assign addr[15051]= 2071310720;
assign addr[15052]= 1969828744;
assign addr[15053]= 1828428082;
assign addr[15054]= 1649974225;
assign addr[15055]= 1438083551;
assign addr[15056]= 1197050035;
assign addr[15057]= 931758235;
assign addr[15058]= 647584304;
assign addr[15059]= 350287041;
assign addr[15060]= 45891193;
assign addr[15061]= -259434643;
assign addr[15062]= -559503022;
assign addr[15063]= -848233042;
assign addr[15064]= -1119773573;
assign addr[15065]= -1368621831;
assign addr[15066]= -1589734894;
assign addr[15067]= -1778631892;
assign addr[15068]= -1931484818;
assign addr[15069]= -2045196100;
assign addr[15070]= -2117461370;
assign addr[15071]= -2146816171;
assign addr[15072]= -2132665626;
assign addr[15073]= -2075296495;
assign addr[15074]= -1975871368;
assign addr[15075]= -1836405100;
assign addr[15076]= -1659723983;
assign addr[15077]= -1449408469;
assign addr[15078]= -1209720613;
assign addr[15079]= -945517704;
assign addr[15080]= -662153826;
assign addr[15081]= -365371365;
assign addr[15082]= -61184634;
assign addr[15083]= 244242007;
assign addr[15084]= 544719071;
assign addr[15085]= 834157373;
assign addr[15086]= 1106691431;
assign addr[15087]= 1356798326;
assign addr[15088]= 1579409630;
assign addr[15089]= 1770014111;
assign addr[15090]= 1924749160;
assign addr[15091]= 2040479063;
assign addr[15092]= 2114858546;
assign addr[15093]= 2146380306;
assign addr[15094]= 2134405552;
assign addr[15095]= 2079176953;
assign addr[15096]= 1981813720;
assign addr[15097]= 1844288924;
assign addr[15098]= 1669389513;
assign addr[15099]= 1460659832;
assign addr[15100]= 1222329801;
assign addr[15101]= 959229189;
assign addr[15102]= 676689746;
assign addr[15103]= 380437148;
assign addr[15104]= 76474970;
assign addr[15105]= -229036977;
assign addr[15106]= -529907477;
assign addr[15107]= -820039373;
assign addr[15108]= -1093553126;
assign addr[15109]= -1344905966;
assign addr[15110]= -1569004214;
assign addr[15111]= -1761306505;
assign addr[15112]= -1917915825;
assign addr[15113]= -2035658475;
assign addr[15114]= -2112148396;
assign addr[15115]= -2145835515;
assign addr[15116]= -2136037160;
assign addr[15117]= -2082951896;
assign addr[15118]= -1987655498;
assign addr[15119]= -1852079154;
assign addr[15120]= -1678970324;
assign addr[15121]= -1471837070;
assign addr[15122]= -1234876957;
assign addr[15123]= -972891995;
assign addr[15124]= -691191324;
assign addr[15125]= -395483624;
assign addr[15126]= -91761426;
assign addr[15127]= 213820322;
assign addr[15128]= 515068990;
assign addr[15129]= 805879757;
assign addr[15130]= 1080359326;
assign addr[15131]= 1332945355;
assign addr[15132]= 1558519173;
assign addr[15133]= 1752509516;
assign addr[15134]= 1910985158;
assign addr[15135]= 2030734582;
assign addr[15136]= 2109331059;
assign addr[15137]= 2145181827;
assign addr[15138]= 2137560369;
assign addr[15139]= 2086621133;
assign addr[15140]= 1993396407;
assign addr[15141]= 1859775393;
assign addr[15142]= 1688465931;
assign addr[15143]= 1482939614;
assign addr[15144]= 1247361445;
assign addr[15145]= 986505429;
assign addr[15146]= 705657826;
assign addr[15147]= 410510029;
assign addr[15148]= 107043224;
assign addr[15149]= -198592817;
assign addr[15150]= -500204365;
assign addr[15151]= -791679244;
assign addr[15152]= -1067110699;
assign addr[15153]= -1320917099;
assign addr[15154]= -1547955041;
assign addr[15155]= -1743623590;
assign addr[15156]= -1903957513;
assign addr[15157]= -2025707632;
assign addr[15158]= -2106406677;
assign addr[15159]= -2144419275;
assign addr[15160]= -2138975100;
assign addr[15161]= -2090184478;
assign addr[15162]= -1999036154;
assign addr[15163]= -1867377253;
assign addr[15164]= -1697875851;
assign addr[15165]= -1493966902;
assign addr[15166]= -1259782632;
assign addr[15167]= -1000068799;
assign addr[15168]= -720088517;
assign addr[15169]= -425515602;
assign addr[15170]= -122319591;
assign addr[15171]= 183355234;
assign addr[15172]= 485314355;
assign addr[15173]= 777438554;
assign addr[15174]= 1053807919;
assign addr[15175]= 1308821808;
assign addr[15176]= 1537312353;
assign addr[15177]= 1734649179;
assign addr[15178]= 1896833245;
assign addr[15179]= 2020577882;
assign addr[15180]= 2103375398;
assign addr[15181]= 2143547897;
assign addr[15182]= 2140281282;
assign addr[15183]= 2093641749;
assign addr[15184]= 2004574453;
assign addr[15185]= 1874884346;
assign addr[15186]= 1707199606;
assign addr[15187]= 1504918373;
assign addr[15188]= 1272139887;
assign addr[15189]= 1013581418;
assign addr[15190]= 734482665;
assign addr[15191]= 440499581;
assign addr[15192]= 137589750;
assign addr[15193]= -168108346;
assign addr[15194]= -470399716;
assign addr[15195]= -763158411;
assign addr[15196]= -1040451659;
assign addr[15197]= -1296660098;
assign addr[15198]= -1526591649;
assign addr[15199]= -1725586737;
assign addr[15200]= -1889612716;
assign addr[15201]= -2015345591;
assign addr[15202]= -2100237377;
assign addr[15203]= -2142567738;
assign addr[15204]= -2141478848;
assign addr[15205]= -2096992772;
assign addr[15206]= -2010011024;
assign addr[15207]= -1882296293;
assign addr[15208]= -1716436725;
assign addr[15209]= -1515793473;
assign addr[15210]= -1284432584;
assign addr[15211]= -1027042599;
assign addr[15212]= -748839539;
assign addr[15213]= -455461206;
assign addr[15214]= -152852926;
assign addr[15215]= 152852926;
assign addr[15216]= 455461206;
assign addr[15217]= 748839539;
assign addr[15218]= 1027042599;
assign addr[15219]= 1284432584;
assign addr[15220]= 1515793473;
assign addr[15221]= 1716436725;
assign addr[15222]= 1882296293;
assign addr[15223]= 2010011024;
assign addr[15224]= 2096992772;
assign addr[15225]= 2141478848;
assign addr[15226]= 2142567738;
assign addr[15227]= 2100237377;
assign addr[15228]= 2015345591;
assign addr[15229]= 1889612716;
assign addr[15230]= 1725586737;
assign addr[15231]= 1526591649;
assign addr[15232]= 1296660098;
assign addr[15233]= 1040451659;
assign addr[15234]= 763158411;
assign addr[15235]= 470399716;
assign addr[15236]= 168108346;
assign addr[15237]= -137589750;
assign addr[15238]= -440499581;
assign addr[15239]= -734482665;
assign addr[15240]= -1013581418;
assign addr[15241]= -1272139887;
assign addr[15242]= -1504918373;
assign addr[15243]= -1707199606;
assign addr[15244]= -1874884346;
assign addr[15245]= -2004574453;
assign addr[15246]= -2093641749;
assign addr[15247]= -2140281282;
assign addr[15248]= -2143547897;
assign addr[15249]= -2103375398;
assign addr[15250]= -2020577882;
assign addr[15251]= -1896833245;
assign addr[15252]= -1734649179;
assign addr[15253]= -1537312353;
assign addr[15254]= -1308821808;
assign addr[15255]= -1053807919;
assign addr[15256]= -777438554;
assign addr[15257]= -485314355;
assign addr[15258]= -183355234;
assign addr[15259]= 122319591;
assign addr[15260]= 425515602;
assign addr[15261]= 720088517;
assign addr[15262]= 1000068799;
assign addr[15263]= 1259782632;
assign addr[15264]= 1493966902;
assign addr[15265]= 1697875851;
assign addr[15266]= 1867377253;
assign addr[15267]= 1999036154;
assign addr[15268]= 2090184478;
assign addr[15269]= 2138975100;
assign addr[15270]= 2144419275;
assign addr[15271]= 2106406677;
assign addr[15272]= 2025707632;
assign addr[15273]= 1903957513;
assign addr[15274]= 1743623590;
assign addr[15275]= 1547955041;
assign addr[15276]= 1320917099;
assign addr[15277]= 1067110699;
assign addr[15278]= 791679244;
assign addr[15279]= 500204365;
assign addr[15280]= 198592817;
assign addr[15281]= -107043224;
assign addr[15282]= -410510029;
assign addr[15283]= -705657826;
assign addr[15284]= -986505429;
assign addr[15285]= -1247361445;
assign addr[15286]= -1482939614;
assign addr[15287]= -1688465931;
assign addr[15288]= -1859775393;
assign addr[15289]= -1993396407;
assign addr[15290]= -2086621133;
assign addr[15291]= -2137560369;
assign addr[15292]= -2145181827;
assign addr[15293]= -2109331059;
assign addr[15294]= -2030734582;
assign addr[15295]= -1910985158;
assign addr[15296]= -1752509516;
assign addr[15297]= -1558519173;
assign addr[15298]= -1332945355;
assign addr[15299]= -1080359326;
assign addr[15300]= -805879757;
assign addr[15301]= -515068990;
assign addr[15302]= -213820322;
assign addr[15303]= 91761426;
assign addr[15304]= 395483624;
assign addr[15305]= 691191324;
assign addr[15306]= 972891995;
assign addr[15307]= 1234876957;
assign addr[15308]= 1471837070;
assign addr[15309]= 1678970324;
assign addr[15310]= 1852079154;
assign addr[15311]= 1987655498;
assign addr[15312]= 2082951896;
assign addr[15313]= 2136037160;
assign addr[15314]= 2145835515;
assign addr[15315]= 2112148396;
assign addr[15316]= 2035658475;
assign addr[15317]= 1917915825;
assign addr[15318]= 1761306505;
assign addr[15319]= 1569004214;
assign addr[15320]= 1344905966;
assign addr[15321]= 1093553126;
assign addr[15322]= 820039373;
assign addr[15323]= 529907477;
assign addr[15324]= 229036977;
assign addr[15325]= -76474970;
assign addr[15326]= -380437148;
assign addr[15327]= -676689746;
assign addr[15328]= -959229189;
assign addr[15329]= -1222329801;
assign addr[15330]= -1460659832;
assign addr[15331]= -1669389513;
assign addr[15332]= -1844288924;
assign addr[15333]= -1981813720;
assign addr[15334]= -2079176953;
assign addr[15335]= -2134405552;
assign addr[15336]= -2146380306;
assign addr[15337]= -2114858546;
assign addr[15338]= -2040479063;
assign addr[15339]= -1924749160;
assign addr[15340]= -1770014111;
assign addr[15341]= -1579409630;
assign addr[15342]= -1356798326;
assign addr[15343]= -1106691431;
assign addr[15344]= -834157373;
assign addr[15345]= -544719071;
assign addr[15346]= -244242007;
assign addr[15347]= 61184634;
assign addr[15348]= 365371365;
assign addr[15349]= 662153826;
assign addr[15350]= 945517704;
assign addr[15351]= 1209720613;
assign addr[15352]= 1449408469;
assign addr[15353]= 1659723983;
assign addr[15354]= 1836405100;
assign addr[15355]= 1975871368;
assign addr[15356]= 2075296495;
assign addr[15357]= 2132665626;
assign addr[15358]= 2146816171;
assign addr[15359]= 2117461370;
assign addr[15360]= 2045196100;
assign addr[15361]= 1931484818;
assign addr[15362]= 1778631892;
assign addr[15363]= 1589734894;
assign addr[15364]= 1368621831;
assign addr[15365]= 1119773573;
assign addr[15366]= 848233042;
assign addr[15367]= 559503022;
assign addr[15368]= 259434643;
assign addr[15369]= -45891193;
assign addr[15370]= -350287041;
assign addr[15371]= -647584304;
assign addr[15372]= -931758235;
assign addr[15373]= -1197050035;
assign addr[15374]= -1438083551;
assign addr[15375]= -1649974225;
assign addr[15376]= -1828428082;
assign addr[15377]= -1969828744;
assign addr[15378]= -2071310720;
assign addr[15379]= -2130817471;
assign addr[15380]= -2147143090;
assign addr[15381]= -2119956737;
assign addr[15382]= -2049809346;
assign addr[15383]= -1938122457;
assign addr[15384]= -1787159411;
assign addr[15385]= -1599979481;
assign addr[15386]= -1380375881;
assign addr[15387]= -1132798888;
assign addr[15388]= -862265664;
assign addr[15389]= -574258580;
assign addr[15390]= -274614114;
assign addr[15391]= 30595422;
assign addr[15392]= 335184940;
assign addr[15393]= 632981917;
assign addr[15394]= 917951481;
assign addr[15395]= 1184318708;
assign addr[15396]= 1426685652;
assign addr[15397]= 1640140734;
assign addr[15398]= 1820358275;
assign addr[15399]= 1963686155;
assign addr[15400]= 2067219829;
assign addr[15401]= 2128861181;
assign addr[15402]= 2147361045;
assign addr[15403]= 2122344521;
assign addr[15404]= 2054318569;
assign addr[15405]= 1944661739;
assign addr[15406]= 1795596234;
assign addr[15407]= 1610142873;
assign addr[15408]= 1392059879;
assign addr[15409]= 1145766716;
assign addr[15410]= 876254528;
assign addr[15411]= 588984994;
assign addr[15412]= 289779648;
assign addr[15413]= -15298099;
assign addr[15414]= -320065829;
assign addr[15415]= -618347408;
assign addr[15416]= -904098143;
assign addr[15417]= -1171527280;
assign addr[15418]= -1415215352;
assign addr[15419]= -1630224009;
assign addr[15420]= -1812196087;
assign addr[15421]= -1957443913;
assign addr[15422]= -2063024031;
assign addr[15423]= -2126796855;
assign addr[15424]= -2147470025;
assign addr[15425]= -2124624598;
assign addr[15426]= -2058723538;
assign addr[15427]= -1951102334;
assign addr[15428]= -1803941934;
assign addr[15429]= -1620224553;
assign addr[15430]= -1403673233;
assign addr[15431]= -1158676398;
assign addr[15432]= -890198924;
assign addr[15433]= -603681519;
assign addr[15434]= -304930476;
assign addr[15435]= 0;
assign addr[15436]= 304930476;
assign addr[15437]= 603681519;
assign addr[15438]= 890198924;
assign addr[15439]= 1158676398;
assign addr[15440]= 1403673233;
assign addr[15441]= 1620224553;
assign addr[15442]= 1803941934;
assign addr[15443]= 1951102334;
assign addr[15444]= 2058723538;
assign addr[15445]= 2124624598;
assign addr[15446]= 2147470025;
assign addr[15447]= 2126796855;
assign addr[15448]= 2063024031;
assign addr[15449]= 1957443913;
assign addr[15450]= 1812196087;
assign addr[15451]= 1630224009;
assign addr[15452]= 1415215352;
assign addr[15453]= 1171527280;
assign addr[15454]= 904098143;
assign addr[15455]= 618347408;
assign addr[15456]= 320065829;
assign addr[15457]= 15298099;
assign addr[15458]= -289779648;
assign addr[15459]= -588984994;
assign addr[15460]= -876254528;
assign addr[15461]= -1145766716;
assign addr[15462]= -1392059879;
assign addr[15463]= -1610142873;
assign addr[15464]= -1795596234;
assign addr[15465]= -1944661739;
assign addr[15466]= -2054318569;
assign addr[15467]= -2122344521;
assign addr[15468]= -2147361045;
assign addr[15469]= -2128861181;
assign addr[15470]= -2067219829;
assign addr[15471]= -1963686155;
assign addr[15472]= -1820358275;
assign addr[15473]= -1640140734;
assign addr[15474]= -1426685652;
assign addr[15475]= -1184318708;
assign addr[15476]= -917951481;
assign addr[15477]= -632981917;
assign addr[15478]= -335184940;
assign addr[15479]= -30595422;
assign addr[15480]= 274614114;
assign addr[15481]= 574258580;
assign addr[15482]= 862265664;
assign addr[15483]= 1132798888;
assign addr[15484]= 1380375881;
assign addr[15485]= 1599979481;
assign addr[15486]= 1787159411;
assign addr[15487]= 1938122457;
assign addr[15488]= 2049809346;
assign addr[15489]= 2119956737;
assign addr[15490]= 2147143090;
assign addr[15491]= 2130817471;
assign addr[15492]= 2071310720;
assign addr[15493]= 1969828744;
assign addr[15494]= 1828428082;
assign addr[15495]= 1649974225;
assign addr[15496]= 1438083551;
assign addr[15497]= 1197050035;
assign addr[15498]= 931758235;
assign addr[15499]= 647584304;
assign addr[15500]= 350287041;
assign addr[15501]= 45891193;
assign addr[15502]= -259434643;
assign addr[15503]= -559503022;
assign addr[15504]= -848233042;
assign addr[15505]= -1119773573;
assign addr[15506]= -1368621831;
assign addr[15507]= -1589734894;
assign addr[15508]= -1778631892;
assign addr[15509]= -1931484818;
assign addr[15510]= -2045196100;
assign addr[15511]= -2117461370;
assign addr[15512]= -2146816171;
assign addr[15513]= -2132665626;
assign addr[15514]= -2075296495;
assign addr[15515]= -1975871368;
assign addr[15516]= -1836405100;
assign addr[15517]= -1659723983;
assign addr[15518]= -1449408469;
assign addr[15519]= -1209720613;
assign addr[15520]= -945517704;
assign addr[15521]= -662153826;
assign addr[15522]= -365371365;
assign addr[15523]= -61184634;
assign addr[15524]= 244242007;
assign addr[15525]= 544719071;
assign addr[15526]= 834157373;
assign addr[15527]= 1106691431;
assign addr[15528]= 1356798326;
assign addr[15529]= 1579409630;
assign addr[15530]= 1770014111;
assign addr[15531]= 1924749160;
assign addr[15532]= 2040479063;
assign addr[15533]= 2114858546;
assign addr[15534]= 2146380306;
assign addr[15535]= 2134405552;
assign addr[15536]= 2079176953;
assign addr[15537]= 1981813720;
assign addr[15538]= 1844288924;
assign addr[15539]= 1669389513;
assign addr[15540]= 1460659832;
assign addr[15541]= 1222329801;
assign addr[15542]= 959229189;
assign addr[15543]= 676689746;
assign addr[15544]= 380437148;
assign addr[15545]= 76474970;
assign addr[15546]= -229036977;
assign addr[15547]= -529907477;
assign addr[15548]= -820039373;
assign addr[15549]= -1093553126;
assign addr[15550]= -1344905966;
assign addr[15551]= -1569004214;
assign addr[15552]= -1761306505;
assign addr[15553]= -1917915825;
assign addr[15554]= -2035658475;
assign addr[15555]= -2112148396;
assign addr[15556]= -2145835515;
assign addr[15557]= -2136037160;
assign addr[15558]= -2082951896;
assign addr[15559]= -1987655498;
assign addr[15560]= -1852079154;
assign addr[15561]= -1678970324;
assign addr[15562]= -1471837070;
assign addr[15563]= -1234876957;
assign addr[15564]= -972891995;
assign addr[15565]= -691191324;
assign addr[15566]= -395483624;
assign addr[15567]= -91761426;
assign addr[15568]= 213820322;
assign addr[15569]= 515068990;
assign addr[15570]= 805879757;
assign addr[15571]= 1080359326;
assign addr[15572]= 1332945355;
assign addr[15573]= 1558519173;
assign addr[15574]= 1752509516;
assign addr[15575]= 1910985158;
assign addr[15576]= 2030734582;
assign addr[15577]= 2109331059;
assign addr[15578]= 2145181827;
assign addr[15579]= 2137560369;
assign addr[15580]= 2086621133;
assign addr[15581]= 1993396407;
assign addr[15582]= 1859775393;
assign addr[15583]= 1688465931;
assign addr[15584]= 1482939614;
assign addr[15585]= 1247361445;
assign addr[15586]= 986505429;
assign addr[15587]= 705657826;
assign addr[15588]= 410510029;
assign addr[15589]= 107043224;
assign addr[15590]= -198592817;
assign addr[15591]= -500204365;
assign addr[15592]= -791679244;
assign addr[15593]= -1067110699;
assign addr[15594]= -1320917099;
assign addr[15595]= -1547955041;
assign addr[15596]= -1743623590;
assign addr[15597]= -1903957513;
assign addr[15598]= -2025707632;
assign addr[15599]= -2106406677;
assign addr[15600]= -2144419275;
assign addr[15601]= -2138975100;
assign addr[15602]= -2090184478;
assign addr[15603]= -1999036154;
assign addr[15604]= -1867377253;
assign addr[15605]= -1697875851;
assign addr[15606]= -1493966902;
assign addr[15607]= -1259782632;
assign addr[15608]= -1000068799;
assign addr[15609]= -720088517;
assign addr[15610]= -425515602;
assign addr[15611]= -122319591;
assign addr[15612]= 183355234;
assign addr[15613]= 485314355;
assign addr[15614]= 777438554;
assign addr[15615]= 1053807919;
assign addr[15616]= 1308821808;
assign addr[15617]= 1537312353;
assign addr[15618]= 1734649179;
assign addr[15619]= 1896833245;
assign addr[15620]= 2020577882;
assign addr[15621]= 2103375398;
assign addr[15622]= 2143547897;
assign addr[15623]= 2140281282;
assign addr[15624]= 2093641749;
assign addr[15625]= 2004574453;
assign addr[15626]= 1874884346;
assign addr[15627]= 1707199606;
assign addr[15628]= 1504918373;
assign addr[15629]= 1272139887;
assign addr[15630]= 1013581418;
assign addr[15631]= 734482665;
assign addr[15632]= 440499581;
assign addr[15633]= 137589750;
assign addr[15634]= -168108346;
assign addr[15635]= -470399716;
assign addr[15636]= -763158411;
assign addr[15637]= -1040451659;
assign addr[15638]= -1296660098;
assign addr[15639]= -1526591649;
assign addr[15640]= -1725586737;
assign addr[15641]= -1889612716;
assign addr[15642]= -2015345591;
assign addr[15643]= -2100237377;
assign addr[15644]= -2142567738;
assign addr[15645]= -2141478848;
assign addr[15646]= -2096992772;
assign addr[15647]= -2010011024;
assign addr[15648]= -1882296293;
assign addr[15649]= -1716436725;
assign addr[15650]= -1515793473;
assign addr[15651]= -1284432584;
assign addr[15652]= -1027042599;
assign addr[15653]= -748839539;
assign addr[15654]= -455461206;
assign addr[15655]= -152852926;
assign addr[15656]= 152852926;
assign addr[15657]= 455461206;
assign addr[15658]= 748839539;
assign addr[15659]= 1027042599;
assign addr[15660]= 1284432584;
assign addr[15661]= 1515793473;
assign addr[15662]= 1716436725;
assign addr[15663]= 1882296293;
assign addr[15664]= 2010011024;
assign addr[15665]= 2096992772;
assign addr[15666]= 2141478848;
assign addr[15667]= 2142567738;
assign addr[15668]= 2100237377;
assign addr[15669]= 2015345591;
assign addr[15670]= 1889612716;
assign addr[15671]= 1725586737;
assign addr[15672]= 1526591649;
assign addr[15673]= 1296660098;
assign addr[15674]= 1040451659;
assign addr[15675]= 763158411;
assign addr[15676]= 470399716;
assign addr[15677]= 168108346;
assign addr[15678]= -137589750;
assign addr[15679]= -440499581;
assign addr[15680]= -734482665;
assign addr[15681]= -1013581418;
assign addr[15682]= -1272139887;
assign addr[15683]= -1504918373;
assign addr[15684]= -1707199606;
assign addr[15685]= -1874884346;
assign addr[15686]= -2004574453;
assign addr[15687]= -2093641749;
assign addr[15688]= -2140281282;
assign addr[15689]= -2143547897;
assign addr[15690]= -2103375398;
assign addr[15691]= -2020577882;
assign addr[15692]= -1896833245;
assign addr[15693]= -1734649179;
assign addr[15694]= -1537312353;
assign addr[15695]= -1308821808;
assign addr[15696]= -1053807919;
assign addr[15697]= -777438554;
assign addr[15698]= -485314355;
assign addr[15699]= -183355234;
assign addr[15700]= 122319591;
assign addr[15701]= 425515602;
assign addr[15702]= 720088517;
assign addr[15703]= 1000068799;
assign addr[15704]= 1259782632;
assign addr[15705]= 1493966902;
assign addr[15706]= 1697875851;
assign addr[15707]= 1867377253;
assign addr[15708]= 1999036154;
assign addr[15709]= 2090184478;
assign addr[15710]= 2138975100;
assign addr[15711]= 2144419275;
assign addr[15712]= 2106406677;
assign addr[15713]= 2025707632;
assign addr[15714]= 1903957513;
assign addr[15715]= 1743623590;
assign addr[15716]= 1547955041;
assign addr[15717]= 1320917099;
assign addr[15718]= 1067110699;
assign addr[15719]= 791679244;
assign addr[15720]= 500204365;
assign addr[15721]= 198592817;
assign addr[15722]= -107043224;
assign addr[15723]= -410510029;
assign addr[15724]= -705657826;
assign addr[15725]= -986505429;
assign addr[15726]= -1247361445;
assign addr[15727]= -1482939614;
assign addr[15728]= -1688465931;
assign addr[15729]= -1859775393;
assign addr[15730]= -1993396407;
assign addr[15731]= -2086621133;
assign addr[15732]= -2137560369;
assign addr[15733]= -2145181827;
assign addr[15734]= -2109331059;
assign addr[15735]= -2030734582;
assign addr[15736]= -1910985158;
assign addr[15737]= -1752509516;
assign addr[15738]= -1558519173;
assign addr[15739]= -1332945355;
assign addr[15740]= -1080359326;
assign addr[15741]= -805879757;
assign addr[15742]= -515068990;
assign addr[15743]= -213820322;
assign addr[15744]= 91761426;
assign addr[15745]= 395483624;
assign addr[15746]= 691191324;
assign addr[15747]= 972891995;
assign addr[15748]= 1234876957;
assign addr[15749]= 1471837070;
assign addr[15750]= 1678970324;
assign addr[15751]= 1852079154;
assign addr[15752]= 1987655498;
assign addr[15753]= 2082951896;
assign addr[15754]= 2136037160;
assign addr[15755]= 2145835515;
assign addr[15756]= 2112148396;
assign addr[15757]= 2035658475;
assign addr[15758]= 1917915825;
assign addr[15759]= 1761306505;
assign addr[15760]= 1569004214;
assign addr[15761]= 1344905966;
assign addr[15762]= 1093553126;
assign addr[15763]= 820039373;
assign addr[15764]= 529907477;
assign addr[15765]= 229036977;
assign addr[15766]= -76474970;
assign addr[15767]= -380437148;
assign addr[15768]= -676689746;
assign addr[15769]= -959229189;
assign addr[15770]= -1222329801;
assign addr[15771]= -1460659832;
assign addr[15772]= -1669389513;
assign addr[15773]= -1844288924;
assign addr[15774]= -1981813720;
assign addr[15775]= -2079176953;
assign addr[15776]= -2134405552;
assign addr[15777]= -2146380306;
assign addr[15778]= -2114858546;
assign addr[15779]= -2040479063;
assign addr[15780]= -1924749160;
assign addr[15781]= -1770014111;
assign addr[15782]= -1579409630;
assign addr[15783]= -1356798326;
assign addr[15784]= -1106691431;
assign addr[15785]= -834157373;
assign addr[15786]= -544719071;
assign addr[15787]= -244242007;
assign addr[15788]= 61184634;
assign addr[15789]= 365371365;
assign addr[15790]= 662153826;
assign addr[15791]= 945517704;
assign addr[15792]= 1209720613;
assign addr[15793]= 1449408469;
assign addr[15794]= 1659723983;
assign addr[15795]= 1836405100;
assign addr[15796]= 1975871368;
assign addr[15797]= 2075296495;
assign addr[15798]= 2132665626;
assign addr[15799]= 2146816171;
assign addr[15800]= 2117461370;
assign addr[15801]= 2045196100;
assign addr[15802]= 1931484818;
assign addr[15803]= 1778631892;
assign addr[15804]= 1589734894;
assign addr[15805]= 1368621831;
assign addr[15806]= 1119773573;
assign addr[15807]= 848233042;
assign addr[15808]= 559503022;
assign addr[15809]= 259434643;
assign addr[15810]= -45891193;
assign addr[15811]= -350287041;
assign addr[15812]= -647584304;
assign addr[15813]= -931758235;
assign addr[15814]= -1197050035;
assign addr[15815]= -1438083551;
assign addr[15816]= -1649974225;
assign addr[15817]= -1828428082;
assign addr[15818]= -1969828744;
assign addr[15819]= -2071310720;
assign addr[15820]= -2130817471;
assign addr[15821]= -2147143090;
assign addr[15822]= -2119956737;
assign addr[15823]= -2049809346;
assign addr[15824]= -1938122457;
assign addr[15825]= -1787159411;
assign addr[15826]= -1599979481;
assign addr[15827]= -1380375881;
assign addr[15828]= -1132798888;
assign addr[15829]= -862265664;
assign addr[15830]= -574258580;
assign addr[15831]= -274614114;
assign addr[15832]= 30595422;
assign addr[15833]= 335184940;
assign addr[15834]= 632981917;
assign addr[15835]= 917951481;
assign addr[15836]= 1184318708;
assign addr[15837]= 1426685652;
assign addr[15838]= 1640140734;
assign addr[15839]= 1820358275;
assign addr[15840]= 1963686155;
assign addr[15841]= 2067219829;
assign addr[15842]= 2128861181;
assign addr[15843]= 2147361045;
assign addr[15844]= 2122344521;
assign addr[15845]= 2054318569;
assign addr[15846]= 1944661739;
assign addr[15847]= 1795596234;
assign addr[15848]= 1610142873;
assign addr[15849]= 1392059879;
assign addr[15850]= 1145766716;
assign addr[15851]= 876254528;
assign addr[15852]= 588984994;
assign addr[15853]= 289779648;
assign addr[15854]= -15298099;
assign addr[15855]= -320065829;
assign addr[15856]= -618347408;
assign addr[15857]= -904098143;
assign addr[15858]= -1171527280;
assign addr[15859]= -1415215352;
assign addr[15860]= -1630224009;
assign addr[15861]= -1812196087;
assign addr[15862]= -1957443913;
assign addr[15863]= -2063024031;
assign addr[15864]= -2126796855;
assign addr[15865]= -2147470025;
assign addr[15866]= -2124624598;
assign addr[15867]= -2058723538;
assign addr[15868]= -1951102334;
assign addr[15869]= -1803941934;
assign addr[15870]= -1620224553;
assign addr[15871]= -1403673233;
assign addr[15872]= -1158676398;
assign addr[15873]= -890198924;
assign addr[15874]= -603681519;
assign addr[15875]= -304930476;
assign addr[15876]= 0;
assign addr[15877]= 304930476;
assign addr[15878]= 603681519;
assign addr[15879]= 890198924;
assign addr[15880]= 1158676398;
assign addr[15881]= 1403673233;
assign addr[15882]= 1620224553;
assign addr[15883]= 1803941934;
assign addr[15884]= 1951102334;
assign addr[15885]= 2058723538;
assign addr[15886]= 2124624598;
assign addr[15887]= 2147470025;
assign addr[15888]= 2126796855;
assign addr[15889]= 2063024031;
assign addr[15890]= 1957443913;
assign addr[15891]= 1812196087;
assign addr[15892]= 1630224009;
assign addr[15893]= 1415215352;
assign addr[15894]= 1171527280;
assign addr[15895]= 904098143;
assign addr[15896]= 618347408;
assign addr[15897]= 320065829;
assign addr[15898]= 15298099;
assign addr[15899]= -289779648;
assign addr[15900]= -588984994;
assign addr[15901]= -876254528;
assign addr[15902]= -1145766716;
assign addr[15903]= -1392059879;
assign addr[15904]= -1610142873;
assign addr[15905]= -1795596234;
assign addr[15906]= -1944661739;
assign addr[15907]= -2054318569;
assign addr[15908]= -2122344521;
assign addr[15909]= -2147361045;
assign addr[15910]= -2128861181;
assign addr[15911]= -2067219829;
assign addr[15912]= -1963686155;
assign addr[15913]= -1820358275;
assign addr[15914]= -1640140734;
assign addr[15915]= -1426685652;
assign addr[15916]= -1184318708;
assign addr[15917]= -917951481;
assign addr[15918]= -632981917;
assign addr[15919]= -335184940;
assign addr[15920]= -30595422;
assign addr[15921]= 274614114;
assign addr[15922]= 574258580;
assign addr[15923]= 862265664;
assign addr[15924]= 1132798888;
assign addr[15925]= 1380375881;
assign addr[15926]= 1599979481;
assign addr[15927]= 1787159411;
assign addr[15928]= 1938122457;
assign addr[15929]= 2049809346;
assign addr[15930]= 2119956737;
assign addr[15931]= 2147143090;
assign addr[15932]= 2130817471;
assign addr[15933]= 2071310720;
assign addr[15934]= 1969828744;
assign addr[15935]= 1828428082;
assign addr[15936]= 1649974225;
assign addr[15937]= 1438083551;
assign addr[15938]= 1197050035;
assign addr[15939]= 931758235;
assign addr[15940]= 647584304;
assign addr[15941]= 350287041;
assign addr[15942]= 45891193;
assign addr[15943]= -259434643;
assign addr[15944]= -559503022;
assign addr[15945]= -848233042;
assign addr[15946]= -1119773573;
assign addr[15947]= -1368621831;
assign addr[15948]= -1589734894;
assign addr[15949]= -1778631892;
assign addr[15950]= -1931484818;
assign addr[15951]= -2045196100;
assign addr[15952]= -2117461370;
assign addr[15953]= -2146816171;
assign addr[15954]= -2132665626;
assign addr[15955]= -2075296495;
assign addr[15956]= -1975871368;
assign addr[15957]= -1836405100;
assign addr[15958]= -1659723983;
assign addr[15959]= -1449408469;
assign addr[15960]= -1209720613;
assign addr[15961]= -945517704;
assign addr[15962]= -662153826;
assign addr[15963]= -365371365;
assign addr[15964]= -61184634;
assign addr[15965]= 244242007;
assign addr[15966]= 544719071;
assign addr[15967]= 834157373;
assign addr[15968]= 1106691431;
assign addr[15969]= 1356798326;
assign addr[15970]= 1579409630;
assign addr[15971]= 1770014111;
assign addr[15972]= 1924749160;
assign addr[15973]= 2040479063;
assign addr[15974]= 2114858546;
assign addr[15975]= 2146380306;
assign addr[15976]= 2134405552;
assign addr[15977]= 2079176953;
assign addr[15978]= 1981813720;
assign addr[15979]= 1844288924;
assign addr[15980]= 1669389513;
assign addr[15981]= 1460659832;
assign addr[15982]= 1222329801;
assign addr[15983]= 959229189;
assign addr[15984]= 676689746;
assign addr[15985]= 380437148;
assign addr[15986]= 76474970;
assign addr[15987]= -229036977;
assign addr[15988]= -529907477;
assign addr[15989]= -820039373;
assign addr[15990]= -1093553126;
assign addr[15991]= -1344905966;
assign addr[15992]= -1569004214;
assign addr[15993]= -1761306505;
assign addr[15994]= -1917915825;
assign addr[15995]= -2035658475;
assign addr[15996]= -2112148396;
assign addr[15997]= -2145835515;
assign addr[15998]= -2136037160;
assign addr[15999]= -2082951896;
assign addr[16000]= -1987655498;
assign addr[16001]= -1852079154;
assign addr[16002]= -1678970324;
assign addr[16003]= -1471837070;
assign addr[16004]= -1234876957;
assign addr[16005]= -972891995;
assign addr[16006]= -691191324;
assign addr[16007]= -395483624;
assign addr[16008]= -91761426;
assign addr[16009]= 213820322;
assign addr[16010]= 515068990;
assign addr[16011]= 805879757;
assign addr[16012]= 1080359326;
assign addr[16013]= 1332945355;
assign addr[16014]= 1558519173;
assign addr[16015]= 1752509516;
assign addr[16016]= 1910985158;
assign addr[16017]= 2030734582;
assign addr[16018]= 2109331059;
assign addr[16019]= 2145181827;
assign addr[16020]= 2137560369;
assign addr[16021]= 2086621133;
assign addr[16022]= 1993396407;
assign addr[16023]= 1859775393;
assign addr[16024]= 1688465931;
assign addr[16025]= 1482939614;
assign addr[16026]= 1247361445;
assign addr[16027]= 986505429;
assign addr[16028]= 705657826;
assign addr[16029]= 410510029;
assign addr[16030]= 107043224;
assign addr[16031]= -198592817;
assign addr[16032]= -500204365;
assign addr[16033]= -791679244;
assign addr[16034]= -1067110699;
assign addr[16035]= -1320917099;
assign addr[16036]= -1547955041;
assign addr[16037]= -1743623590;
assign addr[16038]= -1903957513;
assign addr[16039]= -2025707632;
assign addr[16040]= -2106406677;
assign addr[16041]= -2144419275;
assign addr[16042]= -2138975100;
assign addr[16043]= -2090184478;
assign addr[16044]= -1999036154;
assign addr[16045]= -1867377253;
assign addr[16046]= -1697875851;
assign addr[16047]= -1493966902;
assign addr[16048]= -1259782632;
assign addr[16049]= -1000068799;
assign addr[16050]= -720088517;
assign addr[16051]= -425515602;
assign addr[16052]= -122319591;
assign addr[16053]= 183355234;
assign addr[16054]= 485314355;
assign addr[16055]= 777438554;
assign addr[16056]= 1053807919;
assign addr[16057]= 1308821808;
assign addr[16058]= 1537312353;
assign addr[16059]= 1734649179;
assign addr[16060]= 1896833245;
assign addr[16061]= 2020577882;
assign addr[16062]= 2103375398;
assign addr[16063]= 2143547897;
assign addr[16064]= 2140281282;
assign addr[16065]= 2093641749;
assign addr[16066]= 2004574453;
assign addr[16067]= 1874884346;
assign addr[16068]= 1707199606;
assign addr[16069]= 1504918373;
assign addr[16070]= 1272139887;
assign addr[16071]= 1013581418;
assign addr[16072]= 734482665;
assign addr[16073]= 440499581;
assign addr[16074]= 137589750;
assign addr[16075]= -168108346;
assign addr[16076]= -470399716;
assign addr[16077]= -763158411;
assign addr[16078]= -1040451659;
assign addr[16079]= -1296660098;
assign addr[16080]= -1526591649;
assign addr[16081]= -1725586737;
assign addr[16082]= -1889612716;
assign addr[16083]= -2015345591;
assign addr[16084]= -2100237377;
assign addr[16085]= -2142567738;
assign addr[16086]= -2141478848;
assign addr[16087]= -2096992772;
assign addr[16088]= -2010011024;
assign addr[16089]= -1882296293;
assign addr[16090]= -1716436725;
assign addr[16091]= -1515793473;
assign addr[16092]= -1284432584;
assign addr[16093]= -1027042599;
assign addr[16094]= -748839539;
assign addr[16095]= -455461206;
assign addr[16096]= -152852926;
assign addr[16097]= 152852926;
assign addr[16098]= 455461206;
assign addr[16099]= 748839539;
assign addr[16100]= 1027042599;
assign addr[16101]= 1284432584;
assign addr[16102]= 1515793473;
assign addr[16103]= 1716436725;
assign addr[16104]= 1882296293;
assign addr[16105]= 2010011024;
assign addr[16106]= 2096992772;
assign addr[16107]= 2141478848;
assign addr[16108]= 2142567738;
assign addr[16109]= 2100237377;
assign addr[16110]= 2015345591;
assign addr[16111]= 1889612716;
assign addr[16112]= 1725586737;
assign addr[16113]= 1526591649;
assign addr[16114]= 1296660098;
assign addr[16115]= 1040451659;
assign addr[16116]= 763158411;
assign addr[16117]= 470399716;
assign addr[16118]= 168108346;
assign addr[16119]= -137589750;
assign addr[16120]= -440499581;
assign addr[16121]= -734482665;
assign addr[16122]= -1013581418;
assign addr[16123]= -1272139887;
assign addr[16124]= -1504918373;
assign addr[16125]= -1707199606;
assign addr[16126]= -1874884346;
assign addr[16127]= -2004574453;
assign addr[16128]= -2093641749;
assign addr[16129]= -2140281282;
assign addr[16130]= -2143547897;
assign addr[16131]= -2103375398;
assign addr[16132]= -2020577882;
assign addr[16133]= -1896833245;
assign addr[16134]= -1734649179;
assign addr[16135]= -1537312353;
assign addr[16136]= -1308821808;
assign addr[16137]= -1053807919;
assign addr[16138]= -777438554;
assign addr[16139]= -485314355;
assign addr[16140]= -183355234;
assign addr[16141]= 122319591;
assign addr[16142]= 425515602;
assign addr[16143]= 720088517;
assign addr[16144]= 1000068799;
assign addr[16145]= 1259782632;
assign addr[16146]= 1493966902;
assign addr[16147]= 1697875851;
assign addr[16148]= 1867377253;
assign addr[16149]= 1999036154;
assign addr[16150]= 2090184478;
assign addr[16151]= 2138975100;
assign addr[16152]= 2144419275;
assign addr[16153]= 2106406677;
assign addr[16154]= 2025707632;
assign addr[16155]= 1903957513;
assign addr[16156]= 1743623590;
assign addr[16157]= 1547955041;
assign addr[16158]= 1320917099;
assign addr[16159]= 1067110699;
assign addr[16160]= 791679244;
assign addr[16161]= 500204365;
assign addr[16162]= 198592817;
assign addr[16163]= -107043224;
assign addr[16164]= -410510029;
assign addr[16165]= -705657826;
assign addr[16166]= -986505429;
assign addr[16167]= -1247361445;
assign addr[16168]= -1482939614;
assign addr[16169]= -1688465931;
assign addr[16170]= -1859775393;
assign addr[16171]= -1993396407;
assign addr[16172]= -2086621133;
assign addr[16173]= -2137560369;
assign addr[16174]= -2145181827;
assign addr[16175]= -2109331059;
assign addr[16176]= -2030734582;
assign addr[16177]= -1910985158;
assign addr[16178]= -1752509516;
assign addr[16179]= -1558519173;
assign addr[16180]= -1332945355;
assign addr[16181]= -1080359326;
assign addr[16182]= -805879757;
assign addr[16183]= -515068990;
assign addr[16184]= -213820322;
assign addr[16185]= 91761426;
assign addr[16186]= 395483624;
assign addr[16187]= 691191324;
assign addr[16188]= 972891995;
assign addr[16189]= 1234876957;
assign addr[16190]= 1471837070;
assign addr[16191]= 1678970324;
assign addr[16192]= 1852079154;
assign addr[16193]= 1987655498;
assign addr[16194]= 2082951896;
assign addr[16195]= 2136037160;
assign addr[16196]= 2145835515;
assign addr[16197]= 2112148396;
assign addr[16198]= 2035658475;
assign addr[16199]= 1917915825;
assign addr[16200]= 1761306505;
assign addr[16201]= 1569004214;
assign addr[16202]= 1344905966;
assign addr[16203]= 1093553126;
assign addr[16204]= 820039373;
assign addr[16205]= 529907477;
assign addr[16206]= 229036977;
assign addr[16207]= -76474970;
assign addr[16208]= -380437148;
assign addr[16209]= -676689746;
assign addr[16210]= -959229189;
assign addr[16211]= -1222329801;
assign addr[16212]= -1460659832;
assign addr[16213]= -1669389513;
assign addr[16214]= -1844288924;
assign addr[16215]= -1981813720;
assign addr[16216]= -2079176953;
assign addr[16217]= -2134405552;
assign addr[16218]= -2146380306;
assign addr[16219]= -2114858546;
assign addr[16220]= -2040479063;
assign addr[16221]= -1924749160;
assign addr[16222]= -1770014111;
assign addr[16223]= -1579409630;
assign addr[16224]= -1356798326;
assign addr[16225]= -1106691431;
assign addr[16226]= -834157373;
assign addr[16227]= -544719071;
assign addr[16228]= -244242007;
assign addr[16229]= 61184634;
assign addr[16230]= 365371365;
assign addr[16231]= 662153826;
assign addr[16232]= 945517704;
assign addr[16233]= 1209720613;
assign addr[16234]= 1449408469;
assign addr[16235]= 1659723983;
assign addr[16236]= 1836405100;
assign addr[16237]= 1975871368;
assign addr[16238]= 2075296495;
assign addr[16239]= 2132665626;
assign addr[16240]= 2146816171;
assign addr[16241]= 2117461370;
assign addr[16242]= 2045196100;
assign addr[16243]= 1931484818;
assign addr[16244]= 1778631892;
assign addr[16245]= 1589734894;
assign addr[16246]= 1368621831;
assign addr[16247]= 1119773573;
assign addr[16248]= 848233042;
assign addr[16249]= 559503022;
assign addr[16250]= 259434643;
assign addr[16251]= -45891193;
assign addr[16252]= -350287041;
assign addr[16253]= -647584304;
assign addr[16254]= -931758235;
assign addr[16255]= -1197050035;
assign addr[16256]= -1438083551;
assign addr[16257]= -1649974225;
assign addr[16258]= -1828428082;
assign addr[16259]= -1969828744;
assign addr[16260]= -2071310720;
assign addr[16261]= -2130817471;
assign addr[16262]= -2147143090;
assign addr[16263]= -2119956737;
assign addr[16264]= -2049809346;
assign addr[16265]= -1938122457;
assign addr[16266]= -1787159411;
assign addr[16267]= -1599979481;
assign addr[16268]= -1380375881;
assign addr[16269]= -1132798888;
assign addr[16270]= -862265664;
assign addr[16271]= -574258580;
assign addr[16272]= -274614114;
assign addr[16273]= 30595422;
assign addr[16274]= 335184940;
assign addr[16275]= 632981917;
assign addr[16276]= 917951481;
assign addr[16277]= 1184318708;
assign addr[16278]= 1426685652;
assign addr[16279]= 1640140734;
assign addr[16280]= 1820358275;
assign addr[16281]= 1963686155;
assign addr[16282]= 2067219829;
assign addr[16283]= 2128861181;
assign addr[16284]= 2147361045;
assign addr[16285]= 2122344521;
assign addr[16286]= 2054318569;
assign addr[16287]= 1944661739;
assign addr[16288]= 1795596234;
assign addr[16289]= 1610142873;
assign addr[16290]= 1392059879;
assign addr[16291]= 1145766716;
assign addr[16292]= 876254528;
assign addr[16293]= 588984994;
assign addr[16294]= 289779648;
assign addr[16295]= -15298099;
assign addr[16296]= -320065829;
assign addr[16297]= -618347408;
assign addr[16298]= -904098143;
assign addr[16299]= -1171527280;
assign addr[16300]= -1415215352;
assign addr[16301]= -1630224009;
assign addr[16302]= -1812196087;
assign addr[16303]= -1957443913;
assign addr[16304]= -2063024031;
assign addr[16305]= -2126796855;
assign addr[16306]= -2147470025;
assign addr[16307]= -2124624598;
assign addr[16308]= -2058723538;
assign addr[16309]= -1951102334;
assign addr[16310]= -1803941934;
assign addr[16311]= -1620224553;
assign addr[16312]= -1403673233;
assign addr[16313]= -1158676398;
assign addr[16314]= -890198924;
assign addr[16315]= -603681519;
assign addr[16316]= -304930476;
assign addr[16317]= 0;
assign addr[16318]= 304930476;
assign addr[16319]= 603681519;
assign addr[16320]= 890198924;
assign addr[16321]= 1158676398;
assign addr[16322]= 1403673233;
assign addr[16323]= 1620224553;
assign addr[16324]= 1803941934;
assign addr[16325]= 1951102334;
assign addr[16326]= 2058723538;
assign addr[16327]= 2124624598;
assign addr[16328]= 2147470025;
assign addr[16329]= 2126796855;
assign addr[16330]= 2063024031;
assign addr[16331]= 1957443913;
assign addr[16332]= 1812196087;
assign addr[16333]= 1630224009;
assign addr[16334]= 1415215352;
assign addr[16335]= 1171527280;
assign addr[16336]= 904098143;
assign addr[16337]= 618347408;
assign addr[16338]= 320065829;
assign addr[16339]= 15298099;
assign addr[16340]= -289779648;
assign addr[16341]= -588984994;
assign addr[16342]= -876254528;
assign addr[16343]= -1145766716;
assign addr[16344]= -1392059879;
assign addr[16345]= -1610142873;
assign addr[16346]= -1795596234;
assign addr[16347]= -1944661739;
assign addr[16348]= -2054318569;
assign addr[16349]= -2122344521;
assign addr[16350]= -2147361045;
assign addr[16351]= -2128861181;
assign addr[16352]= -2067219829;
assign addr[16353]= -1963686155;
assign addr[16354]= -1820358275;
assign addr[16355]= -1640140734;
assign addr[16356]= -1426685652;
assign addr[16357]= -1184318708;
assign addr[16358]= -917951481;
assign addr[16359]= -632981917;
assign addr[16360]= -335184940;
assign addr[16361]= -30595422;
assign addr[16362]= 274614114;
assign addr[16363]= 574258580;
assign addr[16364]= 862265664;
assign addr[16365]= 1132798888;
assign addr[16366]= 1380375881;
assign addr[16367]= 1599979481;
assign addr[16368]= 1787159411;
assign addr[16369]= 1938122457;
assign addr[16370]= 2049809346;
assign addr[16371]= 2119956737;
assign addr[16372]= 2147143090;
assign addr[16373]= 2130817471;
assign addr[16374]= 2071310720;
assign addr[16375]= 1969828744;
assign addr[16376]= 1828428082;
assign addr[16377]= 1649974225;
assign addr[16378]= 1438083551;
assign addr[16379]= 1197050035;
assign addr[16380]= 931758235;
assign addr[16381]= 647584304;
assign addr[16382]= 350287041;
assign addr[16383]= 45891193;
assign addr[16384]= -259434643;
assign addr[16385]= -559503022;
assign addr[16386]= -848233042;
assign addr[16387]= -1119773573;
assign addr[16388]= -1368621831;
assign addr[16389]= -1589734894;
assign addr[16390]= -1778631892;
assign addr[16391]= -1931484818;
assign addr[16392]= -2045196100;
assign addr[16393]= -2117461370;
assign addr[16394]= -2146816171;
assign addr[16395]= -2132665626;
assign addr[16396]= -2075296495;
assign addr[16397]= -1975871368;
assign addr[16398]= -1836405100;
assign addr[16399]= -1659723983;
assign addr[16400]= -1449408469;
assign addr[16401]= -1209720613;
assign addr[16402]= -945517704;
assign addr[16403]= -662153826;
assign addr[16404]= -365371365;
assign addr[16405]= -61184634;
assign addr[16406]= 244242007;
assign addr[16407]= 544719071;
assign addr[16408]= 834157373;
assign addr[16409]= 1106691431;
assign addr[16410]= 1356798326;
assign addr[16411]= 1579409630;
assign addr[16412]= 1770014111;
assign addr[16413]= 1924749160;
assign addr[16414]= 2040479063;
assign addr[16415]= 2114858546;
assign addr[16416]= 2146380306;
assign addr[16417]= 2134405552;
assign addr[16418]= 2079176953;
assign addr[16419]= 1981813720;
assign addr[16420]= 1844288924;
assign addr[16421]= 1669389513;
assign addr[16422]= 1460659832;
assign addr[16423]= 1222329801;
assign addr[16424]= 959229189;
assign addr[16425]= 676689746;
assign addr[16426]= 380437148;
assign addr[16427]= 76474970;
assign addr[16428]= -229036977;
assign addr[16429]= -529907477;
assign addr[16430]= -820039373;
assign addr[16431]= -1093553126;
assign addr[16432]= -1344905966;
assign addr[16433]= -1569004214;
assign addr[16434]= -1761306505;
assign addr[16435]= -1917915825;
assign addr[16436]= -2035658475;
assign addr[16437]= -2112148396;
assign addr[16438]= -2145835515;
assign addr[16439]= -2136037160;
assign addr[16440]= -2082951896;
assign addr[16441]= -1987655498;
assign addr[16442]= -1852079154;
assign addr[16443]= -1678970324;
assign addr[16444]= -1471837070;
assign addr[16445]= -1234876957;
assign addr[16446]= -972891995;
assign addr[16447]= -691191324;
assign addr[16448]= -395483624;
assign addr[16449]= -91761426;
assign addr[16450]= 213820322;
assign addr[16451]= 515068990;
assign addr[16452]= 805879757;
assign addr[16453]= 1080359326;
assign addr[16454]= 1332945355;
assign addr[16455]= 1558519173;
assign addr[16456]= 1752509516;
assign addr[16457]= 1910985158;
assign addr[16458]= 2030734582;
assign addr[16459]= 2109331059;
assign addr[16460]= 2145181827;
assign addr[16461]= 2137560369;
assign addr[16462]= 2086621133;
assign addr[16463]= 1993396407;
assign addr[16464]= 1859775393;
assign addr[16465]= 1688465931;
assign addr[16466]= 1482939614;
assign addr[16467]= 1247361445;
assign addr[16468]= 986505429;
assign addr[16469]= 705657826;
assign addr[16470]= 410510029;
assign addr[16471]= 107043224;
assign addr[16472]= -198592817;
assign addr[16473]= -500204365;
assign addr[16474]= -791679244;
assign addr[16475]= -1067110699;
assign addr[16476]= -1320917099;
assign addr[16477]= -1547955041;
assign addr[16478]= -1743623590;
assign addr[16479]= -1903957513;
assign addr[16480]= -2025707632;
assign addr[16481]= -2106406677;
assign addr[16482]= -2144419275;
assign addr[16483]= -2138975100;
assign addr[16484]= -2090184478;
assign addr[16485]= -1999036154;
assign addr[16486]= -1867377253;
assign addr[16487]= -1697875851;
assign addr[16488]= -1493966902;
assign addr[16489]= -1259782632;
assign addr[16490]= -1000068799;
assign addr[16491]= -720088517;
assign addr[16492]= -425515602;
assign addr[16493]= -122319591;
assign addr[16494]= 183355234;
assign addr[16495]= 485314355;
assign addr[16496]= 777438554;
assign addr[16497]= 1053807919;
assign addr[16498]= 1308821808;
assign addr[16499]= 1537312353;
assign addr[16500]= 1734649179;
assign addr[16501]= 1896833245;
assign addr[16502]= 2020577882;
assign addr[16503]= 2103375398;
assign addr[16504]= 2143547897;
assign addr[16505]= 2140281282;
assign addr[16506]= 2093641749;
assign addr[16507]= 2004574453;
assign addr[16508]= 1874884346;
assign addr[16509]= 1707199606;
assign addr[16510]= 1504918373;
assign addr[16511]= 1272139887;
assign addr[16512]= 1013581418;
assign addr[16513]= 734482665;
assign addr[16514]= 440499581;
assign addr[16515]= 137589750;
assign addr[16516]= -168108346;
assign addr[16517]= -470399716;
assign addr[16518]= -763158411;
assign addr[16519]= -1040451659;
assign addr[16520]= -1296660098;
assign addr[16521]= -1526591649;
assign addr[16522]= -1725586737;
assign addr[16523]= -1889612716;
assign addr[16524]= -2015345591;
assign addr[16525]= -2100237377;
assign addr[16526]= -2142567738;
assign addr[16527]= -2141478848;
assign addr[16528]= -2096992772;
assign addr[16529]= -2010011024;
assign addr[16530]= -1882296293;
assign addr[16531]= -1716436725;
assign addr[16532]= -1515793473;
assign addr[16533]= -1284432584;
assign addr[16534]= -1027042599;
assign addr[16535]= -748839539;
assign addr[16536]= -455461206;
assign addr[16537]= -152852926;
assign addr[16538]= 152852926;
assign addr[16539]= 455461206;
assign addr[16540]= 748839539;
assign addr[16541]= 1027042599;
assign addr[16542]= 1284432584;
assign addr[16543]= 1515793473;
assign addr[16544]= 1716436725;
assign addr[16545]= 1882296293;
assign addr[16546]= 2010011024;
assign addr[16547]= 2096992772;
assign addr[16548]= 2141478848;
assign addr[16549]= 2142567738;
assign addr[16550]= 2100237377;
assign addr[16551]= 2015345591;
assign addr[16552]= 1889612716;
assign addr[16553]= 1725586737;
assign addr[16554]= 1526591649;
assign addr[16555]= 1296660098;
assign addr[16556]= 1040451659;
assign addr[16557]= 763158411;
assign addr[16558]= 470399716;
assign addr[16559]= 168108346;
assign addr[16560]= -137589750;
assign addr[16561]= -440499581;
assign addr[16562]= -734482665;
assign addr[16563]= -1013581418;
assign addr[16564]= -1272139887;
assign addr[16565]= -1504918373;
assign addr[16566]= -1707199606;
assign addr[16567]= -1874884346;
assign addr[16568]= -2004574453;
assign addr[16569]= -2093641749;
assign addr[16570]= -2140281282;
assign addr[16571]= -2143547897;
assign addr[16572]= -2103375398;
assign addr[16573]= -2020577882;
assign addr[16574]= -1896833245;
assign addr[16575]= -1734649179;
assign addr[16576]= -1537312353;
assign addr[16577]= -1308821808;
assign addr[16578]= -1053807919;
assign addr[16579]= -777438554;
assign addr[16580]= -485314355;
assign addr[16581]= -183355234;
assign addr[16582]= 122319591;
assign addr[16583]= 425515602;
assign addr[16584]= 720088517;
assign addr[16585]= 1000068799;
assign addr[16586]= 1259782632;
assign addr[16587]= 1493966902;
assign addr[16588]= 1697875851;
assign addr[16589]= 1867377253;
assign addr[16590]= 1999036154;
assign addr[16591]= 2090184478;
assign addr[16592]= 2138975100;
assign addr[16593]= 2144419275;
assign addr[16594]= 2106406677;
assign addr[16595]= 2025707632;
assign addr[16596]= 1903957513;
assign addr[16597]= 1743623590;
assign addr[16598]= 1547955041;
assign addr[16599]= 1320917099;
assign addr[16600]= 1067110699;
assign addr[16601]= 791679244;
assign addr[16602]= 500204365;
assign addr[16603]= 198592817;
assign addr[16604]= -107043224;
assign addr[16605]= -410510029;
assign addr[16606]= -705657826;
assign addr[16607]= -986505429;
assign addr[16608]= -1247361445;
assign addr[16609]= -1482939614;
assign addr[16610]= -1688465931;
assign addr[16611]= -1859775393;
assign addr[16612]= -1993396407;
assign addr[16613]= -2086621133;
assign addr[16614]= -2137560369;
assign addr[16615]= -2145181827;
assign addr[16616]= -2109331059;
assign addr[16617]= -2030734582;
assign addr[16618]= -1910985158;
assign addr[16619]= -1752509516;
assign addr[16620]= -1558519173;
assign addr[16621]= -1332945355;
assign addr[16622]= -1080359326;
assign addr[16623]= -805879757;
assign addr[16624]= -515068990;
assign addr[16625]= -213820322;
assign addr[16626]= 91761426;
assign addr[16627]= 395483624;
assign addr[16628]= 691191324;
assign addr[16629]= 972891995;
assign addr[16630]= 1234876957;
assign addr[16631]= 1471837070;
assign addr[16632]= 1678970324;
assign addr[16633]= 1852079154;
assign addr[16634]= 1987655498;
assign addr[16635]= 2082951896;
assign addr[16636]= 2136037160;
assign addr[16637]= 2145835515;
assign addr[16638]= 2112148396;
assign addr[16639]= 2035658475;
assign addr[16640]= 1917915825;
assign addr[16641]= 1761306505;
assign addr[16642]= 1569004214;
assign addr[16643]= 1344905966;
assign addr[16644]= 1093553126;
assign addr[16645]= 820039373;
assign addr[16646]= 529907477;
assign addr[16647]= 229036977;
assign addr[16648]= -76474970;
assign addr[16649]= -380437148;
assign addr[16650]= -676689746;
assign addr[16651]= -959229189;
assign addr[16652]= -1222329801;
assign addr[16653]= -1460659832;
assign addr[16654]= -1669389513;
assign addr[16655]= -1844288924;
assign addr[16656]= -1981813720;
assign addr[16657]= -2079176953;
assign addr[16658]= -2134405552;
assign addr[16659]= -2146380306;
assign addr[16660]= -2114858546;
assign addr[16661]= -2040479063;
assign addr[16662]= -1924749160;
assign addr[16663]= -1770014111;
assign addr[16664]= -1579409630;
assign addr[16665]= -1356798326;
assign addr[16666]= -1106691431;
assign addr[16667]= -834157373;
assign addr[16668]= -544719071;
assign addr[16669]= -244242007;
assign addr[16670]= 61184634;
assign addr[16671]= 365371365;
assign addr[16672]= 662153826;
assign addr[16673]= 945517704;
assign addr[16674]= 1209720613;
assign addr[16675]= 1449408469;
assign addr[16676]= 1659723983;
assign addr[16677]= 1836405100;
assign addr[16678]= 1975871368;
assign addr[16679]= 2075296495;
assign addr[16680]= 2132665626;
assign addr[16681]= 2146816171;
assign addr[16682]= 2117461370;
assign addr[16683]= 2045196100;
assign addr[16684]= 1931484818;
assign addr[16685]= 1778631892;
assign addr[16686]= 1589734894;
assign addr[16687]= 1368621831;
assign addr[16688]= 1119773573;
assign addr[16689]= 848233042;
assign addr[16690]= 559503022;
assign addr[16691]= 259434643;
assign addr[16692]= -45891193;
assign addr[16693]= -350287041;
assign addr[16694]= -647584304;
assign addr[16695]= -931758235;
assign addr[16696]= -1197050035;
assign addr[16697]= -1438083551;
assign addr[16698]= -1649974225;
assign addr[16699]= -1828428082;
assign addr[16700]= -1969828744;
assign addr[16701]= -2071310720;
assign addr[16702]= -2130817471;
assign addr[16703]= -2147143090;
assign addr[16704]= -2119956737;
assign addr[16705]= -2049809346;
assign addr[16706]= -1938122457;
assign addr[16707]= -1787159411;
assign addr[16708]= -1599979481;
assign addr[16709]= -1380375881;
assign addr[16710]= -1132798888;
assign addr[16711]= -862265664;
assign addr[16712]= -574258580;
assign addr[16713]= -274614114;
assign addr[16714]= 30595422;
assign addr[16715]= 335184940;
assign addr[16716]= 632981917;
assign addr[16717]= 917951481;
assign addr[16718]= 1184318708;
assign addr[16719]= 1426685652;
assign addr[16720]= 1640140734;
assign addr[16721]= 1820358275;
assign addr[16722]= 1963686155;
assign addr[16723]= 2067219829;
assign addr[16724]= 2128861181;
assign addr[16725]= 2147361045;
assign addr[16726]= 2122344521;
assign addr[16727]= 2054318569;
assign addr[16728]= 1944661739;
assign addr[16729]= 1795596234;
assign addr[16730]= 1610142873;
assign addr[16731]= 1392059879;
assign addr[16732]= 1145766716;
assign addr[16733]= 876254528;
assign addr[16734]= 588984994;
assign addr[16735]= 289779648;
assign addr[16736]= -15298099;
assign addr[16737]= -320065829;
assign addr[16738]= -618347408;
assign addr[16739]= -904098143;
assign addr[16740]= -1171527280;
assign addr[16741]= -1415215352;
assign addr[16742]= -1630224009;
assign addr[16743]= -1812196087;
assign addr[16744]= -1957443913;
assign addr[16745]= -2063024031;
assign addr[16746]= -2126796855;
assign addr[16747]= -2147470025;
assign addr[16748]= -2124624598;
assign addr[16749]= -2058723538;
assign addr[16750]= -1951102334;
assign addr[16751]= -1803941934;
assign addr[16752]= -1620224553;
assign addr[16753]= -1403673233;
assign addr[16754]= -1158676398;
assign addr[16755]= -890198924;
assign addr[16756]= -603681519;
assign addr[16757]= -304930476;
assign addr[16758]= 0;
assign addr[16759]= 304930476;
assign addr[16760]= 603681519;
assign addr[16761]= 890198924;
assign addr[16762]= 1158676398;
assign addr[16763]= 1403673233;
assign addr[16764]= 1620224553;
assign addr[16765]= 1803941934;
assign addr[16766]= 1951102334;
assign addr[16767]= 2058723538;
assign addr[16768]= 2124624598;
assign addr[16769]= 2147470025;
assign addr[16770]= 2126796855;
assign addr[16771]= 2063024031;
assign addr[16772]= 1957443913;
assign addr[16773]= 1812196087;
assign addr[16774]= 1630224009;
assign addr[16775]= 1415215352;
assign addr[16776]= 1171527280;
assign addr[16777]= 904098143;
assign addr[16778]= 618347408;
assign addr[16779]= 320065829;
assign addr[16780]= 15298099;
assign addr[16781]= -289779648;
assign addr[16782]= -588984994;
assign addr[16783]= -876254528;
assign addr[16784]= -1145766716;
assign addr[16785]= -1392059879;
assign addr[16786]= -1610142873;
assign addr[16787]= -1795596234;
assign addr[16788]= -1944661739;
assign addr[16789]= -2054318569;
assign addr[16790]= -2122344521;
assign addr[16791]= -2147361045;
assign addr[16792]= -2128861181;
assign addr[16793]= -2067219829;
assign addr[16794]= -1963686155;
assign addr[16795]= -1820358275;
assign addr[16796]= -1640140734;
assign addr[16797]= -1426685652;
assign addr[16798]= -1184318708;
assign addr[16799]= -917951481;
assign addr[16800]= -632981917;
assign addr[16801]= -335184940;
assign addr[16802]= -30595422;
assign addr[16803]= 274614114;
assign addr[16804]= 574258580;
assign addr[16805]= 862265664;
assign addr[16806]= 1132798888;
assign addr[16807]= 1380375881;
assign addr[16808]= 1599979481;
assign addr[16809]= 1787159411;
assign addr[16810]= 1938122457;
assign addr[16811]= 2049809346;
assign addr[16812]= 2119956737;
assign addr[16813]= 2147143090;
assign addr[16814]= 2130817471;
assign addr[16815]= 2071310720;
assign addr[16816]= 1969828744;
assign addr[16817]= 1828428082;
assign addr[16818]= 1649974225;
assign addr[16819]= 1438083551;
assign addr[16820]= 1197050035;
assign addr[16821]= 931758235;
assign addr[16822]= 647584304;
assign addr[16823]= 350287041;
assign addr[16824]= 45891193;
assign addr[16825]= -259434643;
assign addr[16826]= -559503022;
assign addr[16827]= -848233042;
assign addr[16828]= -1119773573;
assign addr[16829]= -1368621831;
assign addr[16830]= -1589734894;
assign addr[16831]= -1778631892;
assign addr[16832]= -1931484818;
assign addr[16833]= -2045196100;
assign addr[16834]= -2117461370;
assign addr[16835]= -2146816171;
assign addr[16836]= -2132665626;
assign addr[16837]= -2075296495;
assign addr[16838]= -1975871368;
assign addr[16839]= -1836405100;
assign addr[16840]= -1659723983;
assign addr[16841]= -1449408469;
assign addr[16842]= -1209720613;
assign addr[16843]= -945517704;
assign addr[16844]= -662153826;
assign addr[16845]= -365371365;
assign addr[16846]= -61184634;
assign addr[16847]= 244242007;
assign addr[16848]= 544719071;
assign addr[16849]= 834157373;
assign addr[16850]= 1106691431;
assign addr[16851]= 1356798326;
assign addr[16852]= 1579409630;
assign addr[16853]= 1770014111;
assign addr[16854]= 1924749160;
assign addr[16855]= 2040479063;
assign addr[16856]= 2114858546;
assign addr[16857]= 2146380306;
assign addr[16858]= 2134405552;
assign addr[16859]= 2079176953;
assign addr[16860]= 1981813720;
assign addr[16861]= 1844288924;
assign addr[16862]= 1669389513;
assign addr[16863]= 1460659832;
assign addr[16864]= 1222329801;
assign addr[16865]= 959229189;
assign addr[16866]= 676689746;
assign addr[16867]= 380437148;
assign addr[16868]= 76474970;
assign addr[16869]= -229036977;
assign addr[16870]= -529907477;
assign addr[16871]= -820039373;
assign addr[16872]= -1093553126;
assign addr[16873]= -1344905966;
assign addr[16874]= -1569004214;
assign addr[16875]= -1761306505;
assign addr[16876]= -1917915825;
assign addr[16877]= -2035658475;
assign addr[16878]= -2112148396;
assign addr[16879]= -2145835515;
assign addr[16880]= -2136037160;
assign addr[16881]= -2082951896;
assign addr[16882]= -1987655498;
assign addr[16883]= -1852079154;
assign addr[16884]= -1678970324;
assign addr[16885]= -1471837070;
assign addr[16886]= -1234876957;
assign addr[16887]= -972891995;
assign addr[16888]= -691191324;
assign addr[16889]= -395483624;
assign addr[16890]= -91761426;
assign addr[16891]= 213820322;
assign addr[16892]= 515068990;
assign addr[16893]= 805879757;
assign addr[16894]= 1080359326;
assign addr[16895]= 1332945355;
assign addr[16896]= 1558519173;
assign addr[16897]= 1752509516;
assign addr[16898]= 1910985158;
assign addr[16899]= 2030734582;
assign addr[16900]= 2109331059;
assign addr[16901]= 2145181827;
assign addr[16902]= 2137560369;
assign addr[16903]= 2086621133;
assign addr[16904]= 1993396407;
assign addr[16905]= 1859775393;
assign addr[16906]= 1688465931;
assign addr[16907]= 1482939614;
assign addr[16908]= 1247361445;
assign addr[16909]= 986505429;
assign addr[16910]= 705657826;
assign addr[16911]= 410510029;
assign addr[16912]= 107043224;
assign addr[16913]= -198592817;
assign addr[16914]= -500204365;
assign addr[16915]= -791679244;
assign addr[16916]= -1067110699;
assign addr[16917]= -1320917099;
assign addr[16918]= -1547955041;
assign addr[16919]= -1743623590;
assign addr[16920]= -1903957513;
assign addr[16921]= -2025707632;
assign addr[16922]= -2106406677;
assign addr[16923]= -2144419275;
assign addr[16924]= -2138975100;
assign addr[16925]= -2090184478;
assign addr[16926]= -1999036154;
assign addr[16927]= -1867377253;
assign addr[16928]= -1697875851;
assign addr[16929]= -1493966902;
assign addr[16930]= -1259782632;
assign addr[16931]= -1000068799;
assign addr[16932]= -720088517;
assign addr[16933]= -425515602;
assign addr[16934]= -122319591;
assign addr[16935]= 183355234;
assign addr[16936]= 485314355;
assign addr[16937]= 777438554;
assign addr[16938]= 1053807919;
assign addr[16939]= 1308821808;
assign addr[16940]= 1537312353;
assign addr[16941]= 1734649179;
assign addr[16942]= 1896833245;
assign addr[16943]= 2020577882;
assign addr[16944]= 2103375398;
assign addr[16945]= 2143547897;
assign addr[16946]= 2140281282;
assign addr[16947]= 2093641749;
assign addr[16948]= 2004574453;
assign addr[16949]= 1874884346;
assign addr[16950]= 1707199606;
assign addr[16951]= 1504918373;
assign addr[16952]= 1272139887;
assign addr[16953]= 1013581418;
assign addr[16954]= 734482665;
assign addr[16955]= 440499581;
assign addr[16956]= 137589750;
assign addr[16957]= -168108346;
assign addr[16958]= -470399716;
assign addr[16959]= -763158411;
assign addr[16960]= -1040451659;
assign addr[16961]= -1296660098;
assign addr[16962]= -1526591649;
assign addr[16963]= -1725586737;
assign addr[16964]= -1889612716;
assign addr[16965]= -2015345591;
assign addr[16966]= -2100237377;
assign addr[16967]= -2142567738;
assign addr[16968]= -2141478848;
assign addr[16969]= -2096992772;
assign addr[16970]= -2010011024;
assign addr[16971]= -1882296293;
assign addr[16972]= -1716436725;
assign addr[16973]= -1515793473;
assign addr[16974]= -1284432584;
assign addr[16975]= -1027042599;
assign addr[16976]= -748839539;
assign addr[16977]= -455461206;
assign addr[16978]= -152852926;
assign addr[16979]= 152852926;
assign addr[16980]= 455461206;
assign addr[16981]= 748839539;
assign addr[16982]= 1027042599;
assign addr[16983]= 1284432584;
assign addr[16984]= 1515793473;
assign addr[16985]= 1716436725;
assign addr[16986]= 1882296293;
assign addr[16987]= 2010011024;
assign addr[16988]= 2096992772;
assign addr[16989]= 2141478848;
assign addr[16990]= 2142567738;
assign addr[16991]= 2100237377;
assign addr[16992]= 2015345591;
assign addr[16993]= 1889612716;
assign addr[16994]= 1725586737;
assign addr[16995]= 1526591649;
assign addr[16996]= 1296660098;
assign addr[16997]= 1040451659;
assign addr[16998]= 763158411;
assign addr[16999]= 470399716;
assign addr[17000]= 168108346;
assign addr[17001]= -137589750;
assign addr[17002]= -440499581;
assign addr[17003]= -734482665;
assign addr[17004]= -1013581418;
assign addr[17005]= -1272139887;
assign addr[17006]= -1504918373;
assign addr[17007]= -1707199606;
assign addr[17008]= -1874884346;
assign addr[17009]= -2004574453;
assign addr[17010]= -2093641749;
assign addr[17011]= -2140281282;
assign addr[17012]= -2143547897;
assign addr[17013]= -2103375398;
assign addr[17014]= -2020577882;
assign addr[17015]= -1896833245;
assign addr[17016]= -1734649179;
assign addr[17017]= -1537312353;
assign addr[17018]= -1308821808;
assign addr[17019]= -1053807919;
assign addr[17020]= -777438554;
assign addr[17021]= -485314355;
assign addr[17022]= -183355234;
assign addr[17023]= 122319591;
assign addr[17024]= 425515602;
assign addr[17025]= 720088517;
assign addr[17026]= 1000068799;
assign addr[17027]= 1259782632;
assign addr[17028]= 1493966902;
assign addr[17029]= 1697875851;
assign addr[17030]= 1867377253;
assign addr[17031]= 1999036154;
assign addr[17032]= 2090184478;
assign addr[17033]= 2138975100;
assign addr[17034]= 2144419275;
assign addr[17035]= 2106406677;
assign addr[17036]= 2025707632;
assign addr[17037]= 1903957513;
assign addr[17038]= 1743623590;
assign addr[17039]= 1547955041;
assign addr[17040]= 1320917099;
assign addr[17041]= 1067110699;
assign addr[17042]= 791679244;
assign addr[17043]= 500204365;
assign addr[17044]= 198592817;
assign addr[17045]= -107043224;
assign addr[17046]= -410510029;
assign addr[17047]= -705657826;
assign addr[17048]= -986505429;
assign addr[17049]= -1247361445;
assign addr[17050]= -1482939614;
assign addr[17051]= -1688465931;
assign addr[17052]= -1859775393;
assign addr[17053]= -1993396407;
assign addr[17054]= -2086621133;
assign addr[17055]= -2137560369;
assign addr[17056]= -2145181827;
assign addr[17057]= -2109331059;
assign addr[17058]= -2030734582;
assign addr[17059]= -1910985158;
assign addr[17060]= -1752509516;
assign addr[17061]= -1558519173;
assign addr[17062]= -1332945355;
assign addr[17063]= -1080359326;
assign addr[17064]= -805879757;
assign addr[17065]= -515068990;
assign addr[17066]= -213820322;
assign addr[17067]= 91761426;
assign addr[17068]= 395483624;
assign addr[17069]= 691191324;
assign addr[17070]= 972891995;
assign addr[17071]= 1234876957;
assign addr[17072]= 1471837070;
assign addr[17073]= 1678970324;
assign addr[17074]= 1852079154;
assign addr[17075]= 1987655498;
assign addr[17076]= 2082951896;
assign addr[17077]= 2136037160;
assign addr[17078]= 2145835515;
assign addr[17079]= 2112148396;
assign addr[17080]= 2035658475;
assign addr[17081]= 1917915825;
assign addr[17082]= 1761306505;
assign addr[17083]= 1569004214;
assign addr[17084]= 1344905966;
assign addr[17085]= 1093553126;
assign addr[17086]= 820039373;
assign addr[17087]= 529907477;
assign addr[17088]= 229036977;
assign addr[17089]= -76474970;
assign addr[17090]= -380437148;
assign addr[17091]= -676689746;
assign addr[17092]= -959229189;
assign addr[17093]= -1222329801;
assign addr[17094]= -1460659832;
assign addr[17095]= -1669389513;
assign addr[17096]= -1844288924;
assign addr[17097]= -1981813720;
assign addr[17098]= -2079176953;
assign addr[17099]= -2134405552;
assign addr[17100]= -2146380306;
assign addr[17101]= -2114858546;
assign addr[17102]= -2040479063;
assign addr[17103]= -1924749160;
assign addr[17104]= -1770014111;
assign addr[17105]= -1579409630;
assign addr[17106]= -1356798326;
assign addr[17107]= -1106691431;
assign addr[17108]= -834157373;
assign addr[17109]= -544719071;
assign addr[17110]= -244242007;
assign addr[17111]= 61184634;
assign addr[17112]= 365371365;
assign addr[17113]= 662153826;
assign addr[17114]= 945517704;
assign addr[17115]= 1209720613;
assign addr[17116]= 1449408469;
assign addr[17117]= 1659723983;
assign addr[17118]= 1836405100;
assign addr[17119]= 1975871368;
assign addr[17120]= 2075296495;
assign addr[17121]= 2132665626;
assign addr[17122]= 2146816171;
assign addr[17123]= 2117461370;
assign addr[17124]= 2045196100;
assign addr[17125]= 1931484818;
assign addr[17126]= 1778631892;
assign addr[17127]= 1589734894;
assign addr[17128]= 1368621831;
assign addr[17129]= 1119773573;
assign addr[17130]= 848233042;
assign addr[17131]= 559503022;
assign addr[17132]= 259434643;
assign addr[17133]= -45891193;
assign addr[17134]= -350287041;
assign addr[17135]= -647584304;
assign addr[17136]= -931758235;
assign addr[17137]= -1197050035;
assign addr[17138]= -1438083551;
assign addr[17139]= -1649974225;
assign addr[17140]= -1828428082;
assign addr[17141]= -1969828744;
assign addr[17142]= -2071310720;
assign addr[17143]= -2130817471;
assign addr[17144]= -2147143090;
assign addr[17145]= -2119956737;
assign addr[17146]= -2049809346;
assign addr[17147]= -1938122457;
assign addr[17148]= -1787159411;
assign addr[17149]= -1599979481;
assign addr[17150]= -1380375881;
assign addr[17151]= -1132798888;
assign addr[17152]= -862265664;
assign addr[17153]= -574258580;
assign addr[17154]= -274614114;
assign addr[17155]= 30595422;
assign addr[17156]= 335184940;
assign addr[17157]= 632981917;
assign addr[17158]= 917951481;
assign addr[17159]= 1184318708;
assign addr[17160]= 1426685652;
assign addr[17161]= 1640140734;
assign addr[17162]= 1820358275;
assign addr[17163]= 1963686155;
assign addr[17164]= 2067219829;
assign addr[17165]= 2128861181;
assign addr[17166]= 2147361045;
assign addr[17167]= 2122344521;
assign addr[17168]= 2054318569;
assign addr[17169]= 1944661739;
assign addr[17170]= 1795596234;
assign addr[17171]= 1610142873;
assign addr[17172]= 1392059879;
assign addr[17173]= 1145766716;
assign addr[17174]= 876254528;
assign addr[17175]= 588984994;
assign addr[17176]= 289779648;
assign addr[17177]= -15298099;
assign addr[17178]= -320065829;
assign addr[17179]= -618347408;
assign addr[17180]= -904098143;
assign addr[17181]= -1171527280;
assign addr[17182]= -1415215352;
assign addr[17183]= -1630224009;
assign addr[17184]= -1812196087;
assign addr[17185]= -1957443913;
assign addr[17186]= -2063024031;
assign addr[17187]= -2126796855;
assign addr[17188]= -2147470025;
assign addr[17189]= -2124624598;
assign addr[17190]= -2058723538;
assign addr[17191]= -1951102334;
assign addr[17192]= -1803941934;
assign addr[17193]= -1620224553;
assign addr[17194]= -1403673233;
assign addr[17195]= -1158676398;
assign addr[17196]= -890198924;
assign addr[17197]= -603681519;
assign addr[17198]= -304930476;
assign addr[17199]= 0;
assign addr[17200]= 304930476;
assign addr[17201]= 603681519;
assign addr[17202]= 890198924;
assign addr[17203]= 1158676398;
assign addr[17204]= 1403673233;
assign addr[17205]= 1620224553;
assign addr[17206]= 1803941934;
assign addr[17207]= 1951102334;
assign addr[17208]= 2058723538;
assign addr[17209]= 2124624598;
assign addr[17210]= 2147470025;
assign addr[17211]= 2126796855;
assign addr[17212]= 2063024031;
assign addr[17213]= 1957443913;
assign addr[17214]= 1812196087;
assign addr[17215]= 1630224009;
assign addr[17216]= 1415215352;
assign addr[17217]= 1171527280;
assign addr[17218]= 904098143;
assign addr[17219]= 618347408;
assign addr[17220]= 320065829;
assign addr[17221]= 15298099;
assign addr[17222]= -289779648;
assign addr[17223]= -588984994;
assign addr[17224]= -876254528;
assign addr[17225]= -1145766716;
assign addr[17226]= -1392059879;
assign addr[17227]= -1610142873;
assign addr[17228]= -1795596234;
assign addr[17229]= -1944661739;
assign addr[17230]= -2054318569;
assign addr[17231]= -2122344521;
assign addr[17232]= -2147361045;
assign addr[17233]= -2128861181;
assign addr[17234]= -2067219829;
assign addr[17235]= -1963686155;
assign addr[17236]= -1820358275;
assign addr[17237]= -1640140734;
assign addr[17238]= -1426685652;
assign addr[17239]= -1184318708;
assign addr[17240]= -917951481;
assign addr[17241]= -632981917;
assign addr[17242]= -335184940;
assign addr[17243]= -30595422;
assign addr[17244]= 274614114;
assign addr[17245]= 574258580;
assign addr[17246]= 862265664;
assign addr[17247]= 1132798888;
assign addr[17248]= 1380375881;
assign addr[17249]= 1599979481;
assign addr[17250]= 1787159411;
assign addr[17251]= 1938122457;
assign addr[17252]= 2049809346;
assign addr[17253]= 2119956737;
assign addr[17254]= 2147143090;
assign addr[17255]= 2130817471;
assign addr[17256]= 2071310720;
assign addr[17257]= 1969828744;
assign addr[17258]= 1828428082;
assign addr[17259]= 1649974225;
assign addr[17260]= 1438083551;
assign addr[17261]= 1197050035;
assign addr[17262]= 931758235;
assign addr[17263]= 647584304;
assign addr[17264]= 350287041;
assign addr[17265]= 45891193;
assign addr[17266]= -259434643;
assign addr[17267]= -559503022;
assign addr[17268]= -848233042;
assign addr[17269]= -1119773573;
assign addr[17270]= -1368621831;
assign addr[17271]= -1589734894;
assign addr[17272]= -1778631892;
assign addr[17273]= -1931484818;
assign addr[17274]= -2045196100;
assign addr[17275]= -2117461370;
assign addr[17276]= -2146816171;
assign addr[17277]= -2132665626;
assign addr[17278]= -2075296495;
assign addr[17279]= -1975871368;
assign addr[17280]= -1836405100;
assign addr[17281]= -1659723983;
assign addr[17282]= -1449408469;
assign addr[17283]= -1209720613;
assign addr[17284]= -945517704;
assign addr[17285]= -662153826;
assign addr[17286]= -365371365;
assign addr[17287]= -61184634;
assign addr[17288]= 244242007;
assign addr[17289]= 544719071;
assign addr[17290]= 834157373;
assign addr[17291]= 1106691431;
assign addr[17292]= 1356798326;
assign addr[17293]= 1579409630;
assign addr[17294]= 1770014111;
assign addr[17295]= 1924749160;
assign addr[17296]= 2040479063;
assign addr[17297]= 2114858546;
assign addr[17298]= 2146380306;
assign addr[17299]= 2134405552;
assign addr[17300]= 2079176953;
assign addr[17301]= 1981813720;
assign addr[17302]= 1844288924;
assign addr[17303]= 1669389513;
assign addr[17304]= 1460659832;
assign addr[17305]= 1222329801;
assign addr[17306]= 959229189;
assign addr[17307]= 676689746;
assign addr[17308]= 380437148;
assign addr[17309]= 76474970;
assign addr[17310]= -229036977;
assign addr[17311]= -529907477;
assign addr[17312]= -820039373;
assign addr[17313]= -1093553126;
assign addr[17314]= -1344905966;
assign addr[17315]= -1569004214;
assign addr[17316]= -1761306505;
assign addr[17317]= -1917915825;
assign addr[17318]= -2035658475;
assign addr[17319]= -2112148396;
assign addr[17320]= -2145835515;
assign addr[17321]= -2136037160;
assign addr[17322]= -2082951896;
assign addr[17323]= -1987655498;
assign addr[17324]= -1852079154;
assign addr[17325]= -1678970324;
assign addr[17326]= -1471837070;
assign addr[17327]= -1234876957;
assign addr[17328]= -972891995;
assign addr[17329]= -691191324;
assign addr[17330]= -395483624;
assign addr[17331]= -91761426;
assign addr[17332]= 213820322;
assign addr[17333]= 515068990;
assign addr[17334]= 805879757;
assign addr[17335]= 1080359326;
assign addr[17336]= 1332945355;
assign addr[17337]= 1558519173;
assign addr[17338]= 1752509516;
assign addr[17339]= 1910985158;
assign addr[17340]= 2030734582;
assign addr[17341]= 2109331059;
assign addr[17342]= 2145181827;
assign addr[17343]= 2137560369;
assign addr[17344]= 2086621133;
assign addr[17345]= 1993396407;
assign addr[17346]= 1859775393;
assign addr[17347]= 1688465931;
assign addr[17348]= 1482939614;
assign addr[17349]= 1247361445;
assign addr[17350]= 986505429;
assign addr[17351]= 705657826;
assign addr[17352]= 410510029;
assign addr[17353]= 107043224;
assign addr[17354]= -198592817;
assign addr[17355]= -500204365;
assign addr[17356]= -791679244;
assign addr[17357]= -1067110699;
assign addr[17358]= -1320917099;
assign addr[17359]= -1547955041;
assign addr[17360]= -1743623590;
assign addr[17361]= -1903957513;
assign addr[17362]= -2025707632;
assign addr[17363]= -2106406677;
assign addr[17364]= -2144419275;
assign addr[17365]= -2138975100;
assign addr[17366]= -2090184478;
assign addr[17367]= -1999036154;
assign addr[17368]= -1867377253;
assign addr[17369]= -1697875851;
assign addr[17370]= -1493966902;
assign addr[17371]= -1259782632;
assign addr[17372]= -1000068799;
assign addr[17373]= -720088517;
assign addr[17374]= -425515602;
assign addr[17375]= -122319591;
assign addr[17376]= 183355234;
assign addr[17377]= 485314355;
assign addr[17378]= 777438554;
assign addr[17379]= 1053807919;
assign addr[17380]= 1308821808;
assign addr[17381]= 1537312353;
assign addr[17382]= 1734649179;
assign addr[17383]= 1896833245;
assign addr[17384]= 2020577882;
assign addr[17385]= 2103375398;
assign addr[17386]= 2143547897;
assign addr[17387]= 2140281282;
assign addr[17388]= 2093641749;
assign addr[17389]= 2004574453;
assign addr[17390]= 1874884346;
assign addr[17391]= 1707199606;
assign addr[17392]= 1504918373;
assign addr[17393]= 1272139887;
assign addr[17394]= 1013581418;
assign addr[17395]= 734482665;
assign addr[17396]= 440499581;
assign addr[17397]= 137589750;
assign addr[17398]= -168108346;
assign addr[17399]= -470399716;
assign addr[17400]= -763158411;
assign addr[17401]= -1040451659;
assign addr[17402]= -1296660098;
assign addr[17403]= -1526591649;
assign addr[17404]= -1725586737;
assign addr[17405]= -1889612716;
assign addr[17406]= -2015345591;
assign addr[17407]= -2100237377;
assign addr[17408]= -2142567738;
assign addr[17409]= -2141478848;
assign addr[17410]= -2096992772;
assign addr[17411]= -2010011024;
assign addr[17412]= -1882296293;
assign addr[17413]= -1716436725;
assign addr[17414]= -1515793473;
assign addr[17415]= -1284432584;
assign addr[17416]= -1027042599;
assign addr[17417]= -748839539;
assign addr[17418]= -455461206;
assign addr[17419]= -152852926;
assign addr[17420]= 152852926;
assign addr[17421]= 455461206;
assign addr[17422]= 748839539;
assign addr[17423]= 1027042599;
assign addr[17424]= 1284432584;
assign addr[17425]= 1515793473;
assign addr[17426]= 1716436725;
assign addr[17427]= 1882296293;
assign addr[17428]= 2010011024;
assign addr[17429]= 2096992772;
assign addr[17430]= 2141478848;
assign addr[17431]= 2142567738;
assign addr[17432]= 2100237377;
assign addr[17433]= 2015345591;
assign addr[17434]= 1889612716;
assign addr[17435]= 1725586737;
assign addr[17436]= 1526591649;
assign addr[17437]= 1296660098;
assign addr[17438]= 1040451659;
assign addr[17439]= 763158411;
assign addr[17440]= 470399716;
assign addr[17441]= 168108346;
assign addr[17442]= -137589750;
assign addr[17443]= -440499581;
assign addr[17444]= -734482665;
assign addr[17445]= -1013581418;
assign addr[17446]= -1272139887;
assign addr[17447]= -1504918373;
assign addr[17448]= -1707199606;
assign addr[17449]= -1874884346;
assign addr[17450]= -2004574453;
assign addr[17451]= -2093641749;
assign addr[17452]= -2140281282;
assign addr[17453]= -2143547897;
assign addr[17454]= -2103375398;
assign addr[17455]= -2020577882;
assign addr[17456]= -1896833245;
assign addr[17457]= -1734649179;
assign addr[17458]= -1537312353;
assign addr[17459]= -1308821808;
assign addr[17460]= -1053807919;
assign addr[17461]= -777438554;
assign addr[17462]= -485314355;
assign addr[17463]= -183355234;
assign addr[17464]= 122319591;
assign addr[17465]= 425515602;
assign addr[17466]= 720088517;
assign addr[17467]= 1000068799;
assign addr[17468]= 1259782632;
assign addr[17469]= 1493966902;
assign addr[17470]= 1697875851;
assign addr[17471]= 1867377253;
assign addr[17472]= 1999036154;
assign addr[17473]= 2090184478;
assign addr[17474]= 2138975100;
assign addr[17475]= 2144419275;
assign addr[17476]= 2106406677;
assign addr[17477]= 2025707632;
assign addr[17478]= 1903957513;
assign addr[17479]= 1743623590;
assign addr[17480]= 1547955041;
assign addr[17481]= 1320917099;
assign addr[17482]= 1067110699;
assign addr[17483]= 791679244;
assign addr[17484]= 500204365;
assign addr[17485]= 198592817;
assign addr[17486]= -107043224;
assign addr[17487]= -410510029;
assign addr[17488]= -705657826;
assign addr[17489]= -986505429;
assign addr[17490]= -1247361445;
assign addr[17491]= -1482939614;
assign addr[17492]= -1688465931;
assign addr[17493]= -1859775393;
assign addr[17494]= -1993396407;
assign addr[17495]= -2086621133;
assign addr[17496]= -2137560369;
assign addr[17497]= -2145181827;
assign addr[17498]= -2109331059;
assign addr[17499]= -2030734582;
assign addr[17500]= -1910985158;
assign addr[17501]= -1752509516;
assign addr[17502]= -1558519173;
assign addr[17503]= -1332945355;
assign addr[17504]= -1080359326;
assign addr[17505]= -805879757;
assign addr[17506]= -515068990;
assign addr[17507]= -213820322;
assign addr[17508]= 91761426;
assign addr[17509]= 395483624;
assign addr[17510]= 691191324;
assign addr[17511]= 972891995;
assign addr[17512]= 1234876957;
assign addr[17513]= 1471837070;
assign addr[17514]= 1678970324;
assign addr[17515]= 1852079154;
assign addr[17516]= 1987655498;
assign addr[17517]= 2082951896;
assign addr[17518]= 2136037160;
assign addr[17519]= 2145835515;
assign addr[17520]= 2112148396;
assign addr[17521]= 2035658475;
assign addr[17522]= 1917915825;
assign addr[17523]= 1761306505;
assign addr[17524]= 1569004214;
assign addr[17525]= 1344905966;
assign addr[17526]= 1093553126;
assign addr[17527]= 820039373;
assign addr[17528]= 529907477;
assign addr[17529]= 229036977;
assign addr[17530]= -76474970;
assign addr[17531]= -380437148;
assign addr[17532]= -676689746;
assign addr[17533]= -959229189;
assign addr[17534]= -1222329801;
assign addr[17535]= -1460659832;
assign addr[17536]= -1669389513;
assign addr[17537]= -1844288924;
assign addr[17538]= -1981813720;
assign addr[17539]= -2079176953;
assign addr[17540]= -2134405552;
assign addr[17541]= -2146380306;
assign addr[17542]= -2114858546;
assign addr[17543]= -2040479063;
assign addr[17544]= -1924749160;
assign addr[17545]= -1770014111;
assign addr[17546]= -1579409630;
assign addr[17547]= -1356798326;
assign addr[17548]= -1106691431;
assign addr[17549]= -834157373;
assign addr[17550]= -544719071;
assign addr[17551]= -244242007;
assign addr[17552]= 61184634;
assign addr[17553]= 365371365;
assign addr[17554]= 662153826;
assign addr[17555]= 945517704;
assign addr[17556]= 1209720613;
assign addr[17557]= 1449408469;
assign addr[17558]= 1659723983;
assign addr[17559]= 1836405100;
assign addr[17560]= 1975871368;
assign addr[17561]= 2075296495;
assign addr[17562]= 2132665626;
assign addr[17563]= 2146816171;
assign addr[17564]= 2117461370;
assign addr[17565]= 2045196100;
assign addr[17566]= 1931484818;
assign addr[17567]= 1778631892;
assign addr[17568]= 1589734894;
assign addr[17569]= 1368621831;
assign addr[17570]= 1119773573;
assign addr[17571]= 848233042;
assign addr[17572]= 559503022;
assign addr[17573]= 259434643;
assign addr[17574]= -45891193;
assign addr[17575]= -350287041;
assign addr[17576]= -647584304;
assign addr[17577]= -931758235;
assign addr[17578]= -1197050035;
assign addr[17579]= -1438083551;
assign addr[17580]= -1649974225;
assign addr[17581]= -1828428082;
assign addr[17582]= -1969828744;
assign addr[17583]= -2071310720;
assign addr[17584]= -2130817471;
assign addr[17585]= -2147143090;
assign addr[17586]= -2119956737;
assign addr[17587]= -2049809346;
assign addr[17588]= -1938122457;
assign addr[17589]= -1787159411;
assign addr[17590]= -1599979481;
assign addr[17591]= -1380375881;
assign addr[17592]= -1132798888;
assign addr[17593]= -862265664;
assign addr[17594]= -574258580;
assign addr[17595]= -274614114;
assign addr[17596]= 30595422;
assign addr[17597]= 335184940;
assign addr[17598]= 632981917;
assign addr[17599]= 917951481;
assign addr[17600]= 1184318708;
assign addr[17601]= 1426685652;
assign addr[17602]= 1640140734;
assign addr[17603]= 1820358275;
assign addr[17604]= 1963686155;
assign addr[17605]= 2067219829;
assign addr[17606]= 2128861181;
assign addr[17607]= 2147361045;
assign addr[17608]= 2122344521;
assign addr[17609]= 2054318569;
assign addr[17610]= 1944661739;
assign addr[17611]= 1795596234;
assign addr[17612]= 1610142873;
assign addr[17613]= 1392059879;
assign addr[17614]= 1145766716;
assign addr[17615]= 876254528;
assign addr[17616]= 588984994;
assign addr[17617]= 289779648;
assign addr[17618]= -15298099;
assign addr[17619]= -320065829;
assign addr[17620]= -618347408;
assign addr[17621]= -904098143;
assign addr[17622]= -1171527280;
assign addr[17623]= -1415215352;
assign addr[17624]= -1630224009;
assign addr[17625]= -1812196087;
assign addr[17626]= -1957443913;
assign addr[17627]= -2063024031;
assign addr[17628]= -2126796855;
assign addr[17629]= -2147470025;
assign addr[17630]= -2124624598;
assign addr[17631]= -2058723538;
assign addr[17632]= -1951102334;
assign addr[17633]= -1803941934;
assign addr[17634]= -1620224553;
assign addr[17635]= -1403673233;
assign addr[17636]= -1158676398;
assign addr[17637]= -890198924;
assign addr[17638]= -603681519;
assign addr[17639]= -304930476;
assign addr[17640]= 0;
assign addr[17641]= 304930476;
assign addr[17642]= 603681519;
assign addr[17643]= 890198924;
assign addr[17644]= 1158676398;
assign addr[17645]= 1403673233;
assign addr[17646]= 1620224553;
assign addr[17647]= 1803941934;
assign addr[17648]= 1951102334;
assign addr[17649]= 2058723538;
assign addr[17650]= 2124624598;
assign addr[17651]= 2147470025;
assign addr[17652]= 2126796855;
assign addr[17653]= 2063024031;
assign addr[17654]= 1957443913;
assign addr[17655]= 1812196087;
assign addr[17656]= 1630224009;
assign addr[17657]= 1415215352;
assign addr[17658]= 1171527280;
assign addr[17659]= 904098143;
assign addr[17660]= 618347408;
assign addr[17661]= 320065829;
assign addr[17662]= 15298099;
assign addr[17663]= -289779648;
assign addr[17664]= -588984994;
assign addr[17665]= -876254528;
assign addr[17666]= -1145766716;
assign addr[17667]= -1392059879;
assign addr[17668]= -1610142873;
assign addr[17669]= -1795596234;
assign addr[17670]= -1944661739;
assign addr[17671]= -2054318569;
assign addr[17672]= -2122344521;
assign addr[17673]= -2147361045;
assign addr[17674]= -2128861181;
assign addr[17675]= -2067219829;
assign addr[17676]= -1963686155;
assign addr[17677]= -1820358275;
assign addr[17678]= -1640140734;
assign addr[17679]= -1426685652;
assign addr[17680]= -1184318708;
assign addr[17681]= -917951481;
assign addr[17682]= -632981917;
assign addr[17683]= -335184940;
assign addr[17684]= -30595422;
assign addr[17685]= 274614114;
assign addr[17686]= 574258580;
assign addr[17687]= 862265664;
assign addr[17688]= 1132798888;
assign addr[17689]= 1380375881;
assign addr[17690]= 1599979481;
assign addr[17691]= 1787159411;
assign addr[17692]= 1938122457;
assign addr[17693]= 2049809346;
assign addr[17694]= 2119956737;
assign addr[17695]= 2147143090;
assign addr[17696]= 2130817471;
assign addr[17697]= 2071310720;
assign addr[17698]= 1969828744;
assign addr[17699]= 1828428082;
assign addr[17700]= 1649974225;
assign addr[17701]= 1438083551;
assign addr[17702]= 1197050035;
assign addr[17703]= 931758235;
assign addr[17704]= 647584304;
assign addr[17705]= 350287041;
assign addr[17706]= 45891193;
assign addr[17707]= -259434643;
assign addr[17708]= -559503022;
assign addr[17709]= -848233042;
assign addr[17710]= -1119773573;
assign addr[17711]= -1368621831;
assign addr[17712]= -1589734894;
assign addr[17713]= -1778631892;
assign addr[17714]= -1931484818;
assign addr[17715]= -2045196100;
assign addr[17716]= -2117461370;
assign addr[17717]= -2146816171;
assign addr[17718]= -2132665626;
assign addr[17719]= -2075296495;
assign addr[17720]= -1975871368;
assign addr[17721]= -1836405100;
assign addr[17722]= -1659723983;
assign addr[17723]= -1449408469;
assign addr[17724]= -1209720613;
assign addr[17725]= -945517704;
assign addr[17726]= -662153826;
assign addr[17727]= -365371365;
assign addr[17728]= -61184634;
assign addr[17729]= 244242007;
assign addr[17730]= 544719071;
assign addr[17731]= 834157373;
assign addr[17732]= 1106691431;
assign addr[17733]= 1356798326;
assign addr[17734]= 1579409630;
assign addr[17735]= 1770014111;
assign addr[17736]= 1924749160;
assign addr[17737]= 2040479063;
assign addr[17738]= 2114858546;
assign addr[17739]= 2146380306;
assign addr[17740]= 2134405552;
assign addr[17741]= 2079176953;
assign addr[17742]= 1981813720;
assign addr[17743]= 1844288924;
assign addr[17744]= 1669389513;
assign addr[17745]= 1460659832;
assign addr[17746]= 1222329801;
assign addr[17747]= 959229189;
assign addr[17748]= 676689746;
assign addr[17749]= 380437148;
assign addr[17750]= 76474970;
assign addr[17751]= -229036977;
assign addr[17752]= -529907477;
assign addr[17753]= -820039373;
assign addr[17754]= -1093553126;
assign addr[17755]= -1344905966;
assign addr[17756]= -1569004214;
assign addr[17757]= -1761306505;
assign addr[17758]= -1917915825;
assign addr[17759]= -2035658475;
assign addr[17760]= -2112148396;
assign addr[17761]= -2145835515;
assign addr[17762]= -2136037160;
assign addr[17763]= -2082951896;
assign addr[17764]= -1987655498;
assign addr[17765]= -1852079154;
assign addr[17766]= -1678970324;
assign addr[17767]= -1471837070;
assign addr[17768]= -1234876957;
assign addr[17769]= -972891995;
assign addr[17770]= -691191324;
assign addr[17771]= -395483624;
assign addr[17772]= -91761426;
assign addr[17773]= 213820322;
assign addr[17774]= 515068990;
assign addr[17775]= 805879757;
assign addr[17776]= 1080359326;
assign addr[17777]= 1332945355;
assign addr[17778]= 1558519173;
assign addr[17779]= 1752509516;
assign addr[17780]= 1910985158;
assign addr[17781]= 2030734582;
assign addr[17782]= 2109331059;
assign addr[17783]= 2145181827;
assign addr[17784]= 2137560369;
assign addr[17785]= 2086621133;
assign addr[17786]= 1993396407;
assign addr[17787]= 1859775393;
assign addr[17788]= 1688465931;
assign addr[17789]= 1482939614;
assign addr[17790]= 1247361445;
assign addr[17791]= 986505429;
assign addr[17792]= 705657826;
assign addr[17793]= 410510029;
assign addr[17794]= 107043224;
assign addr[17795]= -198592817;
assign addr[17796]= -500204365;
assign addr[17797]= -791679244;
assign addr[17798]= -1067110699;
assign addr[17799]= -1320917099;
assign addr[17800]= -1547955041;
assign addr[17801]= -1743623590;
assign addr[17802]= -1903957513;
assign addr[17803]= -2025707632;
assign addr[17804]= -2106406677;
assign addr[17805]= -2144419275;
assign addr[17806]= -2138975100;
assign addr[17807]= -2090184478;
assign addr[17808]= -1999036154;
assign addr[17809]= -1867377253;
assign addr[17810]= -1697875851;
assign addr[17811]= -1493966902;
assign addr[17812]= -1259782632;
assign addr[17813]= -1000068799;
assign addr[17814]= -720088517;
assign addr[17815]= -425515602;
assign addr[17816]= -122319591;
assign addr[17817]= 183355234;
assign addr[17818]= 485314355;
assign addr[17819]= 777438554;
assign addr[17820]= 1053807919;
assign addr[17821]= 1308821808;
assign addr[17822]= 1537312353;
assign addr[17823]= 1734649179;
assign addr[17824]= 1896833245;
assign addr[17825]= 2020577882;
assign addr[17826]= 2103375398;
assign addr[17827]= 2143547897;
assign addr[17828]= 2140281282;
assign addr[17829]= 2093641749;
assign addr[17830]= 2004574453;
assign addr[17831]= 1874884346;
assign addr[17832]= 1707199606;
assign addr[17833]= 1504918373;
assign addr[17834]= 1272139887;
assign addr[17835]= 1013581418;
assign addr[17836]= 734482665;
assign addr[17837]= 440499581;
assign addr[17838]= 137589750;
assign addr[17839]= -168108346;
assign addr[17840]= -470399716;
assign addr[17841]= -763158411;
assign addr[17842]= -1040451659;
assign addr[17843]= -1296660098;
assign addr[17844]= -1526591649;
assign addr[17845]= -1725586737;
assign addr[17846]= -1889612716;
assign addr[17847]= -2015345591;
assign addr[17848]= -2100237377;
assign addr[17849]= -2142567738;
assign addr[17850]= -2141478848;
assign addr[17851]= -2096992772;
assign addr[17852]= -2010011024;
assign addr[17853]= -1882296293;
assign addr[17854]= -1716436725;
assign addr[17855]= -1515793473;
assign addr[17856]= -1284432584;
assign addr[17857]= -1027042599;
assign addr[17858]= -748839539;
assign addr[17859]= -455461206;
assign addr[17860]= -152852926;
assign addr[17861]= 152852926;
assign addr[17862]= 455461206;
assign addr[17863]= 748839539;
assign addr[17864]= 1027042599;
assign addr[17865]= 1284432584;
assign addr[17866]= 1515793473;
assign addr[17867]= 1716436725;
assign addr[17868]= 1882296293;
assign addr[17869]= 2010011024;
assign addr[17870]= 2096992772;
assign addr[17871]= 2141478848;
assign addr[17872]= 2142567738;
assign addr[17873]= 2100237377;
assign addr[17874]= 2015345591;
assign addr[17875]= 1889612716;
assign addr[17876]= 1725586737;
assign addr[17877]= 1526591649;
assign addr[17878]= 1296660098;
assign addr[17879]= 1040451659;
assign addr[17880]= 763158411;
assign addr[17881]= 470399716;
assign addr[17882]= 168108346;
assign addr[17883]= -137589750;
assign addr[17884]= -440499581;
assign addr[17885]= -734482665;
assign addr[17886]= -1013581418;
assign addr[17887]= -1272139887;
assign addr[17888]= -1504918373;
assign addr[17889]= -1707199606;
assign addr[17890]= -1874884346;
assign addr[17891]= -2004574453;
assign addr[17892]= -2093641749;
assign addr[17893]= -2140281282;
assign addr[17894]= -2143547897;
assign addr[17895]= -2103375398;
assign addr[17896]= -2020577882;
assign addr[17897]= -1896833245;
assign addr[17898]= -1734649179;
assign addr[17899]= -1537312353;
assign addr[17900]= -1308821808;
assign addr[17901]= -1053807919;
assign addr[17902]= -777438554;
assign addr[17903]= -485314355;
assign addr[17904]= -183355234;
assign addr[17905]= 122319591;
assign addr[17906]= 425515602;
assign addr[17907]= 720088517;
assign addr[17908]= 1000068799;
assign addr[17909]= 1259782632;
assign addr[17910]= 1493966902;
assign addr[17911]= 1697875851;
assign addr[17912]= 1867377253;
assign addr[17913]= 1999036154;
assign addr[17914]= 2090184478;
assign addr[17915]= 2138975100;
assign addr[17916]= 2144419275;
assign addr[17917]= 2106406677;
assign addr[17918]= 2025707632;
assign addr[17919]= 1903957513;
assign addr[17920]= 1743623590;
assign addr[17921]= 1547955041;
assign addr[17922]= 1320917099;
assign addr[17923]= 1067110699;
assign addr[17924]= 791679244;
assign addr[17925]= 500204365;
assign addr[17926]= 198592817;
assign addr[17927]= -107043224;
assign addr[17928]= -410510029;
assign addr[17929]= -705657826;
assign addr[17930]= -986505429;
assign addr[17931]= -1247361445;
assign addr[17932]= -1482939614;
assign addr[17933]= -1688465931;
assign addr[17934]= -1859775393;
assign addr[17935]= -1993396407;
assign addr[17936]= -2086621133;
assign addr[17937]= -2137560369;
assign addr[17938]= -2145181827;
assign addr[17939]= -2109331059;
assign addr[17940]= -2030734582;
assign addr[17941]= -1910985158;
assign addr[17942]= -1752509516;
assign addr[17943]= -1558519173;
assign addr[17944]= -1332945355;
assign addr[17945]= -1080359326;
assign addr[17946]= -805879757;
assign addr[17947]= -515068990;
assign addr[17948]= -213820322;
assign addr[17949]= 91761426;
assign addr[17950]= 395483624;
assign addr[17951]= 691191324;
assign addr[17952]= 972891995;
assign addr[17953]= 1234876957;
assign addr[17954]= 1471837070;
assign addr[17955]= 1678970324;
assign addr[17956]= 1852079154;
assign addr[17957]= 1987655498;
assign addr[17958]= 2082951896;
assign addr[17959]= 2136037160;
assign addr[17960]= 2145835515;
assign addr[17961]= 2112148396;
assign addr[17962]= 2035658475;
assign addr[17963]= 1917915825;
assign addr[17964]= 1761306505;
assign addr[17965]= 1569004214;
assign addr[17966]= 1344905966;
assign addr[17967]= 1093553126;
assign addr[17968]= 820039373;
assign addr[17969]= 529907477;
assign addr[17970]= 229036977;
assign addr[17971]= -76474970;
assign addr[17972]= -380437148;
assign addr[17973]= -676689746;
assign addr[17974]= -959229189;
assign addr[17975]= -1222329801;
assign addr[17976]= -1460659832;
assign addr[17977]= -1669389513;
assign addr[17978]= -1844288924;
assign addr[17979]= -1981813720;
assign addr[17980]= -2079176953;
assign addr[17981]= -2134405552;
assign addr[17982]= -2146380306;
assign addr[17983]= -2114858546;
assign addr[17984]= -2040479063;
assign addr[17985]= -1924749160;
assign addr[17986]= -1770014111;
assign addr[17987]= -1579409630;
assign addr[17988]= -1356798326;
assign addr[17989]= -1106691431;
assign addr[17990]= -834157373;
assign addr[17991]= -544719071;
assign addr[17992]= -244242007;
assign addr[17993]= 61184634;
assign addr[17994]= 365371365;
assign addr[17995]= 662153826;
assign addr[17996]= 945517704;
assign addr[17997]= 1209720613;
assign addr[17998]= 1449408469;
assign addr[17999]= 1659723983;
assign addr[18000]= 1836405100;
assign addr[18001]= 1975871368;
assign addr[18002]= 2075296495;
assign addr[18003]= 2132665626;
assign addr[18004]= 2146816171;
assign addr[18005]= 2117461370;
assign addr[18006]= 2045196100;
assign addr[18007]= 1931484818;
assign addr[18008]= 1778631892;
assign addr[18009]= 1589734894;
assign addr[18010]= 1368621831;
assign addr[18011]= 1119773573;
assign addr[18012]= 848233042;
assign addr[18013]= 559503022;
assign addr[18014]= 259434643;
assign addr[18015]= -45891193;
assign addr[18016]= -350287041;
assign addr[18017]= -647584304;
assign addr[18018]= -931758235;
assign addr[18019]= -1197050035;
assign addr[18020]= -1438083551;
assign addr[18021]= -1649974225;
assign addr[18022]= -1828428082;
assign addr[18023]= -1969828744;
assign addr[18024]= -2071310720;
assign addr[18025]= -2130817471;
assign addr[18026]= -2147143090;
assign addr[18027]= -2119956737;
assign addr[18028]= -2049809346;
assign addr[18029]= -1938122457;
assign addr[18030]= -1787159411;
assign addr[18031]= -1599979481;
assign addr[18032]= -1380375881;
assign addr[18033]= -1132798888;
assign addr[18034]= -862265664;
assign addr[18035]= -574258580;
assign addr[18036]= -274614114;
assign addr[18037]= 30595422;
assign addr[18038]= 335184940;
assign addr[18039]= 632981917;
assign addr[18040]= 917951481;
assign addr[18041]= 1184318708;
assign addr[18042]= 1426685652;
assign addr[18043]= 1640140734;
assign addr[18044]= 1820358275;
assign addr[18045]= 1963686155;
assign addr[18046]= 2067219829;
assign addr[18047]= 2128861181;
assign addr[18048]= 2147361045;
assign addr[18049]= 2122344521;
assign addr[18050]= 2054318569;
assign addr[18051]= 1944661739;
assign addr[18052]= 1795596234;
assign addr[18053]= 1610142873;
assign addr[18054]= 1392059879;
assign addr[18055]= 1145766716;
assign addr[18056]= 876254528;
assign addr[18057]= 588984994;
assign addr[18058]= 289779648;
assign addr[18059]= -15298099;
assign addr[18060]= -320065829;
assign addr[18061]= -618347408;
assign addr[18062]= -904098143;
assign addr[18063]= -1171527280;
assign addr[18064]= -1415215352;
assign addr[18065]= -1630224009;
assign addr[18066]= -1812196087;
assign addr[18067]= -1957443913;
assign addr[18068]= -2063024031;
assign addr[18069]= -2126796855;
assign addr[18070]= -2147470025;
assign addr[18071]= -2124624598;
assign addr[18072]= -2058723538;
assign addr[18073]= -1951102334;
assign addr[18074]= -1803941934;
assign addr[18075]= -1620224553;
assign addr[18076]= -1403673233;
assign addr[18077]= -1158676398;
assign addr[18078]= -890198924;
assign addr[18079]= -603681519;
assign addr[18080]= -304930476;
assign addr[18081]= 0;
assign addr[18082]= 304930476;
assign addr[18083]= 603681519;
assign addr[18084]= 890198924;
assign addr[18085]= 1158676398;
assign addr[18086]= 1403673233;
assign addr[18087]= 1620224553;
assign addr[18088]= 1803941934;
assign addr[18089]= 1951102334;
assign addr[18090]= 2058723538;
assign addr[18091]= 2124624598;
assign addr[18092]= 2147470025;
assign addr[18093]= 2126796855;
assign addr[18094]= 2063024031;
assign addr[18095]= 1957443913;
assign addr[18096]= 1812196087;
assign addr[18097]= 1630224009;
assign addr[18098]= 1415215352;
assign addr[18099]= 1171527280;
assign addr[18100]= 904098143;
assign addr[18101]= 618347408;
assign addr[18102]= 320065829;
assign addr[18103]= 15298099;
assign addr[18104]= -289779648;
assign addr[18105]= -588984994;
assign addr[18106]= -876254528;
assign addr[18107]= -1145766716;
assign addr[18108]= -1392059879;
assign addr[18109]= -1610142873;
assign addr[18110]= -1795596234;
assign addr[18111]= -1944661739;
assign addr[18112]= -2054318569;
assign addr[18113]= -2122344521;
assign addr[18114]= -2147361045;
assign addr[18115]= -2128861181;
assign addr[18116]= -2067219829;
assign addr[18117]= -1963686155;
assign addr[18118]= -1820358275;
assign addr[18119]= -1640140734;
assign addr[18120]= -1426685652;
assign addr[18121]= -1184318708;
assign addr[18122]= -917951481;
assign addr[18123]= -632981917;
assign addr[18124]= -335184940;
assign addr[18125]= -30595422;
assign addr[18126]= 274614114;
assign addr[18127]= 574258580;
assign addr[18128]= 862265664;
assign addr[18129]= 1132798888;
assign addr[18130]= 1380375881;
assign addr[18131]= 1599979481;
assign addr[18132]= 1787159411;
assign addr[18133]= 1938122457;
assign addr[18134]= 2049809346;
assign addr[18135]= 2119956737;
assign addr[18136]= 2147143090;
assign addr[18137]= 2130817471;
assign addr[18138]= 2071310720;
assign addr[18139]= 1969828744;
assign addr[18140]= 1828428082;
assign addr[18141]= 1649974225;
assign addr[18142]= 1438083551;
assign addr[18143]= 1197050035;
assign addr[18144]= 931758235;
assign addr[18145]= 647584304;
assign addr[18146]= 350287041;
assign addr[18147]= 45891193;
assign addr[18148]= -259434643;
assign addr[18149]= -559503022;
assign addr[18150]= -848233042;
assign addr[18151]= -1119773573;
assign addr[18152]= -1368621831;
assign addr[18153]= -1589734894;
assign addr[18154]= -1778631892;
assign addr[18155]= -1931484818;
assign addr[18156]= -2045196100;
assign addr[18157]= -2117461370;
assign addr[18158]= -2146816171;
assign addr[18159]= -2132665626;
assign addr[18160]= -2075296495;
assign addr[18161]= -1975871368;
assign addr[18162]= -1836405100;
assign addr[18163]= -1659723983;
assign addr[18164]= -1449408469;
assign addr[18165]= -1209720613;
assign addr[18166]= -945517704;
assign addr[18167]= -662153826;
assign addr[18168]= -365371365;
assign addr[18169]= -61184634;
assign addr[18170]= 244242007;
assign addr[18171]= 544719071;
assign addr[18172]= 834157373;
assign addr[18173]= 1106691431;
assign addr[18174]= 1356798326;
assign addr[18175]= 1579409630;
assign addr[18176]= 1770014111;
assign addr[18177]= 1924749160;
assign addr[18178]= 2040479063;
assign addr[18179]= 2114858546;
assign addr[18180]= 2146380306;
assign addr[18181]= 2134405552;
assign addr[18182]= 2079176953;
assign addr[18183]= 1981813720;
assign addr[18184]= 1844288924;
assign addr[18185]= 1669389513;
assign addr[18186]= 1460659832;
assign addr[18187]= 1222329801;
assign addr[18188]= 959229189;
assign addr[18189]= 676689746;
assign addr[18190]= 380437148;
assign addr[18191]= 76474970;
assign addr[18192]= -229036977;
assign addr[18193]= -529907477;
assign addr[18194]= -820039373;
assign addr[18195]= -1093553126;
assign addr[18196]= -1344905966;
assign addr[18197]= -1569004214;
assign addr[18198]= -1761306505;
assign addr[18199]= -1917915825;
assign addr[18200]= -2035658475;
assign addr[18201]= -2112148396;
assign addr[18202]= -2145835515;
assign addr[18203]= -2136037160;
assign addr[18204]= -2082951896;
assign addr[18205]= -1987655498;
assign addr[18206]= -1852079154;
assign addr[18207]= -1678970324;
assign addr[18208]= -1471837070;
assign addr[18209]= -1234876957;
assign addr[18210]= -972891995;
assign addr[18211]= -691191324;
assign addr[18212]= -395483624;
assign addr[18213]= -91761426;
assign addr[18214]= 213820322;
assign addr[18215]= 515068990;
assign addr[18216]= 805879757;
assign addr[18217]= 1080359326;
assign addr[18218]= 1332945355;
assign addr[18219]= 1558519173;
assign addr[18220]= 1752509516;
assign addr[18221]= 1910985158;
assign addr[18222]= 2030734582;
assign addr[18223]= 2109331059;
assign addr[18224]= 2145181827;
assign addr[18225]= 2137560369;
assign addr[18226]= 2086621133;
assign addr[18227]= 1993396407;
assign addr[18228]= 1859775393;
assign addr[18229]= 1688465931;
assign addr[18230]= 1482939614;
assign addr[18231]= 1247361445;
assign addr[18232]= 986505429;
assign addr[18233]= 705657826;
assign addr[18234]= 410510029;
assign addr[18235]= 107043224;
assign addr[18236]= -198592817;
assign addr[18237]= -500204365;
assign addr[18238]= -791679244;
assign addr[18239]= -1067110699;
assign addr[18240]= -1320917099;
assign addr[18241]= -1547955041;
assign addr[18242]= -1743623590;
assign addr[18243]= -1903957513;
assign addr[18244]= -2025707632;
assign addr[18245]= -2106406677;
assign addr[18246]= -2144419275;
assign addr[18247]= -2138975100;
assign addr[18248]= -2090184478;
assign addr[18249]= -1999036154;
assign addr[18250]= -1867377253;
assign addr[18251]= -1697875851;
assign addr[18252]= -1493966902;
assign addr[18253]= -1259782632;
assign addr[18254]= -1000068799;
assign addr[18255]= -720088517;
assign addr[18256]= -425515602;
assign addr[18257]= -122319591;
assign addr[18258]= 183355234;
assign addr[18259]= 485314355;
assign addr[18260]= 777438554;
assign addr[18261]= 1053807919;
assign addr[18262]= 1308821808;
assign addr[18263]= 1537312353;
assign addr[18264]= 1734649179;
assign addr[18265]= 1896833245;
assign addr[18266]= 2020577882;
assign addr[18267]= 2103375398;
assign addr[18268]= 2143547897;
assign addr[18269]= 2140281282;
assign addr[18270]= 2093641749;
assign addr[18271]= 2004574453;
assign addr[18272]= 1874884346;
assign addr[18273]= 1707199606;
assign addr[18274]= 1504918373;
assign addr[18275]= 1272139887;
assign addr[18276]= 1013581418;
assign addr[18277]= 734482665;
assign addr[18278]= 440499581;
assign addr[18279]= 137589750;
assign addr[18280]= -168108346;
assign addr[18281]= -470399716;
assign addr[18282]= -763158411;
assign addr[18283]= -1040451659;
assign addr[18284]= -1296660098;
assign addr[18285]= -1526591649;
assign addr[18286]= -1725586737;
assign addr[18287]= -1889612716;
assign addr[18288]= -2015345591;
assign addr[18289]= -2100237377;
assign addr[18290]= -2142567738;
assign addr[18291]= -2141478848;
assign addr[18292]= -2096992772;
assign addr[18293]= -2010011024;
assign addr[18294]= -1882296293;
assign addr[18295]= -1716436725;
assign addr[18296]= -1515793473;
assign addr[18297]= -1284432584;
assign addr[18298]= -1027042599;
assign addr[18299]= -748839539;
assign addr[18300]= -455461206;
assign addr[18301]= -152852926;
assign addr[18302]= 152852926;
assign addr[18303]= 455461206;
assign addr[18304]= 748839539;
assign addr[18305]= 1027042599;
assign addr[18306]= 1284432584;
assign addr[18307]= 1515793473;
assign addr[18308]= 1716436725;
assign addr[18309]= 1882296293;
assign addr[18310]= 2010011024;
assign addr[18311]= 2096992772;
assign addr[18312]= 2141478848;
assign addr[18313]= 2142567738;
assign addr[18314]= 2100237377;
assign addr[18315]= 2015345591;
assign addr[18316]= 1889612716;
assign addr[18317]= 1725586737;
assign addr[18318]= 1526591649;
assign addr[18319]= 1296660098;
assign addr[18320]= 1040451659;
assign addr[18321]= 763158411;
assign addr[18322]= 470399716;
assign addr[18323]= 168108346;
assign addr[18324]= -137589750;
assign addr[18325]= -440499581;
assign addr[18326]= -734482665;
assign addr[18327]= -1013581418;
assign addr[18328]= -1272139887;
assign addr[18329]= -1504918373;
assign addr[18330]= -1707199606;
assign addr[18331]= -1874884346;
assign addr[18332]= -2004574453;
assign addr[18333]= -2093641749;
assign addr[18334]= -2140281282;
assign addr[18335]= -2143547897;
assign addr[18336]= -2103375398;
assign addr[18337]= -2020577882;
assign addr[18338]= -1896833245;
assign addr[18339]= -1734649179;
assign addr[18340]= -1537312353;
assign addr[18341]= -1308821808;
assign addr[18342]= -1053807919;
assign addr[18343]= -777438554;
assign addr[18344]= -485314355;
assign addr[18345]= -183355234;
assign addr[18346]= 122319591;
assign addr[18347]= 425515602;
assign addr[18348]= 720088517;
assign addr[18349]= 1000068799;
assign addr[18350]= 1259782632;
assign addr[18351]= 1493966902;
assign addr[18352]= 1697875851;
assign addr[18353]= 1867377253;
assign addr[18354]= 1999036154;
assign addr[18355]= 2090184478;
assign addr[18356]= 2138975100;
assign addr[18357]= 2144419275;
assign addr[18358]= 2106406677;
assign addr[18359]= 2025707632;
assign addr[18360]= 1903957513;
assign addr[18361]= 1743623590;
assign addr[18362]= 1547955041;
assign addr[18363]= 1320917099;
assign addr[18364]= 1067110699;
assign addr[18365]= 791679244;
assign addr[18366]= 500204365;
assign addr[18367]= 198592817;
assign addr[18368]= -107043224;
assign addr[18369]= -410510029;
assign addr[18370]= -705657826;
assign addr[18371]= -986505429;
assign addr[18372]= -1247361445;
assign addr[18373]= -1482939614;
assign addr[18374]= -1688465931;
assign addr[18375]= -1859775393;
assign addr[18376]= -1993396407;
assign addr[18377]= -2086621133;
assign addr[18378]= -2137560369;
assign addr[18379]= -2145181827;
assign addr[18380]= -2109331059;
assign addr[18381]= -2030734582;
assign addr[18382]= -1910985158;
assign addr[18383]= -1752509516;
assign addr[18384]= -1558519173;
assign addr[18385]= -1332945355;
assign addr[18386]= -1080359326;
assign addr[18387]= -805879757;
assign addr[18388]= -515068990;
assign addr[18389]= -213820322;
assign addr[18390]= 91761426;
assign addr[18391]= 395483624;
assign addr[18392]= 691191324;
assign addr[18393]= 972891995;
assign addr[18394]= 1234876957;
assign addr[18395]= 1471837070;
assign addr[18396]= 1678970324;
assign addr[18397]= 1852079154;
assign addr[18398]= 1987655498;
assign addr[18399]= 2082951896;
assign addr[18400]= 2136037160;
assign addr[18401]= 2145835515;
assign addr[18402]= 2112148396;
assign addr[18403]= 2035658475;
assign addr[18404]= 1917915825;
assign addr[18405]= 1761306505;
assign addr[18406]= 1569004214;
assign addr[18407]= 1344905966;
assign addr[18408]= 1093553126;
assign addr[18409]= 820039373;
assign addr[18410]= 529907477;
assign addr[18411]= 229036977;
assign addr[18412]= -76474970;
assign addr[18413]= -380437148;
assign addr[18414]= -676689746;
assign addr[18415]= -959229189;
assign addr[18416]= -1222329801;
assign addr[18417]= -1460659832;
assign addr[18418]= -1669389513;
assign addr[18419]= -1844288924;
assign addr[18420]= -1981813720;
assign addr[18421]= -2079176953;
assign addr[18422]= -2134405552;
assign addr[18423]= -2146380306;
assign addr[18424]= -2114858546;
assign addr[18425]= -2040479063;
assign addr[18426]= -1924749160;
assign addr[18427]= -1770014111;
assign addr[18428]= -1579409630;
assign addr[18429]= -1356798326;
assign addr[18430]= -1106691431;
assign addr[18431]= -834157373;
assign addr[18432]= -544719071;
assign addr[18433]= -244242007;
assign addr[18434]= 61184634;
assign addr[18435]= 365371365;
assign addr[18436]= 662153826;
assign addr[18437]= 945517704;
assign addr[18438]= 1209720613;
assign addr[18439]= 1449408469;
assign addr[18440]= 1659723983;
assign addr[18441]= 1836405100;
assign addr[18442]= 1975871368;
assign addr[18443]= 2075296495;
assign addr[18444]= 2132665626;
assign addr[18445]= 2146816171;
assign addr[18446]= 2117461370;
assign addr[18447]= 2045196100;
assign addr[18448]= 1931484818;
assign addr[18449]= 1778631892;
assign addr[18450]= 1589734894;
assign addr[18451]= 1368621831;
assign addr[18452]= 1119773573;
assign addr[18453]= 848233042;
assign addr[18454]= 559503022;
assign addr[18455]= 259434643;
assign addr[18456]= -45891193;
assign addr[18457]= -350287041;
assign addr[18458]= -647584304;
assign addr[18459]= -931758235;
assign addr[18460]= -1197050035;
assign addr[18461]= -1438083551;
assign addr[18462]= -1649974225;
assign addr[18463]= -1828428082;
assign addr[18464]= -1969828744;
assign addr[18465]= -2071310720;
assign addr[18466]= -2130817471;
assign addr[18467]= -2147143090;
assign addr[18468]= -2119956737;
assign addr[18469]= -2049809346;
assign addr[18470]= -1938122457;
assign addr[18471]= -1787159411;
assign addr[18472]= -1599979481;
assign addr[18473]= -1380375881;
assign addr[18474]= -1132798888;
assign addr[18475]= -862265664;
assign addr[18476]= -574258580;
assign addr[18477]= -274614114;
assign addr[18478]= 30595422;
assign addr[18479]= 335184940;
assign addr[18480]= 632981917;
assign addr[18481]= 917951481;
assign addr[18482]= 1184318708;
assign addr[18483]= 1426685652;
assign addr[18484]= 1640140734;
assign addr[18485]= 1820358275;
assign addr[18486]= 1963686155;
assign addr[18487]= 2067219829;
assign addr[18488]= 2128861181;
assign addr[18489]= 2147361045;
assign addr[18490]= 2122344521;
assign addr[18491]= 2054318569;
assign addr[18492]= 1944661739;
assign addr[18493]= 1795596234;
assign addr[18494]= 1610142873;
assign addr[18495]= 1392059879;
assign addr[18496]= 1145766716;
assign addr[18497]= 876254528;
assign addr[18498]= 588984994;
assign addr[18499]= 289779648;
assign addr[18500]= -15298099;
assign addr[18501]= -320065829;
assign addr[18502]= -618347408;
assign addr[18503]= -904098143;
assign addr[18504]= -1171527280;
assign addr[18505]= -1415215352;
assign addr[18506]= -1630224009;
assign addr[18507]= -1812196087;
assign addr[18508]= -1957443913;
assign addr[18509]= -2063024031;
assign addr[18510]= -2126796855;
assign addr[18511]= -2147470025;
assign addr[18512]= -2124624598;
assign addr[18513]= -2058723538;
assign addr[18514]= -1951102334;
assign addr[18515]= -1803941934;
assign addr[18516]= -1620224553;
assign addr[18517]= -1403673233;
assign addr[18518]= -1158676398;
assign addr[18519]= -890198924;
assign addr[18520]= -603681519;
assign addr[18521]= -304930476;
assign addr[18522]= 0;
assign addr[18523]= 304930476;
assign addr[18524]= 603681519;
assign addr[18525]= 890198924;
assign addr[18526]= 1158676398;
assign addr[18527]= 1403673233;
assign addr[18528]= 1620224553;
assign addr[18529]= 1803941934;
assign addr[18530]= 1951102334;
assign addr[18531]= 2058723538;
assign addr[18532]= 2124624598;
assign addr[18533]= 2147470025;
assign addr[18534]= 2126796855;
assign addr[18535]= 2063024031;
assign addr[18536]= 1957443913;
assign addr[18537]= 1812196087;
assign addr[18538]= 1630224009;
assign addr[18539]= 1415215352;
assign addr[18540]= 1171527280;
assign addr[18541]= 904098143;
assign addr[18542]= 618347408;
assign addr[18543]= 320065829;
assign addr[18544]= 15298099;
assign addr[18545]= -289779648;
assign addr[18546]= -588984994;
assign addr[18547]= -876254528;
assign addr[18548]= -1145766716;
assign addr[18549]= -1392059879;
assign addr[18550]= -1610142873;
assign addr[18551]= -1795596234;
assign addr[18552]= -1944661739;
assign addr[18553]= -2054318569;
assign addr[18554]= -2122344521;
assign addr[18555]= -2147361045;
assign addr[18556]= -2128861181;
assign addr[18557]= -2067219829;
assign addr[18558]= -1963686155;
assign addr[18559]= -1820358275;
assign addr[18560]= -1640140734;
assign addr[18561]= -1426685652;
assign addr[18562]= -1184318708;
assign addr[18563]= -917951481;
assign addr[18564]= -632981917;
assign addr[18565]= -335184940;
assign addr[18566]= -30595422;
assign addr[18567]= 274614114;
assign addr[18568]= 574258580;
assign addr[18569]= 862265664;
assign addr[18570]= 1132798888;
assign addr[18571]= 1380375881;
assign addr[18572]= 1599979481;
assign addr[18573]= 1787159411;
assign addr[18574]= 1938122457;
assign addr[18575]= 2049809346;
assign addr[18576]= 2119956737;
assign addr[18577]= 2147143090;
assign addr[18578]= 2130817471;
assign addr[18579]= 2071310720;
assign addr[18580]= 1969828744;
assign addr[18581]= 1828428082;
assign addr[18582]= 1649974225;
assign addr[18583]= 1438083551;
assign addr[18584]= 1197050035;
assign addr[18585]= 931758235;
assign addr[18586]= 647584304;
assign addr[18587]= 350287041;
assign addr[18588]= 45891193;
assign addr[18589]= -259434643;
assign addr[18590]= -559503022;
assign addr[18591]= -848233042;
assign addr[18592]= -1119773573;
assign addr[18593]= -1368621831;
assign addr[18594]= -1589734894;
assign addr[18595]= -1778631892;
assign addr[18596]= -1931484818;
assign addr[18597]= -2045196100;
assign addr[18598]= -2117461370;
assign addr[18599]= -2146816171;
assign addr[18600]= -2132665626;
assign addr[18601]= -2075296495;
assign addr[18602]= -1975871368;
assign addr[18603]= -1836405100;
assign addr[18604]= -1659723983;
assign addr[18605]= -1449408469;
assign addr[18606]= -1209720613;
assign addr[18607]= -945517704;
assign addr[18608]= -662153826;
assign addr[18609]= -365371365;
assign addr[18610]= -61184634;
assign addr[18611]= 244242007;
assign addr[18612]= 544719071;
assign addr[18613]= 834157373;
assign addr[18614]= 1106691431;
assign addr[18615]= 1356798326;
assign addr[18616]= 1579409630;
assign addr[18617]= 1770014111;
assign addr[18618]= 1924749160;
assign addr[18619]= 2040479063;
assign addr[18620]= 2114858546;
assign addr[18621]= 2146380306;
assign addr[18622]= 2134405552;
assign addr[18623]= 2079176953;
assign addr[18624]= 1981813720;
assign addr[18625]= 1844288924;
assign addr[18626]= 1669389513;
assign addr[18627]= 1460659832;
assign addr[18628]= 1222329801;
assign addr[18629]= 959229189;
assign addr[18630]= 676689746;
assign addr[18631]= 380437148;
assign addr[18632]= 76474970;
assign addr[18633]= -229036977;
assign addr[18634]= -529907477;
assign addr[18635]= -820039373;
assign addr[18636]= -1093553126;
assign addr[18637]= -1344905966;
assign addr[18638]= -1569004214;
assign addr[18639]= -1761306505;
assign addr[18640]= -1917915825;
assign addr[18641]= -2035658475;
assign addr[18642]= -2112148396;
assign addr[18643]= -2145835515;
assign addr[18644]= -2136037160;
assign addr[18645]= -2082951896;
assign addr[18646]= -1987655498;
assign addr[18647]= -1852079154;
assign addr[18648]= -1678970324;
assign addr[18649]= -1471837070;
assign addr[18650]= -1234876957;
assign addr[18651]= -972891995;
assign addr[18652]= -691191324;
assign addr[18653]= -395483624;
assign addr[18654]= -91761426;
assign addr[18655]= 213820322;
assign addr[18656]= 515068990;
assign addr[18657]= 805879757;
assign addr[18658]= 1080359326;
assign addr[18659]= 1332945355;
assign addr[18660]= 1558519173;
assign addr[18661]= 1752509516;
assign addr[18662]= 1910985158;
assign addr[18663]= 2030734582;
assign addr[18664]= 2109331059;
assign addr[18665]= 2145181827;
assign addr[18666]= 2137560369;
assign addr[18667]= 2086621133;
assign addr[18668]= 1993396407;
assign addr[18669]= 1859775393;
assign addr[18670]= 1688465931;
assign addr[18671]= 1482939614;
assign addr[18672]= 1247361445;
assign addr[18673]= 986505429;
assign addr[18674]= 705657826;
assign addr[18675]= 410510029;
assign addr[18676]= 107043224;
assign addr[18677]= -198592817;
assign addr[18678]= -500204365;
assign addr[18679]= -791679244;
assign addr[18680]= -1067110699;
assign addr[18681]= -1320917099;
assign addr[18682]= -1547955041;
assign addr[18683]= -1743623590;
assign addr[18684]= -1903957513;
assign addr[18685]= -2025707632;
assign addr[18686]= -2106406677;
assign addr[18687]= -2144419275;
assign addr[18688]= -2138975100;
assign addr[18689]= -2090184478;
assign addr[18690]= -1999036154;
assign addr[18691]= -1867377253;
assign addr[18692]= -1697875851;
assign addr[18693]= -1493966902;
assign addr[18694]= -1259782632;
assign addr[18695]= -1000068799;
assign addr[18696]= -720088517;
assign addr[18697]= -425515602;
assign addr[18698]= -122319591;
assign addr[18699]= 183355234;
assign addr[18700]= 485314355;
assign addr[18701]= 777438554;
assign addr[18702]= 1053807919;
assign addr[18703]= 1308821808;
assign addr[18704]= 1537312353;
assign addr[18705]= 1734649179;
assign addr[18706]= 1896833245;
assign addr[18707]= 2020577882;
assign addr[18708]= 2103375398;
assign addr[18709]= 2143547897;
assign addr[18710]= 2140281282;
assign addr[18711]= 2093641749;
assign addr[18712]= 2004574453;
assign addr[18713]= 1874884346;
assign addr[18714]= 1707199606;
assign addr[18715]= 1504918373;
assign addr[18716]= 1272139887;
assign addr[18717]= 1013581418;
assign addr[18718]= 734482665;
assign addr[18719]= 440499581;
assign addr[18720]= 137589750;
assign addr[18721]= -168108346;
assign addr[18722]= -470399716;
assign addr[18723]= -763158411;
assign addr[18724]= -1040451659;
assign addr[18725]= -1296660098;
assign addr[18726]= -1526591649;
assign addr[18727]= -1725586737;
assign addr[18728]= -1889612716;
assign addr[18729]= -2015345591;
assign addr[18730]= -2100237377;
assign addr[18731]= -2142567738;
assign addr[18732]= -2141478848;
assign addr[18733]= -2096992772;
assign addr[18734]= -2010011024;
assign addr[18735]= -1882296293;
assign addr[18736]= -1716436725;
assign addr[18737]= -1515793473;
assign addr[18738]= -1284432584;
assign addr[18739]= -1027042599;
assign addr[18740]= -748839539;
assign addr[18741]= -455461206;
assign addr[18742]= -152852926;
assign addr[18743]= 152852926;
assign addr[18744]= 455461206;
assign addr[18745]= 748839539;
assign addr[18746]= 1027042599;
assign addr[18747]= 1284432584;
assign addr[18748]= 1515793473;
assign addr[18749]= 1716436725;
assign addr[18750]= 1882296293;
assign addr[18751]= 2010011024;
assign addr[18752]= 2096992772;
assign addr[18753]= 2141478848;
assign addr[18754]= 2142567738;
assign addr[18755]= 2100237377;
assign addr[18756]= 2015345591;
assign addr[18757]= 1889612716;
assign addr[18758]= 1725586737;
assign addr[18759]= 1526591649;
assign addr[18760]= 1296660098;
assign addr[18761]= 1040451659;
assign addr[18762]= 763158411;
assign addr[18763]= 470399716;
assign addr[18764]= 168108346;
assign addr[18765]= -137589750;
assign addr[18766]= -440499581;
assign addr[18767]= -734482665;
assign addr[18768]= -1013581418;
assign addr[18769]= -1272139887;
assign addr[18770]= -1504918373;
assign addr[18771]= -1707199606;
assign addr[18772]= -1874884346;
assign addr[18773]= -2004574453;
assign addr[18774]= -2093641749;
assign addr[18775]= -2140281282;
assign addr[18776]= -2143547897;
assign addr[18777]= -2103375398;
assign addr[18778]= -2020577882;
assign addr[18779]= -1896833245;
assign addr[18780]= -1734649179;
assign addr[18781]= -1537312353;
assign addr[18782]= -1308821808;
assign addr[18783]= -1053807919;
assign addr[18784]= -777438554;
assign addr[18785]= -485314355;
assign addr[18786]= -183355234;
assign addr[18787]= 122319591;
assign addr[18788]= 425515602;
assign addr[18789]= 720088517;
assign addr[18790]= 1000068799;
assign addr[18791]= 1259782632;
assign addr[18792]= 1493966902;
assign addr[18793]= 1697875851;
assign addr[18794]= 1867377253;
assign addr[18795]= 1999036154;
assign addr[18796]= 2090184478;
assign addr[18797]= 2138975100;
assign addr[18798]= 2144419275;
assign addr[18799]= 2106406677;
assign addr[18800]= 2025707632;
assign addr[18801]= 1903957513;
assign addr[18802]= 1743623590;
assign addr[18803]= 1547955041;
assign addr[18804]= 1320917099;
assign addr[18805]= 1067110699;
assign addr[18806]= 791679244;
assign addr[18807]= 500204365;
assign addr[18808]= 198592817;
assign addr[18809]= -107043224;
assign addr[18810]= -410510029;
assign addr[18811]= -705657826;
assign addr[18812]= -986505429;
assign addr[18813]= -1247361445;
assign addr[18814]= -1482939614;
assign addr[18815]= -1688465931;
assign addr[18816]= -1859775393;
assign addr[18817]= -1993396407;
assign addr[18818]= -2086621133;
assign addr[18819]= -2137560369;
assign addr[18820]= -2145181827;
assign addr[18821]= -2109331059;
assign addr[18822]= -2030734582;
assign addr[18823]= -1910985158;
assign addr[18824]= -1752509516;
assign addr[18825]= -1558519173;
assign addr[18826]= -1332945355;
assign addr[18827]= -1080359326;
assign addr[18828]= -805879757;
assign addr[18829]= -515068990;
assign addr[18830]= -213820322;
assign addr[18831]= 91761426;
assign addr[18832]= 395483624;
assign addr[18833]= 691191324;
assign addr[18834]= 972891995;
assign addr[18835]= 1234876957;
assign addr[18836]= 1471837070;
assign addr[18837]= 1678970324;
assign addr[18838]= 1852079154;
assign addr[18839]= 1987655498;
assign addr[18840]= 2082951896;
assign addr[18841]= 2136037160;
assign addr[18842]= 2145835515;
assign addr[18843]= 2112148396;
assign addr[18844]= 2035658475;
assign addr[18845]= 1917915825;
assign addr[18846]= 1761306505;
assign addr[18847]= 1569004214;
assign addr[18848]= 1344905966;
assign addr[18849]= 1093553126;
assign addr[18850]= 820039373;
assign addr[18851]= 529907477;
assign addr[18852]= 229036977;
assign addr[18853]= -76474970;
assign addr[18854]= -380437148;
assign addr[18855]= -676689746;
assign addr[18856]= -959229189;
assign addr[18857]= -1222329801;
assign addr[18858]= -1460659832;
assign addr[18859]= -1669389513;
assign addr[18860]= -1844288924;
assign addr[18861]= -1981813720;
assign addr[18862]= -2079176953;
assign addr[18863]= -2134405552;
assign addr[18864]= -2146380306;
assign addr[18865]= -2114858546;
assign addr[18866]= -2040479063;
assign addr[18867]= -1924749160;
assign addr[18868]= -1770014111;
assign addr[18869]= -1579409630;
assign addr[18870]= -1356798326;
assign addr[18871]= -1106691431;
assign addr[18872]= -834157373;
assign addr[18873]= -544719071;
assign addr[18874]= -244242007;
assign addr[18875]= 61184634;
assign addr[18876]= 365371365;
assign addr[18877]= 662153826;
assign addr[18878]= 945517704;
assign addr[18879]= 1209720613;
assign addr[18880]= 1449408469;
assign addr[18881]= 1659723983;
assign addr[18882]= 1836405100;
assign addr[18883]= 1975871368;
assign addr[18884]= 2075296495;
assign addr[18885]= 2132665626;
assign addr[18886]= 2146816171;
assign addr[18887]= 2117461370;
assign addr[18888]= 2045196100;
assign addr[18889]= 1931484818;
assign addr[18890]= 1778631892;
assign addr[18891]= 1589734894;
assign addr[18892]= 1368621831;
assign addr[18893]= 1119773573;
assign addr[18894]= 848233042;
assign addr[18895]= 559503022;
assign addr[18896]= 259434643;
assign addr[18897]= -45891193;
assign addr[18898]= -350287041;
assign addr[18899]= -647584304;
assign addr[18900]= -931758235;
assign addr[18901]= -1197050035;
assign addr[18902]= -1438083551;
assign addr[18903]= -1649974225;
assign addr[18904]= -1828428082;
assign addr[18905]= -1969828744;
assign addr[18906]= -2071310720;
assign addr[18907]= -2130817471;
assign addr[18908]= -2147143090;
assign addr[18909]= -2119956737;
assign addr[18910]= -2049809346;
assign addr[18911]= -1938122457;
assign addr[18912]= -1787159411;
assign addr[18913]= -1599979481;
assign addr[18914]= -1380375881;
assign addr[18915]= -1132798888;
assign addr[18916]= -862265664;
assign addr[18917]= -574258580;
assign addr[18918]= -274614114;
assign addr[18919]= 30595422;
assign addr[18920]= 335184940;
assign addr[18921]= 632981917;
assign addr[18922]= 917951481;
assign addr[18923]= 1184318708;
assign addr[18924]= 1426685652;
assign addr[18925]= 1640140734;
assign addr[18926]= 1820358275;
assign addr[18927]= 1963686155;
assign addr[18928]= 2067219829;
assign addr[18929]= 2128861181;
assign addr[18930]= 2147361045;
assign addr[18931]= 2122344521;
assign addr[18932]= 2054318569;
assign addr[18933]= 1944661739;
assign addr[18934]= 1795596234;
assign addr[18935]= 1610142873;
assign addr[18936]= 1392059879;
assign addr[18937]= 1145766716;
assign addr[18938]= 876254528;
assign addr[18939]= 588984994;
assign addr[18940]= 289779648;
assign addr[18941]= -15298099;
assign addr[18942]= -320065829;
assign addr[18943]= -618347408;
assign addr[18944]= -904098143;
assign addr[18945]= -1171527280;
assign addr[18946]= -1415215352;
assign addr[18947]= -1630224009;
assign addr[18948]= -1812196087;
assign addr[18949]= -1957443913;
assign addr[18950]= -2063024031;
assign addr[18951]= -2126796855;
assign addr[18952]= -2147470025;
assign addr[18953]= -2124624598;
assign addr[18954]= -2058723538;
assign addr[18955]= -1951102334;
assign addr[18956]= -1803941934;
assign addr[18957]= -1620224553;
assign addr[18958]= -1403673233;
assign addr[18959]= -1158676398;
assign addr[18960]= -890198924;
assign addr[18961]= -603681519;
assign addr[18962]= -304930476;
assign addr[18963]= 0;
assign addr[18964]= 304930476;
assign addr[18965]= 603681519;
assign addr[18966]= 890198924;
assign addr[18967]= 1158676398;
assign addr[18968]= 1403673233;
assign addr[18969]= 1620224553;
assign addr[18970]= 1803941934;
assign addr[18971]= 1951102334;
assign addr[18972]= 2058723538;
assign addr[18973]= 2124624598;
assign addr[18974]= 2147470025;
assign addr[18975]= 2126796855;
assign addr[18976]= 2063024031;
assign addr[18977]= 1957443913;
assign addr[18978]= 1812196087;
assign addr[18979]= 1630224009;
assign addr[18980]= 1415215352;
assign addr[18981]= 1171527280;
assign addr[18982]= 904098143;
assign addr[18983]= 618347408;
assign addr[18984]= 320065829;
assign addr[18985]= 15298099;
assign addr[18986]= -289779648;
assign addr[18987]= -588984994;
assign addr[18988]= -876254528;
assign addr[18989]= -1145766716;
assign addr[18990]= -1392059879;
assign addr[18991]= -1610142873;
assign addr[18992]= -1795596234;
assign addr[18993]= -1944661739;
assign addr[18994]= -2054318569;
assign addr[18995]= -2122344521;
assign addr[18996]= -2147361045;
assign addr[18997]= -2128861181;
assign addr[18998]= -2067219829;
assign addr[18999]= -1963686155;
assign addr[19000]= -1820358275;
assign addr[19001]= -1640140734;
assign addr[19002]= -1426685652;
assign addr[19003]= -1184318708;
assign addr[19004]= -917951481;
assign addr[19005]= -632981917;
assign addr[19006]= -335184940;
assign addr[19007]= -30595422;
assign addr[19008]= 274614114;
assign addr[19009]= 574258580;
assign addr[19010]= 862265664;
assign addr[19011]= 1132798888;
assign addr[19012]= 1380375881;
assign addr[19013]= 1599979481;
assign addr[19014]= 1787159411;
assign addr[19015]= 1938122457;
assign addr[19016]= 2049809346;
assign addr[19017]= 2119956737;
assign addr[19018]= 2147143090;
assign addr[19019]= 2130817471;
assign addr[19020]= 2071310720;
assign addr[19021]= 1969828744;
assign addr[19022]= 1828428082;
assign addr[19023]= 1649974225;
assign addr[19024]= 1438083551;
assign addr[19025]= 1197050035;
assign addr[19026]= 931758235;
assign addr[19027]= 647584304;
assign addr[19028]= 350287041;
assign addr[19029]= 45891193;
assign addr[19030]= -259434643;
assign addr[19031]= -559503022;
assign addr[19032]= -848233042;
assign addr[19033]= -1119773573;
assign addr[19034]= -1368621831;
assign addr[19035]= -1589734894;
assign addr[19036]= -1778631892;
assign addr[19037]= -1931484818;
assign addr[19038]= -2045196100;
assign addr[19039]= -2117461370;
assign addr[19040]= -2146816171;
assign addr[19041]= -2132665626;
assign addr[19042]= -2075296495;
assign addr[19043]= -1975871368;
assign addr[19044]= -1836405100;
assign addr[19045]= -1659723983;
assign addr[19046]= -1449408469;
assign addr[19047]= -1209720613;
assign addr[19048]= -945517704;
assign addr[19049]= -662153826;
assign addr[19050]= -365371365;
assign addr[19051]= -61184634;
assign addr[19052]= 244242007;
assign addr[19053]= 544719071;
assign addr[19054]= 834157373;
assign addr[19055]= 1106691431;
assign addr[19056]= 1356798326;
assign addr[19057]= 1579409630;
assign addr[19058]= 1770014111;
assign addr[19059]= 1924749160;
assign addr[19060]= 2040479063;
assign addr[19061]= 2114858546;
assign addr[19062]= 2146380306;
assign addr[19063]= 2134405552;
assign addr[19064]= 2079176953;
assign addr[19065]= 1981813720;
assign addr[19066]= 1844288924;
assign addr[19067]= 1669389513;
assign addr[19068]= 1460659832;
assign addr[19069]= 1222329801;
assign addr[19070]= 959229189;
assign addr[19071]= 676689746;
assign addr[19072]= 380437148;
assign addr[19073]= 76474970;
assign addr[19074]= -229036977;
assign addr[19075]= -529907477;
assign addr[19076]= -820039373;
assign addr[19077]= -1093553126;
assign addr[19078]= -1344905966;
assign addr[19079]= -1569004214;
assign addr[19080]= -1761306505;
assign addr[19081]= -1917915825;
assign addr[19082]= -2035658475;
assign addr[19083]= -2112148396;
assign addr[19084]= -2145835515;
assign addr[19085]= -2136037160;
assign addr[19086]= -2082951896;
assign addr[19087]= -1987655498;
assign addr[19088]= -1852079154;
assign addr[19089]= -1678970324;
assign addr[19090]= -1471837070;
assign addr[19091]= -1234876957;
assign addr[19092]= -972891995;
assign addr[19093]= -691191324;
assign addr[19094]= -395483624;
assign addr[19095]= -91761426;
assign addr[19096]= 213820322;
assign addr[19097]= 515068990;
assign addr[19098]= 805879757;
assign addr[19099]= 1080359326;
assign addr[19100]= 1332945355;
assign addr[19101]= 1558519173;
assign addr[19102]= 1752509516;
assign addr[19103]= 1910985158;
assign addr[19104]= 2030734582;
assign addr[19105]= 2109331059;
assign addr[19106]= 2145181827;
assign addr[19107]= 2137560369;
assign addr[19108]= 2086621133;
assign addr[19109]= 1993396407;
assign addr[19110]= 1859775393;
assign addr[19111]= 1688465931;
assign addr[19112]= 1482939614;
assign addr[19113]= 1247361445;
assign addr[19114]= 986505429;
assign addr[19115]= 705657826;
assign addr[19116]= 410510029;
assign addr[19117]= 107043224;
assign addr[19118]= -198592817;
assign addr[19119]= -500204365;
assign addr[19120]= -791679244;
assign addr[19121]= -1067110699;
assign addr[19122]= -1320917099;
assign addr[19123]= -1547955041;
assign addr[19124]= -1743623590;
assign addr[19125]= -1903957513;
assign addr[19126]= -2025707632;
assign addr[19127]= -2106406677;
assign addr[19128]= -2144419275;
assign addr[19129]= -2138975100;
assign addr[19130]= -2090184478;
assign addr[19131]= -1999036154;
assign addr[19132]= -1867377253;
assign addr[19133]= -1697875851;
assign addr[19134]= -1493966902;
assign addr[19135]= -1259782632;
assign addr[19136]= -1000068799;
assign addr[19137]= -720088517;
assign addr[19138]= -425515602;
assign addr[19139]= -122319591;
assign addr[19140]= 183355234;
assign addr[19141]= 485314355;
assign addr[19142]= 777438554;
assign addr[19143]= 1053807919;
assign addr[19144]= 1308821808;
assign addr[19145]= 1537312353;
assign addr[19146]= 1734649179;
assign addr[19147]= 1896833245;
assign addr[19148]= 2020577882;
assign addr[19149]= 2103375398;
assign addr[19150]= 2143547897;
assign addr[19151]= 2140281282;
assign addr[19152]= 2093641749;
assign addr[19153]= 2004574453;
assign addr[19154]= 1874884346;
assign addr[19155]= 1707199606;
assign addr[19156]= 1504918373;
assign addr[19157]= 1272139887;
assign addr[19158]= 1013581418;
assign addr[19159]= 734482665;
assign addr[19160]= 440499581;
assign addr[19161]= 137589750;
assign addr[19162]= -168108346;
assign addr[19163]= -470399716;
assign addr[19164]= -763158411;
assign addr[19165]= -1040451659;
assign addr[19166]= -1296660098;
assign addr[19167]= -1526591649;
assign addr[19168]= -1725586737;
assign addr[19169]= -1889612716;
assign addr[19170]= -2015345591;
assign addr[19171]= -2100237377;
assign addr[19172]= -2142567738;
assign addr[19173]= -2141478848;
assign addr[19174]= -2096992772;
assign addr[19175]= -2010011024;
assign addr[19176]= -1882296293;
assign addr[19177]= -1716436725;
assign addr[19178]= -1515793473;
assign addr[19179]= -1284432584;
assign addr[19180]= -1027042599;
assign addr[19181]= -748839539;
assign addr[19182]= -455461206;
assign addr[19183]= -152852926;
assign addr[19184]= 152852926;
assign addr[19185]= 455461206;
assign addr[19186]= 748839539;
assign addr[19187]= 1027042599;
assign addr[19188]= 1284432584;
assign addr[19189]= 1515793473;
assign addr[19190]= 1716436725;
assign addr[19191]= 1882296293;
assign addr[19192]= 2010011024;
assign addr[19193]= 2096992772;
assign addr[19194]= 2141478848;
assign addr[19195]= 2142567738;
assign addr[19196]= 2100237377;
assign addr[19197]= 2015345591;
assign addr[19198]= 1889612716;
assign addr[19199]= 1725586737;
assign addr[19200]= 1526591649;
assign addr[19201]= 1296660098;
assign addr[19202]= 1040451659;
assign addr[19203]= 763158411;
assign addr[19204]= 470399716;
assign addr[19205]= 168108346;
assign addr[19206]= -137589750;
assign addr[19207]= -440499581;
assign addr[19208]= -734482665;
assign addr[19209]= -1013581418;
assign addr[19210]= -1272139887;
assign addr[19211]= -1504918373;
assign addr[19212]= -1707199606;
assign addr[19213]= -1874884346;
assign addr[19214]= -2004574453;
assign addr[19215]= -2093641749;
assign addr[19216]= -2140281282;
assign addr[19217]= -2143547897;
assign addr[19218]= -2103375398;
assign addr[19219]= -2020577882;
assign addr[19220]= -1896833245;
assign addr[19221]= -1734649179;
assign addr[19222]= -1537312353;
assign addr[19223]= -1308821808;
assign addr[19224]= -1053807919;
assign addr[19225]= -777438554;
assign addr[19226]= -485314355;
assign addr[19227]= -183355234;
assign addr[19228]= 122319591;
assign addr[19229]= 425515602;
assign addr[19230]= 720088517;
assign addr[19231]= 1000068799;
assign addr[19232]= 1259782632;
assign addr[19233]= 1493966902;
assign addr[19234]= 1697875851;
assign addr[19235]= 1867377253;
assign addr[19236]= 1999036154;
assign addr[19237]= 2090184478;
assign addr[19238]= 2138975100;
assign addr[19239]= 2144419275;
assign addr[19240]= 2106406677;
assign addr[19241]= 2025707632;
assign addr[19242]= 1903957513;
assign addr[19243]= 1743623590;
assign addr[19244]= 1547955041;
assign addr[19245]= 1320917099;
assign addr[19246]= 1067110699;
assign addr[19247]= 791679244;
assign addr[19248]= 500204365;
assign addr[19249]= 198592817;
assign addr[19250]= -107043224;
assign addr[19251]= -410510029;
assign addr[19252]= -705657826;
assign addr[19253]= -986505429;
assign addr[19254]= -1247361445;
assign addr[19255]= -1482939614;
assign addr[19256]= -1688465931;
assign addr[19257]= -1859775393;
assign addr[19258]= -1993396407;
assign addr[19259]= -2086621133;
assign addr[19260]= -2137560369;
assign addr[19261]= -2145181827;
assign addr[19262]= -2109331059;
assign addr[19263]= -2030734582;
assign addr[19264]= -1910985158;
assign addr[19265]= -1752509516;
assign addr[19266]= -1558519173;
assign addr[19267]= -1332945355;
assign addr[19268]= -1080359326;
assign addr[19269]= -805879757;
assign addr[19270]= -515068990;
assign addr[19271]= -213820322;
assign addr[19272]= 91761426;
assign addr[19273]= 395483624;
assign addr[19274]= 691191324;
assign addr[19275]= 972891995;
assign addr[19276]= 1234876957;
assign addr[19277]= 1471837070;
assign addr[19278]= 1678970324;
assign addr[19279]= 1852079154;
assign addr[19280]= 1987655498;
assign addr[19281]= 2082951896;
assign addr[19282]= 2136037160;
assign addr[19283]= 2145835515;
assign addr[19284]= 2112148396;
assign addr[19285]= 2035658475;
assign addr[19286]= 1917915825;
assign addr[19287]= 1761306505;
assign addr[19288]= 1569004214;
assign addr[19289]= 1344905966;
assign addr[19290]= 1093553126;
assign addr[19291]= 820039373;
assign addr[19292]= 529907477;
assign addr[19293]= 229036977;
assign addr[19294]= -76474970;
assign addr[19295]= -380437148;
assign addr[19296]= -676689746;
assign addr[19297]= -959229189;
assign addr[19298]= -1222329801;
assign addr[19299]= -1460659832;
assign addr[19300]= -1669389513;
assign addr[19301]= -1844288924;
assign addr[19302]= -1981813720;
assign addr[19303]= -2079176953;
assign addr[19304]= -2134405552;
assign addr[19305]= -2146380306;
assign addr[19306]= -2114858546;
assign addr[19307]= -2040479063;
assign addr[19308]= -1924749160;
assign addr[19309]= -1770014111;
assign addr[19310]= -1579409630;
assign addr[19311]= -1356798326;
assign addr[19312]= -1106691431;
assign addr[19313]= -834157373;
assign addr[19314]= -544719071;
assign addr[19315]= -244242007;
assign addr[19316]= 61184634;
assign addr[19317]= 365371365;
assign addr[19318]= 662153826;
assign addr[19319]= 945517704;
assign addr[19320]= 1209720613;
assign addr[19321]= 1449408469;
assign addr[19322]= 1659723983;
assign addr[19323]= 1836405100;
assign addr[19324]= 1975871368;
assign addr[19325]= 2075296495;
assign addr[19326]= 2132665626;
assign addr[19327]= 2146816171;
assign addr[19328]= 2117461370;
assign addr[19329]= 2045196100;
assign addr[19330]= 1931484818;
assign addr[19331]= 1778631892;
assign addr[19332]= 1589734894;
assign addr[19333]= 1368621831;
assign addr[19334]= 1119773573;
assign addr[19335]= 848233042;
assign addr[19336]= 559503022;
assign addr[19337]= 259434643;
assign addr[19338]= -45891193;
assign addr[19339]= -350287041;
assign addr[19340]= -647584304;
assign addr[19341]= -931758235;
assign addr[19342]= -1197050035;
assign addr[19343]= -1438083551;
assign addr[19344]= -1649974225;
assign addr[19345]= -1828428082;
assign addr[19346]= -1969828744;
assign addr[19347]= -2071310720;
assign addr[19348]= -2130817471;
assign addr[19349]= -2147143090;
assign addr[19350]= -2119956737;
assign addr[19351]= -2049809346;
assign addr[19352]= -1938122457;
assign addr[19353]= -1787159411;
assign addr[19354]= -1599979481;
assign addr[19355]= -1380375881;
assign addr[19356]= -1132798888;
assign addr[19357]= -862265664;
assign addr[19358]= -574258580;
assign addr[19359]= -274614114;
assign addr[19360]= 30595422;
assign addr[19361]= 335184940;
assign addr[19362]= 632981917;
assign addr[19363]= 917951481;
assign addr[19364]= 1184318708;
assign addr[19365]= 1426685652;
assign addr[19366]= 1640140734;
assign addr[19367]= 1820358275;
assign addr[19368]= 1963686155;
assign addr[19369]= 2067219829;
assign addr[19370]= 2128861181;
assign addr[19371]= 2147361045;
assign addr[19372]= 2122344521;
assign addr[19373]= 2054318569;
assign addr[19374]= 1944661739;
assign addr[19375]= 1795596234;
assign addr[19376]= 1610142873;
assign addr[19377]= 1392059879;
assign addr[19378]= 1145766716;
assign addr[19379]= 876254528;
assign addr[19380]= 588984994;
assign addr[19381]= 289779648;
assign addr[19382]= -15298099;
assign addr[19383]= -320065829;
assign addr[19384]= -618347408;
assign addr[19385]= -904098143;
assign addr[19386]= -1171527280;
assign addr[19387]= -1415215352;
assign addr[19388]= -1630224009;
assign addr[19389]= -1812196087;
assign addr[19390]= -1957443913;
assign addr[19391]= -2063024031;
assign addr[19392]= -2126796855;
assign addr[19393]= -2147470025;
assign addr[19394]= -2124624598;
assign addr[19395]= -2058723538;
assign addr[19396]= -1951102334;
assign addr[19397]= -1803941934;
assign addr[19398]= -1620224553;
assign addr[19399]= -1403673233;
assign addr[19400]= -1158676398;
assign addr[19401]= -890198924;
assign addr[19402]= -603681519;
assign addr[19403]= -304930476;
assign addr[19404]= 0;
assign addr[19405]= 304930476;
assign addr[19406]= 603681519;
assign addr[19407]= 890198924;
assign addr[19408]= 1158676398;
assign addr[19409]= 1403673233;
assign addr[19410]= 1620224553;
assign addr[19411]= 1803941934;
assign addr[19412]= 1951102334;
assign addr[19413]= 2058723538;
assign addr[19414]= 2124624598;
assign addr[19415]= 2147470025;
assign addr[19416]= 2126796855;
assign addr[19417]= 2063024031;
assign addr[19418]= 1957443913;
assign addr[19419]= 1812196087;
assign addr[19420]= 1630224009;
assign addr[19421]= 1415215352;
assign addr[19422]= 1171527280;
assign addr[19423]= 904098143;
assign addr[19424]= 618347408;
assign addr[19425]= 320065829;
assign addr[19426]= 15298099;
assign addr[19427]= -289779648;
assign addr[19428]= -588984994;
assign addr[19429]= -876254528;
assign addr[19430]= -1145766716;
assign addr[19431]= -1392059879;
assign addr[19432]= -1610142873;
assign addr[19433]= -1795596234;
assign addr[19434]= -1944661739;
assign addr[19435]= -2054318569;
assign addr[19436]= -2122344521;
assign addr[19437]= -2147361045;
assign addr[19438]= -2128861181;
assign addr[19439]= -2067219829;
assign addr[19440]= -1963686155;
assign addr[19441]= -1820358275;
assign addr[19442]= -1640140734;
assign addr[19443]= -1426685652;
assign addr[19444]= -1184318708;
assign addr[19445]= -917951481;
assign addr[19446]= -632981917;
assign addr[19447]= -335184940;
assign addr[19448]= -30595422;
assign addr[19449]= 274614114;
assign addr[19450]= 574258580;
assign addr[19451]= 862265664;
assign addr[19452]= 1132798888;
assign addr[19453]= 1380375881;
assign addr[19454]= 1599979481;
assign addr[19455]= 1787159411;
assign addr[19456]= 1938122457;
assign addr[19457]= 2049809346;
assign addr[19458]= 2119956737;
assign addr[19459]= 2147143090;
assign addr[19460]= 2130817471;
assign addr[19461]= 2071310720;
assign addr[19462]= 1969828744;
assign addr[19463]= 1828428082;
assign addr[19464]= 1649974225;
assign addr[19465]= 1438083551;
assign addr[19466]= 1197050035;
assign addr[19467]= 931758235;
assign addr[19468]= 647584304;
assign addr[19469]= 350287041;
assign addr[19470]= 45891193;
assign addr[19471]= -259434643;
assign addr[19472]= -559503022;
assign addr[19473]= -848233042;
assign addr[19474]= -1119773573;
assign addr[19475]= -1368621831;
assign addr[19476]= -1589734894;
assign addr[19477]= -1778631892;
assign addr[19478]= -1931484818;
assign addr[19479]= -2045196100;
assign addr[19480]= -2117461370;
assign addr[19481]= -2146816171;
assign addr[19482]= -2132665626;
assign addr[19483]= -2075296495;
assign addr[19484]= -1975871368;
assign addr[19485]= -1836405100;
assign addr[19486]= -1659723983;
assign addr[19487]= -1449408469;
assign addr[19488]= -1209720613;
assign addr[19489]= -945517704;
assign addr[19490]= -662153826;
assign addr[19491]= -365371365;
assign addr[19492]= -61184634;
assign addr[19493]= 244242007;
assign addr[19494]= 544719071;
assign addr[19495]= 834157373;
assign addr[19496]= 1106691431;
assign addr[19497]= 1356798326;
assign addr[19498]= 1579409630;
assign addr[19499]= 1770014111;
assign addr[19500]= 1924749160;
assign addr[19501]= 2040479063;
assign addr[19502]= 2114858546;
assign addr[19503]= 2146380306;
assign addr[19504]= 2134405552;
assign addr[19505]= 2079176953;
assign addr[19506]= 1981813720;
assign addr[19507]= 1844288924;
assign addr[19508]= 1669389513;
assign addr[19509]= 1460659832;
assign addr[19510]= 1222329801;
assign addr[19511]= 959229189;
assign addr[19512]= 676689746;
assign addr[19513]= 380437148;
assign addr[19514]= 76474970;
assign addr[19515]= -229036977;
assign addr[19516]= -529907477;
assign addr[19517]= -820039373;
assign addr[19518]= -1093553126;
assign addr[19519]= -1344905966;
assign addr[19520]= -1569004214;
assign addr[19521]= -1761306505;
assign addr[19522]= -1917915825;
assign addr[19523]= -2035658475;
assign addr[19524]= -2112148396;
assign addr[19525]= -2145835515;
assign addr[19526]= -2136037160;
assign addr[19527]= -2082951896;
assign addr[19528]= -1987655498;
assign addr[19529]= -1852079154;
assign addr[19530]= -1678970324;
assign addr[19531]= -1471837070;
assign addr[19532]= -1234876957;
assign addr[19533]= -972891995;
assign addr[19534]= -691191324;
assign addr[19535]= -395483624;
assign addr[19536]= -91761426;
assign addr[19537]= 213820322;
assign addr[19538]= 515068990;
assign addr[19539]= 805879757;
assign addr[19540]= 1080359326;
assign addr[19541]= 1332945355;
assign addr[19542]= 1558519173;
assign addr[19543]= 1752509516;
assign addr[19544]= 1910985158;
assign addr[19545]= 2030734582;
assign addr[19546]= 2109331059;
assign addr[19547]= 2145181827;
assign addr[19548]= 2137560369;
assign addr[19549]= 2086621133;
assign addr[19550]= 1993396407;
assign addr[19551]= 1859775393;
assign addr[19552]= 1688465931;
assign addr[19553]= 1482939614;
assign addr[19554]= 1247361445;
assign addr[19555]= 986505429;
assign addr[19556]= 705657826;
assign addr[19557]= 410510029;
assign addr[19558]= 107043224;
assign addr[19559]= -198592817;
assign addr[19560]= -500204365;
assign addr[19561]= -791679244;
assign addr[19562]= -1067110699;
assign addr[19563]= -1320917099;
assign addr[19564]= -1547955041;
assign addr[19565]= -1743623590;
assign addr[19566]= -1903957513;
assign addr[19567]= -2025707632;
assign addr[19568]= -2106406677;
assign addr[19569]= -2144419275;
assign addr[19570]= -2138975100;
assign addr[19571]= -2090184478;
assign addr[19572]= -1999036154;
assign addr[19573]= -1867377253;
assign addr[19574]= -1697875851;
assign addr[19575]= -1493966902;
assign addr[19576]= -1259782632;
assign addr[19577]= -1000068799;
assign addr[19578]= -720088517;
assign addr[19579]= -425515602;
assign addr[19580]= -122319591;
assign addr[19581]= 183355234;
assign addr[19582]= 485314355;
assign addr[19583]= 777438554;
assign addr[19584]= 1053807919;
assign addr[19585]= 1308821808;
assign addr[19586]= 1537312353;
assign addr[19587]= 1734649179;
assign addr[19588]= 1896833245;
assign addr[19589]= 2020577882;
assign addr[19590]= 2103375398;
assign addr[19591]= 2143547897;
assign addr[19592]= 2140281282;
assign addr[19593]= 2093641749;
assign addr[19594]= 2004574453;
assign addr[19595]= 1874884346;
assign addr[19596]= 1707199606;
assign addr[19597]= 1504918373;
assign addr[19598]= 1272139887;
assign addr[19599]= 1013581418;
assign addr[19600]= 734482665;
assign addr[19601]= 440499581;
assign addr[19602]= 137589750;
assign addr[19603]= -168108346;
assign addr[19604]= -470399716;
assign addr[19605]= -763158411;
assign addr[19606]= -1040451659;
assign addr[19607]= -1296660098;
assign addr[19608]= -1526591649;
assign addr[19609]= -1725586737;
assign addr[19610]= -1889612716;
assign addr[19611]= -2015345591;
assign addr[19612]= -2100237377;
assign addr[19613]= -2142567738;
assign addr[19614]= -2141478848;
assign addr[19615]= -2096992772;
assign addr[19616]= -2010011024;
assign addr[19617]= -1882296293;
assign addr[19618]= -1716436725;
assign addr[19619]= -1515793473;
assign addr[19620]= -1284432584;
assign addr[19621]= -1027042599;
assign addr[19622]= -748839539;
assign addr[19623]= -455461206;
assign addr[19624]= -152852926;
assign addr[19625]= 152852926;
assign addr[19626]= 455461206;
assign addr[19627]= 748839539;
assign addr[19628]= 1027042599;
assign addr[19629]= 1284432584;
assign addr[19630]= 1515793473;
assign addr[19631]= 1716436725;
assign addr[19632]= 1882296293;
assign addr[19633]= 2010011024;
assign addr[19634]= 2096992772;
assign addr[19635]= 2141478848;
assign addr[19636]= 2142567738;
assign addr[19637]= 2100237377;
assign addr[19638]= 2015345591;
assign addr[19639]= 1889612716;
assign addr[19640]= 1725586737;
assign addr[19641]= 1526591649;
assign addr[19642]= 1296660098;
assign addr[19643]= 1040451659;
assign addr[19644]= 763158411;
assign addr[19645]= 470399716;
assign addr[19646]= 168108346;
assign addr[19647]= -137589750;
assign addr[19648]= -440499581;
assign addr[19649]= -734482665;
assign addr[19650]= -1013581418;
assign addr[19651]= -1272139887;
assign addr[19652]= -1504918373;
assign addr[19653]= -1707199606;
assign addr[19654]= -1874884346;
assign addr[19655]= -2004574453;
assign addr[19656]= -2093641749;
assign addr[19657]= -2140281282;
assign addr[19658]= -2143547897;
assign addr[19659]= -2103375398;
assign addr[19660]= -2020577882;
assign addr[19661]= -1896833245;
assign addr[19662]= -1734649179;
assign addr[19663]= -1537312353;
assign addr[19664]= -1308821808;
assign addr[19665]= -1053807919;
assign addr[19666]= -777438554;
assign addr[19667]= -485314355;
assign addr[19668]= -183355234;
assign addr[19669]= 122319591;
assign addr[19670]= 425515602;
assign addr[19671]= 720088517;
assign addr[19672]= 1000068799;
assign addr[19673]= 1259782632;
assign addr[19674]= 1493966902;
assign addr[19675]= 1697875851;
assign addr[19676]= 1867377253;
assign addr[19677]= 1999036154;
assign addr[19678]= 2090184478;
assign addr[19679]= 2138975100;
assign addr[19680]= 2144419275;
assign addr[19681]= 2106406677;
assign addr[19682]= 2025707632;
assign addr[19683]= 1903957513;
assign addr[19684]= 1743623590;
assign addr[19685]= 1547955041;
assign addr[19686]= 1320917099;
assign addr[19687]= 1067110699;
assign addr[19688]= 791679244;
assign addr[19689]= 500204365;
assign addr[19690]= 198592817;
assign addr[19691]= -107043224;
assign addr[19692]= -410510029;
assign addr[19693]= -705657826;
assign addr[19694]= -986505429;
assign addr[19695]= -1247361445;
assign addr[19696]= -1482939614;
assign addr[19697]= -1688465931;
assign addr[19698]= -1859775393;
assign addr[19699]= -1993396407;
assign addr[19700]= -2086621133;
assign addr[19701]= -2137560369;
assign addr[19702]= -2145181827;
assign addr[19703]= -2109331059;
assign addr[19704]= -2030734582;
assign addr[19705]= -1910985158;
assign addr[19706]= -1752509516;
assign addr[19707]= -1558519173;
assign addr[19708]= -1332945355;
assign addr[19709]= -1080359326;
assign addr[19710]= -805879757;
assign addr[19711]= -515068990;
assign addr[19712]= -213820322;
assign addr[19713]= 91761426;
assign addr[19714]= 395483624;
assign addr[19715]= 691191324;
assign addr[19716]= 972891995;
assign addr[19717]= 1234876957;
assign addr[19718]= 1471837070;
assign addr[19719]= 1678970324;
assign addr[19720]= 1852079154;
assign addr[19721]= 1987655498;
assign addr[19722]= 2082951896;
assign addr[19723]= 2136037160;
assign addr[19724]= 2145835515;
assign addr[19725]= 2112148396;
assign addr[19726]= 2035658475;
assign addr[19727]= 1917915825;
assign addr[19728]= 1761306505;
assign addr[19729]= 1569004214;
assign addr[19730]= 1344905966;
assign addr[19731]= 1093553126;
assign addr[19732]= 820039373;
assign addr[19733]= 529907477;
assign addr[19734]= 229036977;
assign addr[19735]= -76474970;
assign addr[19736]= -380437148;
assign addr[19737]= -676689746;
assign addr[19738]= -959229189;
assign addr[19739]= -1222329801;
assign addr[19740]= -1460659832;
assign addr[19741]= -1669389513;
assign addr[19742]= -1844288924;
assign addr[19743]= -1981813720;
assign addr[19744]= -2079176953;
assign addr[19745]= -2134405552;
assign addr[19746]= -2146380306;
assign addr[19747]= -2114858546;
assign addr[19748]= -2040479063;
assign addr[19749]= -1924749160;
assign addr[19750]= -1770014111;
assign addr[19751]= -1579409630;
assign addr[19752]= -1356798326;
assign addr[19753]= -1106691431;
assign addr[19754]= -834157373;
assign addr[19755]= -544719071;
assign addr[19756]= -244242007;
assign addr[19757]= 61184634;
assign addr[19758]= 365371365;
assign addr[19759]= 662153826;
assign addr[19760]= 945517704;
assign addr[19761]= 1209720613;
assign addr[19762]= 1449408469;
assign addr[19763]= 1659723983;
assign addr[19764]= 1836405100;
assign addr[19765]= 1975871368;
assign addr[19766]= 2075296495;
assign addr[19767]= 2132665626;
assign addr[19768]= 2146816171;
assign addr[19769]= 2117461370;
assign addr[19770]= 2045196100;
assign addr[19771]= 1931484818;
assign addr[19772]= 1778631892;
assign addr[19773]= 1589734894;
assign addr[19774]= 1368621831;
assign addr[19775]= 1119773573;
assign addr[19776]= 848233042;
assign addr[19777]= 559503022;
assign addr[19778]= 259434643;
assign addr[19779]= -45891193;
assign addr[19780]= -350287041;
assign addr[19781]= -647584304;
assign addr[19782]= -931758235;
assign addr[19783]= -1197050035;
assign addr[19784]= -1438083551;
assign addr[19785]= -1649974225;
assign addr[19786]= -1828428082;
assign addr[19787]= -1969828744;
assign addr[19788]= -2071310720;
assign addr[19789]= -2130817471;
assign addr[19790]= -2147143090;
assign addr[19791]= -2119956737;
assign addr[19792]= -2049809346;
assign addr[19793]= -1938122457;
assign addr[19794]= -1787159411;
assign addr[19795]= -1599979481;
assign addr[19796]= -1380375881;
assign addr[19797]= -1132798888;
assign addr[19798]= -862265664;
assign addr[19799]= -574258580;
assign addr[19800]= -274614114;
assign addr[19801]= 30595422;
assign addr[19802]= 335184940;
assign addr[19803]= 632981917;
assign addr[19804]= 917951481;
assign addr[19805]= 1184318708;
assign addr[19806]= 1426685652;
assign addr[19807]= 1640140734;
assign addr[19808]= 1820358275;
assign addr[19809]= 1963686155;
assign addr[19810]= 2067219829;
assign addr[19811]= 2128861181;
assign addr[19812]= 2147361045;
assign addr[19813]= 2122344521;
assign addr[19814]= 2054318569;
assign addr[19815]= 1944661739;
assign addr[19816]= 1795596234;
assign addr[19817]= 1610142873;
assign addr[19818]= 1392059879;
assign addr[19819]= 1145766716;
assign addr[19820]= 876254528;
assign addr[19821]= 588984994;
assign addr[19822]= 289779648;
assign addr[19823]= -15298099;
assign addr[19824]= -320065829;
assign addr[19825]= -618347408;
assign addr[19826]= -904098143;
assign addr[19827]= -1171527280;
assign addr[19828]= -1415215352;
assign addr[19829]= -1630224009;
assign addr[19830]= -1812196087;
assign addr[19831]= -1957443913;
assign addr[19832]= -2063024031;
assign addr[19833]= -2126796855;
assign addr[19834]= -2147470025;
assign addr[19835]= -2124624598;
assign addr[19836]= -2058723538;
assign addr[19837]= -1951102334;
assign addr[19838]= -1803941934;
assign addr[19839]= -1620224553;
assign addr[19840]= -1403673233;
assign addr[19841]= -1158676398;
assign addr[19842]= -890198924;
assign addr[19843]= -603681519;
assign addr[19844]= -304930476;
assign addr[19845]= 0;
assign addr[19846]= 304930476;
assign addr[19847]= 603681519;
assign addr[19848]= 890198924;
assign addr[19849]= 1158676398;
assign addr[19850]= 1403673233;
assign addr[19851]= 1620224553;
assign addr[19852]= 1803941934;
assign addr[19853]= 1951102334;
assign addr[19854]= 2058723538;
assign addr[19855]= 2124624598;
assign addr[19856]= 2147470025;
assign addr[19857]= 2126796855;
assign addr[19858]= 2063024031;
assign addr[19859]= 1957443913;
assign addr[19860]= 1812196087;
assign addr[19861]= 1630224009;
assign addr[19862]= 1415215352;
assign addr[19863]= 1171527280;
assign addr[19864]= 904098143;
assign addr[19865]= 618347408;
assign addr[19866]= 320065829;
assign addr[19867]= 15298099;
assign addr[19868]= -289779648;
assign addr[19869]= -588984994;
assign addr[19870]= -876254528;
assign addr[19871]= -1145766716;
assign addr[19872]= -1392059879;
assign addr[19873]= -1610142873;
assign addr[19874]= -1795596234;
assign addr[19875]= -1944661739;
assign addr[19876]= -2054318569;
assign addr[19877]= -2122344521;
assign addr[19878]= -2147361045;
assign addr[19879]= -2128861181;
assign addr[19880]= -2067219829;
assign addr[19881]= -1963686155;
assign addr[19882]= -1820358275;
assign addr[19883]= -1640140734;
assign addr[19884]= -1426685652;
assign addr[19885]= -1184318708;
assign addr[19886]= -917951481;
assign addr[19887]= -632981917;
assign addr[19888]= -335184940;
assign addr[19889]= -30595422;
assign addr[19890]= 274614114;
assign addr[19891]= 574258580;
assign addr[19892]= 862265664;
assign addr[19893]= 1132798888;
assign addr[19894]= 1380375881;
assign addr[19895]= 1599979481;
assign addr[19896]= 1787159411;
assign addr[19897]= 1938122457;
assign addr[19898]= 2049809346;
assign addr[19899]= 2119956737;
assign addr[19900]= 2147143090;
assign addr[19901]= 2130817471;
assign addr[19902]= 2071310720;
assign addr[19903]= 1969828744;
assign addr[19904]= 1828428082;
assign addr[19905]= 1649974225;
assign addr[19906]= 1438083551;
assign addr[19907]= 1197050035;
assign addr[19908]= 931758235;
assign addr[19909]= 647584304;
assign addr[19910]= 350287041;
assign addr[19911]= 45891193;
assign addr[19912]= -259434643;
assign addr[19913]= -559503022;
assign addr[19914]= -848233042;
assign addr[19915]= -1119773573;
assign addr[19916]= -1368621831;
assign addr[19917]= -1589734894;
assign addr[19918]= -1778631892;
assign addr[19919]= -1931484818;
assign addr[19920]= -2045196100;
assign addr[19921]= -2117461370;
assign addr[19922]= -2146816171;
assign addr[19923]= -2132665626;
assign addr[19924]= -2075296495;
assign addr[19925]= -1975871368;
assign addr[19926]= -1836405100;
assign addr[19927]= -1659723983;
assign addr[19928]= -1449408469;
assign addr[19929]= -1209720613;
assign addr[19930]= -945517704;
assign addr[19931]= -662153826;
assign addr[19932]= -365371365;
assign addr[19933]= -61184634;
assign addr[19934]= 244242007;
assign addr[19935]= 544719071;
assign addr[19936]= 834157373;
assign addr[19937]= 1106691431;
assign addr[19938]= 1356798326;
assign addr[19939]= 1579409630;
assign addr[19940]= 1770014111;
assign addr[19941]= 1924749160;
assign addr[19942]= 2040479063;
assign addr[19943]= 2114858546;
assign addr[19944]= 2146380306;
assign addr[19945]= 2134405552;
assign addr[19946]= 2079176953;
assign addr[19947]= 1981813720;
assign addr[19948]= 1844288924;
assign addr[19949]= 1669389513;
assign addr[19950]= 1460659832;
assign addr[19951]= 1222329801;
assign addr[19952]= 959229189;
assign addr[19953]= 676689746;
assign addr[19954]= 380437148;
assign addr[19955]= 76474970;
assign addr[19956]= -229036977;
assign addr[19957]= -529907477;
assign addr[19958]= -820039373;
assign addr[19959]= -1093553126;
assign addr[19960]= -1344905966;
assign addr[19961]= -1569004214;
assign addr[19962]= -1761306505;
assign addr[19963]= -1917915825;
assign addr[19964]= -2035658475;
assign addr[19965]= -2112148396;
assign addr[19966]= -2145835515;
assign addr[19967]= -2136037160;
assign addr[19968]= -2082951896;
assign addr[19969]= -1987655498;
assign addr[19970]= -1852079154;
assign addr[19971]= -1678970324;
assign addr[19972]= -1471837070;
assign addr[19973]= -1234876957;
assign addr[19974]= -972891995;
assign addr[19975]= -691191324;
assign addr[19976]= -395483624;
assign addr[19977]= -91761426;
assign addr[19978]= 213820322;
assign addr[19979]= 515068990;
assign addr[19980]= 805879757;
assign addr[19981]= 1080359326;
assign addr[19982]= 1332945355;
assign addr[19983]= 1558519173;
assign addr[19984]= 1752509516;
assign addr[19985]= 1910985158;
assign addr[19986]= 2030734582;
assign addr[19987]= 2109331059;
assign addr[19988]= 2145181827;
assign addr[19989]= 2137560369;
assign addr[19990]= 2086621133;
assign addr[19991]= 1993396407;
assign addr[19992]= 1859775393;
assign addr[19993]= 1688465931;
assign addr[19994]= 1482939614;
assign addr[19995]= 1247361445;
assign addr[19996]= 986505429;
assign addr[19997]= 705657826;
assign addr[19998]= 410510029;
assign addr[19999]= 107043224;
assign addr[20000]= -198592817;
assign addr[20001]= -500204365;
assign addr[20002]= -791679244;
assign addr[20003]= -1067110699;
assign addr[20004]= -1320917099;
assign addr[20005]= -1547955041;
assign addr[20006]= -1743623590;
assign addr[20007]= -1903957513;
assign addr[20008]= -2025707632;
assign addr[20009]= -2106406677;
assign addr[20010]= -2144419275;
assign addr[20011]= -2138975100;
assign addr[20012]= -2090184478;
assign addr[20013]= -1999036154;
assign addr[20014]= -1867377253;
assign addr[20015]= -1697875851;
assign addr[20016]= -1493966902;
assign addr[20017]= -1259782632;
assign addr[20018]= -1000068799;
assign addr[20019]= -720088517;
assign addr[20020]= -425515602;
assign addr[20021]= -122319591;
assign addr[20022]= 183355234;
assign addr[20023]= 485314355;
assign addr[20024]= 777438554;
assign addr[20025]= 1053807919;
assign addr[20026]= 1308821808;
assign addr[20027]= 1537312353;
assign addr[20028]= 1734649179;
assign addr[20029]= 1896833245;
assign addr[20030]= 2020577882;
assign addr[20031]= 2103375398;
assign addr[20032]= 2143547897;
assign addr[20033]= 2140281282;
assign addr[20034]= 2093641749;
assign addr[20035]= 2004574453;
assign addr[20036]= 1874884346;
assign addr[20037]= 1707199606;
assign addr[20038]= 1504918373;
assign addr[20039]= 1272139887;
assign addr[20040]= 1013581418;
assign addr[20041]= 734482665;
assign addr[20042]= 440499581;
assign addr[20043]= 137589750;
assign addr[20044]= -168108346;
assign addr[20045]= -470399716;
assign addr[20046]= -763158411;
assign addr[20047]= -1040451659;
assign addr[20048]= -1296660098;
assign addr[20049]= -1526591649;
assign addr[20050]= -1725586737;
assign addr[20051]= -1889612716;
assign addr[20052]= -2015345591;
assign addr[20053]= -2100237377;
assign addr[20054]= -2142567738;
assign addr[20055]= -2141478848;
assign addr[20056]= -2096992772;
assign addr[20057]= -2010011024;
assign addr[20058]= -1882296293;
assign addr[20059]= -1716436725;
assign addr[20060]= -1515793473;
assign addr[20061]= -1284432584;
assign addr[20062]= -1027042599;
assign addr[20063]= -748839539;
assign addr[20064]= -455461206;
assign addr[20065]= -152852926;
assign addr[20066]= 152852926;
assign addr[20067]= 455461206;
assign addr[20068]= 748839539;
assign addr[20069]= 1027042599;
assign addr[20070]= 1284432584;
assign addr[20071]= 1515793473;
assign addr[20072]= 1716436725;
assign addr[20073]= 1882296293;
assign addr[20074]= 2010011024;
assign addr[20075]= 2096992772;
assign addr[20076]= 2141478848;
assign addr[20077]= 2142567738;
assign addr[20078]= 2100237377;
assign addr[20079]= 2015345591;
assign addr[20080]= 1889612716;
assign addr[20081]= 1725586737;
assign addr[20082]= 1526591649;
assign addr[20083]= 1296660098;
assign addr[20084]= 1040451659;
assign addr[20085]= 763158411;
assign addr[20086]= 470399716;
assign addr[20087]= 168108346;
assign addr[20088]= -137589750;
assign addr[20089]= -440499581;
assign addr[20090]= -734482665;
assign addr[20091]= -1013581418;
assign addr[20092]= -1272139887;
assign addr[20093]= -1504918373;
assign addr[20094]= -1707199606;
assign addr[20095]= -1874884346;
assign addr[20096]= -2004574453;
assign addr[20097]= -2093641749;
assign addr[20098]= -2140281282;
assign addr[20099]= -2143547897;
assign addr[20100]= -2103375398;
assign addr[20101]= -2020577882;
assign addr[20102]= -1896833245;
assign addr[20103]= -1734649179;
assign addr[20104]= -1537312353;
assign addr[20105]= -1308821808;
assign addr[20106]= -1053807919;
assign addr[20107]= -777438554;
assign addr[20108]= -485314355;
assign addr[20109]= -183355234;
assign addr[20110]= 122319591;
assign addr[20111]= 425515602;
assign addr[20112]= 720088517;
assign addr[20113]= 1000068799;
assign addr[20114]= 1259782632;
assign addr[20115]= 1493966902;
assign addr[20116]= 1697875851;
assign addr[20117]= 1867377253;
assign addr[20118]= 1999036154;
assign addr[20119]= 2090184478;
assign addr[20120]= 2138975100;
assign addr[20121]= 2144419275;
assign addr[20122]= 2106406677;
assign addr[20123]= 2025707632;
assign addr[20124]= 1903957513;
assign addr[20125]= 1743623590;
assign addr[20126]= 1547955041;
assign addr[20127]= 1320917099;
assign addr[20128]= 1067110699;
assign addr[20129]= 791679244;
assign addr[20130]= 500204365;
assign addr[20131]= 198592817;
assign addr[20132]= -107043224;
assign addr[20133]= -410510029;
assign addr[20134]= -705657826;
assign addr[20135]= -986505429;
assign addr[20136]= -1247361445;
assign addr[20137]= -1482939614;
assign addr[20138]= -1688465931;
assign addr[20139]= -1859775393;
assign addr[20140]= -1993396407;
assign addr[20141]= -2086621133;
assign addr[20142]= -2137560369;
assign addr[20143]= -2145181827;
assign addr[20144]= -2109331059;
assign addr[20145]= -2030734582;
assign addr[20146]= -1910985158;
assign addr[20147]= -1752509516;
assign addr[20148]= -1558519173;
assign addr[20149]= -1332945355;
assign addr[20150]= -1080359326;
assign addr[20151]= -805879757;
assign addr[20152]= -515068990;
assign addr[20153]= -213820322;
assign addr[20154]= 91761426;
assign addr[20155]= 395483624;
assign addr[20156]= 691191324;
assign addr[20157]= 972891995;
assign addr[20158]= 1234876957;
assign addr[20159]= 1471837070;
assign addr[20160]= 1678970324;
assign addr[20161]= 1852079154;
assign addr[20162]= 1987655498;
assign addr[20163]= 2082951896;
assign addr[20164]= 2136037160;
assign addr[20165]= 2145835515;
assign addr[20166]= 2112148396;
assign addr[20167]= 2035658475;
assign addr[20168]= 1917915825;
assign addr[20169]= 1761306505;
assign addr[20170]= 1569004214;
assign addr[20171]= 1344905966;
assign addr[20172]= 1093553126;
assign addr[20173]= 820039373;
assign addr[20174]= 529907477;
assign addr[20175]= 229036977;
assign addr[20176]= -76474970;
assign addr[20177]= -380437148;
assign addr[20178]= -676689746;
assign addr[20179]= -959229189;
assign addr[20180]= -1222329801;
assign addr[20181]= -1460659832;
assign addr[20182]= -1669389513;
assign addr[20183]= -1844288924;
assign addr[20184]= -1981813720;
assign addr[20185]= -2079176953;
assign addr[20186]= -2134405552;
assign addr[20187]= -2146380306;
assign addr[20188]= -2114858546;
assign addr[20189]= -2040479063;
assign addr[20190]= -1924749160;
assign addr[20191]= -1770014111;
assign addr[20192]= -1579409630;
assign addr[20193]= -1356798326;
assign addr[20194]= -1106691431;
assign addr[20195]= -834157373;
assign addr[20196]= -544719071;
assign addr[20197]= -244242007;
assign addr[20198]= 61184634;
assign addr[20199]= 365371365;
assign addr[20200]= 662153826;
assign addr[20201]= 945517704;
assign addr[20202]= 1209720613;
assign addr[20203]= 1449408469;
assign addr[20204]= 1659723983;
assign addr[20205]= 1836405100;
assign addr[20206]= 1975871368;
assign addr[20207]= 2075296495;
assign addr[20208]= 2132665626;
assign addr[20209]= 2146816171;
assign addr[20210]= 2117461370;
assign addr[20211]= 2045196100;
assign addr[20212]= 1931484818;
assign addr[20213]= 1778631892;
assign addr[20214]= 1589734894;
assign addr[20215]= 1368621831;
assign addr[20216]= 1119773573;
assign addr[20217]= 848233042;
assign addr[20218]= 559503022;
assign addr[20219]= 259434643;
assign addr[20220]= -45891193;
assign addr[20221]= -350287041;
assign addr[20222]= -647584304;
assign addr[20223]= -931758235;
assign addr[20224]= -1197050035;
assign addr[20225]= -1438083551;
assign addr[20226]= -1649974225;
assign addr[20227]= -1828428082;
assign addr[20228]= -1969828744;
assign addr[20229]= -2071310720;
assign addr[20230]= -2130817471;
assign addr[20231]= -2147143090;
assign addr[20232]= -2119956737;
assign addr[20233]= -2049809346;
assign addr[20234]= -1938122457;
assign addr[20235]= -1787159411;
assign addr[20236]= -1599979481;
assign addr[20237]= -1380375881;
assign addr[20238]= -1132798888;
assign addr[20239]= -862265664;
assign addr[20240]= -574258580;
assign addr[20241]= -274614114;
assign addr[20242]= 30595422;
assign addr[20243]= 335184940;
assign addr[20244]= 632981917;
assign addr[20245]= 917951481;
assign addr[20246]= 1184318708;
assign addr[20247]= 1426685652;
assign addr[20248]= 1640140734;
assign addr[20249]= 1820358275;
assign addr[20250]= 1963686155;
assign addr[20251]= 2067219829;
assign addr[20252]= 2128861181;
assign addr[20253]= 2147361045;
assign addr[20254]= 2122344521;
assign addr[20255]= 2054318569;
assign addr[20256]= 1944661739;
assign addr[20257]= 1795596234;
assign addr[20258]= 1610142873;
assign addr[20259]= 1392059879;
assign addr[20260]= 1145766716;
assign addr[20261]= 876254528;
assign addr[20262]= 588984994;
assign addr[20263]= 289779648;
assign addr[20264]= -15298099;
assign addr[20265]= -320065829;
assign addr[20266]= -618347408;
assign addr[20267]= -904098143;
assign addr[20268]= -1171527280;
assign addr[20269]= -1415215352;
assign addr[20270]= -1630224009;
assign addr[20271]= -1812196087;
assign addr[20272]= -1957443913;
assign addr[20273]= -2063024031;
assign addr[20274]= -2126796855;
assign addr[20275]= -2147470025;
assign addr[20276]= -2124624598;
assign addr[20277]= -2058723538;
assign addr[20278]= -1951102334;
assign addr[20279]= -1803941934;
assign addr[20280]= -1620224553;
assign addr[20281]= -1403673233;
assign addr[20282]= -1158676398;
assign addr[20283]= -890198924;
assign addr[20284]= -603681519;
assign addr[20285]= -304930476;
assign addr[20286]= 0;
assign addr[20287]= 304930476;
assign addr[20288]= 603681519;
assign addr[20289]= 890198924;
assign addr[20290]= 1158676398;
assign addr[20291]= 1403673233;
assign addr[20292]= 1620224553;
assign addr[20293]= 1803941934;
assign addr[20294]= 1951102334;
assign addr[20295]= 2058723538;
assign addr[20296]= 2124624598;
assign addr[20297]= 2147470025;
assign addr[20298]= 2126796855;
assign addr[20299]= 2063024031;
assign addr[20300]= 1957443913;
assign addr[20301]= 1812196087;
assign addr[20302]= 1630224009;
assign addr[20303]= 1415215352;
assign addr[20304]= 1171527280;
assign addr[20305]= 904098143;
assign addr[20306]= 618347408;
assign addr[20307]= 320065829;
assign addr[20308]= 15298099;
assign addr[20309]= -289779648;
assign addr[20310]= -588984994;
assign addr[20311]= -876254528;
assign addr[20312]= -1145766716;
assign addr[20313]= -1392059879;
assign addr[20314]= -1610142873;
assign addr[20315]= -1795596234;
assign addr[20316]= -1944661739;
assign addr[20317]= -2054318569;
assign addr[20318]= -2122344521;
assign addr[20319]= -2147361045;
assign addr[20320]= -2128861181;
assign addr[20321]= -2067219829;
assign addr[20322]= -1963686155;
assign addr[20323]= -1820358275;
assign addr[20324]= -1640140734;
assign addr[20325]= -1426685652;
assign addr[20326]= -1184318708;
assign addr[20327]= -917951481;
assign addr[20328]= -632981917;
assign addr[20329]= -335184940;
assign addr[20330]= -30595422;
assign addr[20331]= 274614114;
assign addr[20332]= 574258580;
assign addr[20333]= 862265664;
assign addr[20334]= 1132798888;
assign addr[20335]= 1380375881;
assign addr[20336]= 1599979481;
assign addr[20337]= 1787159411;
assign addr[20338]= 1938122457;
assign addr[20339]= 2049809346;
assign addr[20340]= 2119956737;
assign addr[20341]= 2147143090;
assign addr[20342]= 2130817471;
assign addr[20343]= 2071310720;
assign addr[20344]= 1969828744;
assign addr[20345]= 1828428082;
assign addr[20346]= 1649974225;
assign addr[20347]= 1438083551;
assign addr[20348]= 1197050035;
assign addr[20349]= 931758235;
assign addr[20350]= 647584304;
assign addr[20351]= 350287041;
assign addr[20352]= 45891193;
assign addr[20353]= -259434643;
assign addr[20354]= -559503022;
assign addr[20355]= -848233042;
assign addr[20356]= -1119773573;
assign addr[20357]= -1368621831;
assign addr[20358]= -1589734894;
assign addr[20359]= -1778631892;
assign addr[20360]= -1931484818;
assign addr[20361]= -2045196100;
assign addr[20362]= -2117461370;
assign addr[20363]= -2146816171;
assign addr[20364]= -2132665626;
assign addr[20365]= -2075296495;
assign addr[20366]= -1975871368;
assign addr[20367]= -1836405100;
assign addr[20368]= -1659723983;
assign addr[20369]= -1449408469;
assign addr[20370]= -1209720613;
assign addr[20371]= -945517704;
assign addr[20372]= -662153826;
assign addr[20373]= -365371365;
assign addr[20374]= -61184634;
assign addr[20375]= 244242007;
assign addr[20376]= 544719071;
assign addr[20377]= 834157373;
assign addr[20378]= 1106691431;
assign addr[20379]= 1356798326;
assign addr[20380]= 1579409630;
assign addr[20381]= 1770014111;
assign addr[20382]= 1924749160;
assign addr[20383]= 2040479063;
assign addr[20384]= 2114858546;
assign addr[20385]= 2146380306;
assign addr[20386]= 2134405552;
assign addr[20387]= 2079176953;
assign addr[20388]= 1981813720;
assign addr[20389]= 1844288924;
assign addr[20390]= 1669389513;
assign addr[20391]= 1460659832;
assign addr[20392]= 1222329801;
assign addr[20393]= 959229189;
assign addr[20394]= 676689746;
assign addr[20395]= 380437148;
assign addr[20396]= 76474970;
assign addr[20397]= -229036977;
assign addr[20398]= -529907477;
assign addr[20399]= -820039373;
assign addr[20400]= -1093553126;
assign addr[20401]= -1344905966;
assign addr[20402]= -1569004214;
assign addr[20403]= -1761306505;
assign addr[20404]= -1917915825;
assign addr[20405]= -2035658475;
assign addr[20406]= -2112148396;
assign addr[20407]= -2145835515;
assign addr[20408]= -2136037160;
assign addr[20409]= -2082951896;
assign addr[20410]= -1987655498;
assign addr[20411]= -1852079154;
assign addr[20412]= -1678970324;
assign addr[20413]= -1471837070;
assign addr[20414]= -1234876957;
assign addr[20415]= -972891995;
assign addr[20416]= -691191324;
assign addr[20417]= -395483624;
assign addr[20418]= -91761426;
assign addr[20419]= 213820322;
assign addr[20420]= 515068990;
assign addr[20421]= 805879757;
assign addr[20422]= 1080359326;
assign addr[20423]= 1332945355;
assign addr[20424]= 1558519173;
assign addr[20425]= 1752509516;
assign addr[20426]= 1910985158;
assign addr[20427]= 2030734582;
assign addr[20428]= 2109331059;
assign addr[20429]= 2145181827;
assign addr[20430]= 2137560369;
assign addr[20431]= 2086621133;
assign addr[20432]= 1993396407;
assign addr[20433]= 1859775393;
assign addr[20434]= 1688465931;
assign addr[20435]= 1482939614;
assign addr[20436]= 1247361445;
assign addr[20437]= 986505429;
assign addr[20438]= 705657826;
assign addr[20439]= 410510029;
assign addr[20440]= 107043224;
assign addr[20441]= -198592817;
assign addr[20442]= -500204365;
assign addr[20443]= -791679244;
assign addr[20444]= -1067110699;
assign addr[20445]= -1320917099;
assign addr[20446]= -1547955041;
assign addr[20447]= -1743623590;
assign addr[20448]= -1903957513;
assign addr[20449]= -2025707632;
assign addr[20450]= -2106406677;
assign addr[20451]= -2144419275;
assign addr[20452]= -2138975100;
assign addr[20453]= -2090184478;
assign addr[20454]= -1999036154;
assign addr[20455]= -1867377253;
assign addr[20456]= -1697875851;
assign addr[20457]= -1493966902;
assign addr[20458]= -1259782632;
assign addr[20459]= -1000068799;
assign addr[20460]= -720088517;
assign addr[20461]= -425515602;
assign addr[20462]= -122319591;
assign addr[20463]= 183355234;
assign addr[20464]= 485314355;
assign addr[20465]= 777438554;
assign addr[20466]= 1053807919;
assign addr[20467]= 1308821808;
assign addr[20468]= 1537312353;
assign addr[20469]= 1734649179;
assign addr[20470]= 1896833245;
assign addr[20471]= 2020577882;
assign addr[20472]= 2103375398;
assign addr[20473]= 2143547897;
assign addr[20474]= 2140281282;
assign addr[20475]= 2093641749;
assign addr[20476]= 2004574453;
assign addr[20477]= 1874884346;
assign addr[20478]= 1707199606;
assign addr[20479]= 1504918373;
assign addr[20480]= 1272139887;
assign addr[20481]= 1013581418;
assign addr[20482]= 734482665;
assign addr[20483]= 440499581;
assign addr[20484]= 137589750;
assign addr[20485]= -168108346;
assign addr[20486]= -470399716;
assign addr[20487]= -763158411;
assign addr[20488]= -1040451659;
assign addr[20489]= -1296660098;
assign addr[20490]= -1526591649;
assign addr[20491]= -1725586737;
assign addr[20492]= -1889612716;
assign addr[20493]= -2015345591;
assign addr[20494]= -2100237377;
assign addr[20495]= -2142567738;
assign addr[20496]= -2141478848;
assign addr[20497]= -2096992772;
assign addr[20498]= -2010011024;
assign addr[20499]= -1882296293;
assign addr[20500]= -1716436725;
assign addr[20501]= -1515793473;
assign addr[20502]= -1284432584;
assign addr[20503]= -1027042599;
assign addr[20504]= -748839539;
assign addr[20505]= -455461206;
assign addr[20506]= -152852926;
assign addr[20507]= 152852926;
assign addr[20508]= 455461206;
assign addr[20509]= 748839539;
assign addr[20510]= 1027042599;
assign addr[20511]= 1284432584;
assign addr[20512]= 1515793473;
assign addr[20513]= 1716436725;
assign addr[20514]= 1882296293;
assign addr[20515]= 2010011024;
assign addr[20516]= 2096992772;
assign addr[20517]= 2141478848;
assign addr[20518]= 2142567738;
assign addr[20519]= 2100237377;
assign addr[20520]= 2015345591;
assign addr[20521]= 1889612716;
assign addr[20522]= 1725586737;
assign addr[20523]= 1526591649;
assign addr[20524]= 1296660098;
assign addr[20525]= 1040451659;
assign addr[20526]= 763158411;
assign addr[20527]= 470399716;
assign addr[20528]= 168108346;
assign addr[20529]= -137589750;
assign addr[20530]= -440499581;
assign addr[20531]= -734482665;
assign addr[20532]= -1013581418;
assign addr[20533]= -1272139887;
assign addr[20534]= -1504918373;
assign addr[20535]= -1707199606;
assign addr[20536]= -1874884346;
assign addr[20537]= -2004574453;
assign addr[20538]= -2093641749;
assign addr[20539]= -2140281282;
assign addr[20540]= -2143547897;
assign addr[20541]= -2103375398;
assign addr[20542]= -2020577882;
assign addr[20543]= -1896833245;
assign addr[20544]= -1734649179;
assign addr[20545]= -1537312353;
assign addr[20546]= -1308821808;
assign addr[20547]= -1053807919;
assign addr[20548]= -777438554;
assign addr[20549]= -485314355;
assign addr[20550]= -183355234;
assign addr[20551]= 122319591;
assign addr[20552]= 425515602;
assign addr[20553]= 720088517;
assign addr[20554]= 1000068799;
assign addr[20555]= 1259782632;
assign addr[20556]= 1493966902;
assign addr[20557]= 1697875851;
assign addr[20558]= 1867377253;
assign addr[20559]= 1999036154;
assign addr[20560]= 2090184478;
assign addr[20561]= 2138975100;
assign addr[20562]= 2144419275;
assign addr[20563]= 2106406677;
assign addr[20564]= 2025707632;
assign addr[20565]= 1903957513;
assign addr[20566]= 1743623590;
assign addr[20567]= 1547955041;
assign addr[20568]= 1320917099;
assign addr[20569]= 1067110699;
assign addr[20570]= 791679244;
assign addr[20571]= 500204365;
assign addr[20572]= 198592817;
assign addr[20573]= -107043224;
assign addr[20574]= -410510029;
assign addr[20575]= -705657826;
assign addr[20576]= -986505429;
assign addr[20577]= -1247361445;
assign addr[20578]= -1482939614;
assign addr[20579]= -1688465931;
assign addr[20580]= -1859775393;
assign addr[20581]= -1993396407;
assign addr[20582]= -2086621133;
assign addr[20583]= -2137560369;
assign addr[20584]= -2145181827;
assign addr[20585]= -2109331059;
assign addr[20586]= -2030734582;
assign addr[20587]= -1910985158;
assign addr[20588]= -1752509516;
assign addr[20589]= -1558519173;
assign addr[20590]= -1332945355;
assign addr[20591]= -1080359326;
assign addr[20592]= -805879757;
assign addr[20593]= -515068990;
assign addr[20594]= -213820322;
assign addr[20595]= 91761426;
assign addr[20596]= 395483624;
assign addr[20597]= 691191324;
assign addr[20598]= 972891995;
assign addr[20599]= 1234876957;
assign addr[20600]= 1471837070;
assign addr[20601]= 1678970324;
assign addr[20602]= 1852079154;
assign addr[20603]= 1987655498;
assign addr[20604]= 2082951896;
assign addr[20605]= 2136037160;
assign addr[20606]= 2145835515;
assign addr[20607]= 2112148396;
assign addr[20608]= 2035658475;
assign addr[20609]= 1917915825;
assign addr[20610]= 1761306505;
assign addr[20611]= 1569004214;
assign addr[20612]= 1344905966;
assign addr[20613]= 1093553126;
assign addr[20614]= 820039373;
assign addr[20615]= 529907477;
assign addr[20616]= 229036977;
assign addr[20617]= -76474970;
assign addr[20618]= -380437148;
assign addr[20619]= -676689746;
assign addr[20620]= -959229189;
assign addr[20621]= -1222329801;
assign addr[20622]= -1460659832;
assign addr[20623]= -1669389513;
assign addr[20624]= -1844288924;
assign addr[20625]= -1981813720;
assign addr[20626]= -2079176953;
assign addr[20627]= -2134405552;
assign addr[20628]= -2146380306;
assign addr[20629]= -2114858546;
assign addr[20630]= -2040479063;
assign addr[20631]= -1924749160;
assign addr[20632]= -1770014111;
assign addr[20633]= -1579409630;
assign addr[20634]= -1356798326;
assign addr[20635]= -1106691431;
assign addr[20636]= -834157373;
assign addr[20637]= -544719071;
assign addr[20638]= -244242007;
assign addr[20639]= 61184634;
assign addr[20640]= 365371365;
assign addr[20641]= 662153826;
assign addr[20642]= 945517704;
assign addr[20643]= 1209720613;
assign addr[20644]= 1449408469;
assign addr[20645]= 1659723983;
assign addr[20646]= 1836405100;
assign addr[20647]= 1975871368;
assign addr[20648]= 2075296495;
assign addr[20649]= 2132665626;
assign addr[20650]= 2146816171;
assign addr[20651]= 2117461370;
assign addr[20652]= 2045196100;
assign addr[20653]= 1931484818;
assign addr[20654]= 1778631892;
assign addr[20655]= 1589734894;
assign addr[20656]= 1368621831;
assign addr[20657]= 1119773573;
assign addr[20658]= 848233042;
assign addr[20659]= 559503022;
assign addr[20660]= 259434643;
assign addr[20661]= -45891193;
assign addr[20662]= -350287041;
assign addr[20663]= -647584304;
assign addr[20664]= -931758235;
assign addr[20665]= -1197050035;
assign addr[20666]= -1438083551;
assign addr[20667]= -1649974225;
assign addr[20668]= -1828428082;
assign addr[20669]= -1969828744;
assign addr[20670]= -2071310720;
assign addr[20671]= -2130817471;
assign addr[20672]= -2147143090;
assign addr[20673]= -2119956737;
assign addr[20674]= -2049809346;
assign addr[20675]= -1938122457;
assign addr[20676]= -1787159411;
assign addr[20677]= -1599979481;
assign addr[20678]= -1380375881;
assign addr[20679]= -1132798888;
assign addr[20680]= -862265664;
assign addr[20681]= -574258580;
assign addr[20682]= -274614114;
assign addr[20683]= 30595422;
assign addr[20684]= 335184940;
assign addr[20685]= 632981917;
assign addr[20686]= 917951481;
assign addr[20687]= 1184318708;
assign addr[20688]= 1426685652;
assign addr[20689]= 1640140734;
assign addr[20690]= 1820358275;
assign addr[20691]= 1963686155;
assign addr[20692]= 2067219829;
assign addr[20693]= 2128861181;
assign addr[20694]= 2147361045;
assign addr[20695]= 2122344521;
assign addr[20696]= 2054318569;
assign addr[20697]= 1944661739;
assign addr[20698]= 1795596234;
assign addr[20699]= 1610142873;
assign addr[20700]= 1392059879;
assign addr[20701]= 1145766716;
assign addr[20702]= 876254528;
assign addr[20703]= 588984994;
assign addr[20704]= 289779648;
assign addr[20705]= -15298099;
assign addr[20706]= -320065829;
assign addr[20707]= -618347408;
assign addr[20708]= -904098143;
assign addr[20709]= -1171527280;
assign addr[20710]= -1415215352;
assign addr[20711]= -1630224009;
assign addr[20712]= -1812196087;
assign addr[20713]= -1957443913;
assign addr[20714]= -2063024031;
assign addr[20715]= -2126796855;
assign addr[20716]= -2147470025;
assign addr[20717]= -2124624598;
assign addr[20718]= -2058723538;
assign addr[20719]= -1951102334;
assign addr[20720]= -1803941934;
assign addr[20721]= -1620224553;
assign addr[20722]= -1403673233;
assign addr[20723]= -1158676398;
assign addr[20724]= -890198924;
assign addr[20725]= -603681519;
assign addr[20726]= -304930476;
assign addr[20727]= 0;
assign addr[20728]= 304930476;
assign addr[20729]= 603681519;
assign addr[20730]= 890198924;
assign addr[20731]= 1158676398;
assign addr[20732]= 1403673233;
assign addr[20733]= 1620224553;
assign addr[20734]= 1803941934;
assign addr[20735]= 1951102334;
assign addr[20736]= 2058723538;
assign addr[20737]= 2124624598;
assign addr[20738]= 2147470025;
assign addr[20739]= 2126796855;
assign addr[20740]= 2063024031;
assign addr[20741]= 1957443913;
assign addr[20742]= 1812196087;
assign addr[20743]= 1630224009;
assign addr[20744]= 1415215352;
assign addr[20745]= 1171527280;
assign addr[20746]= 904098143;
assign addr[20747]= 618347408;
assign addr[20748]= 320065829;
assign addr[20749]= 15298099;
assign addr[20750]= -289779648;
assign addr[20751]= -588984994;
assign addr[20752]= -876254528;
assign addr[20753]= -1145766716;
assign addr[20754]= -1392059879;
assign addr[20755]= -1610142873;
assign addr[20756]= -1795596234;
assign addr[20757]= -1944661739;
assign addr[20758]= -2054318569;
assign addr[20759]= -2122344521;
assign addr[20760]= -2147361045;
assign addr[20761]= -2128861181;
assign addr[20762]= -2067219829;
assign addr[20763]= -1963686155;
assign addr[20764]= -1820358275;
assign addr[20765]= -1640140734;
assign addr[20766]= -1426685652;
assign addr[20767]= -1184318708;
assign addr[20768]= -917951481;
assign addr[20769]= -632981917;
assign addr[20770]= -335184940;
assign addr[20771]= -30595422;
assign addr[20772]= 274614114;
assign addr[20773]= 574258580;
assign addr[20774]= 862265664;
assign addr[20775]= 1132798888;
assign addr[20776]= 1380375881;
assign addr[20777]= 1599979481;
assign addr[20778]= 1787159411;
assign addr[20779]= 1938122457;
assign addr[20780]= 2049809346;
assign addr[20781]= 2119956737;
assign addr[20782]= 2147143090;
assign addr[20783]= 2130817471;
assign addr[20784]= 2071310720;
assign addr[20785]= 1969828744;
assign addr[20786]= 1828428082;
assign addr[20787]= 1649974225;
assign addr[20788]= 1438083551;
assign addr[20789]= 1197050035;
assign addr[20790]= 931758235;
assign addr[20791]= 647584304;
assign addr[20792]= 350287041;
assign addr[20793]= 45891193;
assign addr[20794]= -259434643;
assign addr[20795]= -559503022;
assign addr[20796]= -848233042;
assign addr[20797]= -1119773573;
assign addr[20798]= -1368621831;
assign addr[20799]= -1589734894;
assign addr[20800]= -1778631892;
assign addr[20801]= -1931484818;
assign addr[20802]= -2045196100;
assign addr[20803]= -2117461370;
assign addr[20804]= -2146816171;
assign addr[20805]= -2132665626;
assign addr[20806]= -2075296495;
assign addr[20807]= -1975871368;
assign addr[20808]= -1836405100;
assign addr[20809]= -1659723983;
assign addr[20810]= -1449408469;
assign addr[20811]= -1209720613;
assign addr[20812]= -945517704;
assign addr[20813]= -662153826;
assign addr[20814]= -365371365;
assign addr[20815]= -61184634;
assign addr[20816]= 244242007;
assign addr[20817]= 544719071;
assign addr[20818]= 834157373;
assign addr[20819]= 1106691431;
assign addr[20820]= 1356798326;
assign addr[20821]= 1579409630;
assign addr[20822]= 1770014111;
assign addr[20823]= 1924749160;
assign addr[20824]= 2040479063;
assign addr[20825]= 2114858546;
assign addr[20826]= 2146380306;
assign addr[20827]= 2134405552;
assign addr[20828]= 2079176953;
assign addr[20829]= 1981813720;
assign addr[20830]= 1844288924;
assign addr[20831]= 1669389513;
assign addr[20832]= 1460659832;
assign addr[20833]= 1222329801;
assign addr[20834]= 959229189;
assign addr[20835]= 676689746;
assign addr[20836]= 380437148;
assign addr[20837]= 76474970;
assign addr[20838]= -229036977;
assign addr[20839]= -529907477;
assign addr[20840]= -820039373;
assign addr[20841]= -1093553126;
assign addr[20842]= -1344905966;
assign addr[20843]= -1569004214;
assign addr[20844]= -1761306505;
assign addr[20845]= -1917915825;
assign addr[20846]= -2035658475;
assign addr[20847]= -2112148396;
assign addr[20848]= -2145835515;
assign addr[20849]= -2136037160;
assign addr[20850]= -2082951896;
assign addr[20851]= -1987655498;
assign addr[20852]= -1852079154;
assign addr[20853]= -1678970324;
assign addr[20854]= -1471837070;
assign addr[20855]= -1234876957;
assign addr[20856]= -972891995;
assign addr[20857]= -691191324;
assign addr[20858]= -395483624;
assign addr[20859]= -91761426;
assign addr[20860]= 213820322;
assign addr[20861]= 515068990;
assign addr[20862]= 805879757;
assign addr[20863]= 1080359326;
assign addr[20864]= 1332945355;
assign addr[20865]= 1558519173;
assign addr[20866]= 1752509516;
assign addr[20867]= 1910985158;
assign addr[20868]= 2030734582;
assign addr[20869]= 2109331059;
assign addr[20870]= 2145181827;
assign addr[20871]= 2137560369;
assign addr[20872]= 2086621133;
assign addr[20873]= 1993396407;
assign addr[20874]= 1859775393;
assign addr[20875]= 1688465931;
assign addr[20876]= 1482939614;
assign addr[20877]= 1247361445;
assign addr[20878]= 986505429;
assign addr[20879]= 705657826;
assign addr[20880]= 410510029;
assign addr[20881]= 107043224;
assign addr[20882]= -198592817;
assign addr[20883]= -500204365;
assign addr[20884]= -791679244;
assign addr[20885]= -1067110699;
assign addr[20886]= -1320917099;
assign addr[20887]= -1547955041;
assign addr[20888]= -1743623590;
assign addr[20889]= -1903957513;
assign addr[20890]= -2025707632;
assign addr[20891]= -2106406677;
assign addr[20892]= -2144419275;
assign addr[20893]= -2138975100;
assign addr[20894]= -2090184478;
assign addr[20895]= -1999036154;
assign addr[20896]= -1867377253;
assign addr[20897]= -1697875851;
assign addr[20898]= -1493966902;
assign addr[20899]= -1259782632;
assign addr[20900]= -1000068799;
assign addr[20901]= -720088517;
assign addr[20902]= -425515602;
assign addr[20903]= -122319591;
assign addr[20904]= 183355234;
assign addr[20905]= 485314355;
assign addr[20906]= 777438554;
assign addr[20907]= 1053807919;
assign addr[20908]= 1308821808;
assign addr[20909]= 1537312353;
assign addr[20910]= 1734649179;
assign addr[20911]= 1896833245;
assign addr[20912]= 2020577882;
assign addr[20913]= 2103375398;
assign addr[20914]= 2143547897;
assign addr[20915]= 2140281282;
assign addr[20916]= 2093641749;
assign addr[20917]= 2004574453;
assign addr[20918]= 1874884346;
assign addr[20919]= 1707199606;
assign addr[20920]= 1504918373;
assign addr[20921]= 1272139887;
assign addr[20922]= 1013581418;
assign addr[20923]= 734482665;
assign addr[20924]= 440499581;
assign addr[20925]= 137589750;
assign addr[20926]= -168108346;
assign addr[20927]= -470399716;
assign addr[20928]= -763158411;
assign addr[20929]= -1040451659;
assign addr[20930]= -1296660098;
assign addr[20931]= -1526591649;
assign addr[20932]= -1725586737;
assign addr[20933]= -1889612716;
assign addr[20934]= -2015345591;
assign addr[20935]= -2100237377;
assign addr[20936]= -2142567738;
assign addr[20937]= -2141478848;
assign addr[20938]= -2096992772;
assign addr[20939]= -2010011024;
assign addr[20940]= -1882296293;
assign addr[20941]= -1716436725;
assign addr[20942]= -1515793473;
assign addr[20943]= -1284432584;
assign addr[20944]= -1027042599;
assign addr[20945]= -748839539;
assign addr[20946]= -455461206;
assign addr[20947]= -152852926;
assign addr[20948]= 152852926;
assign addr[20949]= 455461206;
assign addr[20950]= 748839539;
assign addr[20951]= 1027042599;
assign addr[20952]= 1284432584;
assign addr[20953]= 1515793473;
assign addr[20954]= 1716436725;
assign addr[20955]= 1882296293;
assign addr[20956]= 2010011024;
assign addr[20957]= 2096992772;
assign addr[20958]= 2141478848;
assign addr[20959]= 2142567738;
assign addr[20960]= 2100237377;
assign addr[20961]= 2015345591;
assign addr[20962]= 1889612716;
assign addr[20963]= 1725586737;
assign addr[20964]= 1526591649;
assign addr[20965]= 1296660098;
assign addr[20966]= 1040451659;
assign addr[20967]= 763158411;
assign addr[20968]= 470399716;
assign addr[20969]= 168108346;
assign addr[20970]= -137589750;
assign addr[20971]= -440499581;
assign addr[20972]= -734482665;
assign addr[20973]= -1013581418;
assign addr[20974]= -1272139887;
assign addr[20975]= -1504918373;
assign addr[20976]= -1707199606;
assign addr[20977]= -1874884346;
assign addr[20978]= -2004574453;
assign addr[20979]= -2093641749;
assign addr[20980]= -2140281282;
assign addr[20981]= -2143547897;
assign addr[20982]= -2103375398;
assign addr[20983]= -2020577882;
assign addr[20984]= -1896833245;
assign addr[20985]= -1734649179;
assign addr[20986]= -1537312353;
assign addr[20987]= -1308821808;
assign addr[20988]= -1053807919;
assign addr[20989]= -777438554;
assign addr[20990]= -485314355;
assign addr[20991]= -183355234;
assign addr[20992]= 122319591;
assign addr[20993]= 425515602;
assign addr[20994]= 720088517;
assign addr[20995]= 1000068799;
assign addr[20996]= 1259782632;
assign addr[20997]= 1493966902;
assign addr[20998]= 1697875851;
assign addr[20999]= 1867377253;
assign addr[21000]= 1999036154;
assign addr[21001]= 2090184478;
assign addr[21002]= 2138975100;
assign addr[21003]= 2144419275;
assign addr[21004]= 2106406677;
assign addr[21005]= 2025707632;
assign addr[21006]= 1903957513;
assign addr[21007]= 1743623590;
assign addr[21008]= 1547955041;
assign addr[21009]= 1320917099;
assign addr[21010]= 1067110699;
assign addr[21011]= 791679244;
assign addr[21012]= 500204365;
assign addr[21013]= 198592817;
assign addr[21014]= -107043224;
assign addr[21015]= -410510029;
assign addr[21016]= -705657826;
assign addr[21017]= -986505429;
assign addr[21018]= -1247361445;
assign addr[21019]= -1482939614;
assign addr[21020]= -1688465931;
assign addr[21021]= -1859775393;
assign addr[21022]= -1993396407;
assign addr[21023]= -2086621133;
assign addr[21024]= -2137560369;
assign addr[21025]= -2145181827;
assign addr[21026]= -2109331059;
assign addr[21027]= -2030734582;
assign addr[21028]= -1910985158;
assign addr[21029]= -1752509516;
assign addr[21030]= -1558519173;
assign addr[21031]= -1332945355;
assign addr[21032]= -1080359326;
assign addr[21033]= -805879757;
assign addr[21034]= -515068990;
assign addr[21035]= -213820322;
assign addr[21036]= 91761426;
assign addr[21037]= 395483624;
assign addr[21038]= 691191324;
assign addr[21039]= 972891995;
assign addr[21040]= 1234876957;
assign addr[21041]= 1471837070;
assign addr[21042]= 1678970324;
assign addr[21043]= 1852079154;
assign addr[21044]= 1987655498;
assign addr[21045]= 2082951896;
assign addr[21046]= 2136037160;
assign addr[21047]= 2145835515;
assign addr[21048]= 2112148396;
assign addr[21049]= 2035658475;
assign addr[21050]= 1917915825;
assign addr[21051]= 1761306505;
assign addr[21052]= 1569004214;
assign addr[21053]= 1344905966;
assign addr[21054]= 1093553126;
assign addr[21055]= 820039373;
assign addr[21056]= 529907477;
assign addr[21057]= 229036977;
assign addr[21058]= -76474970;
assign addr[21059]= -380437148;
assign addr[21060]= -676689746;
assign addr[21061]= -959229189;
assign addr[21062]= -1222329801;
assign addr[21063]= -1460659832;
assign addr[21064]= -1669389513;
assign addr[21065]= -1844288924;
assign addr[21066]= -1981813720;
assign addr[21067]= -2079176953;
assign addr[21068]= -2134405552;
assign addr[21069]= -2146380306;
assign addr[21070]= -2114858546;
assign addr[21071]= -2040479063;
assign addr[21072]= -1924749160;
assign addr[21073]= -1770014111;
assign addr[21074]= -1579409630;
assign addr[21075]= -1356798326;
assign addr[21076]= -1106691431;
assign addr[21077]= -834157373;
assign addr[21078]= -544719071;
assign addr[21079]= -244242007;
assign addr[21080]= 61184634;
assign addr[21081]= 365371365;
assign addr[21082]= 662153826;
assign addr[21083]= 945517704;
assign addr[21084]= 1209720613;
assign addr[21085]= 1449408469;
assign addr[21086]= 1659723983;
assign addr[21087]= 1836405100;
assign addr[21088]= 1975871368;
assign addr[21089]= 2075296495;
assign addr[21090]= 2132665626;
assign addr[21091]= 2146816171;
assign addr[21092]= 2117461370;
assign addr[21093]= 2045196100;
assign addr[21094]= 1931484818;
assign addr[21095]= 1778631892;
assign addr[21096]= 1589734894;
assign addr[21097]= 1368621831;
assign addr[21098]= 1119773573;
assign addr[21099]= 848233042;
assign addr[21100]= 559503022;
assign addr[21101]= 259434643;
assign addr[21102]= -45891193;
assign addr[21103]= -350287041;
assign addr[21104]= -647584304;
assign addr[21105]= -931758235;
assign addr[21106]= -1197050035;
assign addr[21107]= -1438083551;
assign addr[21108]= -1649974225;
assign addr[21109]= -1828428082;
assign addr[21110]= -1969828744;
assign addr[21111]= -2071310720;
assign addr[21112]= -2130817471;
assign addr[21113]= -2147143090;
assign addr[21114]= -2119956737;
assign addr[21115]= -2049809346;
assign addr[21116]= -1938122457;
assign addr[21117]= -1787159411;
assign addr[21118]= -1599979481;
assign addr[21119]= -1380375881;
assign addr[21120]= -1132798888;
assign addr[21121]= -862265664;
assign addr[21122]= -574258580;
assign addr[21123]= -274614114;
assign addr[21124]= 30595422;
assign addr[21125]= 335184940;
assign addr[21126]= 632981917;
assign addr[21127]= 917951481;
assign addr[21128]= 1184318708;
assign addr[21129]= 1426685652;
assign addr[21130]= 1640140734;
assign addr[21131]= 1820358275;
assign addr[21132]= 1963686155;
assign addr[21133]= 2067219829;
assign addr[21134]= 2128861181;
assign addr[21135]= 2147361045;
assign addr[21136]= 2122344521;
assign addr[21137]= 2054318569;
assign addr[21138]= 1944661739;
assign addr[21139]= 1795596234;
assign addr[21140]= 1610142873;
assign addr[21141]= 1392059879;
assign addr[21142]= 1145766716;
assign addr[21143]= 876254528;
assign addr[21144]= 588984994;
assign addr[21145]= 289779648;
assign addr[21146]= -15298099;
assign addr[21147]= -320065829;
assign addr[21148]= -618347408;
assign addr[21149]= -904098143;
assign addr[21150]= -1171527280;
assign addr[21151]= -1415215352;
assign addr[21152]= -1630224009;
assign addr[21153]= -1812196087;
assign addr[21154]= -1957443913;
assign addr[21155]= -2063024031;
assign addr[21156]= -2126796855;
assign addr[21157]= -2147470025;
assign addr[21158]= -2124624598;
assign addr[21159]= -2058723538;
assign addr[21160]= -1951102334;
assign addr[21161]= -1803941934;
assign addr[21162]= -1620224553;
assign addr[21163]= -1403673233;
assign addr[21164]= -1158676398;
assign addr[21165]= -890198924;
assign addr[21166]= -603681519;
assign addr[21167]= -304930476;
assign addr[21168]= 0;
assign addr[21169]= 304930476;
assign addr[21170]= 603681519;
assign addr[21171]= 890198924;
assign addr[21172]= 1158676398;
assign addr[21173]= 1403673233;
assign addr[21174]= 1620224553;
assign addr[21175]= 1803941934;
assign addr[21176]= 1951102334;
assign addr[21177]= 2058723538;
assign addr[21178]= 2124624598;
assign addr[21179]= 2147470025;
assign addr[21180]= 2126796855;
assign addr[21181]= 2063024031;
assign addr[21182]= 1957443913;
assign addr[21183]= 1812196087;
assign addr[21184]= 1630224009;
assign addr[21185]= 1415215352;
assign addr[21186]= 1171527280;
assign addr[21187]= 904098143;
assign addr[21188]= 618347408;
assign addr[21189]= 320065829;
assign addr[21190]= 15298099;
assign addr[21191]= -289779648;
assign addr[21192]= -588984994;
assign addr[21193]= -876254528;
assign addr[21194]= -1145766716;
assign addr[21195]= -1392059879;
assign addr[21196]= -1610142873;
assign addr[21197]= -1795596234;
assign addr[21198]= -1944661739;
assign addr[21199]= -2054318569;
assign addr[21200]= -2122344521;
assign addr[21201]= -2147361045;
assign addr[21202]= -2128861181;
assign addr[21203]= -2067219829;
assign addr[21204]= -1963686155;
assign addr[21205]= -1820358275;
assign addr[21206]= -1640140734;
assign addr[21207]= -1426685652;
assign addr[21208]= -1184318708;
assign addr[21209]= -917951481;
assign addr[21210]= -632981917;
assign addr[21211]= -335184940;
assign addr[21212]= -30595422;
assign addr[21213]= 274614114;
assign addr[21214]= 574258580;
assign addr[21215]= 862265664;
assign addr[21216]= 1132798888;
assign addr[21217]= 1380375881;
assign addr[21218]= 1599979481;
assign addr[21219]= 1787159411;
assign addr[21220]= 1938122457;
assign addr[21221]= 2049809346;
assign addr[21222]= 2119956737;
assign addr[21223]= 2147143090;
assign addr[21224]= 2130817471;
assign addr[21225]= 2071310720;
assign addr[21226]= 1969828744;
assign addr[21227]= 1828428082;
assign addr[21228]= 1649974225;
assign addr[21229]= 1438083551;
assign addr[21230]= 1197050035;
assign addr[21231]= 931758235;
assign addr[21232]= 647584304;
assign addr[21233]= 350287041;
assign addr[21234]= 45891193;
assign addr[21235]= -259434643;
assign addr[21236]= -559503022;
assign addr[21237]= -848233042;
assign addr[21238]= -1119773573;
assign addr[21239]= -1368621831;
assign addr[21240]= -1589734894;
assign addr[21241]= -1778631892;
assign addr[21242]= -1931484818;
assign addr[21243]= -2045196100;
assign addr[21244]= -2117461370;
assign addr[21245]= -2146816171;
assign addr[21246]= -2132665626;
assign addr[21247]= -2075296495;
assign addr[21248]= -1975871368;
assign addr[21249]= -1836405100;
assign addr[21250]= -1659723983;
assign addr[21251]= -1449408469;
assign addr[21252]= -1209720613;
assign addr[21253]= -945517704;
assign addr[21254]= -662153826;
assign addr[21255]= -365371365;
assign addr[21256]= -61184634;
assign addr[21257]= 244242007;
assign addr[21258]= 544719071;
assign addr[21259]= 834157373;
assign addr[21260]= 1106691431;
assign addr[21261]= 1356798326;
assign addr[21262]= 1579409630;
assign addr[21263]= 1770014111;
assign addr[21264]= 1924749160;
assign addr[21265]= 2040479063;
assign addr[21266]= 2114858546;
assign addr[21267]= 2146380306;
assign addr[21268]= 2134405552;
assign addr[21269]= 2079176953;
assign addr[21270]= 1981813720;
assign addr[21271]= 1844288924;
assign addr[21272]= 1669389513;
assign addr[21273]= 1460659832;
assign addr[21274]= 1222329801;
assign addr[21275]= 959229189;
assign addr[21276]= 676689746;
assign addr[21277]= 380437148;
assign addr[21278]= 76474970;
assign addr[21279]= -229036977;
assign addr[21280]= -529907477;
assign addr[21281]= -820039373;
assign addr[21282]= -1093553126;
assign addr[21283]= -1344905966;
assign addr[21284]= -1569004214;
assign addr[21285]= -1761306505;
assign addr[21286]= -1917915825;
assign addr[21287]= -2035658475;
assign addr[21288]= -2112148396;
assign addr[21289]= -2145835515;
assign addr[21290]= -2136037160;
assign addr[21291]= -2082951896;
assign addr[21292]= -1987655498;
assign addr[21293]= -1852079154;
assign addr[21294]= -1678970324;
assign addr[21295]= -1471837070;
assign addr[21296]= -1234876957;
assign addr[21297]= -972891995;
assign addr[21298]= -691191324;
assign addr[21299]= -395483624;
assign addr[21300]= -91761426;
assign addr[21301]= 213820322;
assign addr[21302]= 515068990;
assign addr[21303]= 805879757;
assign addr[21304]= 1080359326;
assign addr[21305]= 1332945355;
assign addr[21306]= 1558519173;
assign addr[21307]= 1752509516;
assign addr[21308]= 1910985158;
assign addr[21309]= 2030734582;
assign addr[21310]= 2109331059;
assign addr[21311]= 2145181827;
assign addr[21312]= 2137560369;
assign addr[21313]= 2086621133;
assign addr[21314]= 1993396407;
assign addr[21315]= 1859775393;
assign addr[21316]= 1688465931;
assign addr[21317]= 1482939614;
assign addr[21318]= 1247361445;
assign addr[21319]= 986505429;
assign addr[21320]= 705657826;
assign addr[21321]= 410510029;
assign addr[21322]= 107043224;
assign addr[21323]= -198592817;
assign addr[21324]= -500204365;
assign addr[21325]= -791679244;
assign addr[21326]= -1067110699;
assign addr[21327]= -1320917099;
assign addr[21328]= -1547955041;
assign addr[21329]= -1743623590;
assign addr[21330]= -1903957513;
assign addr[21331]= -2025707632;
assign addr[21332]= -2106406677;
assign addr[21333]= -2144419275;
assign addr[21334]= -2138975100;
assign addr[21335]= -2090184478;
assign addr[21336]= -1999036154;
assign addr[21337]= -1867377253;
assign addr[21338]= -1697875851;
assign addr[21339]= -1493966902;
assign addr[21340]= -1259782632;
assign addr[21341]= -1000068799;
assign addr[21342]= -720088517;
assign addr[21343]= -425515602;
assign addr[21344]= -122319591;
assign addr[21345]= 183355234;
assign addr[21346]= 485314355;
assign addr[21347]= 777438554;
assign addr[21348]= 1053807919;
assign addr[21349]= 1308821808;
assign addr[21350]= 1537312353;
assign addr[21351]= 1734649179;
assign addr[21352]= 1896833245;
assign addr[21353]= 2020577882;
assign addr[21354]= 2103375398;
assign addr[21355]= 2143547897;
assign addr[21356]= 2140281282;
assign addr[21357]= 2093641749;
assign addr[21358]= 2004574453;
assign addr[21359]= 1874884346;
assign addr[21360]= 1707199606;
assign addr[21361]= 1504918373;
assign addr[21362]= 1272139887;
assign addr[21363]= 1013581418;
assign addr[21364]= 734482665;
assign addr[21365]= 440499581;
assign addr[21366]= 137589750;
assign addr[21367]= -168108346;
assign addr[21368]= -470399716;
assign addr[21369]= -763158411;
assign addr[21370]= -1040451659;
assign addr[21371]= -1296660098;
assign addr[21372]= -1526591649;
assign addr[21373]= -1725586737;
assign addr[21374]= -1889612716;
assign addr[21375]= -2015345591;
assign addr[21376]= -2100237377;
assign addr[21377]= -2142567738;
assign addr[21378]= -2141478848;
assign addr[21379]= -2096992772;
assign addr[21380]= -2010011024;
assign addr[21381]= -1882296293;
assign addr[21382]= -1716436725;
assign addr[21383]= -1515793473;
assign addr[21384]= -1284432584;
assign addr[21385]= -1027042599;
assign addr[21386]= -748839539;
assign addr[21387]= -455461206;
assign addr[21388]= -152852926;
assign addr[21389]= 152852926;
assign addr[21390]= 455461206;
assign addr[21391]= 748839539;
assign addr[21392]= 1027042599;
assign addr[21393]= 1284432584;
assign addr[21394]= 1515793473;
assign addr[21395]= 1716436725;
assign addr[21396]= 1882296293;
assign addr[21397]= 2010011024;
assign addr[21398]= 2096992772;
assign addr[21399]= 2141478848;
assign addr[21400]= 2142567738;
assign addr[21401]= 2100237377;
assign addr[21402]= 2015345591;
assign addr[21403]= 1889612716;
assign addr[21404]= 1725586737;
assign addr[21405]= 1526591649;
assign addr[21406]= 1296660098;
assign addr[21407]= 1040451659;
assign addr[21408]= 763158411;
assign addr[21409]= 470399716;
assign addr[21410]= 168108346;
assign addr[21411]= -137589750;
assign addr[21412]= -440499581;
assign addr[21413]= -734482665;
assign addr[21414]= -1013581418;
assign addr[21415]= -1272139887;
assign addr[21416]= -1504918373;
assign addr[21417]= -1707199606;
assign addr[21418]= -1874884346;
assign addr[21419]= -2004574453;
assign addr[21420]= -2093641749;
assign addr[21421]= -2140281282;
assign addr[21422]= -2143547897;
assign addr[21423]= -2103375398;
assign addr[21424]= -2020577882;
assign addr[21425]= -1896833245;
assign addr[21426]= -1734649179;
assign addr[21427]= -1537312353;
assign addr[21428]= -1308821808;
assign addr[21429]= -1053807919;
assign addr[21430]= -777438554;
assign addr[21431]= -485314355;
assign addr[21432]= -183355234;
assign addr[21433]= 122319591;
assign addr[21434]= 425515602;
assign addr[21435]= 720088517;
assign addr[21436]= 1000068799;
assign addr[21437]= 1259782632;
assign addr[21438]= 1493966902;
assign addr[21439]= 1697875851;
assign addr[21440]= 1867377253;
assign addr[21441]= 1999036154;
assign addr[21442]= 2090184478;
assign addr[21443]= 2138975100;
assign addr[21444]= 2144419275;
assign addr[21445]= 2106406677;
assign addr[21446]= 2025707632;
assign addr[21447]= 1903957513;
assign addr[21448]= 1743623590;
assign addr[21449]= 1547955041;
assign addr[21450]= 1320917099;
assign addr[21451]= 1067110699;
assign addr[21452]= 791679244;
assign addr[21453]= 500204365;
assign addr[21454]= 198592817;
assign addr[21455]= -107043224;
assign addr[21456]= -410510029;
assign addr[21457]= -705657826;
assign addr[21458]= -986505429;
assign addr[21459]= -1247361445;
assign addr[21460]= -1482939614;
assign addr[21461]= -1688465931;
assign addr[21462]= -1859775393;
assign addr[21463]= -1993396407;
assign addr[21464]= -2086621133;
assign addr[21465]= -2137560369;
assign addr[21466]= -2145181827;
assign addr[21467]= -2109331059;
assign addr[21468]= -2030734582;
assign addr[21469]= -1910985158;
assign addr[21470]= -1752509516;
assign addr[21471]= -1558519173;
assign addr[21472]= -1332945355;
assign addr[21473]= -1080359326;
assign addr[21474]= -805879757;
assign addr[21475]= -515068990;
assign addr[21476]= -213820322;
assign addr[21477]= 91761426;
assign addr[21478]= 395483624;
assign addr[21479]= 691191324;
assign addr[21480]= 972891995;
assign addr[21481]= 1234876957;
assign addr[21482]= 1471837070;
assign addr[21483]= 1678970324;
assign addr[21484]= 1852079154;
assign addr[21485]= 1987655498;
assign addr[21486]= 2082951896;
assign addr[21487]= 2136037160;
assign addr[21488]= 2145835515;
assign addr[21489]= 2112148396;
assign addr[21490]= 2035658475;
assign addr[21491]= 1917915825;
assign addr[21492]= 1761306505;
assign addr[21493]= 1569004214;
assign addr[21494]= 1344905966;
assign addr[21495]= 1093553126;
assign addr[21496]= 820039373;
assign addr[21497]= 529907477;
assign addr[21498]= 229036977;
assign addr[21499]= -76474970;
assign addr[21500]= -380437148;
assign addr[21501]= -676689746;
assign addr[21502]= -959229189;
assign addr[21503]= -1222329801;
assign addr[21504]= -1460659832;
assign addr[21505]= -1669389513;
assign addr[21506]= -1844288924;
assign addr[21507]= -1981813720;
assign addr[21508]= -2079176953;
assign addr[21509]= -2134405552;
assign addr[21510]= -2146380306;
assign addr[21511]= -2114858546;
assign addr[21512]= -2040479063;
assign addr[21513]= -1924749160;
assign addr[21514]= -1770014111;
assign addr[21515]= -1579409630;
assign addr[21516]= -1356798326;
assign addr[21517]= -1106691431;
assign addr[21518]= -834157373;
assign addr[21519]= -544719071;
assign addr[21520]= -244242007;
assign addr[21521]= 61184634;
assign addr[21522]= 365371365;
assign addr[21523]= 662153826;
assign addr[21524]= 945517704;
assign addr[21525]= 1209720613;
assign addr[21526]= 1449408469;
assign addr[21527]= 1659723983;
assign addr[21528]= 1836405100;
assign addr[21529]= 1975871368;
assign addr[21530]= 2075296495;
assign addr[21531]= 2132665626;
assign addr[21532]= 2146816171;
assign addr[21533]= 2117461370;
assign addr[21534]= 2045196100;
assign addr[21535]= 1931484818;
assign addr[21536]= 1778631892;
assign addr[21537]= 1589734894;
assign addr[21538]= 1368621831;
assign addr[21539]= 1119773573;
assign addr[21540]= 848233042;
assign addr[21541]= 559503022;
assign addr[21542]= 259434643;
assign addr[21543]= -45891193;
assign addr[21544]= -350287041;
assign addr[21545]= -647584304;
assign addr[21546]= -931758235;
assign addr[21547]= -1197050035;
assign addr[21548]= -1438083551;
assign addr[21549]= -1649974225;
assign addr[21550]= -1828428082;
assign addr[21551]= -1969828744;
assign addr[21552]= -2071310720;
assign addr[21553]= -2130817471;
assign addr[21554]= -2147143090;
assign addr[21555]= -2119956737;
assign addr[21556]= -2049809346;
assign addr[21557]= -1938122457;
assign addr[21558]= -1787159411;
assign addr[21559]= -1599979481;
assign addr[21560]= -1380375881;
assign addr[21561]= -1132798888;
assign addr[21562]= -862265664;
assign addr[21563]= -574258580;
assign addr[21564]= -274614114;
assign addr[21565]= 30595422;
assign addr[21566]= 335184940;
assign addr[21567]= 632981917;
assign addr[21568]= 917951481;
assign addr[21569]= 1184318708;
assign addr[21570]= 1426685652;
assign addr[21571]= 1640140734;
assign addr[21572]= 1820358275;
assign addr[21573]= 1963686155;
assign addr[21574]= 2067219829;
assign addr[21575]= 2128861181;
assign addr[21576]= 2147361045;
assign addr[21577]= 2122344521;
assign addr[21578]= 2054318569;
assign addr[21579]= 1944661739;
assign addr[21580]= 1795596234;
assign addr[21581]= 1610142873;
assign addr[21582]= 1392059879;
assign addr[21583]= 1145766716;
assign addr[21584]= 876254528;
assign addr[21585]= 588984994;
assign addr[21586]= 289779648;
assign addr[21587]= -15298099;
assign addr[21588]= -320065829;
assign addr[21589]= -618347408;
assign addr[21590]= -904098143;
assign addr[21591]= -1171527280;
assign addr[21592]= -1415215352;
assign addr[21593]= -1630224009;
assign addr[21594]= -1812196087;
assign addr[21595]= -1957443913;
assign addr[21596]= -2063024031;
assign addr[21597]= -2126796855;
assign addr[21598]= -2147470025;
assign addr[21599]= -2124624598;
assign addr[21600]= -2058723538;
assign addr[21601]= -1951102334;
assign addr[21602]= -1803941934;
assign addr[21603]= -1620224553;
assign addr[21604]= -1403673233;
assign addr[21605]= -1158676398;
assign addr[21606]= -890198924;
assign addr[21607]= -603681519;
assign addr[21608]= -304930476;
assign addr[21609]= 0;
assign addr[21610]= 304930476;
assign addr[21611]= 603681519;
assign addr[21612]= 890198924;
assign addr[21613]= 1158676398;
assign addr[21614]= 1403673233;
assign addr[21615]= 1620224553;
assign addr[21616]= 1803941934;
assign addr[21617]= 1951102334;
assign addr[21618]= 2058723538;
assign addr[21619]= 2124624598;
assign addr[21620]= 2147470025;
assign addr[21621]= 2126796855;
assign addr[21622]= 2063024031;
assign addr[21623]= 1957443913;
assign addr[21624]= 1812196087;
assign addr[21625]= 1630224009;
assign addr[21626]= 1415215352;
assign addr[21627]= 1171527280;
assign addr[21628]= 904098143;
assign addr[21629]= 618347408;
assign addr[21630]= 320065829;
assign addr[21631]= 15298099;
assign addr[21632]= -289779648;
assign addr[21633]= -588984994;
assign addr[21634]= -876254528;
assign addr[21635]= -1145766716;
assign addr[21636]= -1392059879;
assign addr[21637]= -1610142873;
assign addr[21638]= -1795596234;
assign addr[21639]= -1944661739;
assign addr[21640]= -2054318569;
assign addr[21641]= -2122344521;
assign addr[21642]= -2147361045;
assign addr[21643]= -2128861181;
assign addr[21644]= -2067219829;
assign addr[21645]= -1963686155;
assign addr[21646]= -1820358275;
assign addr[21647]= -1640140734;
assign addr[21648]= -1426685652;
assign addr[21649]= -1184318708;
assign addr[21650]= -917951481;
assign addr[21651]= -632981917;
assign addr[21652]= -335184940;
assign addr[21653]= -30595422;
assign addr[21654]= 274614114;
assign addr[21655]= 574258580;
assign addr[21656]= 862265664;
assign addr[21657]= 1132798888;
assign addr[21658]= 1380375881;
assign addr[21659]= 1599979481;
assign addr[21660]= 1787159411;
assign addr[21661]= 1938122457;
assign addr[21662]= 2049809346;
assign addr[21663]= 2119956737;
assign addr[21664]= 2147143090;
assign addr[21665]= 2130817471;
assign addr[21666]= 2071310720;
assign addr[21667]= 1969828744;
assign addr[21668]= 1828428082;
assign addr[21669]= 1649974225;
assign addr[21670]= 1438083551;
assign addr[21671]= 1197050035;
assign addr[21672]= 931758235;
assign addr[21673]= 647584304;
assign addr[21674]= 350287041;
assign addr[21675]= 45891193;
assign addr[21676]= -259434643;
assign addr[21677]= -559503022;
assign addr[21678]= -848233042;
assign addr[21679]= -1119773573;
assign addr[21680]= -1368621831;
assign addr[21681]= -1589734894;
assign addr[21682]= -1778631892;
assign addr[21683]= -1931484818;
assign addr[21684]= -2045196100;
assign addr[21685]= -2117461370;
assign addr[21686]= -2146816171;
assign addr[21687]= -2132665626;
assign addr[21688]= -2075296495;
assign addr[21689]= -1975871368;
assign addr[21690]= -1836405100;
assign addr[21691]= -1659723983;
assign addr[21692]= -1449408469;
assign addr[21693]= -1209720613;
assign addr[21694]= -945517704;
assign addr[21695]= -662153826;
assign addr[21696]= -365371365;
assign addr[21697]= -61184634;
assign addr[21698]= 244242007;
assign addr[21699]= 544719071;
assign addr[21700]= 834157373;
assign addr[21701]= 1106691431;
assign addr[21702]= 1356798326;
assign addr[21703]= 1579409630;
assign addr[21704]= 1770014111;
assign addr[21705]= 1924749160;
assign addr[21706]= 2040479063;
assign addr[21707]= 2114858546;
assign addr[21708]= 2146380306;
assign addr[21709]= 2134405552;
assign addr[21710]= 2079176953;
assign addr[21711]= 1981813720;
assign addr[21712]= 1844288924;
assign addr[21713]= 1669389513;
assign addr[21714]= 1460659832;
assign addr[21715]= 1222329801;
assign addr[21716]= 959229189;
assign addr[21717]= 676689746;
assign addr[21718]= 380437148;
assign addr[21719]= 76474970;
assign addr[21720]= -229036977;
assign addr[21721]= -529907477;
assign addr[21722]= -820039373;
assign addr[21723]= -1093553126;
assign addr[21724]= -1344905966;
assign addr[21725]= -1569004214;
assign addr[21726]= -1761306505;
assign addr[21727]= -1917915825;
assign addr[21728]= -2035658475;
assign addr[21729]= -2112148396;
assign addr[21730]= -2145835515;
assign addr[21731]= -2136037160;
assign addr[21732]= -2082951896;
assign addr[21733]= -1987655498;
assign addr[21734]= -1852079154;
assign addr[21735]= -1678970324;
assign addr[21736]= -1471837070;
assign addr[21737]= -1234876957;
assign addr[21738]= -972891995;
assign addr[21739]= -691191324;
assign addr[21740]= -395483624;
assign addr[21741]= -91761426;
assign addr[21742]= 213820322;
assign addr[21743]= 515068990;
assign addr[21744]= 805879757;
assign addr[21745]= 1080359326;
assign addr[21746]= 1332945355;
assign addr[21747]= 1558519173;
assign addr[21748]= 1752509516;
assign addr[21749]= 1910985158;
assign addr[21750]= 2030734582;
assign addr[21751]= 2109331059;
assign addr[21752]= 2145181827;
assign addr[21753]= 2137560369;
assign addr[21754]= 2086621133;
assign addr[21755]= 1993396407;
assign addr[21756]= 1859775393;
assign addr[21757]= 1688465931;
assign addr[21758]= 1482939614;
assign addr[21759]= 1247361445;
assign addr[21760]= 986505429;
assign addr[21761]= 705657826;
assign addr[21762]= 410510029;
assign addr[21763]= 107043224;
assign addr[21764]= -198592817;
assign addr[21765]= -500204365;
assign addr[21766]= -791679244;
assign addr[21767]= -1067110699;
assign addr[21768]= -1320917099;
assign addr[21769]= -1547955041;
assign addr[21770]= -1743623590;
assign addr[21771]= -1903957513;
assign addr[21772]= -2025707632;
assign addr[21773]= -2106406677;
assign addr[21774]= -2144419275;
assign addr[21775]= -2138975100;
assign addr[21776]= -2090184478;
assign addr[21777]= -1999036154;
assign addr[21778]= -1867377253;
assign addr[21779]= -1697875851;
assign addr[21780]= -1493966902;
assign addr[21781]= -1259782632;
assign addr[21782]= -1000068799;
assign addr[21783]= -720088517;
assign addr[21784]= -425515602;
assign addr[21785]= -122319591;
assign addr[21786]= 183355234;
assign addr[21787]= 485314355;
assign addr[21788]= 777438554;
assign addr[21789]= 1053807919;
assign addr[21790]= 1308821808;
assign addr[21791]= 1537312353;
assign addr[21792]= 1734649179;
assign addr[21793]= 1896833245;
assign addr[21794]= 2020577882;
assign addr[21795]= 2103375398;
assign addr[21796]= 2143547897;
assign addr[21797]= 2140281282;
assign addr[21798]= 2093641749;
assign addr[21799]= 2004574453;
assign addr[21800]= 1874884346;
assign addr[21801]= 1707199606;
assign addr[21802]= 1504918373;
assign addr[21803]= 1272139887;
assign addr[21804]= 1013581418;
assign addr[21805]= 734482665;
assign addr[21806]= 440499581;
assign addr[21807]= 137589750;
assign addr[21808]= -168108346;
assign addr[21809]= -470399716;
assign addr[21810]= -763158411;
assign addr[21811]= -1040451659;
assign addr[21812]= -1296660098;
assign addr[21813]= -1526591649;
assign addr[21814]= -1725586737;
assign addr[21815]= -1889612716;
assign addr[21816]= -2015345591;
assign addr[21817]= -2100237377;
assign addr[21818]= -2142567738;
assign addr[21819]= -2141478848;
assign addr[21820]= -2096992772;
assign addr[21821]= -2010011024;
assign addr[21822]= -1882296293;
assign addr[21823]= -1716436725;
assign addr[21824]= -1515793473;
assign addr[21825]= -1284432584;
assign addr[21826]= -1027042599;
assign addr[21827]= -748839539;
assign addr[21828]= -455461206;
assign addr[21829]= -152852926;
assign addr[21830]= 152852926;
assign addr[21831]= 455461206;
assign addr[21832]= 748839539;
assign addr[21833]= 1027042599;
assign addr[21834]= 1284432584;
assign addr[21835]= 1515793473;
assign addr[21836]= 1716436725;
assign addr[21837]= 1882296293;
assign addr[21838]= 2010011024;
assign addr[21839]= 2096992772;
assign addr[21840]= 2141478848;
assign addr[21841]= 2142567738;
assign addr[21842]= 2100237377;
assign addr[21843]= 2015345591;
assign addr[21844]= 1889612716;
assign addr[21845]= 1725586737;
assign addr[21846]= 1526591649;
assign addr[21847]= 1296660098;
assign addr[21848]= 1040451659;
assign addr[21849]= 763158411;
assign addr[21850]= 470399716;
assign addr[21851]= 168108346;
assign addr[21852]= -137589750;
assign addr[21853]= -440499581;
assign addr[21854]= -734482665;
assign addr[21855]= -1013581418;
assign addr[21856]= -1272139887;
assign addr[21857]= -1504918373;
assign addr[21858]= -1707199606;
assign addr[21859]= -1874884346;
assign addr[21860]= -2004574453;
assign addr[21861]= -2093641749;
assign addr[21862]= -2140281282;
assign addr[21863]= -2143547897;
assign addr[21864]= -2103375398;
assign addr[21865]= -2020577882;
assign addr[21866]= -1896833245;
assign addr[21867]= -1734649179;
assign addr[21868]= -1537312353;
assign addr[21869]= -1308821808;
assign addr[21870]= -1053807919;
assign addr[21871]= -777438554;
assign addr[21872]= -485314355;
assign addr[21873]= -183355234;
assign addr[21874]= 122319591;
assign addr[21875]= 425515602;
assign addr[21876]= 720088517;
assign addr[21877]= 1000068799;
assign addr[21878]= 1259782632;
assign addr[21879]= 1493966902;
assign addr[21880]= 1697875851;
assign addr[21881]= 1867377253;
assign addr[21882]= 1999036154;
assign addr[21883]= 2090184478;
assign addr[21884]= 2138975100;
assign addr[21885]= 2144419275;
assign addr[21886]= 2106406677;
assign addr[21887]= 2025707632;
assign addr[21888]= 1903957513;
assign addr[21889]= 1743623590;
assign addr[21890]= 1547955041;
assign addr[21891]= 1320917099;
assign addr[21892]= 1067110699;
assign addr[21893]= 791679244;
assign addr[21894]= 500204365;
assign addr[21895]= 198592817;
assign addr[21896]= -107043224;
assign addr[21897]= -410510029;
assign addr[21898]= -705657826;
assign addr[21899]= -986505429;
assign addr[21900]= -1247361445;
assign addr[21901]= -1482939614;
assign addr[21902]= -1688465931;
assign addr[21903]= -1859775393;
assign addr[21904]= -1993396407;
assign addr[21905]= -2086621133;
assign addr[21906]= -2137560369;
assign addr[21907]= -2145181827;
assign addr[21908]= -2109331059;
assign addr[21909]= -2030734582;
assign addr[21910]= -1910985158;
assign addr[21911]= -1752509516;
assign addr[21912]= -1558519173;
assign addr[21913]= -1332945355;
assign addr[21914]= -1080359326;
assign addr[21915]= -805879757;
assign addr[21916]= -515068990;
assign addr[21917]= -213820322;
assign addr[21918]= 91761426;
assign addr[21919]= 395483624;
assign addr[21920]= 691191324;
assign addr[21921]= 972891995;
assign addr[21922]= 1234876957;
assign addr[21923]= 1471837070;
assign addr[21924]= 1678970324;
assign addr[21925]= 1852079154;
assign addr[21926]= 1987655498;
assign addr[21927]= 2082951896;
assign addr[21928]= 2136037160;
assign addr[21929]= 2145835515;
assign addr[21930]= 2112148396;
assign addr[21931]= 2035658475;
assign addr[21932]= 1917915825;
assign addr[21933]= 1761306505;
assign addr[21934]= 1569004214;
assign addr[21935]= 1344905966;
assign addr[21936]= 1093553126;
assign addr[21937]= 820039373;
assign addr[21938]= 529907477;
assign addr[21939]= 229036977;
assign addr[21940]= -76474970;
assign addr[21941]= -380437148;
assign addr[21942]= -676689746;
assign addr[21943]= -959229189;
assign addr[21944]= -1222329801;
assign addr[21945]= -1460659832;
assign addr[21946]= -1669389513;
assign addr[21947]= -1844288924;
assign addr[21948]= -1981813720;
assign addr[21949]= -2079176953;
assign addr[21950]= -2134405552;
assign addr[21951]= -2146380306;
assign addr[21952]= -2114858546;
assign addr[21953]= -2040479063;
assign addr[21954]= -1924749160;
assign addr[21955]= -1770014111;
assign addr[21956]= -1579409630;
assign addr[21957]= -1356798326;
assign addr[21958]= -1106691431;
assign addr[21959]= -834157373;
assign addr[21960]= -544719071;
assign addr[21961]= -244242007;
assign addr[21962]= 61184634;
assign addr[21963]= 365371365;
assign addr[21964]= 662153826;
assign addr[21965]= 945517704;
assign addr[21966]= 1209720613;
assign addr[21967]= 1449408469;
assign addr[21968]= 1659723983;
assign addr[21969]= 1836405100;
assign addr[21970]= 1975871368;
assign addr[21971]= 2075296495;
assign addr[21972]= 2132665626;
assign addr[21973]= 2146816171;
assign addr[21974]= 2117461370;
assign addr[21975]= 2045196100;
assign addr[21976]= 1931484818;
assign addr[21977]= 1778631892;
assign addr[21978]= 1589734894;
assign addr[21979]= 1368621831;
assign addr[21980]= 1119773573;
assign addr[21981]= 848233042;
assign addr[21982]= 559503022;
assign addr[21983]= 259434643;
assign addr[21984]= -45891193;
assign addr[21985]= -350287041;
assign addr[21986]= -647584304;
assign addr[21987]= -931758235;
assign addr[21988]= -1197050035;
assign addr[21989]= -1438083551;
assign addr[21990]= -1649974225;
assign addr[21991]= -1828428082;
assign addr[21992]= -1969828744;
assign addr[21993]= -2071310720;
assign addr[21994]= -2130817471;
assign addr[21995]= -2147143090;
assign addr[21996]= -2119956737;
assign addr[21997]= -2049809346;
assign addr[21998]= -1938122457;
assign addr[21999]= -1787159411;
assign addr[22000]= -1599979481;
assign addr[22001]= -1380375881;
assign addr[22002]= -1132798888;
assign addr[22003]= -862265664;
assign addr[22004]= -574258580;
assign addr[22005]= -274614114;
assign addr[22006]= 30595422;
assign addr[22007]= 335184940;
assign addr[22008]= 632981917;
assign addr[22009]= 917951481;
assign addr[22010]= 1184318708;
assign addr[22011]= 1426685652;
assign addr[22012]= 1640140734;
assign addr[22013]= 1820358275;
assign addr[22014]= 1963686155;
assign addr[22015]= 2067219829;
assign addr[22016]= 2128861181;
assign addr[22017]= 2147361045;
assign addr[22018]= 2122344521;
assign addr[22019]= 2054318569;
assign addr[22020]= 1944661739;
assign addr[22021]= 1795596234;
assign addr[22022]= 1610142873;
assign addr[22023]= 1392059879;
assign addr[22024]= 1145766716;
assign addr[22025]= 876254528;
assign addr[22026]= 588984994;
assign addr[22027]= 289779648;
assign addr[22028]= -15298099;
assign addr[22029]= -320065829;
assign addr[22030]= -618347408;
assign addr[22031]= -904098143;
assign addr[22032]= -1171527280;
assign addr[22033]= -1415215352;
assign addr[22034]= -1630224009;
assign addr[22035]= -1812196087;
assign addr[22036]= -1957443913;
assign addr[22037]= -2063024031;
assign addr[22038]= -2126796855;
assign addr[22039]= -2147470025;
assign addr[22040]= -2124624598;
assign addr[22041]= -2058723538;
assign addr[22042]= -1951102334;
assign addr[22043]= -1803941934;
assign addr[22044]= -1620224553;
assign addr[22045]= -1403673233;
assign addr[22046]= -1158676398;
assign addr[22047]= -890198924;
assign addr[22048]= -603681519;
assign addr[22049]= -304930476;
assign addr[22050]= 0;
assign addr[22051]= 304930476;
assign addr[22052]= 603681519;
assign addr[22053]= 890198924;
assign addr[22054]= 1158676398;
assign addr[22055]= 1403673233;
assign addr[22056]= 1620224553;
assign addr[22057]= 1803941934;
assign addr[22058]= 1951102334;
assign addr[22059]= 2058723538;
assign addr[22060]= 2124624598;
assign addr[22061]= 2147470025;
assign addr[22062]= 2126796855;
assign addr[22063]= 2063024031;
assign addr[22064]= 1957443913;
assign addr[22065]= 1812196087;
assign addr[22066]= 1630224009;
assign addr[22067]= 1415215352;
assign addr[22068]= 1171527280;
assign addr[22069]= 904098143;
assign addr[22070]= 618347408;
assign addr[22071]= 320065829;
assign addr[22072]= 15298099;
assign addr[22073]= -289779648;
assign addr[22074]= -588984994;
assign addr[22075]= -876254528;
assign addr[22076]= -1145766716;
assign addr[22077]= -1392059879;
assign addr[22078]= -1610142873;
assign addr[22079]= -1795596234;
assign addr[22080]= -1944661739;
assign addr[22081]= -2054318569;
assign addr[22082]= -2122344521;
assign addr[22083]= -2147361045;
assign addr[22084]= -2128861181;
assign addr[22085]= -2067219829;
assign addr[22086]= -1963686155;
assign addr[22087]= -1820358275;
assign addr[22088]= -1640140734;
assign addr[22089]= -1426685652;
assign addr[22090]= -1184318708;
assign addr[22091]= -917951481;
assign addr[22092]= -632981917;
assign addr[22093]= -335184940;
assign addr[22094]= -30595422;
assign addr[22095]= 274614114;
assign addr[22096]= 574258580;
assign addr[22097]= 862265664;
assign addr[22098]= 1132798888;
assign addr[22099]= 1380375881;
assign addr[22100]= 1599979481;
assign addr[22101]= 1787159411;
assign addr[22102]= 1938122457;
assign addr[22103]= 2049809346;
assign addr[22104]= 2119956737;
assign addr[22105]= 2147143090;
assign addr[22106]= 2130817471;
assign addr[22107]= 2071310720;
assign addr[22108]= 1969828744;
assign addr[22109]= 1828428082;
assign addr[22110]= 1649974225;
assign addr[22111]= 1438083551;
assign addr[22112]= 1197050035;
assign addr[22113]= 931758235;
assign addr[22114]= 647584304;
assign addr[22115]= 350287041;
assign addr[22116]= 45891193;
assign addr[22117]= -259434643;
assign addr[22118]= -559503022;
assign addr[22119]= -848233042;
assign addr[22120]= -1119773573;
assign addr[22121]= -1368621831;
assign addr[22122]= -1589734894;
assign addr[22123]= -1778631892;
assign addr[22124]= -1931484818;
assign addr[22125]= -2045196100;
assign addr[22126]= -2117461370;
assign addr[22127]= -2146816171;
assign addr[22128]= -2132665626;
assign addr[22129]= -2075296495;
assign addr[22130]= -1975871368;
assign addr[22131]= -1836405100;
assign addr[22132]= -1659723983;
assign addr[22133]= -1449408469;
assign addr[22134]= -1209720613;
assign addr[22135]= -945517704;
assign addr[22136]= -662153826;
assign addr[22137]= -365371365;
assign addr[22138]= -61184634;
assign addr[22139]= 244242007;
assign addr[22140]= 544719071;
assign addr[22141]= 834157373;
assign addr[22142]= 1106691431;
assign addr[22143]= 1356798326;
assign addr[22144]= 1579409630;
assign addr[22145]= 1770014111;
assign addr[22146]= 1924749160;
assign addr[22147]= 2040479063;
assign addr[22148]= 2114858546;
assign addr[22149]= 2146380306;
assign addr[22150]= 2134405552;
assign addr[22151]= 2079176953;
assign addr[22152]= 1981813720;
assign addr[22153]= 1844288924;
assign addr[22154]= 1669389513;
assign addr[22155]= 1460659832;
assign addr[22156]= 1222329801;
assign addr[22157]= 959229189;
assign addr[22158]= 676689746;
assign addr[22159]= 380437148;
assign addr[22160]= 76474970;
assign addr[22161]= -229036977;
assign addr[22162]= -529907477;
assign addr[22163]= -820039373;
assign addr[22164]= -1093553126;
assign addr[22165]= -1344905966;
assign addr[22166]= -1569004214;
assign addr[22167]= -1761306505;
assign addr[22168]= -1917915825;
assign addr[22169]= -2035658475;
assign addr[22170]= -2112148396;
assign addr[22171]= -2145835515;
assign addr[22172]= -2136037160;
assign addr[22173]= -2082951896;
assign addr[22174]= -1987655498;
assign addr[22175]= -1852079154;
assign addr[22176]= -1678970324;
assign addr[22177]= -1471837070;
assign addr[22178]= -1234876957;
assign addr[22179]= -972891995;
assign addr[22180]= -691191324;
assign addr[22181]= -395483624;
assign addr[22182]= -91761426;
assign addr[22183]= 213820322;
assign addr[22184]= 515068990;
assign addr[22185]= 805879757;
assign addr[22186]= 1080359326;
assign addr[22187]= 1332945355;
assign addr[22188]= 1558519173;
assign addr[22189]= 1752509516;
assign addr[22190]= 1910985158;
assign addr[22191]= 2030734582;
assign addr[22192]= 2109331059;
assign addr[22193]= 2145181827;
assign addr[22194]= 2137560369;
assign addr[22195]= 2086621133;
assign addr[22196]= 1993396407;
assign addr[22197]= 1859775393;
assign addr[22198]= 1688465931;
assign addr[22199]= 1482939614;
assign addr[22200]= 1247361445;
assign addr[22201]= 986505429;
assign addr[22202]= 705657826;
assign addr[22203]= 410510029;
assign addr[22204]= 107043224;
assign addr[22205]= -198592817;
assign addr[22206]= -500204365;
assign addr[22207]= -791679244;
assign addr[22208]= -1067110699;
assign addr[22209]= -1320917099;
assign addr[22210]= -1547955041;
assign addr[22211]= -1743623590;
assign addr[22212]= -1903957513;
assign addr[22213]= -2025707632;
assign addr[22214]= -2106406677;
assign addr[22215]= -2144419275;
assign addr[22216]= -2138975100;
assign addr[22217]= -2090184478;
assign addr[22218]= -1999036154;
assign addr[22219]= -1867377253;
assign addr[22220]= -1697875851;
assign addr[22221]= -1493966902;
assign addr[22222]= -1259782632;
assign addr[22223]= -1000068799;
assign addr[22224]= -720088517;
assign addr[22225]= -425515602;
assign addr[22226]= -122319591;
assign addr[22227]= 183355234;
assign addr[22228]= 485314355;
assign addr[22229]= 777438554;
assign addr[22230]= 1053807919;
assign addr[22231]= 1308821808;
assign addr[22232]= 1537312353;
assign addr[22233]= 1734649179;
assign addr[22234]= 1896833245;
assign addr[22235]= 2020577882;
assign addr[22236]= 2103375398;
assign addr[22237]= 2143547897;
assign addr[22238]= 2140281282;
assign addr[22239]= 2093641749;
assign addr[22240]= 2004574453;
assign addr[22241]= 1874884346;
assign addr[22242]= 1707199606;
assign addr[22243]= 1504918373;
assign addr[22244]= 1272139887;
assign addr[22245]= 1013581418;
assign addr[22246]= 734482665;
assign addr[22247]= 440499581;
assign addr[22248]= 137589750;
assign addr[22249]= -168108346;
assign addr[22250]= -470399716;
assign addr[22251]= -763158411;
assign addr[22252]= -1040451659;
assign addr[22253]= -1296660098;
assign addr[22254]= -1526591649;
assign addr[22255]= -1725586737;
assign addr[22256]= -1889612716;
assign addr[22257]= -2015345591;
assign addr[22258]= -2100237377;
assign addr[22259]= -2142567738;
assign addr[22260]= -2141478848;
assign addr[22261]= -2096992772;
assign addr[22262]= -2010011024;
assign addr[22263]= -1882296293;
assign addr[22264]= -1716436725;
assign addr[22265]= -1515793473;
assign addr[22266]= -1284432584;
assign addr[22267]= -1027042599;
assign addr[22268]= -748839539;
assign addr[22269]= -455461206;
assign addr[22270]= -152852926;
assign addr[22271]= 152852926;
assign addr[22272]= 455461206;
assign addr[22273]= 748839539;
assign addr[22274]= 1027042599;
assign addr[22275]= 1284432584;
assign addr[22276]= 1515793473;
assign addr[22277]= 1716436725;
assign addr[22278]= 1882296293;
assign addr[22279]= 2010011024;
assign addr[22280]= 2096992772;
assign addr[22281]= 2141478848;
assign addr[22282]= 2142567738;
assign addr[22283]= 2100237377;
assign addr[22284]= 2015345591;
assign addr[22285]= 1889612716;
assign addr[22286]= 1725586737;
assign addr[22287]= 1526591649;
assign addr[22288]= 1296660098;
assign addr[22289]= 1040451659;
assign addr[22290]= 763158411;
assign addr[22291]= 470399716;
assign addr[22292]= 168108346;
assign addr[22293]= -137589750;
assign addr[22294]= -440499581;
assign addr[22295]= -734482665;
assign addr[22296]= -1013581418;
assign addr[22297]= -1272139887;
assign addr[22298]= -1504918373;
assign addr[22299]= -1707199606;
assign addr[22300]= -1874884346;
assign addr[22301]= -2004574453;
assign addr[22302]= -2093641749;
assign addr[22303]= -2140281282;
assign addr[22304]= -2143547897;
assign addr[22305]= -2103375398;
assign addr[22306]= -2020577882;
assign addr[22307]= -1896833245;
assign addr[22308]= -1734649179;
assign addr[22309]= -1537312353;
assign addr[22310]= -1308821808;
assign addr[22311]= -1053807919;
assign addr[22312]= -777438554;
assign addr[22313]= -485314355;
assign addr[22314]= -183355234;
assign addr[22315]= 122319591;
assign addr[22316]= 425515602;
assign addr[22317]= 720088517;
assign addr[22318]= 1000068799;
assign addr[22319]= 1259782632;
assign addr[22320]= 1493966902;
assign addr[22321]= 1697875851;
assign addr[22322]= 1867377253;
assign addr[22323]= 1999036154;
assign addr[22324]= 2090184478;
assign addr[22325]= 2138975100;
assign addr[22326]= 2144419275;
assign addr[22327]= 2106406677;
assign addr[22328]= 2025707632;
assign addr[22329]= 1903957513;
assign addr[22330]= 1743623590;
assign addr[22331]= 1547955041;
assign addr[22332]= 1320917099;
assign addr[22333]= 1067110699;
assign addr[22334]= 791679244;
assign addr[22335]= 500204365;
assign addr[22336]= 198592817;
assign addr[22337]= -107043224;
assign addr[22338]= -410510029;
assign addr[22339]= -705657826;
assign addr[22340]= -986505429;
assign addr[22341]= -1247361445;
assign addr[22342]= -1482939614;
assign addr[22343]= -1688465931;
assign addr[22344]= -1859775393;
assign addr[22345]= -1993396407;
assign addr[22346]= -2086621133;
assign addr[22347]= -2137560369;
assign addr[22348]= -2145181827;
assign addr[22349]= -2109331059;
assign addr[22350]= -2030734582;
assign addr[22351]= -1910985158;
assign addr[22352]= -1752509516;
assign addr[22353]= -1558519173;
assign addr[22354]= -1332945355;
assign addr[22355]= -1080359326;
assign addr[22356]= -805879757;
assign addr[22357]= -515068990;
assign addr[22358]= -213820322;
assign addr[22359]= 91761426;
assign addr[22360]= 395483624;
assign addr[22361]= 691191324;
assign addr[22362]= 972891995;
assign addr[22363]= 1234876957;
assign addr[22364]= 1471837070;
assign addr[22365]= 1678970324;
assign addr[22366]= 1852079154;
assign addr[22367]= 1987655498;
assign addr[22368]= 2082951896;
assign addr[22369]= 2136037160;
assign addr[22370]= 2145835515;
assign addr[22371]= 2112148396;
assign addr[22372]= 2035658475;
assign addr[22373]= 1917915825;
assign addr[22374]= 1761306505;
assign addr[22375]= 1569004214;
assign addr[22376]= 1344905966;
assign addr[22377]= 1093553126;
assign addr[22378]= 820039373;
assign addr[22379]= 529907477;
assign addr[22380]= 229036977;
assign addr[22381]= -76474970;
assign addr[22382]= -380437148;
assign addr[22383]= -676689746;
assign addr[22384]= -959229189;
assign addr[22385]= -1222329801;
assign addr[22386]= -1460659832;
assign addr[22387]= -1669389513;
assign addr[22388]= -1844288924;
assign addr[22389]= -1981813720;
assign addr[22390]= -2079176953;
assign addr[22391]= -2134405552;
assign addr[22392]= -2146380306;
assign addr[22393]= -2114858546;
assign addr[22394]= -2040479063;
assign addr[22395]= -1924749160;
assign addr[22396]= -1770014111;
assign addr[22397]= -1579409630;
assign addr[22398]= -1356798326;
assign addr[22399]= -1106691431;
assign addr[22400]= -834157373;
assign addr[22401]= -544719071;
assign addr[22402]= -244242007;
assign addr[22403]= 61184634;
assign addr[22404]= 365371365;
assign addr[22405]= 662153826;
assign addr[22406]= 945517704;
assign addr[22407]= 1209720613;
assign addr[22408]= 1449408469;
assign addr[22409]= 1659723983;
assign addr[22410]= 1836405100;
assign addr[22411]= 1975871368;
assign addr[22412]= 2075296495;
assign addr[22413]= 2132665626;
assign addr[22414]= 2146816171;
assign addr[22415]= 2117461370;
assign addr[22416]= 2045196100;
assign addr[22417]= 1931484818;
assign addr[22418]= 1778631892;
assign addr[22419]= 1589734894;
assign addr[22420]= 1368621831;
assign addr[22421]= 1119773573;
assign addr[22422]= 848233042;
assign addr[22423]= 559503022;
assign addr[22424]= 259434643;
assign addr[22425]= -45891193;
assign addr[22426]= -350287041;
assign addr[22427]= -647584304;
assign addr[22428]= -931758235;
assign addr[22429]= -1197050035;
assign addr[22430]= -1438083551;
assign addr[22431]= -1649974225;
assign addr[22432]= -1828428082;
assign addr[22433]= -1969828744;
assign addr[22434]= -2071310720;
assign addr[22435]= -2130817471;
assign addr[22436]= -2147143090;
assign addr[22437]= -2119956737;
assign addr[22438]= -2049809346;
assign addr[22439]= -1938122457;
assign addr[22440]= -1787159411;
assign addr[22441]= -1599979481;
assign addr[22442]= -1380375881;
assign addr[22443]= -1132798888;
assign addr[22444]= -862265664;
assign addr[22445]= -574258580;
assign addr[22446]= -274614114;
assign addr[22447]= 30595422;
assign addr[22448]= 335184940;
assign addr[22449]= 632981917;
assign addr[22450]= 917951481;
assign addr[22451]= 1184318708;
assign addr[22452]= 1426685652;
assign addr[22453]= 1640140734;
assign addr[22454]= 1820358275;
assign addr[22455]= 1963686155;
assign addr[22456]= 2067219829;
assign addr[22457]= 2128861181;
assign addr[22458]= 2147361045;
assign addr[22459]= 2122344521;
assign addr[22460]= 2054318569;
assign addr[22461]= 1944661739;
assign addr[22462]= 1795596234;
assign addr[22463]= 1610142873;
assign addr[22464]= 1392059879;
assign addr[22465]= 1145766716;
assign addr[22466]= 876254528;
assign addr[22467]= 588984994;
assign addr[22468]= 289779648;
assign addr[22469]= -15298099;
assign addr[22470]= -320065829;
assign addr[22471]= -618347408;
assign addr[22472]= -904098143;
assign addr[22473]= -1171527280;
assign addr[22474]= -1415215352;
assign addr[22475]= -1630224009;
assign addr[22476]= -1812196087;
assign addr[22477]= -1957443913;
assign addr[22478]= -2063024031;
assign addr[22479]= -2126796855;
assign addr[22480]= -2147470025;
assign addr[22481]= -2124624598;
assign addr[22482]= -2058723538;
assign addr[22483]= -1951102334;
assign addr[22484]= -1803941934;
assign addr[22485]= -1620224553;
assign addr[22486]= -1403673233;
assign addr[22487]= -1158676398;
assign addr[22488]= -890198924;
assign addr[22489]= -603681519;
assign addr[22490]= -304930476;
assign addr[22491]= 0;
assign addr[22492]= 304930476;
assign addr[22493]= 603681519;
assign addr[22494]= 890198924;
assign addr[22495]= 1158676398;
assign addr[22496]= 1403673233;
assign addr[22497]= 1620224553;
assign addr[22498]= 1803941934;
assign addr[22499]= 1951102334;
assign addr[22500]= 2058723538;
assign addr[22501]= 2124624598;
assign addr[22502]= 2147470025;
assign addr[22503]= 2126796855;
assign addr[22504]= 2063024031;
assign addr[22505]= 1957443913;
assign addr[22506]= 1812196087;
assign addr[22507]= 1630224009;
assign addr[22508]= 1415215352;
assign addr[22509]= 1171527280;
assign addr[22510]= 904098143;
assign addr[22511]= 618347408;
assign addr[22512]= 320065829;
assign addr[22513]= 15298099;
assign addr[22514]= -289779648;
assign addr[22515]= -588984994;
assign addr[22516]= -876254528;
assign addr[22517]= -1145766716;
assign addr[22518]= -1392059879;
assign addr[22519]= -1610142873;
assign addr[22520]= -1795596234;
assign addr[22521]= -1944661739;
assign addr[22522]= -2054318569;
assign addr[22523]= -2122344521;
assign addr[22524]= -2147361045;
assign addr[22525]= -2128861181;
assign addr[22526]= -2067219829;
assign addr[22527]= -1963686155;
assign addr[22528]= -1820358275;
assign addr[22529]= -1640140734;
assign addr[22530]= -1426685652;
assign addr[22531]= -1184318708;
assign addr[22532]= -917951481;
assign addr[22533]= -632981917;
assign addr[22534]= -335184940;
assign addr[22535]= -30595422;
assign addr[22536]= 274614114;
assign addr[22537]= 574258580;
assign addr[22538]= 862265664;
assign addr[22539]= 1132798888;
assign addr[22540]= 1380375881;
assign addr[22541]= 1599979481;
assign addr[22542]= 1787159411;
assign addr[22543]= 1938122457;
assign addr[22544]= 2049809346;
assign addr[22545]= 2119956737;
assign addr[22546]= 2147143090;
assign addr[22547]= 2130817471;
assign addr[22548]= 2071310720;
assign addr[22549]= 1969828744;
assign addr[22550]= 1828428082;
assign addr[22551]= 1649974225;
assign addr[22552]= 1438083551;
assign addr[22553]= 1197050035;
assign addr[22554]= 931758235;
assign addr[22555]= 647584304;
assign addr[22556]= 350287041;
assign addr[22557]= 45891193;
assign addr[22558]= -259434643;
assign addr[22559]= -559503022;
assign addr[22560]= -848233042;
assign addr[22561]= -1119773573;
assign addr[22562]= -1368621831;
assign addr[22563]= -1589734894;
assign addr[22564]= -1778631892;
assign addr[22565]= -1931484818;
assign addr[22566]= -2045196100;
assign addr[22567]= -2117461370;
assign addr[22568]= -2146816171;
assign addr[22569]= -2132665626;
assign addr[22570]= -2075296495;
assign addr[22571]= -1975871368;
assign addr[22572]= -1836405100;
assign addr[22573]= -1659723983;
assign addr[22574]= -1449408469;
assign addr[22575]= -1209720613;
assign addr[22576]= -945517704;
assign addr[22577]= -662153826;
assign addr[22578]= -365371365;
assign addr[22579]= -61184634;
assign addr[22580]= 244242007;
assign addr[22581]= 544719071;
assign addr[22582]= 834157373;
assign addr[22583]= 1106691431;
assign addr[22584]= 1356798326;
assign addr[22585]= 1579409630;
assign addr[22586]= 1770014111;
assign addr[22587]= 1924749160;
assign addr[22588]= 2040479063;
assign addr[22589]= 2114858546;
assign addr[22590]= 2146380306;
assign addr[22591]= 2134405552;
assign addr[22592]= 2079176953;
assign addr[22593]= 1981813720;
assign addr[22594]= 1844288924;
assign addr[22595]= 1669389513;
assign addr[22596]= 1460659832;
assign addr[22597]= 1222329801;
assign addr[22598]= 959229189;
assign addr[22599]= 676689746;
assign addr[22600]= 380437148;
assign addr[22601]= 76474970;
assign addr[22602]= -229036977;
assign addr[22603]= -529907477;
assign addr[22604]= -820039373;
assign addr[22605]= -1093553126;
assign addr[22606]= -1344905966;
assign addr[22607]= -1569004214;
assign addr[22608]= -1761306505;
assign addr[22609]= -1917915825;
assign addr[22610]= -2035658475;
assign addr[22611]= -2112148396;
assign addr[22612]= -2145835515;
assign addr[22613]= -2136037160;
assign addr[22614]= -2082951896;
assign addr[22615]= -1987655498;
assign addr[22616]= -1852079154;
assign addr[22617]= -1678970324;
assign addr[22618]= -1471837070;
assign addr[22619]= -1234876957;
assign addr[22620]= -972891995;
assign addr[22621]= -691191324;
assign addr[22622]= -395483624;
assign addr[22623]= -91761426;
assign addr[22624]= 213820322;
assign addr[22625]= 515068990;
assign addr[22626]= 805879757;
assign addr[22627]= 1080359326;
assign addr[22628]= 1332945355;
assign addr[22629]= 1558519173;
assign addr[22630]= 1752509516;
assign addr[22631]= 1910985158;
assign addr[22632]= 2030734582;
assign addr[22633]= 2109331059;
assign addr[22634]= 2145181827;
assign addr[22635]= 2137560369;
assign addr[22636]= 2086621133;
assign addr[22637]= 1993396407;
assign addr[22638]= 1859775393;
assign addr[22639]= 1688465931;
assign addr[22640]= 1482939614;
assign addr[22641]= 1247361445;
assign addr[22642]= 986505429;
assign addr[22643]= 705657826;
assign addr[22644]= 410510029;
assign addr[22645]= 107043224;
assign addr[22646]= -198592817;
assign addr[22647]= -500204365;
assign addr[22648]= -791679244;
assign addr[22649]= -1067110699;
assign addr[22650]= -1320917099;
assign addr[22651]= -1547955041;
assign addr[22652]= -1743623590;
assign addr[22653]= -1903957513;
assign addr[22654]= -2025707632;
assign addr[22655]= -2106406677;
assign addr[22656]= -2144419275;
assign addr[22657]= -2138975100;
assign addr[22658]= -2090184478;
assign addr[22659]= -1999036154;
assign addr[22660]= -1867377253;
assign addr[22661]= -1697875851;
assign addr[22662]= -1493966902;
assign addr[22663]= -1259782632;
assign addr[22664]= -1000068799;
assign addr[22665]= -720088517;
assign addr[22666]= -425515602;
assign addr[22667]= -122319591;
assign addr[22668]= 183355234;
assign addr[22669]= 485314355;
assign addr[22670]= 777438554;
assign addr[22671]= 1053807919;
assign addr[22672]= 1308821808;
assign addr[22673]= 1537312353;
assign addr[22674]= 1734649179;
assign addr[22675]= 1896833245;
assign addr[22676]= 2020577882;
assign addr[22677]= 2103375398;
assign addr[22678]= 2143547897;
assign addr[22679]= 2140281282;
assign addr[22680]= 2093641749;
assign addr[22681]= 2004574453;
assign addr[22682]= 1874884346;
assign addr[22683]= 1707199606;
assign addr[22684]= 1504918373;
assign addr[22685]= 1272139887;
assign addr[22686]= 1013581418;
assign addr[22687]= 734482665;
assign addr[22688]= 440499581;
assign addr[22689]= 137589750;
assign addr[22690]= -168108346;
assign addr[22691]= -470399716;
assign addr[22692]= -763158411;
assign addr[22693]= -1040451659;
assign addr[22694]= -1296660098;
assign addr[22695]= -1526591649;
assign addr[22696]= -1725586737;
assign addr[22697]= -1889612716;
assign addr[22698]= -2015345591;
assign addr[22699]= -2100237377;
assign addr[22700]= -2142567738;
assign addr[22701]= -2141478848;
assign addr[22702]= -2096992772;
assign addr[22703]= -2010011024;
assign addr[22704]= -1882296293;
assign addr[22705]= -1716436725;
assign addr[22706]= -1515793473;
assign addr[22707]= -1284432584;
assign addr[22708]= -1027042599;
assign addr[22709]= -748839539;
assign addr[22710]= -455461206;
assign addr[22711]= -152852926;
assign addr[22712]= 152852926;
assign addr[22713]= 455461206;
assign addr[22714]= 748839539;
assign addr[22715]= 1027042599;
assign addr[22716]= 1284432584;
assign addr[22717]= 1515793473;
assign addr[22718]= 1716436725;
assign addr[22719]= 1882296293;
assign addr[22720]= 2010011024;
assign addr[22721]= 2096992772;
assign addr[22722]= 2141478848;
assign addr[22723]= 2142567738;
assign addr[22724]= 2100237377;
assign addr[22725]= 2015345591;
assign addr[22726]= 1889612716;
assign addr[22727]= 1725586737;
assign addr[22728]= 1526591649;
assign addr[22729]= 1296660098;
assign addr[22730]= 1040451659;
assign addr[22731]= 763158411;
assign addr[22732]= 470399716;
assign addr[22733]= 168108346;
assign addr[22734]= -137589750;
assign addr[22735]= -440499581;
assign addr[22736]= -734482665;
assign addr[22737]= -1013581418;
assign addr[22738]= -1272139887;
assign addr[22739]= -1504918373;
assign addr[22740]= -1707199606;
assign addr[22741]= -1874884346;
assign addr[22742]= -2004574453;
assign addr[22743]= -2093641749;
assign addr[22744]= -2140281282;
assign addr[22745]= -2143547897;
assign addr[22746]= -2103375398;
assign addr[22747]= -2020577882;
assign addr[22748]= -1896833245;
assign addr[22749]= -1734649179;
assign addr[22750]= -1537312353;
assign addr[22751]= -1308821808;
assign addr[22752]= -1053807919;
assign addr[22753]= -777438554;
assign addr[22754]= -485314355;
assign addr[22755]= -183355234;
assign addr[22756]= 122319591;
assign addr[22757]= 425515602;
assign addr[22758]= 720088517;
assign addr[22759]= 1000068799;
assign addr[22760]= 1259782632;
assign addr[22761]= 1493966902;
assign addr[22762]= 1697875851;
assign addr[22763]= 1867377253;
assign addr[22764]= 1999036154;
assign addr[22765]= 2090184478;
assign addr[22766]= 2138975100;
assign addr[22767]= 2144419275;
assign addr[22768]= 2106406677;
assign addr[22769]= 2025707632;
assign addr[22770]= 1903957513;
assign addr[22771]= 1743623590;
assign addr[22772]= 1547955041;
assign addr[22773]= 1320917099;
assign addr[22774]= 1067110699;
assign addr[22775]= 791679244;
assign addr[22776]= 500204365;
assign addr[22777]= 198592817;
assign addr[22778]= -107043224;
assign addr[22779]= -410510029;
assign addr[22780]= -705657826;
assign addr[22781]= -986505429;
assign addr[22782]= -1247361445;
assign addr[22783]= -1482939614;
assign addr[22784]= -1688465931;
assign addr[22785]= -1859775393;
assign addr[22786]= -1993396407;
assign addr[22787]= -2086621133;
assign addr[22788]= -2137560369;
assign addr[22789]= -2145181827;
assign addr[22790]= -2109331059;
assign addr[22791]= -2030734582;
assign addr[22792]= -1910985158;
assign addr[22793]= -1752509516;
assign addr[22794]= -1558519173;
assign addr[22795]= -1332945355;
assign addr[22796]= -1080359326;
assign addr[22797]= -805879757;
assign addr[22798]= -515068990;
assign addr[22799]= -213820322;
assign addr[22800]= 91761426;
assign addr[22801]= 395483624;
assign addr[22802]= 691191324;
assign addr[22803]= 972891995;
assign addr[22804]= 1234876957;
assign addr[22805]= 1471837070;
assign addr[22806]= 1678970324;
assign addr[22807]= 1852079154;
assign addr[22808]= 1987655498;
assign addr[22809]= 2082951896;
assign addr[22810]= 2136037160;
assign addr[22811]= 2145835515;
assign addr[22812]= 2112148396;
assign addr[22813]= 2035658475;
assign addr[22814]= 1917915825;
assign addr[22815]= 1761306505;
assign addr[22816]= 1569004214;
assign addr[22817]= 1344905966;
assign addr[22818]= 1093553126;
assign addr[22819]= 820039373;
assign addr[22820]= 529907477;
assign addr[22821]= 229036977;
assign addr[22822]= -76474970;
assign addr[22823]= -380437148;
assign addr[22824]= -676689746;
assign addr[22825]= -959229189;
assign addr[22826]= -1222329801;
assign addr[22827]= -1460659832;
assign addr[22828]= -1669389513;
assign addr[22829]= -1844288924;
assign addr[22830]= -1981813720;
assign addr[22831]= -2079176953;
assign addr[22832]= -2134405552;
assign addr[22833]= -2146380306;
assign addr[22834]= -2114858546;
assign addr[22835]= -2040479063;
assign addr[22836]= -1924749160;
assign addr[22837]= -1770014111;
assign addr[22838]= -1579409630;
assign addr[22839]= -1356798326;
assign addr[22840]= -1106691431;
assign addr[22841]= -834157373;
assign addr[22842]= -544719071;
assign addr[22843]= -244242007;
assign addr[22844]= 61184634;
assign addr[22845]= 365371365;
assign addr[22846]= 662153826;
assign addr[22847]= 945517704;
assign addr[22848]= 1209720613;
assign addr[22849]= 1449408469;
assign addr[22850]= 1659723983;
assign addr[22851]= 1836405100;
assign addr[22852]= 1975871368;
assign addr[22853]= 2075296495;
assign addr[22854]= 2132665626;
assign addr[22855]= 2146816171;
assign addr[22856]= 2117461370;
assign addr[22857]= 2045196100;
assign addr[22858]= 1931484818;
assign addr[22859]= 1778631892;
assign addr[22860]= 1589734894;
assign addr[22861]= 1368621831;
assign addr[22862]= 1119773573;
assign addr[22863]= 848233042;
assign addr[22864]= 559503022;
assign addr[22865]= 259434643;
assign addr[22866]= -45891193;
assign addr[22867]= -350287041;
assign addr[22868]= -647584304;
assign addr[22869]= -931758235;
assign addr[22870]= -1197050035;
assign addr[22871]= -1438083551;
assign addr[22872]= -1649974225;
assign addr[22873]= -1828428082;
assign addr[22874]= -1969828744;
assign addr[22875]= -2071310720;
assign addr[22876]= -2130817471;
assign addr[22877]= -2147143090;
assign addr[22878]= -2119956737;
assign addr[22879]= -2049809346;
assign addr[22880]= -1938122457;
assign addr[22881]= -1787159411;
assign addr[22882]= -1599979481;
assign addr[22883]= -1380375881;
assign addr[22884]= -1132798888;
assign addr[22885]= -862265664;
assign addr[22886]= -574258580;
assign addr[22887]= -274614114;
assign addr[22888]= 30595422;
assign addr[22889]= 335184940;
assign addr[22890]= 632981917;
assign addr[22891]= 917951481;
assign addr[22892]= 1184318708;
assign addr[22893]= 1426685652;
assign addr[22894]= 1640140734;
assign addr[22895]= 1820358275;
assign addr[22896]= 1963686155;
assign addr[22897]= 2067219829;
assign addr[22898]= 2128861181;
assign addr[22899]= 2147361045;
assign addr[22900]= 2122344521;
assign addr[22901]= 2054318569;
assign addr[22902]= 1944661739;
assign addr[22903]= 1795596234;
assign addr[22904]= 1610142873;
assign addr[22905]= 1392059879;
assign addr[22906]= 1145766716;
assign addr[22907]= 876254528;
assign addr[22908]= 588984994;
assign addr[22909]= 289779648;
assign addr[22910]= -15298099;
assign addr[22911]= -320065829;
assign addr[22912]= -618347408;
assign addr[22913]= -904098143;
assign addr[22914]= -1171527280;
assign addr[22915]= -1415215352;
assign addr[22916]= -1630224009;
assign addr[22917]= -1812196087;
assign addr[22918]= -1957443913;
assign addr[22919]= -2063024031;
assign addr[22920]= -2126796855;
assign addr[22921]= -2147470025;
assign addr[22922]= -2124624598;
assign addr[22923]= -2058723538;
assign addr[22924]= -1951102334;
assign addr[22925]= -1803941934;
assign addr[22926]= -1620224553;
assign addr[22927]= -1403673233;
assign addr[22928]= -1158676398;
assign addr[22929]= -890198924;
assign addr[22930]= -603681519;
assign addr[22931]= -304930476;
assign addr[22932]= 0;
assign addr[22933]= 304930476;
assign addr[22934]= 603681519;
assign addr[22935]= 890198924;
assign addr[22936]= 1158676398;
assign addr[22937]= 1403673233;
assign addr[22938]= 1620224553;
assign addr[22939]= 1803941934;
assign addr[22940]= 1951102334;
assign addr[22941]= 2058723538;
assign addr[22942]= 2124624598;
assign addr[22943]= 2147470025;
assign addr[22944]= 2126796855;
assign addr[22945]= 2063024031;
assign addr[22946]= 1957443913;
assign addr[22947]= 1812196087;
assign addr[22948]= 1630224009;
assign addr[22949]= 1415215352;
assign addr[22950]= 1171527280;
assign addr[22951]= 904098143;
assign addr[22952]= 618347408;
assign addr[22953]= 320065829;
assign addr[22954]= 15298099;
assign addr[22955]= -289779648;
assign addr[22956]= -588984994;
assign addr[22957]= -876254528;
assign addr[22958]= -1145766716;
assign addr[22959]= -1392059879;
assign addr[22960]= -1610142873;
assign addr[22961]= -1795596234;
assign addr[22962]= -1944661739;
assign addr[22963]= -2054318569;
assign addr[22964]= -2122344521;
assign addr[22965]= -2147361045;
assign addr[22966]= -2128861181;
assign addr[22967]= -2067219829;
assign addr[22968]= -1963686155;
assign addr[22969]= -1820358275;
assign addr[22970]= -1640140734;
assign addr[22971]= -1426685652;
assign addr[22972]= -1184318708;
assign addr[22973]= -917951481;
assign addr[22974]= -632981917;
assign addr[22975]= -335184940;
assign addr[22976]= -30595422;
assign addr[22977]= 274614114;
assign addr[22978]= 574258580;
assign addr[22979]= 862265664;
assign addr[22980]= 1132798888;
assign addr[22981]= 1380375881;
assign addr[22982]= 1599979481;
assign addr[22983]= 1787159411;
assign addr[22984]= 1938122457;
assign addr[22985]= 2049809346;
assign addr[22986]= 2119956737;
assign addr[22987]= 2147143090;
assign addr[22988]= 2130817471;
assign addr[22989]= 2071310720;
assign addr[22990]= 1969828744;
assign addr[22991]= 1828428082;
assign addr[22992]= 1649974225;
assign addr[22993]= 1438083551;
assign addr[22994]= 1197050035;
assign addr[22995]= 931758235;
assign addr[22996]= 647584304;
assign addr[22997]= 350287041;
assign addr[22998]= 45891193;
assign addr[22999]= -259434643;
assign addr[23000]= -559503022;
assign addr[23001]= -848233042;
assign addr[23002]= -1119773573;
assign addr[23003]= -1368621831;
assign addr[23004]= -1589734894;
assign addr[23005]= -1778631892;
assign addr[23006]= -1931484818;
assign addr[23007]= -2045196100;
assign addr[23008]= -2117461370;
assign addr[23009]= -2146816171;
assign addr[23010]= -2132665626;
assign addr[23011]= -2075296495;
assign addr[23012]= -1975871368;
assign addr[23013]= -1836405100;
assign addr[23014]= -1659723983;
assign addr[23015]= -1449408469;
assign addr[23016]= -1209720613;
assign addr[23017]= -945517704;
assign addr[23018]= -662153826;
assign addr[23019]= -365371365;
assign addr[23020]= -61184634;
assign addr[23021]= 244242007;
assign addr[23022]= 544719071;
assign addr[23023]= 834157373;
assign addr[23024]= 1106691431;
assign addr[23025]= 1356798326;
assign addr[23026]= 1579409630;
assign addr[23027]= 1770014111;
assign addr[23028]= 1924749160;
assign addr[23029]= 2040479063;
assign addr[23030]= 2114858546;
assign addr[23031]= 2146380306;
assign addr[23032]= 2134405552;
assign addr[23033]= 2079176953;
assign addr[23034]= 1981813720;
assign addr[23035]= 1844288924;
assign addr[23036]= 1669389513;
assign addr[23037]= 1460659832;
assign addr[23038]= 1222329801;
assign addr[23039]= 959229189;
assign addr[23040]= 676689746;
assign addr[23041]= 380437148;
assign addr[23042]= 76474970;
assign addr[23043]= -229036977;
assign addr[23044]= -529907477;
assign addr[23045]= -820039373;
assign addr[23046]= -1093553126;
assign addr[23047]= -1344905966;
assign addr[23048]= -1569004214;
assign addr[23049]= -1761306505;
assign addr[23050]= -1917915825;
assign addr[23051]= -2035658475;
assign addr[23052]= -2112148396;
assign addr[23053]= -2145835515;
assign addr[23054]= -2136037160;
assign addr[23055]= -2082951896;
assign addr[23056]= -1987655498;
assign addr[23057]= -1852079154;
assign addr[23058]= -1678970324;
assign addr[23059]= -1471837070;
assign addr[23060]= -1234876957;
assign addr[23061]= -972891995;
assign addr[23062]= -691191324;
assign addr[23063]= -395483624;
assign addr[23064]= -91761426;
assign addr[23065]= 213820322;
assign addr[23066]= 515068990;
assign addr[23067]= 805879757;
assign addr[23068]= 1080359326;
assign addr[23069]= 1332945355;
assign addr[23070]= 1558519173;
assign addr[23071]= 1752509516;
assign addr[23072]= 1910985158;
assign addr[23073]= 2030734582;
assign addr[23074]= 2109331059;
assign addr[23075]= 2145181827;
assign addr[23076]= 2137560369;
assign addr[23077]= 2086621133;
assign addr[23078]= 1993396407;
assign addr[23079]= 1859775393;
assign addr[23080]= 1688465931;
assign addr[23081]= 1482939614;
assign addr[23082]= 1247361445;
assign addr[23083]= 986505429;
assign addr[23084]= 705657826;
assign addr[23085]= 410510029;
assign addr[23086]= 107043224;
assign addr[23087]= -198592817;
assign addr[23088]= -500204365;
assign addr[23089]= -791679244;
assign addr[23090]= -1067110699;
assign addr[23091]= -1320917099;
assign addr[23092]= -1547955041;
assign addr[23093]= -1743623590;
assign addr[23094]= -1903957513;
assign addr[23095]= -2025707632;
assign addr[23096]= -2106406677;
assign addr[23097]= -2144419275;
assign addr[23098]= -2138975100;
assign addr[23099]= -2090184478;
assign addr[23100]= -1999036154;
assign addr[23101]= -1867377253;
assign addr[23102]= -1697875851;
assign addr[23103]= -1493966902;
assign addr[23104]= -1259782632;
assign addr[23105]= -1000068799;
assign addr[23106]= -720088517;
assign addr[23107]= -425515602;
assign addr[23108]= -122319591;
assign addr[23109]= 183355234;
assign addr[23110]= 485314355;
assign addr[23111]= 777438554;
assign addr[23112]= 1053807919;
assign addr[23113]= 1308821808;
assign addr[23114]= 1537312353;
assign addr[23115]= 1734649179;
assign addr[23116]= 1896833245;
assign addr[23117]= 2020577882;
assign addr[23118]= 2103375398;
assign addr[23119]= 2143547897;
assign addr[23120]= 2140281282;
assign addr[23121]= 2093641749;
assign addr[23122]= 2004574453;
assign addr[23123]= 1874884346;
assign addr[23124]= 1707199606;
assign addr[23125]= 1504918373;
assign addr[23126]= 1272139887;
assign addr[23127]= 1013581418;
assign addr[23128]= 734482665;
assign addr[23129]= 440499581;
assign addr[23130]= 137589750;
assign addr[23131]= -168108346;
assign addr[23132]= -470399716;
assign addr[23133]= -763158411;
assign addr[23134]= -1040451659;
assign addr[23135]= -1296660098;
assign addr[23136]= -1526591649;
assign addr[23137]= -1725586737;
assign addr[23138]= -1889612716;
assign addr[23139]= -2015345591;
assign addr[23140]= -2100237377;
assign addr[23141]= -2142567738;
assign addr[23142]= -2141478848;
assign addr[23143]= -2096992772;
assign addr[23144]= -2010011024;
assign addr[23145]= -1882296293;
assign addr[23146]= -1716436725;
assign addr[23147]= -1515793473;
assign addr[23148]= -1284432584;
assign addr[23149]= -1027042599;
assign addr[23150]= -748839539;
assign addr[23151]= -455461206;
assign addr[23152]= -152852926;
assign addr[23153]= 152852926;
assign addr[23154]= 455461206;
assign addr[23155]= 748839539;
assign addr[23156]= 1027042599;
assign addr[23157]= 1284432584;
assign addr[23158]= 1515793473;
assign addr[23159]= 1716436725;
assign addr[23160]= 1882296293;
assign addr[23161]= 2010011024;
assign addr[23162]= 2096992772;
assign addr[23163]= 2141478848;
assign addr[23164]= 2142567738;
assign addr[23165]= 2100237377;
assign addr[23166]= 2015345591;
assign addr[23167]= 1889612716;
assign addr[23168]= 1725586737;
assign addr[23169]= 1526591649;
assign addr[23170]= 1296660098;
assign addr[23171]= 1040451659;
assign addr[23172]= 763158411;
assign addr[23173]= 470399716;
assign addr[23174]= 168108346;
assign addr[23175]= -137589750;
assign addr[23176]= -440499581;
assign addr[23177]= -734482665;
assign addr[23178]= -1013581418;
assign addr[23179]= -1272139887;
assign addr[23180]= -1504918373;
assign addr[23181]= -1707199606;
assign addr[23182]= -1874884346;
assign addr[23183]= -2004574453;
assign addr[23184]= -2093641749;
assign addr[23185]= -2140281282;
assign addr[23186]= -2143547897;
assign addr[23187]= -2103375398;
assign addr[23188]= -2020577882;
assign addr[23189]= -1896833245;
assign addr[23190]= -1734649179;
assign addr[23191]= -1537312353;
assign addr[23192]= -1308821808;
assign addr[23193]= -1053807919;
assign addr[23194]= -777438554;
assign addr[23195]= -485314355;
assign addr[23196]= -183355234;
assign addr[23197]= 122319591;
assign addr[23198]= 425515602;
assign addr[23199]= 720088517;
assign addr[23200]= 1000068799;
assign addr[23201]= 1259782632;
assign addr[23202]= 1493966902;
assign addr[23203]= 1697875851;
assign addr[23204]= 1867377253;
assign addr[23205]= 1999036154;
assign addr[23206]= 2090184478;
assign addr[23207]= 2138975100;
assign addr[23208]= 2144419275;
assign addr[23209]= 2106406677;
assign addr[23210]= 2025707632;
assign addr[23211]= 1903957513;
assign addr[23212]= 1743623590;
assign addr[23213]= 1547955041;
assign addr[23214]= 1320917099;
assign addr[23215]= 1067110699;
assign addr[23216]= 791679244;
assign addr[23217]= 500204365;
assign addr[23218]= 198592817;
assign addr[23219]= -107043224;
assign addr[23220]= -410510029;
assign addr[23221]= -705657826;
assign addr[23222]= -986505429;
assign addr[23223]= -1247361445;
assign addr[23224]= -1482939614;
assign addr[23225]= -1688465931;
assign addr[23226]= -1859775393;
assign addr[23227]= -1993396407;
assign addr[23228]= -2086621133;
assign addr[23229]= -2137560369;
assign addr[23230]= -2145181827;
assign addr[23231]= -2109331059;
assign addr[23232]= -2030734582;
assign addr[23233]= -1910985158;
assign addr[23234]= -1752509516;
assign addr[23235]= -1558519173;
assign addr[23236]= -1332945355;
assign addr[23237]= -1080359326;
assign addr[23238]= -805879757;
assign addr[23239]= -515068990;
assign addr[23240]= -213820322;
assign addr[23241]= 91761426;
assign addr[23242]= 395483624;
assign addr[23243]= 691191324;
assign addr[23244]= 972891995;
assign addr[23245]= 1234876957;
assign addr[23246]= 1471837070;
assign addr[23247]= 1678970324;
assign addr[23248]= 1852079154;
assign addr[23249]= 1987655498;
assign addr[23250]= 2082951896;
assign addr[23251]= 2136037160;
assign addr[23252]= 2145835515;
assign addr[23253]= 2112148396;
assign addr[23254]= 2035658475;
assign addr[23255]= 1917915825;
assign addr[23256]= 1761306505;
assign addr[23257]= 1569004214;
assign addr[23258]= 1344905966;
assign addr[23259]= 1093553126;
assign addr[23260]= 820039373;
assign addr[23261]= 529907477;
assign addr[23262]= 229036977;
assign addr[23263]= -76474970;
assign addr[23264]= -380437148;
assign addr[23265]= -676689746;
assign addr[23266]= -959229189;
assign addr[23267]= -1222329801;
assign addr[23268]= -1460659832;
assign addr[23269]= -1669389513;
assign addr[23270]= -1844288924;
assign addr[23271]= -1981813720;
assign addr[23272]= -2079176953;
assign addr[23273]= -2134405552;
assign addr[23274]= -2146380306;
assign addr[23275]= -2114858546;
assign addr[23276]= -2040479063;
assign addr[23277]= -1924749160;
assign addr[23278]= -1770014111;
assign addr[23279]= -1579409630;
assign addr[23280]= -1356798326;
assign addr[23281]= -1106691431;
assign addr[23282]= -834157373;
assign addr[23283]= -544719071;
assign addr[23284]= -244242007;
assign addr[23285]= 61184634;
assign addr[23286]= 365371365;
assign addr[23287]= 662153826;
assign addr[23288]= 945517704;
assign addr[23289]= 1209720613;
assign addr[23290]= 1449408469;
assign addr[23291]= 1659723983;
assign addr[23292]= 1836405100;
assign addr[23293]= 1975871368;
assign addr[23294]= 2075296495;
assign addr[23295]= 2132665626;
assign addr[23296]= 2146816171;
assign addr[23297]= 2117461370;
assign addr[23298]= 2045196100;
assign addr[23299]= 1931484818;
assign addr[23300]= 1778631892;
assign addr[23301]= 1589734894;
assign addr[23302]= 1368621831;
assign addr[23303]= 1119773573;
assign addr[23304]= 848233042;
assign addr[23305]= 559503022;
assign addr[23306]= 259434643;
assign addr[23307]= -45891193;
assign addr[23308]= -350287041;
assign addr[23309]= -647584304;
assign addr[23310]= -931758235;
assign addr[23311]= -1197050035;
assign addr[23312]= -1438083551;
assign addr[23313]= -1649974225;
assign addr[23314]= -1828428082;
assign addr[23315]= -1969828744;
assign addr[23316]= -2071310720;
assign addr[23317]= -2130817471;
assign addr[23318]= -2147143090;
assign addr[23319]= -2119956737;
assign addr[23320]= -2049809346;
assign addr[23321]= -1938122457;
assign addr[23322]= -1787159411;
assign addr[23323]= -1599979481;
assign addr[23324]= -1380375881;
assign addr[23325]= -1132798888;
assign addr[23326]= -862265664;
assign addr[23327]= -574258580;
assign addr[23328]= -274614114;
assign addr[23329]= 30595422;
assign addr[23330]= 335184940;
assign addr[23331]= 632981917;
assign addr[23332]= 917951481;
assign addr[23333]= 1184318708;
assign addr[23334]= 1426685652;
assign addr[23335]= 1640140734;
assign addr[23336]= 1820358275;
assign addr[23337]= 1963686155;
assign addr[23338]= 2067219829;
assign addr[23339]= 2128861181;
assign addr[23340]= 2147361045;
assign addr[23341]= 2122344521;
assign addr[23342]= 2054318569;
assign addr[23343]= 1944661739;
assign addr[23344]= 1795596234;
assign addr[23345]= 1610142873;
assign addr[23346]= 1392059879;
assign addr[23347]= 1145766716;
assign addr[23348]= 876254528;
assign addr[23349]= 588984994;
assign addr[23350]= 289779648;
assign addr[23351]= -15298099;
assign addr[23352]= -320065829;
assign addr[23353]= -618347408;
assign addr[23354]= -904098143;
assign addr[23355]= -1171527280;
assign addr[23356]= -1415215352;
assign addr[23357]= -1630224009;
assign addr[23358]= -1812196087;
assign addr[23359]= -1957443913;
assign addr[23360]= -2063024031;
assign addr[23361]= -2126796855;
assign addr[23362]= -2147470025;
assign addr[23363]= -2124624598;
assign addr[23364]= -2058723538;
assign addr[23365]= -1951102334;
assign addr[23366]= -1803941934;
assign addr[23367]= -1620224553;
assign addr[23368]= -1403673233;
assign addr[23369]= -1158676398;
assign addr[23370]= -890198924;
assign addr[23371]= -603681519;
assign addr[23372]= -304930476;
assign addr[23373]= 0;
assign addr[23374]= 304930476;
assign addr[23375]= 603681519;
assign addr[23376]= 890198924;
assign addr[23377]= 1158676398;
assign addr[23378]= 1403673233;
assign addr[23379]= 1620224553;
assign addr[23380]= 1803941934;
assign addr[23381]= 1951102334;
assign addr[23382]= 2058723538;
assign addr[23383]= 2124624598;
assign addr[23384]= 2147470025;
assign addr[23385]= 2126796855;
assign addr[23386]= 2063024031;
assign addr[23387]= 1957443913;
assign addr[23388]= 1812196087;
assign addr[23389]= 1630224009;
assign addr[23390]= 1415215352;
assign addr[23391]= 1171527280;
assign addr[23392]= 904098143;
assign addr[23393]= 618347408;
assign addr[23394]= 320065829;
assign addr[23395]= 15298099;
assign addr[23396]= -289779648;
assign addr[23397]= -588984994;
assign addr[23398]= -876254528;
assign addr[23399]= -1145766716;
assign addr[23400]= -1392059879;
assign addr[23401]= -1610142873;
assign addr[23402]= -1795596234;
assign addr[23403]= -1944661739;
assign addr[23404]= -2054318569;
assign addr[23405]= -2122344521;
assign addr[23406]= -2147361045;
assign addr[23407]= -2128861181;
assign addr[23408]= -2067219829;
assign addr[23409]= -1963686155;
assign addr[23410]= -1820358275;
assign addr[23411]= -1640140734;
assign addr[23412]= -1426685652;
assign addr[23413]= -1184318708;
assign addr[23414]= -917951481;
assign addr[23415]= -632981917;
assign addr[23416]= -335184940;
assign addr[23417]= -30595422;
assign addr[23418]= 274614114;
assign addr[23419]= 574258580;
assign addr[23420]= 862265664;
assign addr[23421]= 1132798888;
assign addr[23422]= 1380375881;
assign addr[23423]= 1599979481;
assign addr[23424]= 1787159411;
assign addr[23425]= 1938122457;
assign addr[23426]= 2049809346;
assign addr[23427]= 2119956737;
assign addr[23428]= 2147143090;
assign addr[23429]= 2130817471;
assign addr[23430]= 2071310720;
assign addr[23431]= 1969828744;
assign addr[23432]= 1828428082;
assign addr[23433]= 1649974225;
assign addr[23434]= 1438083551;
assign addr[23435]= 1197050035;
assign addr[23436]= 931758235;
assign addr[23437]= 647584304;
assign addr[23438]= 350287041;
assign addr[23439]= 45891193;
assign addr[23440]= -259434643;
assign addr[23441]= -559503022;
assign addr[23442]= -848233042;
assign addr[23443]= -1119773573;
assign addr[23444]= -1368621831;
assign addr[23445]= -1589734894;
assign addr[23446]= -1778631892;
assign addr[23447]= -1931484818;
assign addr[23448]= -2045196100;
assign addr[23449]= -2117461370;
assign addr[23450]= -2146816171;
assign addr[23451]= -2132665626;
assign addr[23452]= -2075296495;
assign addr[23453]= -1975871368;
assign addr[23454]= -1836405100;
assign addr[23455]= -1659723983;
assign addr[23456]= -1449408469;
assign addr[23457]= -1209720613;
assign addr[23458]= -945517704;
assign addr[23459]= -662153826;
assign addr[23460]= -365371365;
assign addr[23461]= -61184634;
assign addr[23462]= 244242007;
assign addr[23463]= 544719071;
assign addr[23464]= 834157373;
assign addr[23465]= 1106691431;
assign addr[23466]= 1356798326;
assign addr[23467]= 1579409630;
assign addr[23468]= 1770014111;
assign addr[23469]= 1924749160;
assign addr[23470]= 2040479063;
assign addr[23471]= 2114858546;
assign addr[23472]= 2146380306;
assign addr[23473]= 2134405552;
assign addr[23474]= 2079176953;
assign addr[23475]= 1981813720;
assign addr[23476]= 1844288924;
assign addr[23477]= 1669389513;
assign addr[23478]= 1460659832;
assign addr[23479]= 1222329801;
assign addr[23480]= 959229189;
assign addr[23481]= 676689746;
assign addr[23482]= 380437148;
assign addr[23483]= 76474970;
assign addr[23484]= -229036977;
assign addr[23485]= -529907477;
assign addr[23486]= -820039373;
assign addr[23487]= -1093553126;
assign addr[23488]= -1344905966;
assign addr[23489]= -1569004214;
assign addr[23490]= -1761306505;
assign addr[23491]= -1917915825;
assign addr[23492]= -2035658475;
assign addr[23493]= -2112148396;
assign addr[23494]= -2145835515;
assign addr[23495]= -2136037160;
assign addr[23496]= -2082951896;
assign addr[23497]= -1987655498;
assign addr[23498]= -1852079154;
assign addr[23499]= -1678970324;
assign addr[23500]= -1471837070;
assign addr[23501]= -1234876957;
assign addr[23502]= -972891995;
assign addr[23503]= -691191324;
assign addr[23504]= -395483624;
assign addr[23505]= -91761426;
assign addr[23506]= 213820322;
assign addr[23507]= 515068990;
assign addr[23508]= 805879757;
assign addr[23509]= 1080359326;
assign addr[23510]= 1332945355;
assign addr[23511]= 1558519173;
assign addr[23512]= 1752509516;
assign addr[23513]= 1910985158;
assign addr[23514]= 2030734582;
assign addr[23515]= 2109331059;
assign addr[23516]= 2145181827;
assign addr[23517]= 2137560369;
assign addr[23518]= 2086621133;
assign addr[23519]= 1993396407;
assign addr[23520]= 1859775393;
assign addr[23521]= 1688465931;
assign addr[23522]= 1482939614;
assign addr[23523]= 1247361445;
assign addr[23524]= 986505429;
assign addr[23525]= 705657826;
assign addr[23526]= 410510029;
assign addr[23527]= 107043224;
assign addr[23528]= -198592817;
assign addr[23529]= -500204365;
assign addr[23530]= -791679244;
assign addr[23531]= -1067110699;
assign addr[23532]= -1320917099;
assign addr[23533]= -1547955041;
assign addr[23534]= -1743623590;
assign addr[23535]= -1903957513;
assign addr[23536]= -2025707632;
assign addr[23537]= -2106406677;
assign addr[23538]= -2144419275;
assign addr[23539]= -2138975100;
assign addr[23540]= -2090184478;
assign addr[23541]= -1999036154;
assign addr[23542]= -1867377253;
assign addr[23543]= -1697875851;
assign addr[23544]= -1493966902;
assign addr[23545]= -1259782632;
assign addr[23546]= -1000068799;
assign addr[23547]= -720088517;
assign addr[23548]= -425515602;
assign addr[23549]= -122319591;
assign addr[23550]= 183355234;
assign addr[23551]= 485314355;
assign addr[23552]= 777438554;
assign addr[23553]= 1053807919;
assign addr[23554]= 1308821808;
assign addr[23555]= 1537312353;
assign addr[23556]= 1734649179;
assign addr[23557]= 1896833245;
assign addr[23558]= 2020577882;
assign addr[23559]= 2103375398;
assign addr[23560]= 2143547897;
assign addr[23561]= 2140281282;
assign addr[23562]= 2093641749;
assign addr[23563]= 2004574453;
assign addr[23564]= 1874884346;
assign addr[23565]= 1707199606;
assign addr[23566]= 1504918373;
assign addr[23567]= 1272139887;
assign addr[23568]= 1013581418;
assign addr[23569]= 734482665;
assign addr[23570]= 440499581;
assign addr[23571]= 137589750;
assign addr[23572]= -168108346;
assign addr[23573]= -470399716;
assign addr[23574]= -763158411;
assign addr[23575]= -1040451659;
assign addr[23576]= -1296660098;
assign addr[23577]= -1526591649;
assign addr[23578]= -1725586737;
assign addr[23579]= -1889612716;
assign addr[23580]= -2015345591;
assign addr[23581]= -2100237377;
assign addr[23582]= -2142567738;
assign addr[23583]= -2141478848;
assign addr[23584]= -2096992772;
assign addr[23585]= -2010011024;
assign addr[23586]= -1882296293;
assign addr[23587]= -1716436725;
assign addr[23588]= -1515793473;
assign addr[23589]= -1284432584;
assign addr[23590]= -1027042599;
assign addr[23591]= -748839539;
assign addr[23592]= -455461206;
assign addr[23593]= -152852926;
assign addr[23594]= 152852926;
assign addr[23595]= 455461206;
assign addr[23596]= 748839539;
assign addr[23597]= 1027042599;
assign addr[23598]= 1284432584;
assign addr[23599]= 1515793473;
assign addr[23600]= 1716436725;
assign addr[23601]= 1882296293;
assign addr[23602]= 2010011024;
assign addr[23603]= 2096992772;
assign addr[23604]= 2141478848;
assign addr[23605]= 2142567738;
assign addr[23606]= 2100237377;
assign addr[23607]= 2015345591;
assign addr[23608]= 1889612716;
assign addr[23609]= 1725586737;
assign addr[23610]= 1526591649;
assign addr[23611]= 1296660098;
assign addr[23612]= 1040451659;
assign addr[23613]= 763158411;
assign addr[23614]= 470399716;
assign addr[23615]= 168108346;
assign addr[23616]= -137589750;
assign addr[23617]= -440499581;
assign addr[23618]= -734482665;
assign addr[23619]= -1013581418;
assign addr[23620]= -1272139887;
assign addr[23621]= -1504918373;
assign addr[23622]= -1707199606;
assign addr[23623]= -1874884346;
assign addr[23624]= -2004574453;
assign addr[23625]= -2093641749;
assign addr[23626]= -2140281282;
assign addr[23627]= -2143547897;
assign addr[23628]= -2103375398;
assign addr[23629]= -2020577882;
assign addr[23630]= -1896833245;
assign addr[23631]= -1734649179;
assign addr[23632]= -1537312353;
assign addr[23633]= -1308821808;
assign addr[23634]= -1053807919;
assign addr[23635]= -777438554;
assign addr[23636]= -485314355;
assign addr[23637]= -183355234;
assign addr[23638]= 122319591;
assign addr[23639]= 425515602;
assign addr[23640]= 720088517;
assign addr[23641]= 1000068799;
assign addr[23642]= 1259782632;
assign addr[23643]= 1493966902;
assign addr[23644]= 1697875851;
assign addr[23645]= 1867377253;
assign addr[23646]= 1999036154;
assign addr[23647]= 2090184478;
assign addr[23648]= 2138975100;
assign addr[23649]= 2144419275;
assign addr[23650]= 2106406677;
assign addr[23651]= 2025707632;
assign addr[23652]= 1903957513;
assign addr[23653]= 1743623590;
assign addr[23654]= 1547955041;
assign addr[23655]= 1320917099;
assign addr[23656]= 1067110699;
assign addr[23657]= 791679244;
assign addr[23658]= 500204365;
assign addr[23659]= 198592817;
assign addr[23660]= -107043224;
assign addr[23661]= -410510029;
assign addr[23662]= -705657826;
assign addr[23663]= -986505429;
assign addr[23664]= -1247361445;
assign addr[23665]= -1482939614;
assign addr[23666]= -1688465931;
assign addr[23667]= -1859775393;
assign addr[23668]= -1993396407;
assign addr[23669]= -2086621133;
assign addr[23670]= -2137560369;
assign addr[23671]= -2145181827;
assign addr[23672]= -2109331059;
assign addr[23673]= -2030734582;
assign addr[23674]= -1910985158;
assign addr[23675]= -1752509516;
assign addr[23676]= -1558519173;
assign addr[23677]= -1332945355;
assign addr[23678]= -1080359326;
assign addr[23679]= -805879757;
assign addr[23680]= -515068990;
assign addr[23681]= -213820322;
assign addr[23682]= 91761426;
assign addr[23683]= 395483624;
assign addr[23684]= 691191324;
assign addr[23685]= 972891995;
assign addr[23686]= 1234876957;
assign addr[23687]= 1471837070;
assign addr[23688]= 1678970324;
assign addr[23689]= 1852079154;
assign addr[23690]= 1987655498;
assign addr[23691]= 2082951896;
assign addr[23692]= 2136037160;
assign addr[23693]= 2145835515;
assign addr[23694]= 2112148396;
assign addr[23695]= 2035658475;
assign addr[23696]= 1917915825;
assign addr[23697]= 1761306505;
assign addr[23698]= 1569004214;
assign addr[23699]= 1344905966;
assign addr[23700]= 1093553126;
assign addr[23701]= 820039373;
assign addr[23702]= 529907477;
assign addr[23703]= 229036977;
assign addr[23704]= -76474970;
assign addr[23705]= -380437148;
assign addr[23706]= -676689746;
assign addr[23707]= -959229189;
assign addr[23708]= -1222329801;
assign addr[23709]= -1460659832;
assign addr[23710]= -1669389513;
assign addr[23711]= -1844288924;
assign addr[23712]= -1981813720;
assign addr[23713]= -2079176953;
assign addr[23714]= -2134405552;
assign addr[23715]= -2146380306;
assign addr[23716]= -2114858546;
assign addr[23717]= -2040479063;
assign addr[23718]= -1924749160;
assign addr[23719]= -1770014111;
assign addr[23720]= -1579409630;
assign addr[23721]= -1356798326;
assign addr[23722]= -1106691431;
assign addr[23723]= -834157373;
assign addr[23724]= -544719071;
assign addr[23725]= -244242007;
assign addr[23726]= 61184634;
assign addr[23727]= 365371365;
assign addr[23728]= 662153826;
assign addr[23729]= 945517704;
assign addr[23730]= 1209720613;
assign addr[23731]= 1449408469;
assign addr[23732]= 1659723983;
assign addr[23733]= 1836405100;
assign addr[23734]= 1975871368;
assign addr[23735]= 2075296495;
assign addr[23736]= 2132665626;
assign addr[23737]= 2146816171;
assign addr[23738]= 2117461370;
assign addr[23739]= 2045196100;
assign addr[23740]= 1931484818;
assign addr[23741]= 1778631892;
assign addr[23742]= 1589734894;
assign addr[23743]= 1368621831;
assign addr[23744]= 1119773573;
assign addr[23745]= 848233042;
assign addr[23746]= 559503022;
assign addr[23747]= 259434643;
assign addr[23748]= -45891193;
assign addr[23749]= -350287041;
assign addr[23750]= -647584304;
assign addr[23751]= -931758235;
assign addr[23752]= -1197050035;
assign addr[23753]= -1438083551;
assign addr[23754]= -1649974225;
assign addr[23755]= -1828428082;
assign addr[23756]= -1969828744;
assign addr[23757]= -2071310720;
assign addr[23758]= -2130817471;
assign addr[23759]= -2147143090;
assign addr[23760]= -2119956737;
assign addr[23761]= -2049809346;
assign addr[23762]= -1938122457;
assign addr[23763]= -1787159411;
assign addr[23764]= -1599979481;
assign addr[23765]= -1380375881;
assign addr[23766]= -1132798888;
assign addr[23767]= -862265664;
assign addr[23768]= -574258580;
assign addr[23769]= -274614114;
assign addr[23770]= 30595422;
assign addr[23771]= 335184940;
assign addr[23772]= 632981917;
assign addr[23773]= 917951481;
assign addr[23774]= 1184318708;
assign addr[23775]= 1426685652;
assign addr[23776]= 1640140734;
assign addr[23777]= 1820358275;
assign addr[23778]= 1963686155;
assign addr[23779]= 2067219829;
assign addr[23780]= 2128861181;
assign addr[23781]= 2147361045;
assign addr[23782]= 2122344521;
assign addr[23783]= 2054318569;
assign addr[23784]= 1944661739;
assign addr[23785]= 1795596234;
assign addr[23786]= 1610142873;
assign addr[23787]= 1392059879;
assign addr[23788]= 1145766716;
assign addr[23789]= 876254528;
assign addr[23790]= 588984994;
assign addr[23791]= 289779648;
assign addr[23792]= -15298099;
assign addr[23793]= -320065829;
assign addr[23794]= -618347408;
assign addr[23795]= -904098143;
assign addr[23796]= -1171527280;
assign addr[23797]= -1415215352;
assign addr[23798]= -1630224009;
assign addr[23799]= -1812196087;
assign addr[23800]= -1957443913;
assign addr[23801]= -2063024031;
assign addr[23802]= -2126796855;
assign addr[23803]= -2147470025;
assign addr[23804]= -2124624598;
assign addr[23805]= -2058723538;
assign addr[23806]= -1951102334;
assign addr[23807]= -1803941934;
assign addr[23808]= -1620224553;
assign addr[23809]= -1403673233;
assign addr[23810]= -1158676398;
assign addr[23811]= -890198924;
assign addr[23812]= -603681519;
assign addr[23813]= -304930476;
assign addr[23814]= 0;
assign addr[23815]= 304930476;
assign addr[23816]= 603681519;
assign addr[23817]= 890198924;
assign addr[23818]= 1158676398;
assign addr[23819]= 1403673233;
assign addr[23820]= 1620224553;
assign addr[23821]= 1803941934;
assign addr[23822]= 1951102334;
assign addr[23823]= 2058723538;
assign addr[23824]= 2124624598;
assign addr[23825]= 2147470025;
assign addr[23826]= 2126796855;
assign addr[23827]= 2063024031;
assign addr[23828]= 1957443913;
assign addr[23829]= 1812196087;
assign addr[23830]= 1630224009;
assign addr[23831]= 1415215352;
assign addr[23832]= 1171527280;
assign addr[23833]= 904098143;
assign addr[23834]= 618347408;
assign addr[23835]= 320065829;
assign addr[23836]= 15298099;
assign addr[23837]= -289779648;
assign addr[23838]= -588984994;
assign addr[23839]= -876254528;
assign addr[23840]= -1145766716;
assign addr[23841]= -1392059879;
assign addr[23842]= -1610142873;
assign addr[23843]= -1795596234;
assign addr[23844]= -1944661739;
assign addr[23845]= -2054318569;
assign addr[23846]= -2122344521;
assign addr[23847]= -2147361045;
assign addr[23848]= -2128861181;
assign addr[23849]= -2067219829;
assign addr[23850]= -1963686155;
assign addr[23851]= -1820358275;
assign addr[23852]= -1640140734;
assign addr[23853]= -1426685652;
assign addr[23854]= -1184318708;
assign addr[23855]= -917951481;
assign addr[23856]= -632981917;
assign addr[23857]= -335184940;
assign addr[23858]= -30595422;
assign addr[23859]= 274614114;
assign addr[23860]= 574258580;
assign addr[23861]= 862265664;
assign addr[23862]= 1132798888;
assign addr[23863]= 1380375881;
assign addr[23864]= 1599979481;
assign addr[23865]= 1787159411;
assign addr[23866]= 1938122457;
assign addr[23867]= 2049809346;
assign addr[23868]= 2119956737;
assign addr[23869]= 2147143090;
assign addr[23870]= 2130817471;
assign addr[23871]= 2071310720;
assign addr[23872]= 1969828744;
assign addr[23873]= 1828428082;
assign addr[23874]= 1649974225;
assign addr[23875]= 1438083551;
assign addr[23876]= 1197050035;
assign addr[23877]= 931758235;
assign addr[23878]= 647584304;
assign addr[23879]= 350287041;
assign addr[23880]= 45891193;
assign addr[23881]= -259434643;
assign addr[23882]= -559503022;
assign addr[23883]= -848233042;
assign addr[23884]= -1119773573;
assign addr[23885]= -1368621831;
assign addr[23886]= -1589734894;
assign addr[23887]= -1778631892;
assign addr[23888]= -1931484818;
assign addr[23889]= -2045196100;
assign addr[23890]= -2117461370;
assign addr[23891]= -2146816171;
assign addr[23892]= -2132665626;
assign addr[23893]= -2075296495;
assign addr[23894]= -1975871368;
assign addr[23895]= -1836405100;
assign addr[23896]= -1659723983;
assign addr[23897]= -1449408469;
assign addr[23898]= -1209720613;
assign addr[23899]= -945517704;
assign addr[23900]= -662153826;
assign addr[23901]= -365371365;
assign addr[23902]= -61184634;
assign addr[23903]= 244242007;
assign addr[23904]= 544719071;
assign addr[23905]= 834157373;
assign addr[23906]= 1106691431;
assign addr[23907]= 1356798326;
assign addr[23908]= 1579409630;
assign addr[23909]= 1770014111;
assign addr[23910]= 1924749160;
assign addr[23911]= 2040479063;
assign addr[23912]= 2114858546;
assign addr[23913]= 2146380306;
assign addr[23914]= 2134405552;
assign addr[23915]= 2079176953;
assign addr[23916]= 1981813720;
assign addr[23917]= 1844288924;
assign addr[23918]= 1669389513;
assign addr[23919]= 1460659832;
assign addr[23920]= 1222329801;
assign addr[23921]= 959229189;
assign addr[23922]= 676689746;
assign addr[23923]= 380437148;
assign addr[23924]= 76474970;
assign addr[23925]= -229036977;
assign addr[23926]= -529907477;
assign addr[23927]= -820039373;
assign addr[23928]= -1093553126;
assign addr[23929]= -1344905966;
assign addr[23930]= -1569004214;
assign addr[23931]= -1761306505;
assign addr[23932]= -1917915825;
assign addr[23933]= -2035658475;
assign addr[23934]= -2112148396;
assign addr[23935]= -2145835515;
assign addr[23936]= -2136037160;
assign addr[23937]= -2082951896;
assign addr[23938]= -1987655498;
assign addr[23939]= -1852079154;
assign addr[23940]= -1678970324;
assign addr[23941]= -1471837070;
assign addr[23942]= -1234876957;
assign addr[23943]= -972891995;
assign addr[23944]= -691191324;
assign addr[23945]= -395483624;
assign addr[23946]= -91761426;
assign addr[23947]= 213820322;
assign addr[23948]= 515068990;
assign addr[23949]= 805879757;
assign addr[23950]= 1080359326;
assign addr[23951]= 1332945355;
assign addr[23952]= 1558519173;
assign addr[23953]= 1752509516;
assign addr[23954]= 1910985158;
assign addr[23955]= 2030734582;
assign addr[23956]= 2109331059;
assign addr[23957]= 2145181827;
assign addr[23958]= 2137560369;
assign addr[23959]= 2086621133;
assign addr[23960]= 1993396407;
assign addr[23961]= 1859775393;
assign addr[23962]= 1688465931;
assign addr[23963]= 1482939614;
assign addr[23964]= 1247361445;
assign addr[23965]= 986505429;
assign addr[23966]= 705657826;
assign addr[23967]= 410510029;
assign addr[23968]= 107043224;
assign addr[23969]= -198592817;
assign addr[23970]= -500204365;
assign addr[23971]= -791679244;
assign addr[23972]= -1067110699;
assign addr[23973]= -1320917099;
assign addr[23974]= -1547955041;
assign addr[23975]= -1743623590;
assign addr[23976]= -1903957513;
assign addr[23977]= -2025707632;
assign addr[23978]= -2106406677;
assign addr[23979]= -2144419275;
assign addr[23980]= -2138975100;
assign addr[23981]= -2090184478;
assign addr[23982]= -1999036154;
assign addr[23983]= -1867377253;
assign addr[23984]= -1697875851;
assign addr[23985]= -1493966902;
assign addr[23986]= -1259782632;
assign addr[23987]= -1000068799;
assign addr[23988]= -720088517;
assign addr[23989]= -425515602;
assign addr[23990]= -122319591;
assign addr[23991]= 183355234;
assign addr[23992]= 485314355;
assign addr[23993]= 777438554;
assign addr[23994]= 1053807919;
assign addr[23995]= 1308821808;
assign addr[23996]= 1537312353;
assign addr[23997]= 1734649179;
assign addr[23998]= 1896833245;
assign addr[23999]= 2020577882;
assign addr[24000]= 2103375398;
assign addr[24001]= 2143547897;
assign addr[24002]= 2140281282;
assign addr[24003]= 2093641749;
assign addr[24004]= 2004574453;
assign addr[24005]= 1874884346;
assign addr[24006]= 1707199606;
assign addr[24007]= 1504918373;
assign addr[24008]= 1272139887;
assign addr[24009]= 1013581418;
assign addr[24010]= 734482665;
assign addr[24011]= 440499581;
assign addr[24012]= 137589750;
assign addr[24013]= -168108346;
assign addr[24014]= -470399716;
assign addr[24015]= -763158411;
assign addr[24016]= -1040451659;
assign addr[24017]= -1296660098;
assign addr[24018]= -1526591649;
assign addr[24019]= -1725586737;
assign addr[24020]= -1889612716;
assign addr[24021]= -2015345591;
assign addr[24022]= -2100237377;
assign addr[24023]= -2142567738;
assign addr[24024]= -2141478848;
assign addr[24025]= -2096992772;
assign addr[24026]= -2010011024;
assign addr[24027]= -1882296293;
assign addr[24028]= -1716436725;
assign addr[24029]= -1515793473;
assign addr[24030]= -1284432584;
assign addr[24031]= -1027042599;
assign addr[24032]= -748839539;
assign addr[24033]= -455461206;
assign addr[24034]= -152852926;
assign addr[24035]= 152852926;
assign addr[24036]= 455461206;
assign addr[24037]= 748839539;
assign addr[24038]= 1027042599;
assign addr[24039]= 1284432584;
assign addr[24040]= 1515793473;
assign addr[24041]= 1716436725;
assign addr[24042]= 1882296293;
assign addr[24043]= 2010011024;
assign addr[24044]= 2096992772;
assign addr[24045]= 2141478848;
assign addr[24046]= 2142567738;
assign addr[24047]= 2100237377;
assign addr[24048]= 2015345591;
assign addr[24049]= 1889612716;
assign addr[24050]= 1725586737;
assign addr[24051]= 1526591649;
assign addr[24052]= 1296660098;
assign addr[24053]= 1040451659;
assign addr[24054]= 763158411;
assign addr[24055]= 470399716;
assign addr[24056]= 168108346;
assign addr[24057]= -137589750;
assign addr[24058]= -440499581;
assign addr[24059]= -734482665;
assign addr[24060]= -1013581418;
assign addr[24061]= -1272139887;
assign addr[24062]= -1504918373;
assign addr[24063]= -1707199606;
assign addr[24064]= -1874884346;
assign addr[24065]= -2004574453;
assign addr[24066]= -2093641749;
assign addr[24067]= -2140281282;
assign addr[24068]= -2143547897;
assign addr[24069]= -2103375398;
assign addr[24070]= -2020577882;
assign addr[24071]= -1896833245;
assign addr[24072]= -1734649179;
assign addr[24073]= -1537312353;
assign addr[24074]= -1308821808;
assign addr[24075]= -1053807919;
assign addr[24076]= -777438554;
assign addr[24077]= -485314355;
assign addr[24078]= -183355234;
assign addr[24079]= 122319591;
assign addr[24080]= 425515602;
assign addr[24081]= 720088517;
assign addr[24082]= 1000068799;
assign addr[24083]= 1259782632;
assign addr[24084]= 1493966902;
assign addr[24085]= 1697875851;
assign addr[24086]= 1867377253;
assign addr[24087]= 1999036154;
assign addr[24088]= 2090184478;
assign addr[24089]= 2138975100;
assign addr[24090]= 2144419275;
assign addr[24091]= 2106406677;
assign addr[24092]= 2025707632;
assign addr[24093]= 1903957513;
assign addr[24094]= 1743623590;
assign addr[24095]= 1547955041;
assign addr[24096]= 1320917099;
assign addr[24097]= 1067110699;
assign addr[24098]= 791679244;
assign addr[24099]= 500204365;
assign addr[24100]= 198592817;
assign addr[24101]= -107043224;
assign addr[24102]= -410510029;
assign addr[24103]= -705657826;
assign addr[24104]= -986505429;
assign addr[24105]= -1247361445;
assign addr[24106]= -1482939614;
assign addr[24107]= -1688465931;
assign addr[24108]= -1859775393;
assign addr[24109]= -1993396407;
assign addr[24110]= -2086621133;
assign addr[24111]= -2137560369;
assign addr[24112]= -2145181827;
assign addr[24113]= -2109331059;
assign addr[24114]= -2030734582;
assign addr[24115]= -1910985158;
assign addr[24116]= -1752509516;
assign addr[24117]= -1558519173;
assign addr[24118]= -1332945355;
assign addr[24119]= -1080359326;
assign addr[24120]= -805879757;
assign addr[24121]= -515068990;
assign addr[24122]= -213820322;
assign addr[24123]= 91761426;
assign addr[24124]= 395483624;
assign addr[24125]= 691191324;
assign addr[24126]= 972891995;
assign addr[24127]= 1234876957;
assign addr[24128]= 1471837070;
assign addr[24129]= 1678970324;
assign addr[24130]= 1852079154;
assign addr[24131]= 1987655498;
assign addr[24132]= 2082951896;
assign addr[24133]= 2136037160;
assign addr[24134]= 2145835515;
assign addr[24135]= 2112148396;
assign addr[24136]= 2035658475;
assign addr[24137]= 1917915825;
assign addr[24138]= 1761306505;
assign addr[24139]= 1569004214;
assign addr[24140]= 1344905966;
assign addr[24141]= 1093553126;
assign addr[24142]= 820039373;
assign addr[24143]= 529907477;
assign addr[24144]= 229036977;
assign addr[24145]= -76474970;
assign addr[24146]= -380437148;
assign addr[24147]= -676689746;
assign addr[24148]= -959229189;
assign addr[24149]= -1222329801;
assign addr[24150]= -1460659832;
assign addr[24151]= -1669389513;
assign addr[24152]= -1844288924;
assign addr[24153]= -1981813720;
assign addr[24154]= -2079176953;
assign addr[24155]= -2134405552;
assign addr[24156]= -2146380306;
assign addr[24157]= -2114858546;
assign addr[24158]= -2040479063;
assign addr[24159]= -1924749160;
assign addr[24160]= -1770014111;
assign addr[24161]= -1579409630;
assign addr[24162]= -1356798326;
assign addr[24163]= -1106691431;
assign addr[24164]= -834157373;
assign addr[24165]= -544719071;
assign addr[24166]= -244242007;
assign addr[24167]= 61184634;
assign addr[24168]= 365371365;
assign addr[24169]= 662153826;
assign addr[24170]= 945517704;
assign addr[24171]= 1209720613;
assign addr[24172]= 1449408469;
assign addr[24173]= 1659723983;
assign addr[24174]= 1836405100;
assign addr[24175]= 1975871368;
assign addr[24176]= 2075296495;
assign addr[24177]= 2132665626;
assign addr[24178]= 2146816171;
assign addr[24179]= 2117461370;
assign addr[24180]= 2045196100;
assign addr[24181]= 1931484818;
assign addr[24182]= 1778631892;
assign addr[24183]= 1589734894;
assign addr[24184]= 1368621831;
assign addr[24185]= 1119773573;
assign addr[24186]= 848233042;
assign addr[24187]= 559503022;
assign addr[24188]= 259434643;
assign addr[24189]= -45891193;
assign addr[24190]= -350287041;
assign addr[24191]= -647584304;
assign addr[24192]= -931758235;
assign addr[24193]= -1197050035;
assign addr[24194]= -1438083551;
assign addr[24195]= -1649974225;
assign addr[24196]= -1828428082;
assign addr[24197]= -1969828744;
assign addr[24198]= -2071310720;
assign addr[24199]= -2130817471;
assign addr[24200]= -2147143090;
assign addr[24201]= -2119956737;
assign addr[24202]= -2049809346;
assign addr[24203]= -1938122457;
assign addr[24204]= -1787159411;
assign addr[24205]= -1599979481;
assign addr[24206]= -1380375881;
assign addr[24207]= -1132798888;
assign addr[24208]= -862265664;
assign addr[24209]= -574258580;
assign addr[24210]= -274614114;
assign addr[24211]= 30595422;
assign addr[24212]= 335184940;
assign addr[24213]= 632981917;
assign addr[24214]= 917951481;
assign addr[24215]= 1184318708;
assign addr[24216]= 1426685652;
assign addr[24217]= 1640140734;
assign addr[24218]= 1820358275;
assign addr[24219]= 1963686155;
assign addr[24220]= 2067219829;
assign addr[24221]= 2128861181;
assign addr[24222]= 2147361045;
assign addr[24223]= 2122344521;
assign addr[24224]= 2054318569;
assign addr[24225]= 1944661739;
assign addr[24226]= 1795596234;
assign addr[24227]= 1610142873;
assign addr[24228]= 1392059879;
assign addr[24229]= 1145766716;
assign addr[24230]= 876254528;
assign addr[24231]= 588984994;
assign addr[24232]= 289779648;
assign addr[24233]= -15298099;
assign addr[24234]= -320065829;
assign addr[24235]= -618347408;
assign addr[24236]= -904098143;
assign addr[24237]= -1171527280;
assign addr[24238]= -1415215352;
assign addr[24239]= -1630224009;
assign addr[24240]= -1812196087;
assign addr[24241]= -1957443913;
assign addr[24242]= -2063024031;
assign addr[24243]= -2126796855;
assign addr[24244]= -2147470025;
assign addr[24245]= -2124624598;
assign addr[24246]= -2058723538;
assign addr[24247]= -1951102334;
assign addr[24248]= -1803941934;
assign addr[24249]= -1620224553;
assign addr[24250]= -1403673233;
assign addr[24251]= -1158676398;
assign addr[24252]= -890198924;
assign addr[24253]= -603681519;
assign addr[24254]= -304930476;
assign addr[24255]= 0;
assign addr[24256]= 304930476;
assign addr[24257]= 603681519;
assign addr[24258]= 890198924;
assign addr[24259]= 1158676398;
assign addr[24260]= 1403673233;
assign addr[24261]= 1620224553;
assign addr[24262]= 1803941934;
assign addr[24263]= 1951102334;
assign addr[24264]= 2058723538;
assign addr[24265]= 2124624598;
assign addr[24266]= 2147470025;
assign addr[24267]= 2126796855;
assign addr[24268]= 2063024031;
assign addr[24269]= 1957443913;
assign addr[24270]= 1812196087;
assign addr[24271]= 1630224009;
assign addr[24272]= 1415215352;
assign addr[24273]= 1171527280;
assign addr[24274]= 904098143;
assign addr[24275]= 618347408;
assign addr[24276]= 320065829;
assign addr[24277]= 15298099;
assign addr[24278]= -289779648;
assign addr[24279]= -588984994;
assign addr[24280]= -876254528;
assign addr[24281]= -1145766716;
assign addr[24282]= -1392059879;
assign addr[24283]= -1610142873;
assign addr[24284]= -1795596234;
assign addr[24285]= -1944661739;
assign addr[24286]= -2054318569;
assign addr[24287]= -2122344521;
assign addr[24288]= -2147361045;
assign addr[24289]= -2128861181;
assign addr[24290]= -2067219829;
assign addr[24291]= -1963686155;
assign addr[24292]= -1820358275;
assign addr[24293]= -1640140734;
assign addr[24294]= -1426685652;
assign addr[24295]= -1184318708;
assign addr[24296]= -917951481;
assign addr[24297]= -632981917;
assign addr[24298]= -335184940;
assign addr[24299]= -30595422;
assign addr[24300]= 274614114;
assign addr[24301]= 574258580;
assign addr[24302]= 862265664;
assign addr[24303]= 1132798888;
assign addr[24304]= 1380375881;
assign addr[24305]= 1599979481;
assign addr[24306]= 1787159411;
assign addr[24307]= 1938122457;
assign addr[24308]= 2049809346;
assign addr[24309]= 2119956737;
assign addr[24310]= 2147143090;
assign addr[24311]= 2130817471;
assign addr[24312]= 2071310720;
assign addr[24313]= 1969828744;
assign addr[24314]= 1828428082;
assign addr[24315]= 1649974225;
assign addr[24316]= 1438083551;
assign addr[24317]= 1197050035;
assign addr[24318]= 931758235;
assign addr[24319]= 647584304;
assign addr[24320]= 350287041;
assign addr[24321]= 45891193;
assign addr[24322]= -259434643;
assign addr[24323]= -559503022;
assign addr[24324]= -848233042;
assign addr[24325]= -1119773573;
assign addr[24326]= -1368621831;
assign addr[24327]= -1589734894;
assign addr[24328]= -1778631892;
assign addr[24329]= -1931484818;
assign addr[24330]= -2045196100;
assign addr[24331]= -2117461370;
assign addr[24332]= -2146816171;
assign addr[24333]= -2132665626;
assign addr[24334]= -2075296495;
assign addr[24335]= -1975871368;
assign addr[24336]= -1836405100;
assign addr[24337]= -1659723983;
assign addr[24338]= -1449408469;
assign addr[24339]= -1209720613;
assign addr[24340]= -945517704;
assign addr[24341]= -662153826;
assign addr[24342]= -365371365;
assign addr[24343]= -61184634;
assign addr[24344]= 244242007;
assign addr[24345]= 544719071;
assign addr[24346]= 834157373;
assign addr[24347]= 1106691431;
assign addr[24348]= 1356798326;
assign addr[24349]= 1579409630;
assign addr[24350]= 1770014111;
assign addr[24351]= 1924749160;
assign addr[24352]= 2040479063;
assign addr[24353]= 2114858546;
assign addr[24354]= 2146380306;
assign addr[24355]= 2134405552;
assign addr[24356]= 2079176953;
assign addr[24357]= 1981813720;
assign addr[24358]= 1844288924;
assign addr[24359]= 1669389513;
assign addr[24360]= 1460659832;
assign addr[24361]= 1222329801;
assign addr[24362]= 959229189;
assign addr[24363]= 676689746;
assign addr[24364]= 380437148;
assign addr[24365]= 76474970;
assign addr[24366]= -229036977;
assign addr[24367]= -529907477;
assign addr[24368]= -820039373;
assign addr[24369]= -1093553126;
assign addr[24370]= -1344905966;
assign addr[24371]= -1569004214;
assign addr[24372]= -1761306505;
assign addr[24373]= -1917915825;
assign addr[24374]= -2035658475;
assign addr[24375]= -2112148396;
assign addr[24376]= -2145835515;
assign addr[24377]= -2136037160;
assign addr[24378]= -2082951896;
assign addr[24379]= -1987655498;
assign addr[24380]= -1852079154;
assign addr[24381]= -1678970324;
assign addr[24382]= -1471837070;
assign addr[24383]= -1234876957;
assign addr[24384]= -972891995;
assign addr[24385]= -691191324;
assign addr[24386]= -395483624;
assign addr[24387]= -91761426;
assign addr[24388]= 213820322;
assign addr[24389]= 515068990;
assign addr[24390]= 805879757;
assign addr[24391]= 1080359326;
assign addr[24392]= 1332945355;
assign addr[24393]= 1558519173;
assign addr[24394]= 1752509516;
assign addr[24395]= 1910985158;
assign addr[24396]= 2030734582;
assign addr[24397]= 2109331059;
assign addr[24398]= 2145181827;
assign addr[24399]= 2137560369;
assign addr[24400]= 2086621133;
assign addr[24401]= 1993396407;
assign addr[24402]= 1859775393;
assign addr[24403]= 1688465931;
assign addr[24404]= 1482939614;
assign addr[24405]= 1247361445;
assign addr[24406]= 986505429;
assign addr[24407]= 705657826;
assign addr[24408]= 410510029;
assign addr[24409]= 107043224;
assign addr[24410]= -198592817;
assign addr[24411]= -500204365;
assign addr[24412]= -791679244;
assign addr[24413]= -1067110699;
assign addr[24414]= -1320917099;
assign addr[24415]= -1547955041;
assign addr[24416]= -1743623590;
assign addr[24417]= -1903957513;
assign addr[24418]= -2025707632;
assign addr[24419]= -2106406677;
assign addr[24420]= -2144419275;
assign addr[24421]= -2138975100;
assign addr[24422]= -2090184478;
assign addr[24423]= -1999036154;
assign addr[24424]= -1867377253;
assign addr[24425]= -1697875851;
assign addr[24426]= -1493966902;
assign addr[24427]= -1259782632;
assign addr[24428]= -1000068799;
assign addr[24429]= -720088517;
assign addr[24430]= -425515602;
assign addr[24431]= -122319591;
assign addr[24432]= 183355234;
assign addr[24433]= 485314355;
assign addr[24434]= 777438554;
assign addr[24435]= 1053807919;
assign addr[24436]= 1308821808;
assign addr[24437]= 1537312353;
assign addr[24438]= 1734649179;
assign addr[24439]= 1896833245;
assign addr[24440]= 2020577882;
assign addr[24441]= 2103375398;
assign addr[24442]= 2143547897;
assign addr[24443]= 2140281282;
assign addr[24444]= 2093641749;
assign addr[24445]= 2004574453;
assign addr[24446]= 1874884346;
assign addr[24447]= 1707199606;
assign addr[24448]= 1504918373;
assign addr[24449]= 1272139887;
assign addr[24450]= 1013581418;
assign addr[24451]= 734482665;
assign addr[24452]= 440499581;
assign addr[24453]= 137589750;
assign addr[24454]= -168108346;
assign addr[24455]= -470399716;
assign addr[24456]= -763158411;
assign addr[24457]= -1040451659;
assign addr[24458]= -1296660098;
assign addr[24459]= -1526591649;
assign addr[24460]= -1725586737;
assign addr[24461]= -1889612716;
assign addr[24462]= -2015345591;
assign addr[24463]= -2100237377;
assign addr[24464]= -2142567738;
assign addr[24465]= -2141478848;
assign addr[24466]= -2096992772;
assign addr[24467]= -2010011024;
assign addr[24468]= -1882296293;
assign addr[24469]= -1716436725;
assign addr[24470]= -1515793473;
assign addr[24471]= -1284432584;
assign addr[24472]= -1027042599;
assign addr[24473]= -748839539;
assign addr[24474]= -455461206;
assign addr[24475]= -152852926;
assign addr[24476]= 152852926;
assign addr[24477]= 455461206;
assign addr[24478]= 748839539;
assign addr[24479]= 1027042599;
assign addr[24480]= 1284432584;
assign addr[24481]= 1515793473;
assign addr[24482]= 1716436725;
assign addr[24483]= 1882296293;
assign addr[24484]= 2010011024;
assign addr[24485]= 2096992772;
assign addr[24486]= 2141478848;
assign addr[24487]= 2142567738;
assign addr[24488]= 2100237377;
assign addr[24489]= 2015345591;
assign addr[24490]= 1889612716;
assign addr[24491]= 1725586737;
assign addr[24492]= 1526591649;
assign addr[24493]= 1296660098;
assign addr[24494]= 1040451659;
assign addr[24495]= 763158411;
assign addr[24496]= 470399716;
assign addr[24497]= 168108346;
assign addr[24498]= -137589750;
assign addr[24499]= -440499581;
assign addr[24500]= -734482665;
assign addr[24501]= -1013581418;
assign addr[24502]= -1272139887;
assign addr[24503]= -1504918373;
assign addr[24504]= -1707199606;
assign addr[24505]= -1874884346;
assign addr[24506]= -2004574453;
assign addr[24507]= -2093641749;
assign addr[24508]= -2140281282;
assign addr[24509]= -2143547897;
assign addr[24510]= -2103375398;
assign addr[24511]= -2020577882;
assign addr[24512]= -1896833245;
assign addr[24513]= -1734649179;
assign addr[24514]= -1537312353;
assign addr[24515]= -1308821808;
assign addr[24516]= -1053807919;
assign addr[24517]= -777438554;
assign addr[24518]= -485314355;
assign addr[24519]= -183355234;
assign addr[24520]= 122319591;
assign addr[24521]= 425515602;
assign addr[24522]= 720088517;
assign addr[24523]= 1000068799;
assign addr[24524]= 1259782632;
assign addr[24525]= 1493966902;
assign addr[24526]= 1697875851;
assign addr[24527]= 1867377253;
assign addr[24528]= 1999036154;
assign addr[24529]= 2090184478;
assign addr[24530]= 2138975100;
assign addr[24531]= 2144419275;
assign addr[24532]= 2106406677;
assign addr[24533]= 2025707632;
assign addr[24534]= 1903957513;
assign addr[24535]= 1743623590;
assign addr[24536]= 1547955041;
assign addr[24537]= 1320917099;
assign addr[24538]= 1067110699;
assign addr[24539]= 791679244;
assign addr[24540]= 500204365;
assign addr[24541]= 198592817;
assign addr[24542]= -107043224;
assign addr[24543]= -410510029;
assign addr[24544]= -705657826;
assign addr[24545]= -986505429;
assign addr[24546]= -1247361445;
assign addr[24547]= -1482939614;
assign addr[24548]= -1688465931;
assign addr[24549]= -1859775393;
assign addr[24550]= -1993396407;
assign addr[24551]= -2086621133;
assign addr[24552]= -2137560369;
assign addr[24553]= -2145181827;
assign addr[24554]= -2109331059;
assign addr[24555]= -2030734582;
assign addr[24556]= -1910985158;
assign addr[24557]= -1752509516;
assign addr[24558]= -1558519173;
assign addr[24559]= -1332945355;
assign addr[24560]= -1080359326;
assign addr[24561]= -805879757;
assign addr[24562]= -515068990;
assign addr[24563]= -213820322;
assign addr[24564]= 91761426;
assign addr[24565]= 395483624;
assign addr[24566]= 691191324;
assign addr[24567]= 972891995;
assign addr[24568]= 1234876957;
assign addr[24569]= 1471837070;
assign addr[24570]= 1678970324;
assign addr[24571]= 1852079154;
assign addr[24572]= 1987655498;
assign addr[24573]= 2082951896;
assign addr[24574]= 2136037160;
assign addr[24575]= 2145835515;
assign addr[24576]= 2112148396;
assign addr[24577]= 2035658475;
assign addr[24578]= 1917915825;
assign addr[24579]= 1761306505;
assign addr[24580]= 1569004214;
assign addr[24581]= 1344905966;
assign addr[24582]= 1093553126;
assign addr[24583]= 820039373;
assign addr[24584]= 529907477;
assign addr[24585]= 229036977;
assign addr[24586]= -76474970;
assign addr[24587]= -380437148;
assign addr[24588]= -676689746;
assign addr[24589]= -959229189;
assign addr[24590]= -1222329801;
assign addr[24591]= -1460659832;
assign addr[24592]= -1669389513;
assign addr[24593]= -1844288924;
assign addr[24594]= -1981813720;
assign addr[24595]= -2079176953;
assign addr[24596]= -2134405552;
assign addr[24597]= -2146380306;
assign addr[24598]= -2114858546;
assign addr[24599]= -2040479063;
assign addr[24600]= -1924749160;
assign addr[24601]= -1770014111;
assign addr[24602]= -1579409630;
assign addr[24603]= -1356798326;
assign addr[24604]= -1106691431;
assign addr[24605]= -834157373;
assign addr[24606]= -544719071;
assign addr[24607]= -244242007;
assign addr[24608]= 61184634;
assign addr[24609]= 365371365;
assign addr[24610]= 662153826;
assign addr[24611]= 945517704;
assign addr[24612]= 1209720613;
assign addr[24613]= 1449408469;
assign addr[24614]= 1659723983;
assign addr[24615]= 1836405100;
assign addr[24616]= 1975871368;
assign addr[24617]= 2075296495;
assign addr[24618]= 2132665626;
assign addr[24619]= 2146816171;
assign addr[24620]= 2117461370;
assign addr[24621]= 2045196100;
assign addr[24622]= 1931484818;
assign addr[24623]= 1778631892;
assign addr[24624]= 1589734894;
assign addr[24625]= 1368621831;
assign addr[24626]= 1119773573;
assign addr[24627]= 848233042;
assign addr[24628]= 559503022;
assign addr[24629]= 259434643;
assign addr[24630]= -45891193;
assign addr[24631]= -350287041;
assign addr[24632]= -647584304;
assign addr[24633]= -931758235;
assign addr[24634]= -1197050035;
assign addr[24635]= -1438083551;
assign addr[24636]= -1649974225;
assign addr[24637]= -1828428082;
assign addr[24638]= -1969828744;
assign addr[24639]= -2071310720;
assign addr[24640]= -2130817471;
assign addr[24641]= -2147143090;
assign addr[24642]= -2119956737;
assign addr[24643]= -2049809346;
assign addr[24644]= -1938122457;
assign addr[24645]= -1787159411;
assign addr[24646]= -1599979481;
assign addr[24647]= -1380375881;
assign addr[24648]= -1132798888;
assign addr[24649]= -862265664;
assign addr[24650]= -574258580;
assign addr[24651]= -274614114;
assign addr[24652]= 30595422;
assign addr[24653]= 335184940;
assign addr[24654]= 632981917;
assign addr[24655]= 917951481;
assign addr[24656]= 1184318708;
assign addr[24657]= 1426685652;
assign addr[24658]= 1640140734;
assign addr[24659]= 1820358275;
assign addr[24660]= 1963686155;
assign addr[24661]= 2067219829;
assign addr[24662]= 2128861181;
assign addr[24663]= 2147361045;
assign addr[24664]= 2122344521;
assign addr[24665]= 2054318569;
assign addr[24666]= 1944661739;
assign addr[24667]= 1795596234;
assign addr[24668]= 1610142873;
assign addr[24669]= 1392059879;
assign addr[24670]= 1145766716;
assign addr[24671]= 876254528;
assign addr[24672]= 588984994;
assign addr[24673]= 289779648;
assign addr[24674]= -15298099;
assign addr[24675]= -320065829;
assign addr[24676]= -618347408;
assign addr[24677]= -904098143;
assign addr[24678]= -1171527280;
assign addr[24679]= -1415215352;
assign addr[24680]= -1630224009;
assign addr[24681]= -1812196087;
assign addr[24682]= -1957443913;
assign addr[24683]= -2063024031;
assign addr[24684]= -2126796855;
assign addr[24685]= -2147470025;
assign addr[24686]= -2124624598;
assign addr[24687]= -2058723538;
assign addr[24688]= -1951102334;
assign addr[24689]= -1803941934;
assign addr[24690]= -1620224553;
assign addr[24691]= -1403673233;
assign addr[24692]= -1158676398;
assign addr[24693]= -890198924;
assign addr[24694]= -603681519;
assign addr[24695]= -304930476;
assign addr[24696]= 0;
assign addr[24697]= 304930476;
assign addr[24698]= 603681519;
assign addr[24699]= 890198924;
assign addr[24700]= 1158676398;
assign addr[24701]= 1403673233;
assign addr[24702]= 1620224553;
assign addr[24703]= 1803941934;
assign addr[24704]= 1951102334;
assign addr[24705]= 2058723538;
assign addr[24706]= 2124624598;
assign addr[24707]= 2147470025;
assign addr[24708]= 2126796855;
assign addr[24709]= 2063024031;
assign addr[24710]= 1957443913;
assign addr[24711]= 1812196087;
assign addr[24712]= 1630224009;
assign addr[24713]= 1415215352;
assign addr[24714]= 1171527280;
assign addr[24715]= 904098143;
assign addr[24716]= 618347408;
assign addr[24717]= 320065829;
assign addr[24718]= 15298099;
assign addr[24719]= -289779648;
assign addr[24720]= -588984994;
assign addr[24721]= -876254528;
assign addr[24722]= -1145766716;
assign addr[24723]= -1392059879;
assign addr[24724]= -1610142873;
assign addr[24725]= -1795596234;
assign addr[24726]= -1944661739;
assign addr[24727]= -2054318569;
assign addr[24728]= -2122344521;
assign addr[24729]= -2147361045;
assign addr[24730]= -2128861181;
assign addr[24731]= -2067219829;
assign addr[24732]= -1963686155;
assign addr[24733]= -1820358275;
assign addr[24734]= -1640140734;
assign addr[24735]= -1426685652;
assign addr[24736]= -1184318708;
assign addr[24737]= -917951481;
assign addr[24738]= -632981917;
assign addr[24739]= -335184940;
assign addr[24740]= -30595422;
assign addr[24741]= 274614114;
assign addr[24742]= 574258580;
assign addr[24743]= 862265664;
assign addr[24744]= 1132798888;
assign addr[24745]= 1380375881;
assign addr[24746]= 1599979481;
assign addr[24747]= 1787159411;
assign addr[24748]= 1938122457;
assign addr[24749]= 2049809346;
assign addr[24750]= 2119956737;
assign addr[24751]= 2147143090;
assign addr[24752]= 2130817471;
assign addr[24753]= 2071310720;
assign addr[24754]= 1969828744;
assign addr[24755]= 1828428082;
assign addr[24756]= 1649974225;
assign addr[24757]= 1438083551;
assign addr[24758]= 1197050035;
assign addr[24759]= 931758235;
assign addr[24760]= 647584304;
assign addr[24761]= 350287041;
assign addr[24762]= 45891193;
assign addr[24763]= -259434643;
assign addr[24764]= -559503022;
assign addr[24765]= -848233042;
assign addr[24766]= -1119773573;
assign addr[24767]= -1368621831;
assign addr[24768]= -1589734894;
assign addr[24769]= -1778631892;
assign addr[24770]= -1931484818;
assign addr[24771]= -2045196100;
assign addr[24772]= -2117461370;
assign addr[24773]= -2146816171;
assign addr[24774]= -2132665626;
assign addr[24775]= -2075296495;
assign addr[24776]= -1975871368;
assign addr[24777]= -1836405100;
assign addr[24778]= -1659723983;
assign addr[24779]= -1449408469;
assign addr[24780]= -1209720613;
assign addr[24781]= -945517704;
assign addr[24782]= -662153826;
assign addr[24783]= -365371365;
assign addr[24784]= -61184634;
assign addr[24785]= 244242007;
assign addr[24786]= 544719071;
assign addr[24787]= 834157373;
assign addr[24788]= 1106691431;
assign addr[24789]= 1356798326;
assign addr[24790]= 1579409630;
assign addr[24791]= 1770014111;
assign addr[24792]= 1924749160;
assign addr[24793]= 2040479063;
assign addr[24794]= 2114858546;
assign addr[24795]= 2146380306;
assign addr[24796]= 2134405552;
assign addr[24797]= 2079176953;
assign addr[24798]= 1981813720;
assign addr[24799]= 1844288924;
assign addr[24800]= 1669389513;
assign addr[24801]= 1460659832;
assign addr[24802]= 1222329801;
assign addr[24803]= 959229189;
assign addr[24804]= 676689746;
assign addr[24805]= 380437148;
assign addr[24806]= 76474970;
assign addr[24807]= -229036977;
assign addr[24808]= -529907477;
assign addr[24809]= -820039373;
assign addr[24810]= -1093553126;
assign addr[24811]= -1344905966;
assign addr[24812]= -1569004214;
assign addr[24813]= -1761306505;
assign addr[24814]= -1917915825;
assign addr[24815]= -2035658475;
assign addr[24816]= -2112148396;
assign addr[24817]= -2145835515;
assign addr[24818]= -2136037160;
assign addr[24819]= -2082951896;
assign addr[24820]= -1987655498;
assign addr[24821]= -1852079154;
assign addr[24822]= -1678970324;
assign addr[24823]= -1471837070;
assign addr[24824]= -1234876957;
assign addr[24825]= -972891995;
assign addr[24826]= -691191324;
assign addr[24827]= -395483624;
assign addr[24828]= -91761426;
assign addr[24829]= 213820322;
assign addr[24830]= 515068990;
assign addr[24831]= 805879757;
assign addr[24832]= 1080359326;
assign addr[24833]= 1332945355;
assign addr[24834]= 1558519173;
assign addr[24835]= 1752509516;
assign addr[24836]= 1910985158;
assign addr[24837]= 2030734582;
assign addr[24838]= 2109331059;
assign addr[24839]= 2145181827;
assign addr[24840]= 2137560369;
assign addr[24841]= 2086621133;
assign addr[24842]= 1993396407;
assign addr[24843]= 1859775393;
assign addr[24844]= 1688465931;
assign addr[24845]= 1482939614;
assign addr[24846]= 1247361445;
assign addr[24847]= 986505429;
assign addr[24848]= 705657826;
assign addr[24849]= 410510029;
assign addr[24850]= 107043224;
assign addr[24851]= -198592817;
assign addr[24852]= -500204365;
assign addr[24853]= -791679244;
assign addr[24854]= -1067110699;
assign addr[24855]= -1320917099;
assign addr[24856]= -1547955041;
assign addr[24857]= -1743623590;
assign addr[24858]= -1903957513;
assign addr[24859]= -2025707632;
assign addr[24860]= -2106406677;
assign addr[24861]= -2144419275;
assign addr[24862]= -2138975100;
assign addr[24863]= -2090184478;
assign addr[24864]= -1999036154;
assign addr[24865]= -1867377253;
assign addr[24866]= -1697875851;
assign addr[24867]= -1493966902;
assign addr[24868]= -1259782632;
assign addr[24869]= -1000068799;
assign addr[24870]= -720088517;
assign addr[24871]= -425515602;
assign addr[24872]= -122319591;
assign addr[24873]= 183355234;
assign addr[24874]= 485314355;
assign addr[24875]= 777438554;
assign addr[24876]= 1053807919;
assign addr[24877]= 1308821808;
assign addr[24878]= 1537312353;
assign addr[24879]= 1734649179;
assign addr[24880]= 1896833245;
assign addr[24881]= 2020577882;
assign addr[24882]= 2103375398;
assign addr[24883]= 2143547897;
assign addr[24884]= 2140281282;
assign addr[24885]= 2093641749;
assign addr[24886]= 2004574453;
assign addr[24887]= 1874884346;
assign addr[24888]= 1707199606;
assign addr[24889]= 1504918373;
assign addr[24890]= 1272139887;
assign addr[24891]= 1013581418;
assign addr[24892]= 734482665;
assign addr[24893]= 440499581;
assign addr[24894]= 137589750;
assign addr[24895]= -168108346;
assign addr[24896]= -470399716;
assign addr[24897]= -763158411;
assign addr[24898]= -1040451659;
assign addr[24899]= -1296660098;
assign addr[24900]= -1526591649;
assign addr[24901]= -1725586737;
assign addr[24902]= -1889612716;
assign addr[24903]= -2015345591;
assign addr[24904]= -2100237377;
assign addr[24905]= -2142567738;
assign addr[24906]= -2141478848;
assign addr[24907]= -2096992772;
assign addr[24908]= -2010011024;
assign addr[24909]= -1882296293;
assign addr[24910]= -1716436725;
assign addr[24911]= -1515793473;
assign addr[24912]= -1284432584;
assign addr[24913]= -1027042599;
assign addr[24914]= -748839539;
assign addr[24915]= -455461206;
assign addr[24916]= -152852926;
assign addr[24917]= 152852926;
assign addr[24918]= 455461206;
assign addr[24919]= 748839539;
assign addr[24920]= 1027042599;
assign addr[24921]= 1284432584;
assign addr[24922]= 1515793473;
assign addr[24923]= 1716436725;
assign addr[24924]= 1882296293;
assign addr[24925]= 2010011024;
assign addr[24926]= 2096992772;
assign addr[24927]= 2141478848;
assign addr[24928]= 2142567738;
assign addr[24929]= 2100237377;
assign addr[24930]= 2015345591;
assign addr[24931]= 1889612716;
assign addr[24932]= 1725586737;
assign addr[24933]= 1526591649;
assign addr[24934]= 1296660098;
assign addr[24935]= 1040451659;
assign addr[24936]= 763158411;
assign addr[24937]= 470399716;
assign addr[24938]= 168108346;
assign addr[24939]= -137589750;
assign addr[24940]= -440499581;
assign addr[24941]= -734482665;
assign addr[24942]= -1013581418;
assign addr[24943]= -1272139887;
assign addr[24944]= -1504918373;
assign addr[24945]= -1707199606;
assign addr[24946]= -1874884346;
assign addr[24947]= -2004574453;
assign addr[24948]= -2093641749;
assign addr[24949]= -2140281282;
assign addr[24950]= -2143547897;
assign addr[24951]= -2103375398;
assign addr[24952]= -2020577882;
assign addr[24953]= -1896833245;
assign addr[24954]= -1734649179;
assign addr[24955]= -1537312353;
assign addr[24956]= -1308821808;
assign addr[24957]= -1053807919;
assign addr[24958]= -777438554;
assign addr[24959]= -485314355;
assign addr[24960]= -183355234;
assign addr[24961]= 122319591;
assign addr[24962]= 425515602;
assign addr[24963]= 720088517;
assign addr[24964]= 1000068799;
assign addr[24965]= 1259782632;
assign addr[24966]= 1493966902;
assign addr[24967]= 1697875851;
assign addr[24968]= 1867377253;
assign addr[24969]= 1999036154;
assign addr[24970]= 2090184478;
assign addr[24971]= 2138975100;
assign addr[24972]= 2144419275;
assign addr[24973]= 2106406677;
assign addr[24974]= 2025707632;
assign addr[24975]= 1903957513;
assign addr[24976]= 1743623590;
assign addr[24977]= 1547955041;
assign addr[24978]= 1320917099;
assign addr[24979]= 1067110699;
assign addr[24980]= 791679244;
assign addr[24981]= 500204365;
assign addr[24982]= 198592817;
assign addr[24983]= -107043224;
assign addr[24984]= -410510029;
assign addr[24985]= -705657826;
assign addr[24986]= -986505429;
assign addr[24987]= -1247361445;
assign addr[24988]= -1482939614;
assign addr[24989]= -1688465931;
assign addr[24990]= -1859775393;
assign addr[24991]= -1993396407;
assign addr[24992]= -2086621133;
assign addr[24993]= -2137560369;
assign addr[24994]= -2145181827;
assign addr[24995]= -2109331059;
assign addr[24996]= -2030734582;
assign addr[24997]= -1910985158;
assign addr[24998]= -1752509516;
assign addr[24999]= -1558519173;
assign addr[25000]= -1332945355;
assign addr[25001]= -1080359326;
assign addr[25002]= -805879757;
assign addr[25003]= -515068990;
assign addr[25004]= -213820322;
assign addr[25005]= 91761426;
assign addr[25006]= 395483624;
assign addr[25007]= 691191324;
assign addr[25008]= 972891995;
assign addr[25009]= 1234876957;
assign addr[25010]= 1471837070;
assign addr[25011]= 1678970324;
assign addr[25012]= 1852079154;
assign addr[25013]= 1987655498;
assign addr[25014]= 2082951896;
assign addr[25015]= 2136037160;
assign addr[25016]= 2145835515;
assign addr[25017]= 2112148396;
assign addr[25018]= 2035658475;
assign addr[25019]= 1917915825;
assign addr[25020]= 1761306505;
assign addr[25021]= 1569004214;
assign addr[25022]= 1344905966;
assign addr[25023]= 1093553126;
assign addr[25024]= 820039373;
assign addr[25025]= 529907477;
assign addr[25026]= 229036977;
assign addr[25027]= -76474970;
assign addr[25028]= -380437148;
assign addr[25029]= -676689746;
assign addr[25030]= -959229189;
assign addr[25031]= -1222329801;
assign addr[25032]= -1460659832;
assign addr[25033]= -1669389513;
assign addr[25034]= -1844288924;
assign addr[25035]= -1981813720;
assign addr[25036]= -2079176953;
assign addr[25037]= -2134405552;
assign addr[25038]= -2146380306;
assign addr[25039]= -2114858546;
assign addr[25040]= -2040479063;
assign addr[25041]= -1924749160;
assign addr[25042]= -1770014111;
assign addr[25043]= -1579409630;
assign addr[25044]= -1356798326;
assign addr[25045]= -1106691431;
assign addr[25046]= -834157373;
assign addr[25047]= -544719071;
assign addr[25048]= -244242007;
assign addr[25049]= 61184634;
assign addr[25050]= 365371365;
assign addr[25051]= 662153826;
assign addr[25052]= 945517704;
assign addr[25053]= 1209720613;
assign addr[25054]= 1449408469;
assign addr[25055]= 1659723983;
assign addr[25056]= 1836405100;
assign addr[25057]= 1975871368;
assign addr[25058]= 2075296495;
assign addr[25059]= 2132665626;
assign addr[25060]= 2146816171;
assign addr[25061]= 2117461370;
assign addr[25062]= 2045196100;
assign addr[25063]= 1931484818;
assign addr[25064]= 1778631892;
assign addr[25065]= 1589734894;
assign addr[25066]= 1368621831;
assign addr[25067]= 1119773573;
assign addr[25068]= 848233042;
assign addr[25069]= 559503022;
assign addr[25070]= 259434643;
assign addr[25071]= -45891193;
assign addr[25072]= -350287041;
assign addr[25073]= -647584304;
assign addr[25074]= -931758235;
assign addr[25075]= -1197050035;
assign addr[25076]= -1438083551;
assign addr[25077]= -1649974225;
assign addr[25078]= -1828428082;
assign addr[25079]= -1969828744;
assign addr[25080]= -2071310720;
assign addr[25081]= -2130817471;
assign addr[25082]= -2147143090;
assign addr[25083]= -2119956737;
assign addr[25084]= -2049809346;
assign addr[25085]= -1938122457;
assign addr[25086]= -1787159411;
assign addr[25087]= -1599979481;
assign addr[25088]= -1380375881;
assign addr[25089]= -1132798888;
assign addr[25090]= -862265664;
assign addr[25091]= -574258580;
assign addr[25092]= -274614114;
assign addr[25093]= 30595422;
assign addr[25094]= 335184940;
assign addr[25095]= 632981917;
assign addr[25096]= 917951481;
assign addr[25097]= 1184318708;
assign addr[25098]= 1426685652;
assign addr[25099]= 1640140734;
assign addr[25100]= 1820358275;
assign addr[25101]= 1963686155;
assign addr[25102]= 2067219829;
assign addr[25103]= 2128861181;
assign addr[25104]= 2147361045;
assign addr[25105]= 2122344521;
assign addr[25106]= 2054318569;
assign addr[25107]= 1944661739;
assign addr[25108]= 1795596234;
assign addr[25109]= 1610142873;
assign addr[25110]= 1392059879;
assign addr[25111]= 1145766716;
assign addr[25112]= 876254528;
assign addr[25113]= 588984994;
assign addr[25114]= 289779648;
assign addr[25115]= -15298099;
assign addr[25116]= -320065829;
assign addr[25117]= -618347408;
assign addr[25118]= -904098143;
assign addr[25119]= -1171527280;
assign addr[25120]= -1415215352;
assign addr[25121]= -1630224009;
assign addr[25122]= -1812196087;
assign addr[25123]= -1957443913;
assign addr[25124]= -2063024031;
assign addr[25125]= -2126796855;
assign addr[25126]= -2147470025;
assign addr[25127]= -2124624598;
assign addr[25128]= -2058723538;
assign addr[25129]= -1951102334;
assign addr[25130]= -1803941934;
assign addr[25131]= -1620224553;
assign addr[25132]= -1403673233;
assign addr[25133]= -1158676398;
assign addr[25134]= -890198924;
assign addr[25135]= -603681519;
assign addr[25136]= -304930476;
assign addr[25137]= 0;
assign addr[25138]= 304930476;
assign addr[25139]= 603681519;
assign addr[25140]= 890198924;
assign addr[25141]= 1158676398;
assign addr[25142]= 1403673233;
assign addr[25143]= 1620224553;
assign addr[25144]= 1803941934;
assign addr[25145]= 1951102334;
assign addr[25146]= 2058723538;
assign addr[25147]= 2124624598;
assign addr[25148]= 2147470025;
assign addr[25149]= 2126796855;
assign addr[25150]= 2063024031;
assign addr[25151]= 1957443913;
assign addr[25152]= 1812196087;
assign addr[25153]= 1630224009;
assign addr[25154]= 1415215352;
assign addr[25155]= 1171527280;
assign addr[25156]= 904098143;
assign addr[25157]= 618347408;
assign addr[25158]= 320065829;
assign addr[25159]= 15298099;
assign addr[25160]= -289779648;
assign addr[25161]= -588984994;
assign addr[25162]= -876254528;
assign addr[25163]= -1145766716;
assign addr[25164]= -1392059879;
assign addr[25165]= -1610142873;
assign addr[25166]= -1795596234;
assign addr[25167]= -1944661739;
assign addr[25168]= -2054318569;
assign addr[25169]= -2122344521;
assign addr[25170]= -2147361045;
assign addr[25171]= -2128861181;
assign addr[25172]= -2067219829;
assign addr[25173]= -1963686155;
assign addr[25174]= -1820358275;
assign addr[25175]= -1640140734;
assign addr[25176]= -1426685652;
assign addr[25177]= -1184318708;
assign addr[25178]= -917951481;
assign addr[25179]= -632981917;
assign addr[25180]= -335184940;
assign addr[25181]= -30595422;
assign addr[25182]= 274614114;
assign addr[25183]= 574258580;
assign addr[25184]= 862265664;
assign addr[25185]= 1132798888;
assign addr[25186]= 1380375881;
assign addr[25187]= 1599979481;
assign addr[25188]= 1787159411;
assign addr[25189]= 1938122457;
assign addr[25190]= 2049809346;
assign addr[25191]= 2119956737;
assign addr[25192]= 2147143090;
assign addr[25193]= 2130817471;
assign addr[25194]= 2071310720;
assign addr[25195]= 1969828744;
assign addr[25196]= 1828428082;
assign addr[25197]= 1649974225;
assign addr[25198]= 1438083551;
assign addr[25199]= 1197050035;
assign addr[25200]= 931758235;
assign addr[25201]= 647584304;
assign addr[25202]= 350287041;
assign addr[25203]= 45891193;
assign addr[25204]= -259434643;
assign addr[25205]= -559503022;
assign addr[25206]= -848233042;
assign addr[25207]= -1119773573;
assign addr[25208]= -1368621831;
assign addr[25209]= -1589734894;
assign addr[25210]= -1778631892;
assign addr[25211]= -1931484818;
assign addr[25212]= -2045196100;
assign addr[25213]= -2117461370;
assign addr[25214]= -2146816171;
assign addr[25215]= -2132665626;
assign addr[25216]= -2075296495;
assign addr[25217]= -1975871368;
assign addr[25218]= -1836405100;
assign addr[25219]= -1659723983;
assign addr[25220]= -1449408469;
assign addr[25221]= -1209720613;
assign addr[25222]= -945517704;
assign addr[25223]= -662153826;
assign addr[25224]= -365371365;
assign addr[25225]= -61184634;
assign addr[25226]= 244242007;
assign addr[25227]= 544719071;
assign addr[25228]= 834157373;
assign addr[25229]= 1106691431;
assign addr[25230]= 1356798326;
assign addr[25231]= 1579409630;
assign addr[25232]= 1770014111;
assign addr[25233]= 1924749160;
assign addr[25234]= 2040479063;
assign addr[25235]= 2114858546;
assign addr[25236]= 2146380306;
assign addr[25237]= 2134405552;
assign addr[25238]= 2079176953;
assign addr[25239]= 1981813720;
assign addr[25240]= 1844288924;
assign addr[25241]= 1669389513;
assign addr[25242]= 1460659832;
assign addr[25243]= 1222329801;
assign addr[25244]= 959229189;
assign addr[25245]= 676689746;
assign addr[25246]= 380437148;
assign addr[25247]= 76474970;
assign addr[25248]= -229036977;
assign addr[25249]= -529907477;
assign addr[25250]= -820039373;
assign addr[25251]= -1093553126;
assign addr[25252]= -1344905966;
assign addr[25253]= -1569004214;
assign addr[25254]= -1761306505;
assign addr[25255]= -1917915825;
assign addr[25256]= -2035658475;
assign addr[25257]= -2112148396;
assign addr[25258]= -2145835515;
assign addr[25259]= -2136037160;
assign addr[25260]= -2082951896;
assign addr[25261]= -1987655498;
assign addr[25262]= -1852079154;
assign addr[25263]= -1678970324;
assign addr[25264]= -1471837070;
assign addr[25265]= -1234876957;
assign addr[25266]= -972891995;
assign addr[25267]= -691191324;
assign addr[25268]= -395483624;
assign addr[25269]= -91761426;
assign addr[25270]= 213820322;
assign addr[25271]= 515068990;
assign addr[25272]= 805879757;
assign addr[25273]= 1080359326;
assign addr[25274]= 1332945355;
assign addr[25275]= 1558519173;
assign addr[25276]= 1752509516;
assign addr[25277]= 1910985158;
assign addr[25278]= 2030734582;
assign addr[25279]= 2109331059;
assign addr[25280]= 2145181827;
assign addr[25281]= 2137560369;
assign addr[25282]= 2086621133;
assign addr[25283]= 1993396407;
assign addr[25284]= 1859775393;
assign addr[25285]= 1688465931;
assign addr[25286]= 1482939614;
assign addr[25287]= 1247361445;
assign addr[25288]= 986505429;
assign addr[25289]= 705657826;
assign addr[25290]= 410510029;
assign addr[25291]= 107043224;
assign addr[25292]= -198592817;
assign addr[25293]= -500204365;
assign addr[25294]= -791679244;
assign addr[25295]= -1067110699;
assign addr[25296]= -1320917099;
assign addr[25297]= -1547955041;
assign addr[25298]= -1743623590;
assign addr[25299]= -1903957513;
assign addr[25300]= -2025707632;
assign addr[25301]= -2106406677;
assign addr[25302]= -2144419275;
assign addr[25303]= -2138975100;
assign addr[25304]= -2090184478;
assign addr[25305]= -1999036154;
assign addr[25306]= -1867377253;
assign addr[25307]= -1697875851;
assign addr[25308]= -1493966902;
assign addr[25309]= -1259782632;
assign addr[25310]= -1000068799;
assign addr[25311]= -720088517;
assign addr[25312]= -425515602;
assign addr[25313]= -122319591;
assign addr[25314]= 183355234;
assign addr[25315]= 485314355;
assign addr[25316]= 777438554;
assign addr[25317]= 1053807919;
assign addr[25318]= 1308821808;
assign addr[25319]= 1537312353;
assign addr[25320]= 1734649179;
assign addr[25321]= 1896833245;
assign addr[25322]= 2020577882;
assign addr[25323]= 2103375398;
assign addr[25324]= 2143547897;
assign addr[25325]= 2140281282;
assign addr[25326]= 2093641749;
assign addr[25327]= 2004574453;
assign addr[25328]= 1874884346;
assign addr[25329]= 1707199606;
assign addr[25330]= 1504918373;
assign addr[25331]= 1272139887;
assign addr[25332]= 1013581418;
assign addr[25333]= 734482665;
assign addr[25334]= 440499581;
assign addr[25335]= 137589750;
assign addr[25336]= -168108346;
assign addr[25337]= -470399716;
assign addr[25338]= -763158411;
assign addr[25339]= -1040451659;
assign addr[25340]= -1296660098;
assign addr[25341]= -1526591649;
assign addr[25342]= -1725586737;
assign addr[25343]= -1889612716;
assign addr[25344]= -2015345591;
assign addr[25345]= -2100237377;
assign addr[25346]= -2142567738;
assign addr[25347]= -2141478848;
assign addr[25348]= -2096992772;
assign addr[25349]= -2010011024;
assign addr[25350]= -1882296293;
assign addr[25351]= -1716436725;
assign addr[25352]= -1515793473;
assign addr[25353]= -1284432584;
assign addr[25354]= -1027042599;
assign addr[25355]= -748839539;
assign addr[25356]= -455461206;
assign addr[25357]= -152852926;
assign addr[25358]= 152852926;
assign addr[25359]= 455461206;
assign addr[25360]= 748839539;
assign addr[25361]= 1027042599;
assign addr[25362]= 1284432584;
assign addr[25363]= 1515793473;
assign addr[25364]= 1716436725;
assign addr[25365]= 1882296293;
assign addr[25366]= 2010011024;
assign addr[25367]= 2096992772;
assign addr[25368]= 2141478848;
assign addr[25369]= 2142567738;
assign addr[25370]= 2100237377;
assign addr[25371]= 2015345591;
assign addr[25372]= 1889612716;
assign addr[25373]= 1725586737;
assign addr[25374]= 1526591649;
assign addr[25375]= 1296660098;
assign addr[25376]= 1040451659;
assign addr[25377]= 763158411;
assign addr[25378]= 470399716;
assign addr[25379]= 168108346;
assign addr[25380]= -137589750;
assign addr[25381]= -440499581;
assign addr[25382]= -734482665;
assign addr[25383]= -1013581418;
assign addr[25384]= -1272139887;
assign addr[25385]= -1504918373;
assign addr[25386]= -1707199606;
assign addr[25387]= -1874884346;
assign addr[25388]= -2004574453;
assign addr[25389]= -2093641749;
assign addr[25390]= -2140281282;
assign addr[25391]= -2143547897;
assign addr[25392]= -2103375398;
assign addr[25393]= -2020577882;
assign addr[25394]= -1896833245;
assign addr[25395]= -1734649179;
assign addr[25396]= -1537312353;
assign addr[25397]= -1308821808;
assign addr[25398]= -1053807919;
assign addr[25399]= -777438554;
assign addr[25400]= -485314355;
assign addr[25401]= -183355234;
assign addr[25402]= 122319591;
assign addr[25403]= 425515602;
assign addr[25404]= 720088517;
assign addr[25405]= 1000068799;
assign addr[25406]= 1259782632;
assign addr[25407]= 1493966902;
assign addr[25408]= 1697875851;
assign addr[25409]= 1867377253;
assign addr[25410]= 1999036154;
assign addr[25411]= 2090184478;
assign addr[25412]= 2138975100;
assign addr[25413]= 2144419275;
assign addr[25414]= 2106406677;
assign addr[25415]= 2025707632;
assign addr[25416]= 1903957513;
assign addr[25417]= 1743623590;
assign addr[25418]= 1547955041;
assign addr[25419]= 1320917099;
assign addr[25420]= 1067110699;
assign addr[25421]= 791679244;
assign addr[25422]= 500204365;
assign addr[25423]= 198592817;
assign addr[25424]= -107043224;
assign addr[25425]= -410510029;
assign addr[25426]= -705657826;
assign addr[25427]= -986505429;
assign addr[25428]= -1247361445;
assign addr[25429]= -1482939614;
assign addr[25430]= -1688465931;
assign addr[25431]= -1859775393;
assign addr[25432]= -1993396407;
assign addr[25433]= -2086621133;
assign addr[25434]= -2137560369;
assign addr[25435]= -2145181827;
assign addr[25436]= -2109331059;
assign addr[25437]= -2030734582;
assign addr[25438]= -1910985158;
assign addr[25439]= -1752509516;
assign addr[25440]= -1558519173;
assign addr[25441]= -1332945355;
assign addr[25442]= -1080359326;
assign addr[25443]= -805879757;
assign addr[25444]= -515068990;
assign addr[25445]= -213820322;
assign addr[25446]= 91761426;
assign addr[25447]= 395483624;
assign addr[25448]= 691191324;
assign addr[25449]= 972891995;
assign addr[25450]= 1234876957;
assign addr[25451]= 1471837070;
assign addr[25452]= 1678970324;
assign addr[25453]= 1852079154;
assign addr[25454]= 1987655498;
assign addr[25455]= 2082951896;
assign addr[25456]= 2136037160;
assign addr[25457]= 2145835515;
assign addr[25458]= 2112148396;
assign addr[25459]= 2035658475;
assign addr[25460]= 1917915825;
assign addr[25461]= 1761306505;
assign addr[25462]= 1569004214;
assign addr[25463]= 1344905966;
assign addr[25464]= 1093553126;
assign addr[25465]= 820039373;
assign addr[25466]= 529907477;
assign addr[25467]= 229036977;
assign addr[25468]= -76474970;
assign addr[25469]= -380437148;
assign addr[25470]= -676689746;
assign addr[25471]= -959229189;
assign addr[25472]= -1222329801;
assign addr[25473]= -1460659832;
assign addr[25474]= -1669389513;
assign addr[25475]= -1844288924;
assign addr[25476]= -1981813720;
assign addr[25477]= -2079176953;
assign addr[25478]= -2134405552;
assign addr[25479]= -2146380306;
assign addr[25480]= -2114858546;
assign addr[25481]= -2040479063;
assign addr[25482]= -1924749160;
assign addr[25483]= -1770014111;
assign addr[25484]= -1579409630;
assign addr[25485]= -1356798326;
assign addr[25486]= -1106691431;
assign addr[25487]= -834157373;
assign addr[25488]= -544719071;
assign addr[25489]= -244242007;
assign addr[25490]= 61184634;
assign addr[25491]= 365371365;
assign addr[25492]= 662153826;
assign addr[25493]= 945517704;
assign addr[25494]= 1209720613;
assign addr[25495]= 1449408469;
assign addr[25496]= 1659723983;
assign addr[25497]= 1836405100;
assign addr[25498]= 1975871368;
assign addr[25499]= 2075296495;
assign addr[25500]= 2132665626;
assign addr[25501]= 2146816171;
assign addr[25502]= 2117461370;
assign addr[25503]= 2045196100;
assign addr[25504]= 1931484818;
assign addr[25505]= 1778631892;
assign addr[25506]= 1589734894;
assign addr[25507]= 1368621831;
assign addr[25508]= 1119773573;
assign addr[25509]= 848233042;
assign addr[25510]= 559503022;
assign addr[25511]= 259434643;
assign addr[25512]= -45891193;
assign addr[25513]= -350287041;
assign addr[25514]= -647584304;
assign addr[25515]= -931758235;
assign addr[25516]= -1197050035;
assign addr[25517]= -1438083551;
assign addr[25518]= -1649974225;
assign addr[25519]= -1828428082;
assign addr[25520]= -1969828744;
assign addr[25521]= -2071310720;
assign addr[25522]= -2130817471;
assign addr[25523]= -2147143090;
assign addr[25524]= -2119956737;
assign addr[25525]= -2049809346;
assign addr[25526]= -1938122457;
assign addr[25527]= -1787159411;
assign addr[25528]= -1599979481;
assign addr[25529]= -1380375881;
assign addr[25530]= -1132798888;
assign addr[25531]= -862265664;
assign addr[25532]= -574258580;
assign addr[25533]= -274614114;
assign addr[25534]= 30595422;
assign addr[25535]= 335184940;
assign addr[25536]= 632981917;
assign addr[25537]= 917951481;
assign addr[25538]= 1184318708;
assign addr[25539]= 1426685652;
assign addr[25540]= 1640140734;
assign addr[25541]= 1820358275;
assign addr[25542]= 1963686155;
assign addr[25543]= 2067219829;
assign addr[25544]= 2128861181;
assign addr[25545]= 2147361045;
assign addr[25546]= 2122344521;
assign addr[25547]= 2054318569;
assign addr[25548]= 1944661739;
assign addr[25549]= 1795596234;
assign addr[25550]= 1610142873;
assign addr[25551]= 1392059879;
assign addr[25552]= 1145766716;
assign addr[25553]= 876254528;
assign addr[25554]= 588984994;
assign addr[25555]= 289779648;
assign addr[25556]= -15298099;
assign addr[25557]= -320065829;
assign addr[25558]= -618347408;
assign addr[25559]= -904098143;
assign addr[25560]= -1171527280;
assign addr[25561]= -1415215352;
assign addr[25562]= -1630224009;
assign addr[25563]= -1812196087;
assign addr[25564]= -1957443913;
assign addr[25565]= -2063024031;
assign addr[25566]= -2126796855;
assign addr[25567]= -2147470025;
assign addr[25568]= -2124624598;
assign addr[25569]= -2058723538;
assign addr[25570]= -1951102334;
assign addr[25571]= -1803941934;
assign addr[25572]= -1620224553;
assign addr[25573]= -1403673233;
assign addr[25574]= -1158676398;
assign addr[25575]= -890198924;
assign addr[25576]= -603681519;
assign addr[25577]= -304930476;
assign addr[25578]= 0;
assign addr[25579]= 304930476;
assign addr[25580]= 603681519;
assign addr[25581]= 890198924;
assign addr[25582]= 1158676398;
assign addr[25583]= 1403673233;
assign addr[25584]= 1620224553;
assign addr[25585]= 1803941934;
assign addr[25586]= 1951102334;
assign addr[25587]= 2058723538;
assign addr[25588]= 2124624598;
assign addr[25589]= 2147470025;
assign addr[25590]= 2126796855;
assign addr[25591]= 2063024031;
assign addr[25592]= 1957443913;
assign addr[25593]= 1812196087;
assign addr[25594]= 1630224009;
assign addr[25595]= 1415215352;
assign addr[25596]= 1171527280;
assign addr[25597]= 904098143;
assign addr[25598]= 618347408;
assign addr[25599]= 320065829;
assign addr[25600]= 15298099;
assign addr[25601]= -289779648;
assign addr[25602]= -588984994;
assign addr[25603]= -876254528;
assign addr[25604]= -1145766716;
assign addr[25605]= -1392059879;
assign addr[25606]= -1610142873;
assign addr[25607]= -1795596234;
assign addr[25608]= -1944661739;
assign addr[25609]= -2054318569;
assign addr[25610]= -2122344521;
assign addr[25611]= -2147361045;
assign addr[25612]= -2128861181;
assign addr[25613]= -2067219829;
assign addr[25614]= -1963686155;
assign addr[25615]= -1820358275;
assign addr[25616]= -1640140734;
assign addr[25617]= -1426685652;
assign addr[25618]= -1184318708;
assign addr[25619]= -917951481;
assign addr[25620]= -632981917;
assign addr[25621]= -335184940;
assign addr[25622]= -30595422;
assign addr[25623]= 274614114;
assign addr[25624]= 574258580;
assign addr[25625]= 862265664;
assign addr[25626]= 1132798888;
assign addr[25627]= 1380375881;
assign addr[25628]= 1599979481;
assign addr[25629]= 1787159411;
assign addr[25630]= 1938122457;
assign addr[25631]= 2049809346;
assign addr[25632]= 2119956737;
assign addr[25633]= 2147143090;
assign addr[25634]= 2130817471;
assign addr[25635]= 2071310720;
assign addr[25636]= 1969828744;
assign addr[25637]= 1828428082;
assign addr[25638]= 1649974225;
assign addr[25639]= 1438083551;
assign addr[25640]= 1197050035;
assign addr[25641]= 931758235;
assign addr[25642]= 647584304;
assign addr[25643]= 350287041;
assign addr[25644]= 45891193;
assign addr[25645]= -259434643;
assign addr[25646]= -559503022;
assign addr[25647]= -848233042;
assign addr[25648]= -1119773573;
assign addr[25649]= -1368621831;
assign addr[25650]= -1589734894;
assign addr[25651]= -1778631892;
assign addr[25652]= -1931484818;
assign addr[25653]= -2045196100;
assign addr[25654]= -2117461370;
assign addr[25655]= -2146816171;
assign addr[25656]= -2132665626;
assign addr[25657]= -2075296495;
assign addr[25658]= -1975871368;
assign addr[25659]= -1836405100;
assign addr[25660]= -1659723983;
assign addr[25661]= -1449408469;
assign addr[25662]= -1209720613;
assign addr[25663]= -945517704;
assign addr[25664]= -662153826;
assign addr[25665]= -365371365;
assign addr[25666]= -61184634;
assign addr[25667]= 244242007;
assign addr[25668]= 544719071;
assign addr[25669]= 834157373;
assign addr[25670]= 1106691431;
assign addr[25671]= 1356798326;
assign addr[25672]= 1579409630;
assign addr[25673]= 1770014111;
assign addr[25674]= 1924749160;
assign addr[25675]= 2040479063;
assign addr[25676]= 2114858546;
assign addr[25677]= 2146380306;
assign addr[25678]= 2134405552;
assign addr[25679]= 2079176953;
assign addr[25680]= 1981813720;
assign addr[25681]= 1844288924;
assign addr[25682]= 1669389513;
assign addr[25683]= 1460659832;
assign addr[25684]= 1222329801;
assign addr[25685]= 959229189;
assign addr[25686]= 676689746;
assign addr[25687]= 380437148;
assign addr[25688]= 76474970;
assign addr[25689]= -229036977;
assign addr[25690]= -529907477;
assign addr[25691]= -820039373;
assign addr[25692]= -1093553126;
assign addr[25693]= -1344905966;
assign addr[25694]= -1569004214;
assign addr[25695]= -1761306505;
assign addr[25696]= -1917915825;
assign addr[25697]= -2035658475;
assign addr[25698]= -2112148396;
assign addr[25699]= -2145835515;
assign addr[25700]= -2136037160;
assign addr[25701]= -2082951896;
assign addr[25702]= -1987655498;
assign addr[25703]= -1852079154;
assign addr[25704]= -1678970324;
assign addr[25705]= -1471837070;
assign addr[25706]= -1234876957;
assign addr[25707]= -972891995;
assign addr[25708]= -691191324;
assign addr[25709]= -395483624;
assign addr[25710]= -91761426;
assign addr[25711]= 213820322;
assign addr[25712]= 515068990;
assign addr[25713]= 805879757;
assign addr[25714]= 1080359326;
assign addr[25715]= 1332945355;
assign addr[25716]= 1558519173;
assign addr[25717]= 1752509516;
assign addr[25718]= 1910985158;
assign addr[25719]= 2030734582;
assign addr[25720]= 2109331059;
assign addr[25721]= 2145181827;
assign addr[25722]= 2137560369;
assign addr[25723]= 2086621133;
assign addr[25724]= 1993396407;
assign addr[25725]= 1859775393;
assign addr[25726]= 1688465931;
assign addr[25727]= 1482939614;
assign addr[25728]= 1247361445;
assign addr[25729]= 986505429;
assign addr[25730]= 705657826;
assign addr[25731]= 410510029;
assign addr[25732]= 107043224;
assign addr[25733]= -198592817;
assign addr[25734]= -500204365;
assign addr[25735]= -791679244;
assign addr[25736]= -1067110699;
assign addr[25737]= -1320917099;
assign addr[25738]= -1547955041;
assign addr[25739]= -1743623590;
assign addr[25740]= -1903957513;
assign addr[25741]= -2025707632;
assign addr[25742]= -2106406677;
assign addr[25743]= -2144419275;
assign addr[25744]= -2138975100;
assign addr[25745]= -2090184478;
assign addr[25746]= -1999036154;
assign addr[25747]= -1867377253;
assign addr[25748]= -1697875851;
assign addr[25749]= -1493966902;
assign addr[25750]= -1259782632;
assign addr[25751]= -1000068799;
assign addr[25752]= -720088517;
assign addr[25753]= -425515602;
assign addr[25754]= -122319591;
assign addr[25755]= 183355234;
assign addr[25756]= 485314355;
assign addr[25757]= 777438554;
assign addr[25758]= 1053807919;
assign addr[25759]= 1308821808;
assign addr[25760]= 1537312353;
assign addr[25761]= 1734649179;
assign addr[25762]= 1896833245;
assign addr[25763]= 2020577882;
assign addr[25764]= 2103375398;
assign addr[25765]= 2143547897;
assign addr[25766]= 2140281282;
assign addr[25767]= 2093641749;
assign addr[25768]= 2004574453;
assign addr[25769]= 1874884346;
assign addr[25770]= 1707199606;
assign addr[25771]= 1504918373;
assign addr[25772]= 1272139887;
assign addr[25773]= 1013581418;
assign addr[25774]= 734482665;
assign addr[25775]= 440499581;
assign addr[25776]= 137589750;
assign addr[25777]= -168108346;
assign addr[25778]= -470399716;
assign addr[25779]= -763158411;
assign addr[25780]= -1040451659;
assign addr[25781]= -1296660098;
assign addr[25782]= -1526591649;
assign addr[25783]= -1725586737;
assign addr[25784]= -1889612716;
assign addr[25785]= -2015345591;
assign addr[25786]= -2100237377;
assign addr[25787]= -2142567738;
assign addr[25788]= -2141478848;
assign addr[25789]= -2096992772;
assign addr[25790]= -2010011024;
assign addr[25791]= -1882296293;
assign addr[25792]= -1716436725;
assign addr[25793]= -1515793473;
assign addr[25794]= -1284432584;
assign addr[25795]= -1027042599;
assign addr[25796]= -748839539;
assign addr[25797]= -455461206;
assign addr[25798]= -152852926;
assign addr[25799]= 152852926;
assign addr[25800]= 455461206;
assign addr[25801]= 748839539;
assign addr[25802]= 1027042599;
assign addr[25803]= 1284432584;
assign addr[25804]= 1515793473;
assign addr[25805]= 1716436725;
assign addr[25806]= 1882296293;
assign addr[25807]= 2010011024;
assign addr[25808]= 2096992772;
assign addr[25809]= 2141478848;
assign addr[25810]= 2142567738;
assign addr[25811]= 2100237377;
assign addr[25812]= 2015345591;
assign addr[25813]= 1889612716;
assign addr[25814]= 1725586737;
assign addr[25815]= 1526591649;
assign addr[25816]= 1296660098;
assign addr[25817]= 1040451659;
assign addr[25818]= 763158411;
assign addr[25819]= 470399716;
assign addr[25820]= 168108346;
assign addr[25821]= -137589750;
assign addr[25822]= -440499581;
assign addr[25823]= -734482665;
assign addr[25824]= -1013581418;
assign addr[25825]= -1272139887;
assign addr[25826]= -1504918373;
assign addr[25827]= -1707199606;
assign addr[25828]= -1874884346;
assign addr[25829]= -2004574453;
assign addr[25830]= -2093641749;
assign addr[25831]= -2140281282;
assign addr[25832]= -2143547897;
assign addr[25833]= -2103375398;
assign addr[25834]= -2020577882;
assign addr[25835]= -1896833245;
assign addr[25836]= -1734649179;
assign addr[25837]= -1537312353;
assign addr[25838]= -1308821808;
assign addr[25839]= -1053807919;
assign addr[25840]= -777438554;
assign addr[25841]= -485314355;
assign addr[25842]= -183355234;
assign addr[25843]= 122319591;
assign addr[25844]= 425515602;
assign addr[25845]= 720088517;
assign addr[25846]= 1000068799;
assign addr[25847]= 1259782632;
assign addr[25848]= 1493966902;
assign addr[25849]= 1697875851;
assign addr[25850]= 1867377253;
assign addr[25851]= 1999036154;
assign addr[25852]= 2090184478;
assign addr[25853]= 2138975100;
assign addr[25854]= 2144419275;
assign addr[25855]= 2106406677;
assign addr[25856]= 2025707632;
assign addr[25857]= 1903957513;
assign addr[25858]= 1743623590;
assign addr[25859]= 1547955041;
assign addr[25860]= 1320917099;
assign addr[25861]= 1067110699;
assign addr[25862]= 791679244;
assign addr[25863]= 500204365;
assign addr[25864]= 198592817;
assign addr[25865]= -107043224;
assign addr[25866]= -410510029;
assign addr[25867]= -705657826;
assign addr[25868]= -986505429;
assign addr[25869]= -1247361445;
assign addr[25870]= -1482939614;
assign addr[25871]= -1688465931;
assign addr[25872]= -1859775393;
assign addr[25873]= -1993396407;
assign addr[25874]= -2086621133;
assign addr[25875]= -2137560369;
assign addr[25876]= -2145181827;
assign addr[25877]= -2109331059;
assign addr[25878]= -2030734582;
assign addr[25879]= -1910985158;
assign addr[25880]= -1752509516;
assign addr[25881]= -1558519173;
assign addr[25882]= -1332945355;
assign addr[25883]= -1080359326;
assign addr[25884]= -805879757;
assign addr[25885]= -515068990;
assign addr[25886]= -213820322;
assign addr[25887]= 91761426;
assign addr[25888]= 395483624;
assign addr[25889]= 691191324;
assign addr[25890]= 972891995;
assign addr[25891]= 1234876957;
assign addr[25892]= 1471837070;
assign addr[25893]= 1678970324;
assign addr[25894]= 1852079154;
assign addr[25895]= 1987655498;
assign addr[25896]= 2082951896;
assign addr[25897]= 2136037160;
assign addr[25898]= 2145835515;
assign addr[25899]= 2112148396;
assign addr[25900]= 2035658475;
assign addr[25901]= 1917915825;
assign addr[25902]= 1761306505;
assign addr[25903]= 1569004214;
assign addr[25904]= 1344905966;
assign addr[25905]= 1093553126;
assign addr[25906]= 820039373;
assign addr[25907]= 529907477;
assign addr[25908]= 229036977;
assign addr[25909]= -76474970;
assign addr[25910]= -380437148;
assign addr[25911]= -676689746;
assign addr[25912]= -959229189;
assign addr[25913]= -1222329801;
assign addr[25914]= -1460659832;
assign addr[25915]= -1669389513;
assign addr[25916]= -1844288924;
assign addr[25917]= -1981813720;
assign addr[25918]= -2079176953;
assign addr[25919]= -2134405552;
assign addr[25920]= -2146380306;
assign addr[25921]= -2114858546;
assign addr[25922]= -2040479063;
assign addr[25923]= -1924749160;
assign addr[25924]= -1770014111;
assign addr[25925]= -1579409630;
assign addr[25926]= -1356798326;
assign addr[25927]= -1106691431;
assign addr[25928]= -834157373;
assign addr[25929]= -544719071;
assign addr[25930]= -244242007;
assign addr[25931]= 61184634;
assign addr[25932]= 365371365;
assign addr[25933]= 662153826;
assign addr[25934]= 945517704;
assign addr[25935]= 1209720613;
assign addr[25936]= 1449408469;
assign addr[25937]= 1659723983;
assign addr[25938]= 1836405100;
assign addr[25939]= 1975871368;
assign addr[25940]= 2075296495;
assign addr[25941]= 2132665626;
assign addr[25942]= 2146816171;
assign addr[25943]= 2117461370;
assign addr[25944]= 2045196100;
assign addr[25945]= 1931484818;
assign addr[25946]= 1778631892;
assign addr[25947]= 1589734894;
assign addr[25948]= 1368621831;
assign addr[25949]= 1119773573;
assign addr[25950]= 848233042;
assign addr[25951]= 559503022;
assign addr[25952]= 259434643;
assign addr[25953]= -45891193;
assign addr[25954]= -350287041;
assign addr[25955]= -647584304;
assign addr[25956]= -931758235;
assign addr[25957]= -1197050035;
assign addr[25958]= -1438083551;
assign addr[25959]= -1649974225;
assign addr[25960]= -1828428082;
assign addr[25961]= -1969828744;
assign addr[25962]= -2071310720;
assign addr[25963]= -2130817471;
assign addr[25964]= -2147143090;
assign addr[25965]= -2119956737;
assign addr[25966]= -2049809346;
assign addr[25967]= -1938122457;
assign addr[25968]= -1787159411;
assign addr[25969]= -1599979481;
assign addr[25970]= -1380375881;
assign addr[25971]= -1132798888;
assign addr[25972]= -862265664;
assign addr[25973]= -574258580;
assign addr[25974]= -274614114;
assign addr[25975]= 30595422;
assign addr[25976]= 335184940;
assign addr[25977]= 632981917;
assign addr[25978]= 917951481;
assign addr[25979]= 1184318708;
assign addr[25980]= 1426685652;
assign addr[25981]= 1640140734;
assign addr[25982]= 1820358275;
assign addr[25983]= 1963686155;
assign addr[25984]= 2067219829;
assign addr[25985]= 2128861181;
assign addr[25986]= 2147361045;
assign addr[25987]= 2122344521;
assign addr[25988]= 2054318569;
assign addr[25989]= 1944661739;
assign addr[25990]= 1795596234;
assign addr[25991]= 1610142873;
assign addr[25992]= 1392059879;
assign addr[25993]= 1145766716;
assign addr[25994]= 876254528;
assign addr[25995]= 588984994;
assign addr[25996]= 289779648;
assign addr[25997]= -15298099;
assign addr[25998]= -320065829;
assign addr[25999]= -618347408;
assign addr[26000]= -904098143;
assign addr[26001]= -1171527280;
assign addr[26002]= -1415215352;
assign addr[26003]= -1630224009;
assign addr[26004]= -1812196087;
assign addr[26005]= -1957443913;
assign addr[26006]= -2063024031;
assign addr[26007]= -2126796855;
assign addr[26008]= -2147470025;
assign addr[26009]= -2124624598;
assign addr[26010]= -2058723538;
assign addr[26011]= -1951102334;
assign addr[26012]= -1803941934;
assign addr[26013]= -1620224553;
assign addr[26014]= -1403673233;
assign addr[26015]= -1158676398;
assign addr[26016]= -890198924;
assign addr[26017]= -603681519;
assign addr[26018]= -304930476;
assign addr[26019]= 0;
assign addr[26020]= 304930476;
assign addr[26021]= 603681519;
assign addr[26022]= 890198924;
assign addr[26023]= 1158676398;
assign addr[26024]= 1403673233;
assign addr[26025]= 1620224553;
assign addr[26026]= 1803941934;
assign addr[26027]= 1951102334;
assign addr[26028]= 2058723538;
assign addr[26029]= 2124624598;
assign addr[26030]= 2147470025;
assign addr[26031]= 2126796855;
assign addr[26032]= 2063024031;
assign addr[26033]= 1957443913;
assign addr[26034]= 1812196087;
assign addr[26035]= 1630224009;
assign addr[26036]= 1415215352;
assign addr[26037]= 1171527280;
assign addr[26038]= 904098143;
assign addr[26039]= 618347408;
assign addr[26040]= 320065829;
assign addr[26041]= 15298099;
assign addr[26042]= -289779648;
assign addr[26043]= -588984994;
assign addr[26044]= -876254528;
assign addr[26045]= -1145766716;
assign addr[26046]= -1392059879;
assign addr[26047]= -1610142873;
assign addr[26048]= -1795596234;
assign addr[26049]= -1944661739;
assign addr[26050]= -2054318569;
assign addr[26051]= -2122344521;
assign addr[26052]= -2147361045;
assign addr[26053]= -2128861181;
assign addr[26054]= -2067219829;
assign addr[26055]= -1963686155;
assign addr[26056]= -1820358275;
assign addr[26057]= -1640140734;
assign addr[26058]= -1426685652;
assign addr[26059]= -1184318708;
assign addr[26060]= -917951481;
assign addr[26061]= -632981917;
assign addr[26062]= -335184940;
assign addr[26063]= -30595422;
assign addr[26064]= 274614114;
assign addr[26065]= 574258580;
assign addr[26066]= 862265664;
assign addr[26067]= 1132798888;
assign addr[26068]= 1380375881;
assign addr[26069]= 1599979481;
assign addr[26070]= 1787159411;
assign addr[26071]= 1938122457;
assign addr[26072]= 2049809346;
assign addr[26073]= 2119956737;
assign addr[26074]= 2147143090;
assign addr[26075]= 2130817471;
assign addr[26076]= 2071310720;
assign addr[26077]= 1969828744;
assign addr[26078]= 1828428082;
assign addr[26079]= 1649974225;
assign addr[26080]= 1438083551;
assign addr[26081]= 1197050035;
assign addr[26082]= 931758235;
assign addr[26083]= 647584304;
assign addr[26084]= 350287041;
assign addr[26085]= 45891193;
assign addr[26086]= -259434643;
assign addr[26087]= -559503022;
assign addr[26088]= -848233042;
assign addr[26089]= -1119773573;
assign addr[26090]= -1368621831;
assign addr[26091]= -1589734894;
assign addr[26092]= -1778631892;
assign addr[26093]= -1931484818;
assign addr[26094]= -2045196100;
assign addr[26095]= -2117461370;
assign addr[26096]= -2146816171;
assign addr[26097]= -2132665626;
assign addr[26098]= -2075296495;
assign addr[26099]= -1975871368;
assign addr[26100]= -1836405100;
assign addr[26101]= -1659723983;
assign addr[26102]= -1449408469;
assign addr[26103]= -1209720613;
assign addr[26104]= -945517704;
assign addr[26105]= -662153826;
assign addr[26106]= -365371365;
assign addr[26107]= -61184634;
assign addr[26108]= 244242007;
assign addr[26109]= 544719071;
assign addr[26110]= 834157373;
assign addr[26111]= 1106691431;
assign addr[26112]= 1356798326;
assign addr[26113]= 1579409630;
assign addr[26114]= 1770014111;
assign addr[26115]= 1924749160;
assign addr[26116]= 2040479063;
assign addr[26117]= 2114858546;
assign addr[26118]= 2146380306;
assign addr[26119]= 2134405552;
assign addr[26120]= 2079176953;
assign addr[26121]= 1981813720;
assign addr[26122]= 1844288924;
assign addr[26123]= 1669389513;
assign addr[26124]= 1460659832;
assign addr[26125]= 1222329801;
assign addr[26126]= 959229189;
assign addr[26127]= 676689746;
assign addr[26128]= 380437148;
assign addr[26129]= 76474970;
assign addr[26130]= -229036977;
assign addr[26131]= -529907477;
assign addr[26132]= -820039373;
assign addr[26133]= -1093553126;
assign addr[26134]= -1344905966;
assign addr[26135]= -1569004214;
assign addr[26136]= -1761306505;
assign addr[26137]= -1917915825;
assign addr[26138]= -2035658475;
assign addr[26139]= -2112148396;
assign addr[26140]= -2145835515;
assign addr[26141]= -2136037160;
assign addr[26142]= -2082951896;
assign addr[26143]= -1987655498;
assign addr[26144]= -1852079154;
assign addr[26145]= -1678970324;
assign addr[26146]= -1471837070;
assign addr[26147]= -1234876957;
assign addr[26148]= -972891995;
assign addr[26149]= -691191324;
assign addr[26150]= -395483624;
assign addr[26151]= -91761426;
assign addr[26152]= 213820322;
assign addr[26153]= 515068990;
assign addr[26154]= 805879757;
assign addr[26155]= 1080359326;
assign addr[26156]= 1332945355;
assign addr[26157]= 1558519173;
assign addr[26158]= 1752509516;
assign addr[26159]= 1910985158;
assign addr[26160]= 2030734582;
assign addr[26161]= 2109331059;
assign addr[26162]= 2145181827;
assign addr[26163]= 2137560369;
assign addr[26164]= 2086621133;
assign addr[26165]= 1993396407;
assign addr[26166]= 1859775393;
assign addr[26167]= 1688465931;
assign addr[26168]= 1482939614;
assign addr[26169]= 1247361445;
assign addr[26170]= 986505429;
assign addr[26171]= 705657826;
assign addr[26172]= 410510029;
assign addr[26173]= 107043224;
assign addr[26174]= -198592817;
assign addr[26175]= -500204365;
assign addr[26176]= -791679244;
assign addr[26177]= -1067110699;
assign addr[26178]= -1320917099;
assign addr[26179]= -1547955041;
assign addr[26180]= -1743623590;
assign addr[26181]= -1903957513;
assign addr[26182]= -2025707632;
assign addr[26183]= -2106406677;
assign addr[26184]= -2144419275;
assign addr[26185]= -2138975100;
assign addr[26186]= -2090184478;
assign addr[26187]= -1999036154;
assign addr[26188]= -1867377253;
assign addr[26189]= -1697875851;
assign addr[26190]= -1493966902;
assign addr[26191]= -1259782632;
assign addr[26192]= -1000068799;
assign addr[26193]= -720088517;
assign addr[26194]= -425515602;
assign addr[26195]= -122319591;
assign addr[26196]= 183355234;
assign addr[26197]= 485314355;
assign addr[26198]= 777438554;
assign addr[26199]= 1053807919;
assign addr[26200]= 1308821808;
assign addr[26201]= 1537312353;
assign addr[26202]= 1734649179;
assign addr[26203]= 1896833245;
assign addr[26204]= 2020577882;
assign addr[26205]= 2103375398;
assign addr[26206]= 2143547897;
assign addr[26207]= 2140281282;
assign addr[26208]= 2093641749;
assign addr[26209]= 2004574453;
assign addr[26210]= 1874884346;
assign addr[26211]= 1707199606;
assign addr[26212]= 1504918373;
assign addr[26213]= 1272139887;
assign addr[26214]= 1013581418;
assign addr[26215]= 734482665;
assign addr[26216]= 440499581;
assign addr[26217]= 137589750;
assign addr[26218]= -168108346;
assign addr[26219]= -470399716;
assign addr[26220]= -763158411;
assign addr[26221]= -1040451659;
assign addr[26222]= -1296660098;
assign addr[26223]= -1526591649;
assign addr[26224]= -1725586737;
assign addr[26225]= -1889612716;
assign addr[26226]= -2015345591;
assign addr[26227]= -2100237377;
assign addr[26228]= -2142567738;
assign addr[26229]= -2141478848;
assign addr[26230]= -2096992772;
assign addr[26231]= -2010011024;
assign addr[26232]= -1882296293;
assign addr[26233]= -1716436725;
assign addr[26234]= -1515793473;
assign addr[26235]= -1284432584;
assign addr[26236]= -1027042599;
assign addr[26237]= -748839539;
assign addr[26238]= -455461206;
assign addr[26239]= -152852926;
assign addr[26240]= 152852926;
assign addr[26241]= 455461206;
assign addr[26242]= 748839539;
assign addr[26243]= 1027042599;
assign addr[26244]= 1284432584;
assign addr[26245]= 1515793473;
assign addr[26246]= 1716436725;
assign addr[26247]= 1882296293;
assign addr[26248]= 2010011024;
assign addr[26249]= 2096992772;
assign addr[26250]= 2141478848;
assign addr[26251]= 2142567738;
assign addr[26252]= 2100237377;
assign addr[26253]= 2015345591;
assign addr[26254]= 1889612716;
assign addr[26255]= 1725586737;
assign addr[26256]= 1526591649;
assign addr[26257]= 1296660098;
assign addr[26258]= 1040451659;
assign addr[26259]= 763158411;
assign addr[26260]= 470399716;
assign addr[26261]= 168108346;
assign addr[26262]= -137589750;
assign addr[26263]= -440499581;
assign addr[26264]= -734482665;
assign addr[26265]= -1013581418;
assign addr[26266]= -1272139887;
assign addr[26267]= -1504918373;
assign addr[26268]= -1707199606;
assign addr[26269]= -1874884346;
assign addr[26270]= -2004574453;
assign addr[26271]= -2093641749;
assign addr[26272]= -2140281282;
assign addr[26273]= -2143547897;
assign addr[26274]= -2103375398;
assign addr[26275]= -2020577882;
assign addr[26276]= -1896833245;
assign addr[26277]= -1734649179;
assign addr[26278]= -1537312353;
assign addr[26279]= -1308821808;
assign addr[26280]= -1053807919;
assign addr[26281]= -777438554;
assign addr[26282]= -485314355;
assign addr[26283]= -183355234;
assign addr[26284]= 122319591;
assign addr[26285]= 425515602;
assign addr[26286]= 720088517;
assign addr[26287]= 1000068799;
assign addr[26288]= 1259782632;
assign addr[26289]= 1493966902;
assign addr[26290]= 1697875851;
assign addr[26291]= 1867377253;
assign addr[26292]= 1999036154;
assign addr[26293]= 2090184478;
assign addr[26294]= 2138975100;
assign addr[26295]= 2144419275;
assign addr[26296]= 2106406677;
assign addr[26297]= 2025707632;
assign addr[26298]= 1903957513;
assign addr[26299]= 1743623590;
assign addr[26300]= 1547955041;
assign addr[26301]= 1320917099;
assign addr[26302]= 1067110699;
assign addr[26303]= 791679244;
assign addr[26304]= 500204365;
assign addr[26305]= 198592817;
assign addr[26306]= -107043224;
assign addr[26307]= -410510029;
assign addr[26308]= -705657826;
assign addr[26309]= -986505429;
assign addr[26310]= -1247361445;
assign addr[26311]= -1482939614;
assign addr[26312]= -1688465931;
assign addr[26313]= -1859775393;
assign addr[26314]= -1993396407;
assign addr[26315]= -2086621133;
assign addr[26316]= -2137560369;
assign addr[26317]= -2145181827;
assign addr[26318]= -2109331059;
assign addr[26319]= -2030734582;
assign addr[26320]= -1910985158;
assign addr[26321]= -1752509516;
assign addr[26322]= -1558519173;
assign addr[26323]= -1332945355;
assign addr[26324]= -1080359326;
assign addr[26325]= -805879757;
assign addr[26326]= -515068990;
assign addr[26327]= -213820322;
assign addr[26328]= 91761426;
assign addr[26329]= 395483624;
assign addr[26330]= 691191324;
assign addr[26331]= 972891995;
assign addr[26332]= 1234876957;
assign addr[26333]= 1471837070;
assign addr[26334]= 1678970324;
assign addr[26335]= 1852079154;
assign addr[26336]= 1987655498;
assign addr[26337]= 2082951896;
assign addr[26338]= 2136037160;
assign addr[26339]= 2145835515;
assign addr[26340]= 2112148396;
assign addr[26341]= 2035658475;
assign addr[26342]= 1917915825;
assign addr[26343]= 1761306505;
assign addr[26344]= 1569004214;
assign addr[26345]= 1344905966;
assign addr[26346]= 1093553126;
assign addr[26347]= 820039373;
assign addr[26348]= 529907477;
assign addr[26349]= 229036977;
assign addr[26350]= -76474970;
assign addr[26351]= -380437148;
assign addr[26352]= -676689746;
assign addr[26353]= -959229189;
assign addr[26354]= -1222329801;
assign addr[26355]= -1460659832;
assign addr[26356]= -1669389513;
assign addr[26357]= -1844288924;
assign addr[26358]= -1981813720;
assign addr[26359]= -2079176953;
assign addr[26360]= -2134405552;
assign addr[26361]= -2146380306;
assign addr[26362]= -2114858546;
assign addr[26363]= -2040479063;
assign addr[26364]= -1924749160;
assign addr[26365]= -1770014111;
assign addr[26366]= -1579409630;
assign addr[26367]= -1356798326;
assign addr[26368]= -1106691431;
assign addr[26369]= -834157373;
assign addr[26370]= -544719071;
assign addr[26371]= -244242007;
assign addr[26372]= 61184634;
assign addr[26373]= 365371365;
assign addr[26374]= 662153826;
assign addr[26375]= 945517704;
assign addr[26376]= 1209720613;
assign addr[26377]= 1449408469;
assign addr[26378]= 1659723983;
assign addr[26379]= 1836405100;
assign addr[26380]= 1975871368;
assign addr[26381]= 2075296495;
assign addr[26382]= 2132665626;
assign addr[26383]= 2146816171;
assign addr[26384]= 2117461370;
assign addr[26385]= 2045196100;
assign addr[26386]= 1931484818;
assign addr[26387]= 1778631892;
assign addr[26388]= 1589734894;
assign addr[26389]= 1368621831;
assign addr[26390]= 1119773573;
assign addr[26391]= 848233042;
assign addr[26392]= 559503022;
assign addr[26393]= 259434643;
assign addr[26394]= -45891193;
assign addr[26395]= -350287041;
assign addr[26396]= -647584304;
assign addr[26397]= -931758235;
assign addr[26398]= -1197050035;
assign addr[26399]= -1438083551;
assign addr[26400]= -1649974225;
assign addr[26401]= -1828428082;
assign addr[26402]= -1969828744;
assign addr[26403]= -2071310720;
assign addr[26404]= -2130817471;
assign addr[26405]= -2147143090;
assign addr[26406]= -2119956737;
assign addr[26407]= -2049809346;
assign addr[26408]= -1938122457;
assign addr[26409]= -1787159411;
assign addr[26410]= -1599979481;
assign addr[26411]= -1380375881;
assign addr[26412]= -1132798888;
assign addr[26413]= -862265664;
assign addr[26414]= -574258580;
assign addr[26415]= -274614114;
assign addr[26416]= 30595422;
assign addr[26417]= 335184940;
assign addr[26418]= 632981917;
assign addr[26419]= 917951481;
assign addr[26420]= 1184318708;
assign addr[26421]= 1426685652;
assign addr[26422]= 1640140734;
assign addr[26423]= 1820358275;
assign addr[26424]= 1963686155;
assign addr[26425]= 2067219829;
assign addr[26426]= 2128861181;
assign addr[26427]= 2147361045;
assign addr[26428]= 2122344521;
assign addr[26429]= 2054318569;
assign addr[26430]= 1944661739;
assign addr[26431]= 1795596234;
assign addr[26432]= 1610142873;
assign addr[26433]= 1392059879;
assign addr[26434]= 1145766716;
assign addr[26435]= 876254528;
assign addr[26436]= 588984994;
assign addr[26437]= 289779648;
assign addr[26438]= -15298099;
assign addr[26439]= -320065829;
assign addr[26440]= -618347408;
assign addr[26441]= -904098143;
assign addr[26442]= -1171527280;
assign addr[26443]= -1415215352;
assign addr[26444]= -1630224009;
assign addr[26445]= -1812196087;
assign addr[26446]= -1957443913;
assign addr[26447]= -2063024031;
assign addr[26448]= -2126796855;
assign addr[26449]= -2147470025;
assign addr[26450]= -2124624598;
assign addr[26451]= -2058723538;
assign addr[26452]= -1951102334;
assign addr[26453]= -1803941934;
assign addr[26454]= -1620224553;
assign addr[26455]= -1403673233;
assign addr[26456]= -1158676398;
assign addr[26457]= -890198924;
assign addr[26458]= -603681519;
assign addr[26459]= -304930476;
assign addr[26460]= 0;
assign addr[26461]= 304930476;
assign addr[26462]= 603681519;
assign addr[26463]= 890198924;
assign addr[26464]= 1158676398;
assign addr[26465]= 1403673233;
assign addr[26466]= 1620224553;
assign addr[26467]= 1803941934;
assign addr[26468]= 1951102334;
assign addr[26469]= 2058723538;
assign addr[26470]= 2124624598;
assign addr[26471]= 2147470025;
assign addr[26472]= 2126796855;
assign addr[26473]= 2063024031;
assign addr[26474]= 1957443913;
assign addr[26475]= 1812196087;
assign addr[26476]= 1630224009;
assign addr[26477]= 1415215352;
assign addr[26478]= 1171527280;
assign addr[26479]= 904098143;
assign addr[26480]= 618347408;
assign addr[26481]= 320065829;
assign addr[26482]= 15298099;
assign addr[26483]= -289779648;
assign addr[26484]= -588984994;
assign addr[26485]= -876254528;
assign addr[26486]= -1145766716;
assign addr[26487]= -1392059879;
assign addr[26488]= -1610142873;
assign addr[26489]= -1795596234;
assign addr[26490]= -1944661739;
assign addr[26491]= -2054318569;
assign addr[26492]= -2122344521;
assign addr[26493]= -2147361045;
assign addr[26494]= -2128861181;
assign addr[26495]= -2067219829;
assign addr[26496]= -1963686155;
assign addr[26497]= -1820358275;
assign addr[26498]= -1640140734;
assign addr[26499]= -1426685652;
assign addr[26500]= -1184318708;
assign addr[26501]= -917951481;
assign addr[26502]= -632981917;
assign addr[26503]= -335184940;
assign addr[26504]= -30595422;
assign addr[26505]= 274614114;
assign addr[26506]= 574258580;
assign addr[26507]= 862265664;
assign addr[26508]= 1132798888;
assign addr[26509]= 1380375881;
assign addr[26510]= 1599979481;
assign addr[26511]= 1787159411;
assign addr[26512]= 1938122457;
assign addr[26513]= 2049809346;
assign addr[26514]= 2119956737;
assign addr[26515]= 2147143090;
assign addr[26516]= 2130817471;
assign addr[26517]= 2071310720;
assign addr[26518]= 1969828744;
assign addr[26519]= 1828428082;
assign addr[26520]= 1649974225;
assign addr[26521]= 1438083551;
assign addr[26522]= 1197050035;
assign addr[26523]= 931758235;
assign addr[26524]= 647584304;
assign addr[26525]= 350287041;
assign addr[26526]= 45891193;
assign addr[26527]= -259434643;
assign addr[26528]= -559503022;
assign addr[26529]= -848233042;
assign addr[26530]= -1119773573;
assign addr[26531]= -1368621831;
assign addr[26532]= -1589734894;
assign addr[26533]= -1778631892;
assign addr[26534]= -1931484818;
assign addr[26535]= -2045196100;
assign addr[26536]= -2117461370;
assign addr[26537]= -2146816171;
assign addr[26538]= -2132665626;
assign addr[26539]= -2075296495;
assign addr[26540]= -1975871368;
assign addr[26541]= -1836405100;
assign addr[26542]= -1659723983;
assign addr[26543]= -1449408469;
assign addr[26544]= -1209720613;
assign addr[26545]= -945517704;
assign addr[26546]= -662153826;
assign addr[26547]= -365371365;
assign addr[26548]= -61184634;
assign addr[26549]= 244242007;
assign addr[26550]= 544719071;
assign addr[26551]= 834157373;
assign addr[26552]= 1106691431;
assign addr[26553]= 1356798326;
assign addr[26554]= 1579409630;
assign addr[26555]= 1770014111;
assign addr[26556]= 1924749160;
assign addr[26557]= 2040479063;
assign addr[26558]= 2114858546;
assign addr[26559]= 2146380306;
assign addr[26560]= 2134405552;
assign addr[26561]= 2079176953;
assign addr[26562]= 1981813720;
assign addr[26563]= 1844288924;
assign addr[26564]= 1669389513;
assign addr[26565]= 1460659832;
assign addr[26566]= 1222329801;
assign addr[26567]= 959229189;
assign addr[26568]= 676689746;
assign addr[26569]= 380437148;
assign addr[26570]= 76474970;
assign addr[26571]= -229036977;
assign addr[26572]= -529907477;
assign addr[26573]= -820039373;
assign addr[26574]= -1093553126;
assign addr[26575]= -1344905966;
assign addr[26576]= -1569004214;
assign addr[26577]= -1761306505;
assign addr[26578]= -1917915825;
assign addr[26579]= -2035658475;
assign addr[26580]= -2112148396;
assign addr[26581]= -2145835515;
assign addr[26582]= -2136037160;
assign addr[26583]= -2082951896;
assign addr[26584]= -1987655498;
assign addr[26585]= -1852079154;
assign addr[26586]= -1678970324;
assign addr[26587]= -1471837070;
assign addr[26588]= -1234876957;
assign addr[26589]= -972891995;
assign addr[26590]= -691191324;
assign addr[26591]= -395483624;
assign addr[26592]= -91761426;
assign addr[26593]= 213820322;
assign addr[26594]= 515068990;
assign addr[26595]= 805879757;
assign addr[26596]= 1080359326;
assign addr[26597]= 1332945355;
assign addr[26598]= 1558519173;
assign addr[26599]= 1752509516;
assign addr[26600]= 1910985158;
assign addr[26601]= 2030734582;
assign addr[26602]= 2109331059;
assign addr[26603]= 2145181827;
assign addr[26604]= 2137560369;
assign addr[26605]= 2086621133;
assign addr[26606]= 1993396407;
assign addr[26607]= 1859775393;
assign addr[26608]= 1688465931;
assign addr[26609]= 1482939614;
assign addr[26610]= 1247361445;
assign addr[26611]= 986505429;
assign addr[26612]= 705657826;
assign addr[26613]= 410510029;
assign addr[26614]= 107043224;
assign addr[26615]= -198592817;
assign addr[26616]= -500204365;
assign addr[26617]= -791679244;
assign addr[26618]= -1067110699;
assign addr[26619]= -1320917099;
assign addr[26620]= -1547955041;
assign addr[26621]= -1743623590;
assign addr[26622]= -1903957513;
assign addr[26623]= -2025707632;
assign addr[26624]= -2106406677;
assign addr[26625]= -2144419275;
assign addr[26626]= -2138975100;
assign addr[26627]= -2090184478;
assign addr[26628]= -1999036154;
assign addr[26629]= -1867377253;
assign addr[26630]= -1697875851;
assign addr[26631]= -1493966902;
assign addr[26632]= -1259782632;
assign addr[26633]= -1000068799;
assign addr[26634]= -720088517;
assign addr[26635]= -425515602;
assign addr[26636]= -122319591;
assign addr[26637]= 183355234;
assign addr[26638]= 485314355;
assign addr[26639]= 777438554;
assign addr[26640]= 1053807919;
assign addr[26641]= 1308821808;
assign addr[26642]= 1537312353;
assign addr[26643]= 1734649179;
assign addr[26644]= 1896833245;
assign addr[26645]= 2020577882;
assign addr[26646]= 2103375398;
assign addr[26647]= 2143547897;
assign addr[26648]= 2140281282;
assign addr[26649]= 2093641749;
assign addr[26650]= 2004574453;
assign addr[26651]= 1874884346;
assign addr[26652]= 1707199606;
assign addr[26653]= 1504918373;
assign addr[26654]= 1272139887;
assign addr[26655]= 1013581418;
assign addr[26656]= 734482665;
assign addr[26657]= 440499581;
assign addr[26658]= 137589750;
assign addr[26659]= -168108346;
assign addr[26660]= -470399716;
assign addr[26661]= -763158411;
assign addr[26662]= -1040451659;
assign addr[26663]= -1296660098;
assign addr[26664]= -1526591649;
assign addr[26665]= -1725586737;
assign addr[26666]= -1889612716;
assign addr[26667]= -2015345591;
assign addr[26668]= -2100237377;
assign addr[26669]= -2142567738;
assign addr[26670]= -2141478848;
assign addr[26671]= -2096992772;
assign addr[26672]= -2010011024;
assign addr[26673]= -1882296293;
assign addr[26674]= -1716436725;
assign addr[26675]= -1515793473;
assign addr[26676]= -1284432584;
assign addr[26677]= -1027042599;
assign addr[26678]= -748839539;
assign addr[26679]= -455461206;
assign addr[26680]= -152852926;
assign addr[26681]= 152852926;
assign addr[26682]= 455461206;
assign addr[26683]= 748839539;
assign addr[26684]= 1027042599;
assign addr[26685]= 1284432584;
assign addr[26686]= 1515793473;
assign addr[26687]= 1716436725;
assign addr[26688]= 1882296293;
assign addr[26689]= 2010011024;
assign addr[26690]= 2096992772;
assign addr[26691]= 2141478848;
assign addr[26692]= 2142567738;
assign addr[26693]= 2100237377;
assign addr[26694]= 2015345591;
assign addr[26695]= 1889612716;
assign addr[26696]= 1725586737;
assign addr[26697]= 1526591649;
assign addr[26698]= 1296660098;
assign addr[26699]= 1040451659;
assign addr[26700]= 763158411;
assign addr[26701]= 470399716;
assign addr[26702]= 168108346;
assign addr[26703]= -137589750;
assign addr[26704]= -440499581;
assign addr[26705]= -734482665;
assign addr[26706]= -1013581418;
assign addr[26707]= -1272139887;
assign addr[26708]= -1504918373;
assign addr[26709]= -1707199606;
assign addr[26710]= -1874884346;
assign addr[26711]= -2004574453;
assign addr[26712]= -2093641749;
assign addr[26713]= -2140281282;
assign addr[26714]= -2143547897;
assign addr[26715]= -2103375398;
assign addr[26716]= -2020577882;
assign addr[26717]= -1896833245;
assign addr[26718]= -1734649179;
assign addr[26719]= -1537312353;
assign addr[26720]= -1308821808;
assign addr[26721]= -1053807919;
assign addr[26722]= -777438554;
assign addr[26723]= -485314355;
assign addr[26724]= -183355234;
assign addr[26725]= 122319591;
assign addr[26726]= 425515602;
assign addr[26727]= 720088517;
assign addr[26728]= 1000068799;
assign addr[26729]= 1259782632;
assign addr[26730]= 1493966902;
assign addr[26731]= 1697875851;
assign addr[26732]= 1867377253;
assign addr[26733]= 1999036154;
assign addr[26734]= 2090184478;
assign addr[26735]= 2138975100;
assign addr[26736]= 2144419275;
assign addr[26737]= 2106406677;
assign addr[26738]= 2025707632;
assign addr[26739]= 1903957513;
assign addr[26740]= 1743623590;
assign addr[26741]= 1547955041;
assign addr[26742]= 1320917099;
assign addr[26743]= 1067110699;
assign addr[26744]= 791679244;
assign addr[26745]= 500204365;
assign addr[26746]= 198592817;
assign addr[26747]= -107043224;
assign addr[26748]= -410510029;
assign addr[26749]= -705657826;
assign addr[26750]= -986505429;
assign addr[26751]= -1247361445;
assign addr[26752]= -1482939614;
assign addr[26753]= -1688465931;
assign addr[26754]= -1859775393;
assign addr[26755]= -1993396407;
assign addr[26756]= -2086621133;
assign addr[26757]= -2137560369;
assign addr[26758]= -2145181827;
assign addr[26759]= -2109331059;
assign addr[26760]= -2030734582;
assign addr[26761]= -1910985158;
assign addr[26762]= -1752509516;
assign addr[26763]= -1558519173;
assign addr[26764]= -1332945355;
assign addr[26765]= -1080359326;
assign addr[26766]= -805879757;
assign addr[26767]= -515068990;
assign addr[26768]= -213820322;
assign addr[26769]= 91761426;
assign addr[26770]= 395483624;
assign addr[26771]= 691191324;
assign addr[26772]= 972891995;
assign addr[26773]= 1234876957;
assign addr[26774]= 1471837070;
assign addr[26775]= 1678970324;
assign addr[26776]= 1852079154;
assign addr[26777]= 1987655498;
assign addr[26778]= 2082951896;
assign addr[26779]= 2136037160;
assign addr[26780]= 2145835515;
assign addr[26781]= 2112148396;
assign addr[26782]= 2035658475;
assign addr[26783]= 1917915825;
assign addr[26784]= 1761306505;
assign addr[26785]= 1569004214;
assign addr[26786]= 1344905966;
assign addr[26787]= 1093553126;
assign addr[26788]= 820039373;
assign addr[26789]= 529907477;
assign addr[26790]= 229036977;
assign addr[26791]= -76474970;
assign addr[26792]= -380437148;
assign addr[26793]= -676689746;
assign addr[26794]= -959229189;
assign addr[26795]= -1222329801;
assign addr[26796]= -1460659832;
assign addr[26797]= -1669389513;
assign addr[26798]= -1844288924;
assign addr[26799]= -1981813720;
assign addr[26800]= -2079176953;
assign addr[26801]= -2134405552;
assign addr[26802]= -2146380306;
assign addr[26803]= -2114858546;
assign addr[26804]= -2040479063;
assign addr[26805]= -1924749160;
assign addr[26806]= -1770014111;
assign addr[26807]= -1579409630;
assign addr[26808]= -1356798326;
assign addr[26809]= -1106691431;
assign addr[26810]= -834157373;
assign addr[26811]= -544719071;
assign addr[26812]= -244242007;
assign addr[26813]= 61184634;
assign addr[26814]= 365371365;
assign addr[26815]= 662153826;
assign addr[26816]= 945517704;
assign addr[26817]= 1209720613;
assign addr[26818]= 1449408469;
assign addr[26819]= 1659723983;
assign addr[26820]= 1836405100;
assign addr[26821]= 1975871368;
assign addr[26822]= 2075296495;
assign addr[26823]= 2132665626;
assign addr[26824]= 2146816171;
assign addr[26825]= 2117461370;
assign addr[26826]= 2045196100;
assign addr[26827]= 1931484818;
assign addr[26828]= 1778631892;
assign addr[26829]= 1589734894;
assign addr[26830]= 1368621831;
assign addr[26831]= 1119773573;
assign addr[26832]= 848233042;
assign addr[26833]= 559503022;
assign addr[26834]= 259434643;
assign addr[26835]= -45891193;
assign addr[26836]= -350287041;
assign addr[26837]= -647584304;
assign addr[26838]= -931758235;
assign addr[26839]= -1197050035;
assign addr[26840]= -1438083551;
assign addr[26841]= -1649974225;
assign addr[26842]= -1828428082;
assign addr[26843]= -1969828744;
assign addr[26844]= -2071310720;
assign addr[26845]= -2130817471;
assign addr[26846]= -2147143090;
assign addr[26847]= -2119956737;
assign addr[26848]= -2049809346;
assign addr[26849]= -1938122457;
assign addr[26850]= -1787159411;
assign addr[26851]= -1599979481;
assign addr[26852]= -1380375881;
assign addr[26853]= -1132798888;
assign addr[26854]= -862265664;
assign addr[26855]= -574258580;
assign addr[26856]= -274614114;
assign addr[26857]= 30595422;
assign addr[26858]= 335184940;
assign addr[26859]= 632981917;
assign addr[26860]= 917951481;
assign addr[26861]= 1184318708;
assign addr[26862]= 1426685652;
assign addr[26863]= 1640140734;
assign addr[26864]= 1820358275;
assign addr[26865]= 1963686155;
assign addr[26866]= 2067219829;
assign addr[26867]= 2128861181;
assign addr[26868]= 2147361045;
assign addr[26869]= 2122344521;
assign addr[26870]= 2054318569;
assign addr[26871]= 1944661739;
assign addr[26872]= 1795596234;
assign addr[26873]= 1610142873;
assign addr[26874]= 1392059879;
assign addr[26875]= 1145766716;
assign addr[26876]= 876254528;
assign addr[26877]= 588984994;
assign addr[26878]= 289779648;
assign addr[26879]= -15298099;
assign addr[26880]= -320065829;
assign addr[26881]= -618347408;
assign addr[26882]= -904098143;
assign addr[26883]= -1171527280;
assign addr[26884]= -1415215352;
assign addr[26885]= -1630224009;
assign addr[26886]= -1812196087;
assign addr[26887]= -1957443913;
assign addr[26888]= -2063024031;
assign addr[26889]= -2126796855;
assign addr[26890]= -2147470025;
assign addr[26891]= -2124624598;
assign addr[26892]= -2058723538;
assign addr[26893]= -1951102334;
assign addr[26894]= -1803941934;
assign addr[26895]= -1620224553;
assign addr[26896]= -1403673233;
assign addr[26897]= -1158676398;
assign addr[26898]= -890198924;
assign addr[26899]= -603681519;
assign addr[26900]= -304930476;
assign addr[26901]= 0;
assign addr[26902]= 304930476;
assign addr[26903]= 603681519;
assign addr[26904]= 890198924;
assign addr[26905]= 1158676398;
assign addr[26906]= 1403673233;
assign addr[26907]= 1620224553;
assign addr[26908]= 1803941934;
assign addr[26909]= 1951102334;
assign addr[26910]= 2058723538;
assign addr[26911]= 2124624598;
assign addr[26912]= 2147470025;
assign addr[26913]= 2126796855;
assign addr[26914]= 2063024031;
assign addr[26915]= 1957443913;
assign addr[26916]= 1812196087;
assign addr[26917]= 1630224009;
assign addr[26918]= 1415215352;
assign addr[26919]= 1171527280;
assign addr[26920]= 904098143;
assign addr[26921]= 618347408;
assign addr[26922]= 320065829;
assign addr[26923]= 15298099;
assign addr[26924]= -289779648;
assign addr[26925]= -588984994;
assign addr[26926]= -876254528;
assign addr[26927]= -1145766716;
assign addr[26928]= -1392059879;
assign addr[26929]= -1610142873;
assign addr[26930]= -1795596234;
assign addr[26931]= -1944661739;
assign addr[26932]= -2054318569;
assign addr[26933]= -2122344521;
assign addr[26934]= -2147361045;
assign addr[26935]= -2128861181;
assign addr[26936]= -2067219829;
assign addr[26937]= -1963686155;
assign addr[26938]= -1820358275;
assign addr[26939]= -1640140734;
assign addr[26940]= -1426685652;
assign addr[26941]= -1184318708;
assign addr[26942]= -917951481;
assign addr[26943]= -632981917;
assign addr[26944]= -335184940;
assign addr[26945]= -30595422;
assign addr[26946]= 274614114;
assign addr[26947]= 574258580;
assign addr[26948]= 862265664;
assign addr[26949]= 1132798888;
assign addr[26950]= 1380375881;
assign addr[26951]= 1599979481;
assign addr[26952]= 1787159411;
assign addr[26953]= 1938122457;
assign addr[26954]= 2049809346;
assign addr[26955]= 2119956737;
assign addr[26956]= 2147143090;
assign addr[26957]= 2130817471;
assign addr[26958]= 2071310720;
assign addr[26959]= 1969828744;
assign addr[26960]= 1828428082;
assign addr[26961]= 1649974225;
assign addr[26962]= 1438083551;
assign addr[26963]= 1197050035;
assign addr[26964]= 931758235;
assign addr[26965]= 647584304;
assign addr[26966]= 350287041;
assign addr[26967]= 45891193;
assign addr[26968]= -259434643;
assign addr[26969]= -559503022;
assign addr[26970]= -848233042;
assign addr[26971]= -1119773573;
assign addr[26972]= -1368621831;
assign addr[26973]= -1589734894;
assign addr[26974]= -1778631892;
assign addr[26975]= -1931484818;
assign addr[26976]= -2045196100;
assign addr[26977]= -2117461370;
assign addr[26978]= -2146816171;
assign addr[26979]= -2132665626;
assign addr[26980]= -2075296495;
assign addr[26981]= -1975871368;
assign addr[26982]= -1836405100;
assign addr[26983]= -1659723983;
assign addr[26984]= -1449408469;
assign addr[26985]= -1209720613;
assign addr[26986]= -945517704;
assign addr[26987]= -662153826;
assign addr[26988]= -365371365;
assign addr[26989]= -61184634;
assign addr[26990]= 244242007;
assign addr[26991]= 544719071;
assign addr[26992]= 834157373;
assign addr[26993]= 1106691431;
assign addr[26994]= 1356798326;
assign addr[26995]= 1579409630;
assign addr[26996]= 1770014111;
assign addr[26997]= 1924749160;
assign addr[26998]= 2040479063;
assign addr[26999]= 2114858546;
assign addr[27000]= 2146380306;
assign addr[27001]= 2134405552;
assign addr[27002]= 2079176953;
assign addr[27003]= 1981813720;
assign addr[27004]= 1844288924;
assign addr[27005]= 1669389513;
assign addr[27006]= 1460659832;
assign addr[27007]= 1222329801;
assign addr[27008]= 959229189;
assign addr[27009]= 676689746;
assign addr[27010]= 380437148;
assign addr[27011]= 76474970;
assign addr[27012]= -229036977;
assign addr[27013]= -529907477;
assign addr[27014]= -820039373;
assign addr[27015]= -1093553126;
assign addr[27016]= -1344905966;
assign addr[27017]= -1569004214;
assign addr[27018]= -1761306505;
assign addr[27019]= -1917915825;
assign addr[27020]= -2035658475;
assign addr[27021]= -2112148396;
assign addr[27022]= -2145835515;
assign addr[27023]= -2136037160;
assign addr[27024]= -2082951896;
assign addr[27025]= -1987655498;
assign addr[27026]= -1852079154;
assign addr[27027]= -1678970324;
assign addr[27028]= -1471837070;
assign addr[27029]= -1234876957;
assign addr[27030]= -972891995;
assign addr[27031]= -691191324;
assign addr[27032]= -395483624;
assign addr[27033]= -91761426;
assign addr[27034]= 213820322;
assign addr[27035]= 515068990;
assign addr[27036]= 805879757;
assign addr[27037]= 1080359326;
assign addr[27038]= 1332945355;
assign addr[27039]= 1558519173;
assign addr[27040]= 1752509516;
assign addr[27041]= 1910985158;
assign addr[27042]= 2030734582;
assign addr[27043]= 2109331059;
assign addr[27044]= 2145181827;
assign addr[27045]= 2137560369;
assign addr[27046]= 2086621133;
assign addr[27047]= 1993396407;
assign addr[27048]= 1859775393;
assign addr[27049]= 1688465931;
assign addr[27050]= 1482939614;
assign addr[27051]= 1247361445;
assign addr[27052]= 986505429;
assign addr[27053]= 705657826;
assign addr[27054]= 410510029;
assign addr[27055]= 107043224;
assign addr[27056]= -198592817;
assign addr[27057]= -500204365;
assign addr[27058]= -791679244;
assign addr[27059]= -1067110699;
assign addr[27060]= -1320917099;
assign addr[27061]= -1547955041;
assign addr[27062]= -1743623590;
assign addr[27063]= -1903957513;
assign addr[27064]= -2025707632;
assign addr[27065]= -2106406677;
assign addr[27066]= -2144419275;
assign addr[27067]= -2138975100;
assign addr[27068]= -2090184478;
assign addr[27069]= -1999036154;
assign addr[27070]= -1867377253;
assign addr[27071]= -1697875851;
assign addr[27072]= -1493966902;
assign addr[27073]= -1259782632;
assign addr[27074]= -1000068799;
assign addr[27075]= -720088517;
assign addr[27076]= -425515602;
assign addr[27077]= -122319591;
assign addr[27078]= 183355234;
assign addr[27079]= 485314355;
assign addr[27080]= 777438554;
assign addr[27081]= 1053807919;
assign addr[27082]= 1308821808;
assign addr[27083]= 1537312353;
assign addr[27084]= 1734649179;
assign addr[27085]= 1896833245;
assign addr[27086]= 2020577882;
assign addr[27087]= 2103375398;
assign addr[27088]= 2143547897;
assign addr[27089]= 2140281282;
assign addr[27090]= 2093641749;
assign addr[27091]= 2004574453;
assign addr[27092]= 1874884346;
assign addr[27093]= 1707199606;
assign addr[27094]= 1504918373;
assign addr[27095]= 1272139887;
assign addr[27096]= 1013581418;
assign addr[27097]= 734482665;
assign addr[27098]= 440499581;
assign addr[27099]= 137589750;
assign addr[27100]= -168108346;
assign addr[27101]= -470399716;
assign addr[27102]= -763158411;
assign addr[27103]= -1040451659;
assign addr[27104]= -1296660098;
assign addr[27105]= -1526591649;
assign addr[27106]= -1725586737;
assign addr[27107]= -1889612716;
assign addr[27108]= -2015345591;
assign addr[27109]= -2100237377;
assign addr[27110]= -2142567738;
assign addr[27111]= -2141478848;
assign addr[27112]= -2096992772;
assign addr[27113]= -2010011024;
assign addr[27114]= -1882296293;
assign addr[27115]= -1716436725;
assign addr[27116]= -1515793473;
assign addr[27117]= -1284432584;
assign addr[27118]= -1027042599;
assign addr[27119]= -748839539;
assign addr[27120]= -455461206;
assign addr[27121]= -152852926;
assign addr[27122]= 152852926;
assign addr[27123]= 455461206;
assign addr[27124]= 748839539;
assign addr[27125]= 1027042599;
assign addr[27126]= 1284432584;
assign addr[27127]= 1515793473;
assign addr[27128]= 1716436725;
assign addr[27129]= 1882296293;
assign addr[27130]= 2010011024;
assign addr[27131]= 2096992772;
assign addr[27132]= 2141478848;
assign addr[27133]= 2142567738;
assign addr[27134]= 2100237377;
assign addr[27135]= 2015345591;
assign addr[27136]= 1889612716;
assign addr[27137]= 1725586737;
assign addr[27138]= 1526591649;
assign addr[27139]= 1296660098;
assign addr[27140]= 1040451659;
assign addr[27141]= 763158411;
assign addr[27142]= 470399716;
assign addr[27143]= 168108346;
assign addr[27144]= -137589750;
assign addr[27145]= -440499581;
assign addr[27146]= -734482665;
assign addr[27147]= -1013581418;
assign addr[27148]= -1272139887;
assign addr[27149]= -1504918373;
assign addr[27150]= -1707199606;
assign addr[27151]= -1874884346;
assign addr[27152]= -2004574453;
assign addr[27153]= -2093641749;
assign addr[27154]= -2140281282;
assign addr[27155]= -2143547897;
assign addr[27156]= -2103375398;
assign addr[27157]= -2020577882;
assign addr[27158]= -1896833245;
assign addr[27159]= -1734649179;
assign addr[27160]= -1537312353;
assign addr[27161]= -1308821808;
assign addr[27162]= -1053807919;
assign addr[27163]= -777438554;
assign addr[27164]= -485314355;
assign addr[27165]= -183355234;
assign addr[27166]= 122319591;
assign addr[27167]= 425515602;
assign addr[27168]= 720088517;
assign addr[27169]= 1000068799;
assign addr[27170]= 1259782632;
assign addr[27171]= 1493966902;
assign addr[27172]= 1697875851;
assign addr[27173]= 1867377253;
assign addr[27174]= 1999036154;
assign addr[27175]= 2090184478;
assign addr[27176]= 2138975100;
assign addr[27177]= 2144419275;
assign addr[27178]= 2106406677;
assign addr[27179]= 2025707632;
assign addr[27180]= 1903957513;
assign addr[27181]= 1743623590;
assign addr[27182]= 1547955041;
assign addr[27183]= 1320917099;
assign addr[27184]= 1067110699;
assign addr[27185]= 791679244;
assign addr[27186]= 500204365;
assign addr[27187]= 198592817;
assign addr[27188]= -107043224;
assign addr[27189]= -410510029;
assign addr[27190]= -705657826;
assign addr[27191]= -986505429;
assign addr[27192]= -1247361445;
assign addr[27193]= -1482939614;
assign addr[27194]= -1688465931;
assign addr[27195]= -1859775393;
assign addr[27196]= -1993396407;
assign addr[27197]= -2086621133;
assign addr[27198]= -2137560369;
assign addr[27199]= -2145181827;
assign addr[27200]= -2109331059;
assign addr[27201]= -2030734582;
assign addr[27202]= -1910985158;
assign addr[27203]= -1752509516;
assign addr[27204]= -1558519173;
assign addr[27205]= -1332945355;
assign addr[27206]= -1080359326;
assign addr[27207]= -805879757;
assign addr[27208]= -515068990;
assign addr[27209]= -213820322;
assign addr[27210]= 91761426;
assign addr[27211]= 395483624;
assign addr[27212]= 691191324;
assign addr[27213]= 972891995;
assign addr[27214]= 1234876957;
assign addr[27215]= 1471837070;
assign addr[27216]= 1678970324;
assign addr[27217]= 1852079154;
assign addr[27218]= 1987655498;
assign addr[27219]= 2082951896;
assign addr[27220]= 2136037160;
assign addr[27221]= 2145835515;
assign addr[27222]= 2112148396;
assign addr[27223]= 2035658475;
assign addr[27224]= 1917915825;
assign addr[27225]= 1761306505;
assign addr[27226]= 1569004214;
assign addr[27227]= 1344905966;
assign addr[27228]= 1093553126;
assign addr[27229]= 820039373;
assign addr[27230]= 529907477;
assign addr[27231]= 229036977;
assign addr[27232]= -76474970;
assign addr[27233]= -380437148;
assign addr[27234]= -676689746;
assign addr[27235]= -959229189;
assign addr[27236]= -1222329801;
assign addr[27237]= -1460659832;
assign addr[27238]= -1669389513;
assign addr[27239]= -1844288924;
assign addr[27240]= -1981813720;
assign addr[27241]= -2079176953;
assign addr[27242]= -2134405552;
assign addr[27243]= -2146380306;
assign addr[27244]= -2114858546;
assign addr[27245]= -2040479063;
assign addr[27246]= -1924749160;
assign addr[27247]= -1770014111;
assign addr[27248]= -1579409630;
assign addr[27249]= -1356798326;
assign addr[27250]= -1106691431;
assign addr[27251]= -834157373;
assign addr[27252]= -544719071;
assign addr[27253]= -244242007;
assign addr[27254]= 61184634;
assign addr[27255]= 365371365;
assign addr[27256]= 662153826;
assign addr[27257]= 945517704;
assign addr[27258]= 1209720613;
assign addr[27259]= 1449408469;
assign addr[27260]= 1659723983;
assign addr[27261]= 1836405100;
assign addr[27262]= 1975871368;
assign addr[27263]= 2075296495;
assign addr[27264]= 2132665626;
assign addr[27265]= 2146816171;
assign addr[27266]= 2117461370;
assign addr[27267]= 2045196100;
assign addr[27268]= 1931484818;
assign addr[27269]= 1778631892;
assign addr[27270]= 1589734894;
assign addr[27271]= 1368621831;
assign addr[27272]= 1119773573;
assign addr[27273]= 848233042;
assign addr[27274]= 559503022;
assign addr[27275]= 259434643;
assign addr[27276]= -45891193;
assign addr[27277]= -350287041;
assign addr[27278]= -647584304;
assign addr[27279]= -931758235;
assign addr[27280]= -1197050035;
assign addr[27281]= -1438083551;
assign addr[27282]= -1649974225;
assign addr[27283]= -1828428082;
assign addr[27284]= -1969828744;
assign addr[27285]= -2071310720;
assign addr[27286]= -2130817471;
assign addr[27287]= -2147143090;
assign addr[27288]= -2119956737;
assign addr[27289]= -2049809346;
assign addr[27290]= -1938122457;
assign addr[27291]= -1787159411;
assign addr[27292]= -1599979481;
assign addr[27293]= -1380375881;
assign addr[27294]= -1132798888;
assign addr[27295]= -862265664;
assign addr[27296]= -574258580;
assign addr[27297]= -274614114;
assign addr[27298]= 30595422;
assign addr[27299]= 335184940;
assign addr[27300]= 632981917;
assign addr[27301]= 917951481;
assign addr[27302]= 1184318708;
assign addr[27303]= 1426685652;
assign addr[27304]= 1640140734;
assign addr[27305]= 1820358275;
assign addr[27306]= 1963686155;
assign addr[27307]= 2067219829;
assign addr[27308]= 2128861181;
assign addr[27309]= 2147361045;
assign addr[27310]= 2122344521;
assign addr[27311]= 2054318569;
assign addr[27312]= 1944661739;
assign addr[27313]= 1795596234;
assign addr[27314]= 1610142873;
assign addr[27315]= 1392059879;
assign addr[27316]= 1145766716;
assign addr[27317]= 876254528;
assign addr[27318]= 588984994;
assign addr[27319]= 289779648;
assign addr[27320]= -15298099;
assign addr[27321]= -320065829;
assign addr[27322]= -618347408;
assign addr[27323]= -904098143;
assign addr[27324]= -1171527280;
assign addr[27325]= -1415215352;
assign addr[27326]= -1630224009;
assign addr[27327]= -1812196087;
assign addr[27328]= -1957443913;
assign addr[27329]= -2063024031;
assign addr[27330]= -2126796855;
assign addr[27331]= -2147470025;
assign addr[27332]= -2124624598;
assign addr[27333]= -2058723538;
assign addr[27334]= -1951102334;
assign addr[27335]= -1803941934;
assign addr[27336]= -1620224553;
assign addr[27337]= -1403673233;
assign addr[27338]= -1158676398;
assign addr[27339]= -890198924;
assign addr[27340]= -603681519;
assign addr[27341]= -304930476;
assign addr[27342]= 0;
assign addr[27343]= 304930476;
assign addr[27344]= 603681519;
assign addr[27345]= 890198924;
assign addr[27346]= 1158676398;
assign addr[27347]= 1403673233;
assign addr[27348]= 1620224553;
assign addr[27349]= 1803941934;
assign addr[27350]= 1951102334;
assign addr[27351]= 2058723538;
assign addr[27352]= 2124624598;
assign addr[27353]= 2147470025;
assign addr[27354]= 2126796855;
assign addr[27355]= 2063024031;
assign addr[27356]= 1957443913;
assign addr[27357]= 1812196087;
assign addr[27358]= 1630224009;
assign addr[27359]= 1415215352;
assign addr[27360]= 1171527280;
assign addr[27361]= 904098143;
assign addr[27362]= 618347408;
assign addr[27363]= 320065829;
assign addr[27364]= 15298099;
assign addr[27365]= -289779648;
assign addr[27366]= -588984994;
assign addr[27367]= -876254528;
assign addr[27368]= -1145766716;
assign addr[27369]= -1392059879;
assign addr[27370]= -1610142873;
assign addr[27371]= -1795596234;
assign addr[27372]= -1944661739;
assign addr[27373]= -2054318569;
assign addr[27374]= -2122344521;
assign addr[27375]= -2147361045;
assign addr[27376]= -2128861181;
assign addr[27377]= -2067219829;
assign addr[27378]= -1963686155;
assign addr[27379]= -1820358275;
assign addr[27380]= -1640140734;
assign addr[27381]= -1426685652;
assign addr[27382]= -1184318708;
assign addr[27383]= -917951481;
assign addr[27384]= -632981917;
assign addr[27385]= -335184940;
assign addr[27386]= -30595422;
assign addr[27387]= 274614114;
assign addr[27388]= 574258580;
assign addr[27389]= 862265664;
assign addr[27390]= 1132798888;
assign addr[27391]= 1380375881;
assign addr[27392]= 1599979481;
assign addr[27393]= 1787159411;
assign addr[27394]= 1938122457;
assign addr[27395]= 2049809346;
assign addr[27396]= 2119956737;
assign addr[27397]= 2147143090;
assign addr[27398]= 2130817471;
assign addr[27399]= 2071310720;
assign addr[27400]= 1969828744;
assign addr[27401]= 1828428082;
assign addr[27402]= 1649974225;
assign addr[27403]= 1438083551;
assign addr[27404]= 1197050035;
assign addr[27405]= 931758235;
assign addr[27406]= 647584304;
assign addr[27407]= 350287041;
assign addr[27408]= 45891193;
assign addr[27409]= -259434643;
assign addr[27410]= -559503022;
assign addr[27411]= -848233042;
assign addr[27412]= -1119773573;
assign addr[27413]= -1368621831;
assign addr[27414]= -1589734894;
assign addr[27415]= -1778631892;
assign addr[27416]= -1931484818;
assign addr[27417]= -2045196100;
assign addr[27418]= -2117461370;
assign addr[27419]= -2146816171;
assign addr[27420]= -2132665626;
assign addr[27421]= -2075296495;
assign addr[27422]= -1975871368;
assign addr[27423]= -1836405100;
assign addr[27424]= -1659723983;
assign addr[27425]= -1449408469;
assign addr[27426]= -1209720613;
assign addr[27427]= -945517704;
assign addr[27428]= -662153826;
assign addr[27429]= -365371365;
assign addr[27430]= -61184634;
assign addr[27431]= 244242007;
assign addr[27432]= 544719071;
assign addr[27433]= 834157373;
assign addr[27434]= 1106691431;
assign addr[27435]= 1356798326;
assign addr[27436]= 1579409630;
assign addr[27437]= 1770014111;
assign addr[27438]= 1924749160;
assign addr[27439]= 2040479063;
assign addr[27440]= 2114858546;
assign addr[27441]= 2146380306;
assign addr[27442]= 2134405552;
assign addr[27443]= 2079176953;
assign addr[27444]= 1981813720;
assign addr[27445]= 1844288924;
assign addr[27446]= 1669389513;
assign addr[27447]= 1460659832;
assign addr[27448]= 1222329801;
assign addr[27449]= 959229189;
assign addr[27450]= 676689746;
assign addr[27451]= 380437148;
assign addr[27452]= 76474970;
assign addr[27453]= -229036977;
assign addr[27454]= -529907477;
assign addr[27455]= -820039373;
assign addr[27456]= -1093553126;
assign addr[27457]= -1344905966;
assign addr[27458]= -1569004214;
assign addr[27459]= -1761306505;
assign addr[27460]= -1917915825;
assign addr[27461]= -2035658475;
assign addr[27462]= -2112148396;
assign addr[27463]= -2145835515;
assign addr[27464]= -2136037160;
assign addr[27465]= -2082951896;
assign addr[27466]= -1987655498;
assign addr[27467]= -1852079154;
assign addr[27468]= -1678970324;
assign addr[27469]= -1471837070;
assign addr[27470]= -1234876957;
assign addr[27471]= -972891995;
assign addr[27472]= -691191324;
assign addr[27473]= -395483624;
assign addr[27474]= -91761426;
assign addr[27475]= 213820322;
assign addr[27476]= 515068990;
assign addr[27477]= 805879757;
assign addr[27478]= 1080359326;
assign addr[27479]= 1332945355;
assign addr[27480]= 1558519173;
assign addr[27481]= 1752509516;
assign addr[27482]= 1910985158;
assign addr[27483]= 2030734582;
assign addr[27484]= 2109331059;
assign addr[27485]= 2145181827;
assign addr[27486]= 2137560369;
assign addr[27487]= 2086621133;
assign addr[27488]= 1993396407;
assign addr[27489]= 1859775393;
assign addr[27490]= 1688465931;
assign addr[27491]= 1482939614;
assign addr[27492]= 1247361445;
assign addr[27493]= 986505429;
assign addr[27494]= 705657826;
assign addr[27495]= 410510029;
assign addr[27496]= 107043224;
assign addr[27497]= -198592817;
assign addr[27498]= -500204365;
assign addr[27499]= -791679244;
assign addr[27500]= -1067110699;
assign addr[27501]= -1320917099;
assign addr[27502]= -1547955041;
assign addr[27503]= -1743623590;
assign addr[27504]= -1903957513;
assign addr[27505]= -2025707632;
assign addr[27506]= -2106406677;
assign addr[27507]= -2144419275;
assign addr[27508]= -2138975100;
assign addr[27509]= -2090184478;
assign addr[27510]= -1999036154;
assign addr[27511]= -1867377253;
assign addr[27512]= -1697875851;
assign addr[27513]= -1493966902;
assign addr[27514]= -1259782632;
assign addr[27515]= -1000068799;
assign addr[27516]= -720088517;
assign addr[27517]= -425515602;
assign addr[27518]= -122319591;
assign addr[27519]= 183355234;
assign addr[27520]= 485314355;
assign addr[27521]= 777438554;
assign addr[27522]= 1053807919;
assign addr[27523]= 1308821808;
assign addr[27524]= 1537312353;
assign addr[27525]= 1734649179;
assign addr[27526]= 1896833245;
assign addr[27527]= 2020577882;
assign addr[27528]= 2103375398;
assign addr[27529]= 2143547897;
assign addr[27530]= 2140281282;
assign addr[27531]= 2093641749;
assign addr[27532]= 2004574453;
assign addr[27533]= 1874884346;
assign addr[27534]= 1707199606;
assign addr[27535]= 1504918373;
assign addr[27536]= 1272139887;
assign addr[27537]= 1013581418;
assign addr[27538]= 734482665;
assign addr[27539]= 440499581;
assign addr[27540]= 137589750;
assign addr[27541]= -168108346;
assign addr[27542]= -470399716;
assign addr[27543]= -763158411;
assign addr[27544]= -1040451659;
assign addr[27545]= -1296660098;
assign addr[27546]= -1526591649;
assign addr[27547]= -1725586737;
assign addr[27548]= -1889612716;
assign addr[27549]= -2015345591;
assign addr[27550]= -2100237377;
assign addr[27551]= -2142567738;
assign addr[27552]= -2141478848;
assign addr[27553]= -2096992772;
assign addr[27554]= -2010011024;
assign addr[27555]= -1882296293;
assign addr[27556]= -1716436725;
assign addr[27557]= -1515793473;
assign addr[27558]= -1284432584;
assign addr[27559]= -1027042599;
assign addr[27560]= -748839539;
assign addr[27561]= -455461206;
assign addr[27562]= -152852926;
assign addr[27563]= 152852926;
assign addr[27564]= 455461206;
assign addr[27565]= 748839539;
assign addr[27566]= 1027042599;
assign addr[27567]= 1284432584;
assign addr[27568]= 1515793473;
assign addr[27569]= 1716436725;
assign addr[27570]= 1882296293;
assign addr[27571]= 2010011024;
assign addr[27572]= 2096992772;
assign addr[27573]= 2141478848;
assign addr[27574]= 2142567738;
assign addr[27575]= 2100237377;
assign addr[27576]= 2015345591;
assign addr[27577]= 1889612716;
assign addr[27578]= 1725586737;
assign addr[27579]= 1526591649;
assign addr[27580]= 1296660098;
assign addr[27581]= 1040451659;
assign addr[27582]= 763158411;
assign addr[27583]= 470399716;
assign addr[27584]= 168108346;
assign addr[27585]= -137589750;
assign addr[27586]= -440499581;
assign addr[27587]= -734482665;
assign addr[27588]= -1013581418;
assign addr[27589]= -1272139887;
assign addr[27590]= -1504918373;
assign addr[27591]= -1707199606;
assign addr[27592]= -1874884346;
assign addr[27593]= -2004574453;
assign addr[27594]= -2093641749;
assign addr[27595]= -2140281282;
assign addr[27596]= -2143547897;
assign addr[27597]= -2103375398;
assign addr[27598]= -2020577882;
assign addr[27599]= -1896833245;
assign addr[27600]= -1734649179;
assign addr[27601]= -1537312353;
assign addr[27602]= -1308821808;
assign addr[27603]= -1053807919;
assign addr[27604]= -777438554;
assign addr[27605]= -485314355;
assign addr[27606]= -183355234;
assign addr[27607]= 122319591;
assign addr[27608]= 425515602;
assign addr[27609]= 720088517;
assign addr[27610]= 1000068799;
assign addr[27611]= 1259782632;
assign addr[27612]= 1493966902;
assign addr[27613]= 1697875851;
assign addr[27614]= 1867377253;
assign addr[27615]= 1999036154;
assign addr[27616]= 2090184478;
assign addr[27617]= 2138975100;
assign addr[27618]= 2144419275;
assign addr[27619]= 2106406677;
assign addr[27620]= 2025707632;
assign addr[27621]= 1903957513;
assign addr[27622]= 1743623590;
assign addr[27623]= 1547955041;
assign addr[27624]= 1320917099;
assign addr[27625]= 1067110699;
assign addr[27626]= 791679244;
assign addr[27627]= 500204365;
assign addr[27628]= 198592817;
assign addr[27629]= -107043224;
assign addr[27630]= -410510029;
assign addr[27631]= -705657826;
assign addr[27632]= -986505429;
assign addr[27633]= -1247361445;
assign addr[27634]= -1482939614;
assign addr[27635]= -1688465931;
assign addr[27636]= -1859775393;
assign addr[27637]= -1993396407;
assign addr[27638]= -2086621133;
assign addr[27639]= -2137560369;
assign addr[27640]= -2145181827;
assign addr[27641]= -2109331059;
assign addr[27642]= -2030734582;
assign addr[27643]= -1910985158;
assign addr[27644]= -1752509516;
assign addr[27645]= -1558519173;
assign addr[27646]= -1332945355;
assign addr[27647]= -1080359326;
assign addr[27648]= -805879757;
assign addr[27649]= -515068990;
assign addr[27650]= -213820322;
assign addr[27651]= 91761426;
assign addr[27652]= 395483624;
assign addr[27653]= 691191324;
assign addr[27654]= 972891995;
assign addr[27655]= 1234876957;
assign addr[27656]= 1471837070;
assign addr[27657]= 1678970324;
assign addr[27658]= 1852079154;
assign addr[27659]= 1987655498;
assign addr[27660]= 2082951896;
assign addr[27661]= 2136037160;
assign addr[27662]= 2145835515;
assign addr[27663]= 2112148396;
assign addr[27664]= 2035658475;
assign addr[27665]= 1917915825;
assign addr[27666]= 1761306505;
assign addr[27667]= 1569004214;
assign addr[27668]= 1344905966;
assign addr[27669]= 1093553126;
assign addr[27670]= 820039373;
assign addr[27671]= 529907477;
assign addr[27672]= 229036977;
assign addr[27673]= -76474970;
assign addr[27674]= -380437148;
assign addr[27675]= -676689746;
assign addr[27676]= -959229189;
assign addr[27677]= -1222329801;
assign addr[27678]= -1460659832;
assign addr[27679]= -1669389513;
assign addr[27680]= -1844288924;
assign addr[27681]= -1981813720;
assign addr[27682]= -2079176953;
assign addr[27683]= -2134405552;
assign addr[27684]= -2146380306;
assign addr[27685]= -2114858546;
assign addr[27686]= -2040479063;
assign addr[27687]= -1924749160;
assign addr[27688]= -1770014111;
assign addr[27689]= -1579409630;
assign addr[27690]= -1356798326;
assign addr[27691]= -1106691431;
assign addr[27692]= -834157373;
assign addr[27693]= -544719071;
assign addr[27694]= -244242007;
assign addr[27695]= 61184634;
assign addr[27696]= 365371365;
assign addr[27697]= 662153826;
assign addr[27698]= 945517704;
assign addr[27699]= 1209720613;
assign addr[27700]= 1449408469;
assign addr[27701]= 1659723983;
assign addr[27702]= 1836405100;
assign addr[27703]= 1975871368;
assign addr[27704]= 2075296495;
assign addr[27705]= 2132665626;
assign addr[27706]= 2146816171;
assign addr[27707]= 2117461370;
assign addr[27708]= 2045196100;
assign addr[27709]= 1931484818;
assign addr[27710]= 1778631892;
assign addr[27711]= 1589734894;
assign addr[27712]= 1368621831;
assign addr[27713]= 1119773573;
assign addr[27714]= 848233042;
assign addr[27715]= 559503022;
assign addr[27716]= 259434643;
assign addr[27717]= -45891193;
assign addr[27718]= -350287041;
assign addr[27719]= -647584304;
assign addr[27720]= -931758235;
assign addr[27721]= -1197050035;
assign addr[27722]= -1438083551;
assign addr[27723]= -1649974225;
assign addr[27724]= -1828428082;
assign addr[27725]= -1969828744;
assign addr[27726]= -2071310720;
assign addr[27727]= -2130817471;
assign addr[27728]= -2147143090;
assign addr[27729]= -2119956737;
assign addr[27730]= -2049809346;
assign addr[27731]= -1938122457;
assign addr[27732]= -1787159411;
assign addr[27733]= -1599979481;
assign addr[27734]= -1380375881;
assign addr[27735]= -1132798888;
assign addr[27736]= -862265664;
assign addr[27737]= -574258580;
assign addr[27738]= -274614114;
assign addr[27739]= 30595422;
assign addr[27740]= 335184940;
assign addr[27741]= 632981917;
assign addr[27742]= 917951481;
assign addr[27743]= 1184318708;
assign addr[27744]= 1426685652;
assign addr[27745]= 1640140734;
assign addr[27746]= 1820358275;
assign addr[27747]= 1963686155;
assign addr[27748]= 2067219829;
assign addr[27749]= 2128861181;
assign addr[27750]= 2147361045;
assign addr[27751]= 2122344521;
assign addr[27752]= 2054318569;
assign addr[27753]= 1944661739;
assign addr[27754]= 1795596234;
assign addr[27755]= 1610142873;
assign addr[27756]= 1392059879;
assign addr[27757]= 1145766716;
assign addr[27758]= 876254528;
assign addr[27759]= 588984994;
assign addr[27760]= 289779648;
assign addr[27761]= -15298099;
assign addr[27762]= -320065829;
assign addr[27763]= -618347408;
assign addr[27764]= -904098143;
assign addr[27765]= -1171527280;
assign addr[27766]= -1415215352;
assign addr[27767]= -1630224009;
assign addr[27768]= -1812196087;
assign addr[27769]= -1957443913;
assign addr[27770]= -2063024031;
assign addr[27771]= -2126796855;
assign addr[27772]= -2147470025;
assign addr[27773]= -2124624598;
assign addr[27774]= -2058723538;
assign addr[27775]= -1951102334;
assign addr[27776]= -1803941934;
assign addr[27777]= -1620224553;
assign addr[27778]= -1403673233;
assign addr[27779]= -1158676398;
assign addr[27780]= -890198924;
assign addr[27781]= -603681519;
assign addr[27782]= -304930476;
assign addr[27783]= 0;
assign addr[27784]= 304930476;
assign addr[27785]= 603681519;
assign addr[27786]= 890198924;
assign addr[27787]= 1158676398;
assign addr[27788]= 1403673233;
assign addr[27789]= 1620224553;
assign addr[27790]= 1803941934;
assign addr[27791]= 1951102334;
assign addr[27792]= 2058723538;
assign addr[27793]= 2124624598;
assign addr[27794]= 2147470025;
assign addr[27795]= 2126796855;
assign addr[27796]= 2063024031;
assign addr[27797]= 1957443913;
assign addr[27798]= 1812196087;
assign addr[27799]= 1630224009;
assign addr[27800]= 1415215352;
assign addr[27801]= 1171527280;
assign addr[27802]= 904098143;
assign addr[27803]= 618347408;
assign addr[27804]= 320065829;
assign addr[27805]= 15298099;
assign addr[27806]= -289779648;
assign addr[27807]= -588984994;
assign addr[27808]= -876254528;
assign addr[27809]= -1145766716;
assign addr[27810]= -1392059879;
assign addr[27811]= -1610142873;
assign addr[27812]= -1795596234;
assign addr[27813]= -1944661739;
assign addr[27814]= -2054318569;
assign addr[27815]= -2122344521;
assign addr[27816]= -2147361045;
assign addr[27817]= -2128861181;
assign addr[27818]= -2067219829;
assign addr[27819]= -1963686155;
assign addr[27820]= -1820358275;
assign addr[27821]= -1640140734;
assign addr[27822]= -1426685652;
assign addr[27823]= -1184318708;
assign addr[27824]= -917951481;
assign addr[27825]= -632981917;
assign addr[27826]= -335184940;
assign addr[27827]= -30595422;
assign addr[27828]= 274614114;
assign addr[27829]= 574258580;
assign addr[27830]= 862265664;
assign addr[27831]= 1132798888;
assign addr[27832]= 1380375881;
assign addr[27833]= 1599979481;
assign addr[27834]= 1787159411;
assign addr[27835]= 1938122457;
assign addr[27836]= 2049809346;
assign addr[27837]= 2119956737;
assign addr[27838]= 2147143090;
assign addr[27839]= 2130817471;
assign addr[27840]= 2071310720;
assign addr[27841]= 1969828744;
assign addr[27842]= 1828428082;
assign addr[27843]= 1649974225;
assign addr[27844]= 1438083551;
assign addr[27845]= 1197050035;
assign addr[27846]= 931758235;
assign addr[27847]= 647584304;
assign addr[27848]= 350287041;
assign addr[27849]= 45891193;
assign addr[27850]= -259434643;
assign addr[27851]= -559503022;
assign addr[27852]= -848233042;
assign addr[27853]= -1119773573;
assign addr[27854]= -1368621831;
assign addr[27855]= -1589734894;
assign addr[27856]= -1778631892;
assign addr[27857]= -1931484818;
assign addr[27858]= -2045196100;
assign addr[27859]= -2117461370;
assign addr[27860]= -2146816171;
assign addr[27861]= -2132665626;
assign addr[27862]= -2075296495;
assign addr[27863]= -1975871368;
assign addr[27864]= -1836405100;
assign addr[27865]= -1659723983;
assign addr[27866]= -1449408469;
assign addr[27867]= -1209720613;
assign addr[27868]= -945517704;
assign addr[27869]= -662153826;
assign addr[27870]= -365371365;
assign addr[27871]= -61184634;
assign addr[27872]= 244242007;
assign addr[27873]= 544719071;
assign addr[27874]= 834157373;
assign addr[27875]= 1106691431;
assign addr[27876]= 1356798326;
assign addr[27877]= 1579409630;
assign addr[27878]= 1770014111;
assign addr[27879]= 1924749160;
assign addr[27880]= 2040479063;
assign addr[27881]= 2114858546;
assign addr[27882]= 2146380306;
assign addr[27883]= 2134405552;
assign addr[27884]= 2079176953;
assign addr[27885]= 1981813720;
assign addr[27886]= 1844288924;
assign addr[27887]= 1669389513;
assign addr[27888]= 1460659832;
assign addr[27889]= 1222329801;
assign addr[27890]= 959229189;
assign addr[27891]= 676689746;
assign addr[27892]= 380437148;
assign addr[27893]= 76474970;
assign addr[27894]= -229036977;
assign addr[27895]= -529907477;
assign addr[27896]= -820039373;
assign addr[27897]= -1093553126;
assign addr[27898]= -1344905966;
assign addr[27899]= -1569004214;
assign addr[27900]= -1761306505;
assign addr[27901]= -1917915825;
assign addr[27902]= -2035658475;
assign addr[27903]= -2112148396;
assign addr[27904]= -2145835515;
assign addr[27905]= -2136037160;
assign addr[27906]= -2082951896;
assign addr[27907]= -1987655498;
assign addr[27908]= -1852079154;
assign addr[27909]= -1678970324;
assign addr[27910]= -1471837070;
assign addr[27911]= -1234876957;
assign addr[27912]= -972891995;
assign addr[27913]= -691191324;
assign addr[27914]= -395483624;
assign addr[27915]= -91761426;
assign addr[27916]= 213820322;
assign addr[27917]= 515068990;
assign addr[27918]= 805879757;
assign addr[27919]= 1080359326;
assign addr[27920]= 1332945355;
assign addr[27921]= 1558519173;
assign addr[27922]= 1752509516;
assign addr[27923]= 1910985158;
assign addr[27924]= 2030734582;
assign addr[27925]= 2109331059;
assign addr[27926]= 2145181827;
assign addr[27927]= 2137560369;
assign addr[27928]= 2086621133;
assign addr[27929]= 1993396407;
assign addr[27930]= 1859775393;
assign addr[27931]= 1688465931;
assign addr[27932]= 1482939614;
assign addr[27933]= 1247361445;
assign addr[27934]= 986505429;
assign addr[27935]= 705657826;
assign addr[27936]= 410510029;
assign addr[27937]= 107043224;
assign addr[27938]= -198592817;
assign addr[27939]= -500204365;
assign addr[27940]= -791679244;
assign addr[27941]= -1067110699;
assign addr[27942]= -1320917099;
assign addr[27943]= -1547955041;
assign addr[27944]= -1743623590;
assign addr[27945]= -1903957513;
assign addr[27946]= -2025707632;
assign addr[27947]= -2106406677;
assign addr[27948]= -2144419275;
assign addr[27949]= -2138975100;
assign addr[27950]= -2090184478;
assign addr[27951]= -1999036154;
assign addr[27952]= -1867377253;
assign addr[27953]= -1697875851;
assign addr[27954]= -1493966902;
assign addr[27955]= -1259782632;
assign addr[27956]= -1000068799;
assign addr[27957]= -720088517;
assign addr[27958]= -425515602;
assign addr[27959]= -122319591;
assign addr[27960]= 183355234;
assign addr[27961]= 485314355;
assign addr[27962]= 777438554;
assign addr[27963]= 1053807919;
assign addr[27964]= 1308821808;
assign addr[27965]= 1537312353;
assign addr[27966]= 1734649179;
assign addr[27967]= 1896833245;
assign addr[27968]= 2020577882;
assign addr[27969]= 2103375398;
assign addr[27970]= 2143547897;
assign addr[27971]= 2140281282;
assign addr[27972]= 2093641749;
assign addr[27973]= 2004574453;
assign addr[27974]= 1874884346;
assign addr[27975]= 1707199606;
assign addr[27976]= 1504918373;
assign addr[27977]= 1272139887;
assign addr[27978]= 1013581418;
assign addr[27979]= 734482665;
assign addr[27980]= 440499581;
assign addr[27981]= 137589750;
assign addr[27982]= -168108346;
assign addr[27983]= -470399716;
assign addr[27984]= -763158411;
assign addr[27985]= -1040451659;
assign addr[27986]= -1296660098;
assign addr[27987]= -1526591649;
assign addr[27988]= -1725586737;
assign addr[27989]= -1889612716;
assign addr[27990]= -2015345591;
assign addr[27991]= -2100237377;
assign addr[27992]= -2142567738;
assign addr[27993]= -2141478848;
assign addr[27994]= -2096992772;
assign addr[27995]= -2010011024;
assign addr[27996]= -1882296293;
assign addr[27997]= -1716436725;
assign addr[27998]= -1515793473;
assign addr[27999]= -1284432584;
assign addr[28000]= -1027042599;
assign addr[28001]= -748839539;
assign addr[28002]= -455461206;
assign addr[28003]= -152852926;
assign addr[28004]= 152852926;
assign addr[28005]= 455461206;
assign addr[28006]= 748839539;
assign addr[28007]= 1027042599;
assign addr[28008]= 1284432584;
assign addr[28009]= 1515793473;
assign addr[28010]= 1716436725;
assign addr[28011]= 1882296293;
assign addr[28012]= 2010011024;
assign addr[28013]= 2096992772;
assign addr[28014]= 2141478848;
assign addr[28015]= 2142567738;
assign addr[28016]= 2100237377;
assign addr[28017]= 2015345591;
assign addr[28018]= 1889612716;
assign addr[28019]= 1725586737;
assign addr[28020]= 1526591649;
assign addr[28021]= 1296660098;
assign addr[28022]= 1040451659;
assign addr[28023]= 763158411;
assign addr[28024]= 470399716;
assign addr[28025]= 168108346;
assign addr[28026]= -137589750;
assign addr[28027]= -440499581;
assign addr[28028]= -734482665;
assign addr[28029]= -1013581418;
assign addr[28030]= -1272139887;
assign addr[28031]= -1504918373;
assign addr[28032]= -1707199606;
assign addr[28033]= -1874884346;
assign addr[28034]= -2004574453;
assign addr[28035]= -2093641749;
assign addr[28036]= -2140281282;
assign addr[28037]= -2143547897;
assign addr[28038]= -2103375398;
assign addr[28039]= -2020577882;
assign addr[28040]= -1896833245;
assign addr[28041]= -1734649179;
assign addr[28042]= -1537312353;
assign addr[28043]= -1308821808;
assign addr[28044]= -1053807919;
assign addr[28045]= -777438554;
assign addr[28046]= -485314355;
assign addr[28047]= -183355234;
assign addr[28048]= 122319591;
assign addr[28049]= 425515602;
assign addr[28050]= 720088517;
assign addr[28051]= 1000068799;
assign addr[28052]= 1259782632;
assign addr[28053]= 1493966902;
assign addr[28054]= 1697875851;
assign addr[28055]= 1867377253;
assign addr[28056]= 1999036154;
assign addr[28057]= 2090184478;
assign addr[28058]= 2138975100;
assign addr[28059]= 2144419275;
assign addr[28060]= 2106406677;
assign addr[28061]= 2025707632;
assign addr[28062]= 1903957513;
assign addr[28063]= 1743623590;
assign addr[28064]= 1547955041;
assign addr[28065]= 1320917099;
assign addr[28066]= 1067110699;
assign addr[28067]= 791679244;
assign addr[28068]= 500204365;
assign addr[28069]= 198592817;
assign addr[28070]= -107043224;
assign addr[28071]= -410510029;
assign addr[28072]= -705657826;
assign addr[28073]= -986505429;
assign addr[28074]= -1247361445;
assign addr[28075]= -1482939614;
assign addr[28076]= -1688465931;
assign addr[28077]= -1859775393;
assign addr[28078]= -1993396407;
assign addr[28079]= -2086621133;
assign addr[28080]= -2137560369;
assign addr[28081]= -2145181827;
assign addr[28082]= -2109331059;
assign addr[28083]= -2030734582;
assign addr[28084]= -1910985158;
assign addr[28085]= -1752509516;
assign addr[28086]= -1558519173;
assign addr[28087]= -1332945355;
assign addr[28088]= -1080359326;
assign addr[28089]= -805879757;
assign addr[28090]= -515068990;
assign addr[28091]= -213820322;
assign addr[28092]= 91761426;
assign addr[28093]= 395483624;
assign addr[28094]= 691191324;
assign addr[28095]= 972891995;
assign addr[28096]= 1234876957;
assign addr[28097]= 1471837070;
assign addr[28098]= 1678970324;
assign addr[28099]= 1852079154;
assign addr[28100]= 1987655498;
assign addr[28101]= 2082951896;
assign addr[28102]= 2136037160;
assign addr[28103]= 2145835515;
assign addr[28104]= 2112148396;
assign addr[28105]= 2035658475;
assign addr[28106]= 1917915825;
assign addr[28107]= 1761306505;
assign addr[28108]= 1569004214;
assign addr[28109]= 1344905966;
assign addr[28110]= 1093553126;
assign addr[28111]= 820039373;
assign addr[28112]= 529907477;
assign addr[28113]= 229036977;
assign addr[28114]= -76474970;
assign addr[28115]= -380437148;
assign addr[28116]= -676689746;
assign addr[28117]= -959229189;
assign addr[28118]= -1222329801;
assign addr[28119]= -1460659832;
assign addr[28120]= -1669389513;
assign addr[28121]= -1844288924;
assign addr[28122]= -1981813720;
assign addr[28123]= -2079176953;
assign addr[28124]= -2134405552;
assign addr[28125]= -2146380306;
assign addr[28126]= -2114858546;
assign addr[28127]= -2040479063;
assign addr[28128]= -1924749160;
assign addr[28129]= -1770014111;
assign addr[28130]= -1579409630;
assign addr[28131]= -1356798326;
assign addr[28132]= -1106691431;
assign addr[28133]= -834157373;
assign addr[28134]= -544719071;
assign addr[28135]= -244242007;
assign addr[28136]= 61184634;
assign addr[28137]= 365371365;
assign addr[28138]= 662153826;
assign addr[28139]= 945517704;
assign addr[28140]= 1209720613;
assign addr[28141]= 1449408469;
assign addr[28142]= 1659723983;
assign addr[28143]= 1836405100;
assign addr[28144]= 1975871368;
assign addr[28145]= 2075296495;
assign addr[28146]= 2132665626;
assign addr[28147]= 2146816171;
assign addr[28148]= 2117461370;
assign addr[28149]= 2045196100;
assign addr[28150]= 1931484818;
assign addr[28151]= 1778631892;
assign addr[28152]= 1589734894;
assign addr[28153]= 1368621831;
assign addr[28154]= 1119773573;
assign addr[28155]= 848233042;
assign addr[28156]= 559503022;
assign addr[28157]= 259434643;
assign addr[28158]= -45891193;
assign addr[28159]= -350287041;
assign addr[28160]= -647584304;
assign addr[28161]= -931758235;
assign addr[28162]= -1197050035;
assign addr[28163]= -1438083551;
assign addr[28164]= -1649974225;
assign addr[28165]= -1828428082;
assign addr[28166]= -1969828744;
assign addr[28167]= -2071310720;
assign addr[28168]= -2130817471;
assign addr[28169]= -2147143090;
assign addr[28170]= -2119956737;
assign addr[28171]= -2049809346;
assign addr[28172]= -1938122457;
assign addr[28173]= -1787159411;
assign addr[28174]= -1599979481;
assign addr[28175]= -1380375881;
assign addr[28176]= -1132798888;
assign addr[28177]= -862265664;
assign addr[28178]= -574258580;
assign addr[28179]= -274614114;
assign addr[28180]= 30595422;
assign addr[28181]= 335184940;
assign addr[28182]= 632981917;
assign addr[28183]= 917951481;
assign addr[28184]= 1184318708;
assign addr[28185]= 1426685652;
assign addr[28186]= 1640140734;
assign addr[28187]= 1820358275;
assign addr[28188]= 1963686155;
assign addr[28189]= 2067219829;
assign addr[28190]= 2128861181;
assign addr[28191]= 2147361045;
assign addr[28192]= 2122344521;
assign addr[28193]= 2054318569;
assign addr[28194]= 1944661739;
assign addr[28195]= 1795596234;
assign addr[28196]= 1610142873;
assign addr[28197]= 1392059879;
assign addr[28198]= 1145766716;
assign addr[28199]= 876254528;
assign addr[28200]= 588984994;
assign addr[28201]= 289779648;
assign addr[28202]= -15298099;
assign addr[28203]= -320065829;
assign addr[28204]= -618347408;
assign addr[28205]= -904098143;
assign addr[28206]= -1171527280;
assign addr[28207]= -1415215352;
assign addr[28208]= -1630224009;
assign addr[28209]= -1812196087;
assign addr[28210]= -1957443913;
assign addr[28211]= -2063024031;
assign addr[28212]= -2126796855;
assign addr[28213]= -2147470025;
assign addr[28214]= -2124624598;
assign addr[28215]= -2058723538;
assign addr[28216]= -1951102334;
assign addr[28217]= -1803941934;
assign addr[28218]= -1620224553;
assign addr[28219]= -1403673233;
assign addr[28220]= -1158676398;
assign addr[28221]= -890198924;
assign addr[28222]= -603681519;
assign addr[28223]= -304930476;
assign addr[28224]= 0;
assign addr[28225]= 304930476;
assign addr[28226]= 603681519;
assign addr[28227]= 890198924;
assign addr[28228]= 1158676398;
assign addr[28229]= 1403673233;
assign addr[28230]= 1620224553;
assign addr[28231]= 1803941934;
assign addr[28232]= 1951102334;
assign addr[28233]= 2058723538;
assign addr[28234]= 2124624598;
assign addr[28235]= 2147470025;
assign addr[28236]= 2126796855;
assign addr[28237]= 2063024031;
assign addr[28238]= 1957443913;
assign addr[28239]= 1812196087;
assign addr[28240]= 1630224009;
assign addr[28241]= 1415215352;
assign addr[28242]= 1171527280;
assign addr[28243]= 904098143;
assign addr[28244]= 618347408;
assign addr[28245]= 320065829;
assign addr[28246]= 15298099;
assign addr[28247]= -289779648;
assign addr[28248]= -588984994;
assign addr[28249]= -876254528;
assign addr[28250]= -1145766716;
assign addr[28251]= -1392059879;
assign addr[28252]= -1610142873;
assign addr[28253]= -1795596234;
assign addr[28254]= -1944661739;
assign addr[28255]= -2054318569;
assign addr[28256]= -2122344521;
assign addr[28257]= -2147361045;
assign addr[28258]= -2128861181;
assign addr[28259]= -2067219829;
assign addr[28260]= -1963686155;
assign addr[28261]= -1820358275;
assign addr[28262]= -1640140734;
assign addr[28263]= -1426685652;
assign addr[28264]= -1184318708;
assign addr[28265]= -917951481;
assign addr[28266]= -632981917;
assign addr[28267]= -335184940;
assign addr[28268]= -30595422;
assign addr[28269]= 274614114;
assign addr[28270]= 574258580;
assign addr[28271]= 862265664;
assign addr[28272]= 1132798888;
assign addr[28273]= 1380375881;
assign addr[28274]= 1599979481;
assign addr[28275]= 1787159411;
assign addr[28276]= 1938122457;
assign addr[28277]= 2049809346;
assign addr[28278]= 2119956737;
assign addr[28279]= 2147143090;
assign addr[28280]= 2130817471;
assign addr[28281]= 2071310720;
assign addr[28282]= 1969828744;
assign addr[28283]= 1828428082;
assign addr[28284]= 1649974225;
assign addr[28285]= 1438083551;
assign addr[28286]= 1197050035;
assign addr[28287]= 931758235;
assign addr[28288]= 647584304;
assign addr[28289]= 350287041;
assign addr[28290]= 45891193;
assign addr[28291]= -259434643;
assign addr[28292]= -559503022;
assign addr[28293]= -848233042;
assign addr[28294]= -1119773573;
assign addr[28295]= -1368621831;
assign addr[28296]= -1589734894;
assign addr[28297]= -1778631892;
assign addr[28298]= -1931484818;
assign addr[28299]= -2045196100;
assign addr[28300]= -2117461370;
assign addr[28301]= -2146816171;
assign addr[28302]= -2132665626;
assign addr[28303]= -2075296495;
assign addr[28304]= -1975871368;
assign addr[28305]= -1836405100;
assign addr[28306]= -1659723983;
assign addr[28307]= -1449408469;
assign addr[28308]= -1209720613;
assign addr[28309]= -945517704;
assign addr[28310]= -662153826;
assign addr[28311]= -365371365;
assign addr[28312]= -61184634;
assign addr[28313]= 244242007;
assign addr[28314]= 544719071;
assign addr[28315]= 834157373;
assign addr[28316]= 1106691431;
assign addr[28317]= 1356798326;
assign addr[28318]= 1579409630;
assign addr[28319]= 1770014111;
assign addr[28320]= 1924749160;
assign addr[28321]= 2040479063;
assign addr[28322]= 2114858546;
assign addr[28323]= 2146380306;
assign addr[28324]= 2134405552;
assign addr[28325]= 2079176953;
assign addr[28326]= 1981813720;
assign addr[28327]= 1844288924;
assign addr[28328]= 1669389513;
assign addr[28329]= 1460659832;
assign addr[28330]= 1222329801;
assign addr[28331]= 959229189;
assign addr[28332]= 676689746;
assign addr[28333]= 380437148;
assign addr[28334]= 76474970;
assign addr[28335]= -229036977;
assign addr[28336]= -529907477;
assign addr[28337]= -820039373;
assign addr[28338]= -1093553126;
assign addr[28339]= -1344905966;
assign addr[28340]= -1569004214;
assign addr[28341]= -1761306505;
assign addr[28342]= -1917915825;
assign addr[28343]= -2035658475;
assign addr[28344]= -2112148396;
assign addr[28345]= -2145835515;
assign addr[28346]= -2136037160;
assign addr[28347]= -2082951896;
assign addr[28348]= -1987655498;
assign addr[28349]= -1852079154;
assign addr[28350]= -1678970324;
assign addr[28351]= -1471837070;
assign addr[28352]= -1234876957;
assign addr[28353]= -972891995;
assign addr[28354]= -691191324;
assign addr[28355]= -395483624;
assign addr[28356]= -91761426;
assign addr[28357]= 213820322;
assign addr[28358]= 515068990;
assign addr[28359]= 805879757;
assign addr[28360]= 1080359326;
assign addr[28361]= 1332945355;
assign addr[28362]= 1558519173;
assign addr[28363]= 1752509516;
assign addr[28364]= 1910985158;
assign addr[28365]= 2030734582;
assign addr[28366]= 2109331059;
assign addr[28367]= 2145181827;
assign addr[28368]= 2137560369;
assign addr[28369]= 2086621133;
assign addr[28370]= 1993396407;
assign addr[28371]= 1859775393;
assign addr[28372]= 1688465931;
assign addr[28373]= 1482939614;
assign addr[28374]= 1247361445;
assign addr[28375]= 986505429;
assign addr[28376]= 705657826;
assign addr[28377]= 410510029;
assign addr[28378]= 107043224;
assign addr[28379]= -198592817;
assign addr[28380]= -500204365;
assign addr[28381]= -791679244;
assign addr[28382]= -1067110699;
assign addr[28383]= -1320917099;
assign addr[28384]= -1547955041;
assign addr[28385]= -1743623590;
assign addr[28386]= -1903957513;
assign addr[28387]= -2025707632;
assign addr[28388]= -2106406677;
assign addr[28389]= -2144419275;
assign addr[28390]= -2138975100;
assign addr[28391]= -2090184478;
assign addr[28392]= -1999036154;
assign addr[28393]= -1867377253;
assign addr[28394]= -1697875851;
assign addr[28395]= -1493966902;
assign addr[28396]= -1259782632;
assign addr[28397]= -1000068799;
assign addr[28398]= -720088517;
assign addr[28399]= -425515602;
assign addr[28400]= -122319591;
assign addr[28401]= 183355234;
assign addr[28402]= 485314355;
assign addr[28403]= 777438554;
assign addr[28404]= 1053807919;
assign addr[28405]= 1308821808;
assign addr[28406]= 1537312353;
assign addr[28407]= 1734649179;
assign addr[28408]= 1896833245;
assign addr[28409]= 2020577882;
assign addr[28410]= 2103375398;
assign addr[28411]= 2143547897;
assign addr[28412]= 2140281282;
assign addr[28413]= 2093641749;
assign addr[28414]= 2004574453;
assign addr[28415]= 1874884346;
assign addr[28416]= 1707199606;
assign addr[28417]= 1504918373;
assign addr[28418]= 1272139887;
assign addr[28419]= 1013581418;
assign addr[28420]= 734482665;
assign addr[28421]= 440499581;
assign addr[28422]= 137589750;
assign addr[28423]= -168108346;
assign addr[28424]= -470399716;
assign addr[28425]= -763158411;
assign addr[28426]= -1040451659;
assign addr[28427]= -1296660098;
assign addr[28428]= -1526591649;
assign addr[28429]= -1725586737;
assign addr[28430]= -1889612716;
assign addr[28431]= -2015345591;
assign addr[28432]= -2100237377;
assign addr[28433]= -2142567738;
assign addr[28434]= -2141478848;
assign addr[28435]= -2096992772;
assign addr[28436]= -2010011024;
assign addr[28437]= -1882296293;
assign addr[28438]= -1716436725;
assign addr[28439]= -1515793473;
assign addr[28440]= -1284432584;
assign addr[28441]= -1027042599;
assign addr[28442]= -748839539;
assign addr[28443]= -455461206;
assign addr[28444]= -152852926;
assign addr[28445]= 152852926;
assign addr[28446]= 455461206;
assign addr[28447]= 748839539;
assign addr[28448]= 1027042599;
assign addr[28449]= 1284432584;
assign addr[28450]= 1515793473;
assign addr[28451]= 1716436725;
assign addr[28452]= 1882296293;
assign addr[28453]= 2010011024;
assign addr[28454]= 2096992772;
assign addr[28455]= 2141478848;
assign addr[28456]= 2142567738;
assign addr[28457]= 2100237377;
assign addr[28458]= 2015345591;
assign addr[28459]= 1889612716;
assign addr[28460]= 1725586737;
assign addr[28461]= 1526591649;
assign addr[28462]= 1296660098;
assign addr[28463]= 1040451659;
assign addr[28464]= 763158411;
assign addr[28465]= 470399716;
assign addr[28466]= 168108346;
assign addr[28467]= -137589750;
assign addr[28468]= -440499581;
assign addr[28469]= -734482665;
assign addr[28470]= -1013581418;
assign addr[28471]= -1272139887;
assign addr[28472]= -1504918373;
assign addr[28473]= -1707199606;
assign addr[28474]= -1874884346;
assign addr[28475]= -2004574453;
assign addr[28476]= -2093641749;
assign addr[28477]= -2140281282;
assign addr[28478]= -2143547897;
assign addr[28479]= -2103375398;
assign addr[28480]= -2020577882;
assign addr[28481]= -1896833245;
assign addr[28482]= -1734649179;
assign addr[28483]= -1537312353;
assign addr[28484]= -1308821808;
assign addr[28485]= -1053807919;
assign addr[28486]= -777438554;
assign addr[28487]= -485314355;
assign addr[28488]= -183355234;
assign addr[28489]= 122319591;
assign addr[28490]= 425515602;
assign addr[28491]= 720088517;
assign addr[28492]= 1000068799;
assign addr[28493]= 1259782632;
assign addr[28494]= 1493966902;
assign addr[28495]= 1697875851;
assign addr[28496]= 1867377253;
assign addr[28497]= 1999036154;
assign addr[28498]= 2090184478;
assign addr[28499]= 2138975100;
assign addr[28500]= 2144419275;
assign addr[28501]= 2106406677;
assign addr[28502]= 2025707632;
assign addr[28503]= 1903957513;
assign addr[28504]= 1743623590;
assign addr[28505]= 1547955041;
assign addr[28506]= 1320917099;
assign addr[28507]= 1067110699;
assign addr[28508]= 791679244;
assign addr[28509]= 500204365;
assign addr[28510]= 198592817;
assign addr[28511]= -107043224;
assign addr[28512]= -410510029;
assign addr[28513]= -705657826;
assign addr[28514]= -986505429;
assign addr[28515]= -1247361445;
assign addr[28516]= -1482939614;
assign addr[28517]= -1688465931;
assign addr[28518]= -1859775393;
assign addr[28519]= -1993396407;
assign addr[28520]= -2086621133;
assign addr[28521]= -2137560369;
assign addr[28522]= -2145181827;
assign addr[28523]= -2109331059;
assign addr[28524]= -2030734582;
assign addr[28525]= -1910985158;
assign addr[28526]= -1752509516;
assign addr[28527]= -1558519173;
assign addr[28528]= -1332945355;
assign addr[28529]= -1080359326;
assign addr[28530]= -805879757;
assign addr[28531]= -515068990;
assign addr[28532]= -213820322;
assign addr[28533]= 91761426;
assign addr[28534]= 395483624;
assign addr[28535]= 691191324;
assign addr[28536]= 972891995;
assign addr[28537]= 1234876957;
assign addr[28538]= 1471837070;
assign addr[28539]= 1678970324;
assign addr[28540]= 1852079154;
assign addr[28541]= 1987655498;
assign addr[28542]= 2082951896;
assign addr[28543]= 2136037160;
assign addr[28544]= 2145835515;
assign addr[28545]= 2112148396;
assign addr[28546]= 2035658475;
assign addr[28547]= 1917915825;
assign addr[28548]= 1761306505;
assign addr[28549]= 1569004214;
assign addr[28550]= 1344905966;
assign addr[28551]= 1093553126;
assign addr[28552]= 820039373;
assign addr[28553]= 529907477;
assign addr[28554]= 229036977;
assign addr[28555]= -76474970;
assign addr[28556]= -380437148;
assign addr[28557]= -676689746;
assign addr[28558]= -959229189;
assign addr[28559]= -1222329801;
assign addr[28560]= -1460659832;
assign addr[28561]= -1669389513;
assign addr[28562]= -1844288924;
assign addr[28563]= -1981813720;
assign addr[28564]= -2079176953;
assign addr[28565]= -2134405552;
assign addr[28566]= -2146380306;
assign addr[28567]= -2114858546;
assign addr[28568]= -2040479063;
assign addr[28569]= -1924749160;
assign addr[28570]= -1770014111;
assign addr[28571]= -1579409630;
assign addr[28572]= -1356798326;
assign addr[28573]= -1106691431;
assign addr[28574]= -834157373;
assign addr[28575]= -544719071;
assign addr[28576]= -244242007;
assign addr[28577]= 61184634;
assign addr[28578]= 365371365;
assign addr[28579]= 662153826;
assign addr[28580]= 945517704;
assign addr[28581]= 1209720613;
assign addr[28582]= 1449408469;
assign addr[28583]= 1659723983;
assign addr[28584]= 1836405100;
assign addr[28585]= 1975871368;
assign addr[28586]= 2075296495;
assign addr[28587]= 2132665626;
assign addr[28588]= 2146816171;
assign addr[28589]= 2117461370;
assign addr[28590]= 2045196100;
assign addr[28591]= 1931484818;
assign addr[28592]= 1778631892;
assign addr[28593]= 1589734894;
assign addr[28594]= 1368621831;
assign addr[28595]= 1119773573;
assign addr[28596]= 848233042;
assign addr[28597]= 559503022;
assign addr[28598]= 259434643;
assign addr[28599]= -45891193;
assign addr[28600]= -350287041;
assign addr[28601]= -647584304;
assign addr[28602]= -931758235;
assign addr[28603]= -1197050035;
assign addr[28604]= -1438083551;
assign addr[28605]= -1649974225;
assign addr[28606]= -1828428082;
assign addr[28607]= -1969828744;
assign addr[28608]= -2071310720;
assign addr[28609]= -2130817471;
assign addr[28610]= -2147143090;
assign addr[28611]= -2119956737;
assign addr[28612]= -2049809346;
assign addr[28613]= -1938122457;
assign addr[28614]= -1787159411;
assign addr[28615]= -1599979481;
assign addr[28616]= -1380375881;
assign addr[28617]= -1132798888;
assign addr[28618]= -862265664;
assign addr[28619]= -574258580;
assign addr[28620]= -274614114;
assign addr[28621]= 30595422;
assign addr[28622]= 335184940;
assign addr[28623]= 632981917;
assign addr[28624]= 917951481;
assign addr[28625]= 1184318708;
assign addr[28626]= 1426685652;
assign addr[28627]= 1640140734;
assign addr[28628]= 1820358275;
assign addr[28629]= 1963686155;
assign addr[28630]= 2067219829;
assign addr[28631]= 2128861181;
assign addr[28632]= 2147361045;
assign addr[28633]= 2122344521;
assign addr[28634]= 2054318569;
assign addr[28635]= 1944661739;
assign addr[28636]= 1795596234;
assign addr[28637]= 1610142873;
assign addr[28638]= 1392059879;
assign addr[28639]= 1145766716;
assign addr[28640]= 876254528;
assign addr[28641]= 588984994;
assign addr[28642]= 289779648;
assign addr[28643]= -15298099;
assign addr[28644]= -320065829;
assign addr[28645]= -618347408;
assign addr[28646]= -904098143;
assign addr[28647]= -1171527280;
assign addr[28648]= -1415215352;
assign addr[28649]= -1630224009;
assign addr[28650]= -1812196087;
assign addr[28651]= -1957443913;
assign addr[28652]= -2063024031;
assign addr[28653]= -2126796855;
assign addr[28654]= -2147470025;
assign addr[28655]= -2124624598;
assign addr[28656]= -2058723538;
assign addr[28657]= -1951102334;
assign addr[28658]= -1803941934;
assign addr[28659]= -1620224553;
assign addr[28660]= -1403673233;
assign addr[28661]= -1158676398;
assign addr[28662]= -890198924;
assign addr[28663]= -603681519;
assign addr[28664]= -304930476;
assign addr[28665]= 0;
assign addr[28666]= 304930476;
assign addr[28667]= 603681519;
assign addr[28668]= 890198924;
assign addr[28669]= 1158676398;
assign addr[28670]= 1403673233;
assign addr[28671]= 1620224553;
assign addr[28672]= 1803941934;
assign addr[28673]= 1951102334;
assign addr[28674]= 2058723538;
assign addr[28675]= 2124624598;
assign addr[28676]= 2147470025;
assign addr[28677]= 2126796855;
assign addr[28678]= 2063024031;
assign addr[28679]= 1957443913;
assign addr[28680]= 1812196087;
assign addr[28681]= 1630224009;
assign addr[28682]= 1415215352;
assign addr[28683]= 1171527280;
assign addr[28684]= 904098143;
assign addr[28685]= 618347408;
assign addr[28686]= 320065829;
assign addr[28687]= 15298099;
assign addr[28688]= -289779648;
assign addr[28689]= -588984994;
assign addr[28690]= -876254528;
assign addr[28691]= -1145766716;
assign addr[28692]= -1392059879;
assign addr[28693]= -1610142873;
assign addr[28694]= -1795596234;
assign addr[28695]= -1944661739;
assign addr[28696]= -2054318569;
assign addr[28697]= -2122344521;
assign addr[28698]= -2147361045;
assign addr[28699]= -2128861181;
assign addr[28700]= -2067219829;
assign addr[28701]= -1963686155;
assign addr[28702]= -1820358275;
assign addr[28703]= -1640140734;
assign addr[28704]= -1426685652;
assign addr[28705]= -1184318708;
assign addr[28706]= -917951481;
assign addr[28707]= -632981917;
assign addr[28708]= -335184940;
assign addr[28709]= -30595422;
assign addr[28710]= 274614114;
assign addr[28711]= 574258580;
assign addr[28712]= 862265664;
assign addr[28713]= 1132798888;
assign addr[28714]= 1380375881;
assign addr[28715]= 1599979481;
assign addr[28716]= 1787159411;
assign addr[28717]= 1938122457;
assign addr[28718]= 2049809346;
assign addr[28719]= 2119956737;
assign addr[28720]= 2147143090;
assign addr[28721]= 2130817471;
assign addr[28722]= 2071310720;
assign addr[28723]= 1969828744;
assign addr[28724]= 1828428082;
assign addr[28725]= 1649974225;
assign addr[28726]= 1438083551;
assign addr[28727]= 1197050035;
assign addr[28728]= 931758235;
assign addr[28729]= 647584304;
assign addr[28730]= 350287041;
assign addr[28731]= 45891193;
assign addr[28732]= -259434643;
assign addr[28733]= -559503022;
assign addr[28734]= -848233042;
assign addr[28735]= -1119773573;
assign addr[28736]= -1368621831;
assign addr[28737]= -1589734894;
assign addr[28738]= -1778631892;
assign addr[28739]= -1931484818;
assign addr[28740]= -2045196100;
assign addr[28741]= -2117461370;
assign addr[28742]= -2146816171;
assign addr[28743]= -2132665626;
assign addr[28744]= -2075296495;
assign addr[28745]= -1975871368;
assign addr[28746]= -1836405100;
assign addr[28747]= -1659723983;
assign addr[28748]= -1449408469;
assign addr[28749]= -1209720613;
assign addr[28750]= -945517704;
assign addr[28751]= -662153826;
assign addr[28752]= -365371365;
assign addr[28753]= -61184634;
assign addr[28754]= 244242007;
assign addr[28755]= 544719071;
assign addr[28756]= 834157373;
assign addr[28757]= 1106691431;
assign addr[28758]= 1356798326;
assign addr[28759]= 1579409630;
assign addr[28760]= 1770014111;
assign addr[28761]= 1924749160;
assign addr[28762]= 2040479063;
assign addr[28763]= 2114858546;
assign addr[28764]= 2146380306;
assign addr[28765]= 2134405552;
assign addr[28766]= 2079176953;
assign addr[28767]= 1981813720;
assign addr[28768]= 1844288924;
assign addr[28769]= 1669389513;
assign addr[28770]= 1460659832;
assign addr[28771]= 1222329801;
assign addr[28772]= 959229189;
assign addr[28773]= 676689746;
assign addr[28774]= 380437148;
assign addr[28775]= 76474970;
assign addr[28776]= -229036977;
assign addr[28777]= -529907477;
assign addr[28778]= -820039373;
assign addr[28779]= -1093553126;
assign addr[28780]= -1344905966;
assign addr[28781]= -1569004214;
assign addr[28782]= -1761306505;
assign addr[28783]= -1917915825;
assign addr[28784]= -2035658475;
assign addr[28785]= -2112148396;
assign addr[28786]= -2145835515;
assign addr[28787]= -2136037160;
assign addr[28788]= -2082951896;
assign addr[28789]= -1987655498;
assign addr[28790]= -1852079154;
assign addr[28791]= -1678970324;
assign addr[28792]= -1471837070;
assign addr[28793]= -1234876957;
assign addr[28794]= -972891995;
assign addr[28795]= -691191324;
assign addr[28796]= -395483624;
assign addr[28797]= -91761426;
assign addr[28798]= 213820322;
assign addr[28799]= 515068990;
assign addr[28800]= 805879757;
assign addr[28801]= 1080359326;
assign addr[28802]= 1332945355;
assign addr[28803]= 1558519173;
assign addr[28804]= 1752509516;
assign addr[28805]= 1910985158;
assign addr[28806]= 2030734582;
assign addr[28807]= 2109331059;
assign addr[28808]= 2145181827;
assign addr[28809]= 2137560369;
assign addr[28810]= 2086621133;
assign addr[28811]= 1993396407;
assign addr[28812]= 1859775393;
assign addr[28813]= 1688465931;
assign addr[28814]= 1482939614;
assign addr[28815]= 1247361445;
assign addr[28816]= 986505429;
assign addr[28817]= 705657826;
assign addr[28818]= 410510029;
assign addr[28819]= 107043224;
assign addr[28820]= -198592817;
assign addr[28821]= -500204365;
assign addr[28822]= -791679244;
assign addr[28823]= -1067110699;
assign addr[28824]= -1320917099;
assign addr[28825]= -1547955041;
assign addr[28826]= -1743623590;
assign addr[28827]= -1903957513;
assign addr[28828]= -2025707632;
assign addr[28829]= -2106406677;
assign addr[28830]= -2144419275;
assign addr[28831]= -2138975100;
assign addr[28832]= -2090184478;
assign addr[28833]= -1999036154;
assign addr[28834]= -1867377253;
assign addr[28835]= -1697875851;
assign addr[28836]= -1493966902;
assign addr[28837]= -1259782632;
assign addr[28838]= -1000068799;
assign addr[28839]= -720088517;
assign addr[28840]= -425515602;
assign addr[28841]= -122319591;
assign addr[28842]= 183355234;
assign addr[28843]= 485314355;
assign addr[28844]= 777438554;
assign addr[28845]= 1053807919;
assign addr[28846]= 1308821808;
assign addr[28847]= 1537312353;
assign addr[28848]= 1734649179;
assign addr[28849]= 1896833245;
assign addr[28850]= 2020577882;
assign addr[28851]= 2103375398;
assign addr[28852]= 2143547897;
assign addr[28853]= 2140281282;
assign addr[28854]= 2093641749;
assign addr[28855]= 2004574453;
assign addr[28856]= 1874884346;
assign addr[28857]= 1707199606;
assign addr[28858]= 1504918373;
assign addr[28859]= 1272139887;
assign addr[28860]= 1013581418;
assign addr[28861]= 734482665;
assign addr[28862]= 440499581;
assign addr[28863]= 137589750;
assign addr[28864]= -168108346;
assign addr[28865]= -470399716;
assign addr[28866]= -763158411;
assign addr[28867]= -1040451659;
assign addr[28868]= -1296660098;
assign addr[28869]= -1526591649;
assign addr[28870]= -1725586737;
assign addr[28871]= -1889612716;
assign addr[28872]= -2015345591;
assign addr[28873]= -2100237377;
assign addr[28874]= -2142567738;
assign addr[28875]= -2141478848;
assign addr[28876]= -2096992772;
assign addr[28877]= -2010011024;
assign addr[28878]= -1882296293;
assign addr[28879]= -1716436725;
assign addr[28880]= -1515793473;
assign addr[28881]= -1284432584;
assign addr[28882]= -1027042599;
assign addr[28883]= -748839539;
assign addr[28884]= -455461206;
assign addr[28885]= -152852926;
assign addr[28886]= 152852926;
assign addr[28887]= 455461206;
assign addr[28888]= 748839539;
assign addr[28889]= 1027042599;
assign addr[28890]= 1284432584;
assign addr[28891]= 1515793473;
assign addr[28892]= 1716436725;
assign addr[28893]= 1882296293;
assign addr[28894]= 2010011024;
assign addr[28895]= 2096992772;
assign addr[28896]= 2141478848;
assign addr[28897]= 2142567738;
assign addr[28898]= 2100237377;
assign addr[28899]= 2015345591;
assign addr[28900]= 1889612716;
assign addr[28901]= 1725586737;
assign addr[28902]= 1526591649;
assign addr[28903]= 1296660098;
assign addr[28904]= 1040451659;
assign addr[28905]= 763158411;
assign addr[28906]= 470399716;
assign addr[28907]= 168108346;
assign addr[28908]= -137589750;
assign addr[28909]= -440499581;
assign addr[28910]= -734482665;
assign addr[28911]= -1013581418;
assign addr[28912]= -1272139887;
assign addr[28913]= -1504918373;
assign addr[28914]= -1707199606;
assign addr[28915]= -1874884346;
assign addr[28916]= -2004574453;
assign addr[28917]= -2093641749;
assign addr[28918]= -2140281282;
assign addr[28919]= -2143547897;
assign addr[28920]= -2103375398;
assign addr[28921]= -2020577882;
assign addr[28922]= -1896833245;
assign addr[28923]= -1734649179;
assign addr[28924]= -1537312353;
assign addr[28925]= -1308821808;
assign addr[28926]= -1053807919;
assign addr[28927]= -777438554;
assign addr[28928]= -485314355;
assign addr[28929]= -183355234;
assign addr[28930]= 122319591;
assign addr[28931]= 425515602;
assign addr[28932]= 720088517;
assign addr[28933]= 1000068799;
assign addr[28934]= 1259782632;
assign addr[28935]= 1493966902;
assign addr[28936]= 1697875851;
assign addr[28937]= 1867377253;
assign addr[28938]= 1999036154;
assign addr[28939]= 2090184478;
assign addr[28940]= 2138975100;
assign addr[28941]= 2144419275;
assign addr[28942]= 2106406677;
assign addr[28943]= 2025707632;
assign addr[28944]= 1903957513;
assign addr[28945]= 1743623590;
assign addr[28946]= 1547955041;
assign addr[28947]= 1320917099;
assign addr[28948]= 1067110699;
assign addr[28949]= 791679244;
assign addr[28950]= 500204365;
assign addr[28951]= 198592817;
assign addr[28952]= -107043224;
assign addr[28953]= -410510029;
assign addr[28954]= -705657826;
assign addr[28955]= -986505429;
assign addr[28956]= -1247361445;
assign addr[28957]= -1482939614;
assign addr[28958]= -1688465931;
assign addr[28959]= -1859775393;
assign addr[28960]= -1993396407;
assign addr[28961]= -2086621133;
assign addr[28962]= -2137560369;
assign addr[28963]= -2145181827;
assign addr[28964]= -2109331059;
assign addr[28965]= -2030734582;
assign addr[28966]= -1910985158;
assign addr[28967]= -1752509516;
assign addr[28968]= -1558519173;
assign addr[28969]= -1332945355;
assign addr[28970]= -1080359326;
assign addr[28971]= -805879757;
assign addr[28972]= -515068990;
assign addr[28973]= -213820322;
assign addr[28974]= 91761426;
assign addr[28975]= 395483624;
assign addr[28976]= 691191324;
assign addr[28977]= 972891995;
assign addr[28978]= 1234876957;
assign addr[28979]= 1471837070;
assign addr[28980]= 1678970324;
assign addr[28981]= 1852079154;
assign addr[28982]= 1987655498;
assign addr[28983]= 2082951896;
assign addr[28984]= 2136037160;
assign addr[28985]= 2145835515;
assign addr[28986]= 2112148396;
assign addr[28987]= 2035658475;
assign addr[28988]= 1917915825;
assign addr[28989]= 1761306505;
assign addr[28990]= 1569004214;
assign addr[28991]= 1344905966;
assign addr[28992]= 1093553126;
assign addr[28993]= 820039373;
assign addr[28994]= 529907477;
assign addr[28995]= 229036977;
assign addr[28996]= -76474970;
assign addr[28997]= -380437148;
assign addr[28998]= -676689746;
assign addr[28999]= -959229189;
assign addr[29000]= -1222329801;
assign addr[29001]= -1460659832;
assign addr[29002]= -1669389513;
assign addr[29003]= -1844288924;
assign addr[29004]= -1981813720;
assign addr[29005]= -2079176953;
assign addr[29006]= -2134405552;
assign addr[29007]= -2146380306;
assign addr[29008]= -2114858546;
assign addr[29009]= -2040479063;
assign addr[29010]= -1924749160;
assign addr[29011]= -1770014111;
assign addr[29012]= -1579409630;
assign addr[29013]= -1356798326;
assign addr[29014]= -1106691431;
assign addr[29015]= -834157373;
assign addr[29016]= -544719071;
assign addr[29017]= -244242007;
assign addr[29018]= 61184634;
assign addr[29019]= 365371365;
assign addr[29020]= 662153826;
assign addr[29021]= 945517704;
assign addr[29022]= 1209720613;
assign addr[29023]= 1449408469;
assign addr[29024]= 1659723983;
assign addr[29025]= 1836405100;
assign addr[29026]= 1975871368;
assign addr[29027]= 2075296495;
assign addr[29028]= 2132665626;
assign addr[29029]= 2146816171;
assign addr[29030]= 2117461370;
assign addr[29031]= 2045196100;
assign addr[29032]= 1931484818;
assign addr[29033]= 1778631892;
assign addr[29034]= 1589734894;
assign addr[29035]= 1368621831;
assign addr[29036]= 1119773573;
assign addr[29037]= 848233042;
assign addr[29038]= 559503022;
assign addr[29039]= 259434643;
assign addr[29040]= -45891193;
assign addr[29041]= -350287041;
assign addr[29042]= -647584304;
assign addr[29043]= -931758235;
assign addr[29044]= -1197050035;
assign addr[29045]= -1438083551;
assign addr[29046]= -1649974225;
assign addr[29047]= -1828428082;
assign addr[29048]= -1969828744;
assign addr[29049]= -2071310720;
assign addr[29050]= -2130817471;
assign addr[29051]= -2147143090;
assign addr[29052]= -2119956737;
assign addr[29053]= -2049809346;
assign addr[29054]= -1938122457;
assign addr[29055]= -1787159411;
assign addr[29056]= -1599979481;
assign addr[29057]= -1380375881;
assign addr[29058]= -1132798888;
assign addr[29059]= -862265664;
assign addr[29060]= -574258580;
assign addr[29061]= -274614114;
assign addr[29062]= 30595422;
assign addr[29063]= 335184940;
assign addr[29064]= 632981917;
assign addr[29065]= 917951481;
assign addr[29066]= 1184318708;
assign addr[29067]= 1426685652;
assign addr[29068]= 1640140734;
assign addr[29069]= 1820358275;
assign addr[29070]= 1963686155;
assign addr[29071]= 2067219829;
assign addr[29072]= 2128861181;
assign addr[29073]= 2147361045;
assign addr[29074]= 2122344521;
assign addr[29075]= 2054318569;
assign addr[29076]= 1944661739;
assign addr[29077]= 1795596234;
assign addr[29078]= 1610142873;
assign addr[29079]= 1392059879;
assign addr[29080]= 1145766716;
assign addr[29081]= 876254528;
assign addr[29082]= 588984994;
assign addr[29083]= 289779648;
assign addr[29084]= -15298099;
assign addr[29085]= -320065829;
assign addr[29086]= -618347408;
assign addr[29087]= -904098143;
assign addr[29088]= -1171527280;
assign addr[29089]= -1415215352;
assign addr[29090]= -1630224009;
assign addr[29091]= -1812196087;
assign addr[29092]= -1957443913;
assign addr[29093]= -2063024031;
assign addr[29094]= -2126796855;
assign addr[29095]= -2147470025;
assign addr[29096]= -2124624598;
assign addr[29097]= -2058723538;
assign addr[29098]= -1951102334;
assign addr[29099]= -1803941934;
assign addr[29100]= -1620224553;
assign addr[29101]= -1403673233;
assign addr[29102]= -1158676398;
assign addr[29103]= -890198924;
assign addr[29104]= -603681519;
assign addr[29105]= -304930476;
assign addr[29106]= 0;
assign addr[29107]= 304930476;
assign addr[29108]= 603681519;
assign addr[29109]= 890198924;
assign addr[29110]= 1158676398;
assign addr[29111]= 1403673233;
assign addr[29112]= 1620224553;
assign addr[29113]= 1803941934;
assign addr[29114]= 1951102334;
assign addr[29115]= 2058723538;
assign addr[29116]= 2124624598;
assign addr[29117]= 2147470025;
assign addr[29118]= 2126796855;
assign addr[29119]= 2063024031;
assign addr[29120]= 1957443913;
assign addr[29121]= 1812196087;
assign addr[29122]= 1630224009;
assign addr[29123]= 1415215352;
assign addr[29124]= 1171527280;
assign addr[29125]= 904098143;
assign addr[29126]= 618347408;
assign addr[29127]= 320065829;
assign addr[29128]= 15298099;
assign addr[29129]= -289779648;
assign addr[29130]= -588984994;
assign addr[29131]= -876254528;
assign addr[29132]= -1145766716;
assign addr[29133]= -1392059879;
assign addr[29134]= -1610142873;
assign addr[29135]= -1795596234;
assign addr[29136]= -1944661739;
assign addr[29137]= -2054318569;
assign addr[29138]= -2122344521;
assign addr[29139]= -2147361045;
assign addr[29140]= -2128861181;
assign addr[29141]= -2067219829;
assign addr[29142]= -1963686155;
assign addr[29143]= -1820358275;
assign addr[29144]= -1640140734;
assign addr[29145]= -1426685652;
assign addr[29146]= -1184318708;
assign addr[29147]= -917951481;
assign addr[29148]= -632981917;
assign addr[29149]= -335184940;
assign addr[29150]= -30595422;
assign addr[29151]= 274614114;
assign addr[29152]= 574258580;
assign addr[29153]= 862265664;
assign addr[29154]= 1132798888;
assign addr[29155]= 1380375881;
assign addr[29156]= 1599979481;
assign addr[29157]= 1787159411;
assign addr[29158]= 1938122457;
assign addr[29159]= 2049809346;
assign addr[29160]= 2119956737;
assign addr[29161]= 2147143090;
assign addr[29162]= 2130817471;
assign addr[29163]= 2071310720;
assign addr[29164]= 1969828744;
assign addr[29165]= 1828428082;
assign addr[29166]= 1649974225;
assign addr[29167]= 1438083551;
assign addr[29168]= 1197050035;
assign addr[29169]= 931758235;
assign addr[29170]= 647584304;
assign addr[29171]= 350287041;
assign addr[29172]= 45891193;
assign addr[29173]= -259434643;
assign addr[29174]= -559503022;
assign addr[29175]= -848233042;
assign addr[29176]= -1119773573;
assign addr[29177]= -1368621831;
assign addr[29178]= -1589734894;
assign addr[29179]= -1778631892;
assign addr[29180]= -1931484818;
assign addr[29181]= -2045196100;
assign addr[29182]= -2117461370;
assign addr[29183]= -2146816171;
assign addr[29184]= -2132665626;
assign addr[29185]= -2075296495;
assign addr[29186]= -1975871368;
assign addr[29187]= -1836405100;
assign addr[29188]= -1659723983;
assign addr[29189]= -1449408469;
assign addr[29190]= -1209720613;
assign addr[29191]= -945517704;
assign addr[29192]= -662153826;
assign addr[29193]= -365371365;
assign addr[29194]= -61184634;
assign addr[29195]= 244242007;
assign addr[29196]= 544719071;
assign addr[29197]= 834157373;
assign addr[29198]= 1106691431;
assign addr[29199]= 1356798326;
assign addr[29200]= 1579409630;
assign addr[29201]= 1770014111;
assign addr[29202]= 1924749160;
assign addr[29203]= 2040479063;
assign addr[29204]= 2114858546;
assign addr[29205]= 2146380306;
assign addr[29206]= 2134405552;
assign addr[29207]= 2079176953;
assign addr[29208]= 1981813720;
assign addr[29209]= 1844288924;
assign addr[29210]= 1669389513;
assign addr[29211]= 1460659832;
assign addr[29212]= 1222329801;
assign addr[29213]= 959229189;
assign addr[29214]= 676689746;
assign addr[29215]= 380437148;
assign addr[29216]= 76474970;
assign addr[29217]= -229036977;
assign addr[29218]= -529907477;
assign addr[29219]= -820039373;
assign addr[29220]= -1093553126;
assign addr[29221]= -1344905966;
assign addr[29222]= -1569004214;
assign addr[29223]= -1761306505;
assign addr[29224]= -1917915825;
assign addr[29225]= -2035658475;
assign addr[29226]= -2112148396;
assign addr[29227]= -2145835515;
assign addr[29228]= -2136037160;
assign addr[29229]= -2082951896;
assign addr[29230]= -1987655498;
assign addr[29231]= -1852079154;
assign addr[29232]= -1678970324;
assign addr[29233]= -1471837070;
assign addr[29234]= -1234876957;
assign addr[29235]= -972891995;
assign addr[29236]= -691191324;
assign addr[29237]= -395483624;
assign addr[29238]= -91761426;
assign addr[29239]= 213820322;
assign addr[29240]= 515068990;
assign addr[29241]= 805879757;
assign addr[29242]= 1080359326;
assign addr[29243]= 1332945355;
assign addr[29244]= 1558519173;
assign addr[29245]= 1752509516;
assign addr[29246]= 1910985158;
assign addr[29247]= 2030734582;
assign addr[29248]= 2109331059;
assign addr[29249]= 2145181827;
assign addr[29250]= 2137560369;
assign addr[29251]= 2086621133;
assign addr[29252]= 1993396407;
assign addr[29253]= 1859775393;
assign addr[29254]= 1688465931;
assign addr[29255]= 1482939614;
assign addr[29256]= 1247361445;
assign addr[29257]= 986505429;
assign addr[29258]= 705657826;
assign addr[29259]= 410510029;
assign addr[29260]= 107043224;
assign addr[29261]= -198592817;
assign addr[29262]= -500204365;
assign addr[29263]= -791679244;
assign addr[29264]= -1067110699;
assign addr[29265]= -1320917099;
assign addr[29266]= -1547955041;
assign addr[29267]= -1743623590;
assign addr[29268]= -1903957513;
assign addr[29269]= -2025707632;
assign addr[29270]= -2106406677;
assign addr[29271]= -2144419275;
assign addr[29272]= -2138975100;
assign addr[29273]= -2090184478;
assign addr[29274]= -1999036154;
assign addr[29275]= -1867377253;
assign addr[29276]= -1697875851;
assign addr[29277]= -1493966902;
assign addr[29278]= -1259782632;
assign addr[29279]= -1000068799;
assign addr[29280]= -720088517;
assign addr[29281]= -425515602;
assign addr[29282]= -122319591;
assign addr[29283]= 183355234;
assign addr[29284]= 485314355;
assign addr[29285]= 777438554;
assign addr[29286]= 1053807919;
assign addr[29287]= 1308821808;
assign addr[29288]= 1537312353;
assign addr[29289]= 1734649179;
assign addr[29290]= 1896833245;
assign addr[29291]= 2020577882;
assign addr[29292]= 2103375398;
assign addr[29293]= 2143547897;
assign addr[29294]= 2140281282;
assign addr[29295]= 2093641749;
assign addr[29296]= 2004574453;
assign addr[29297]= 1874884346;
assign addr[29298]= 1707199606;
assign addr[29299]= 1504918373;
assign addr[29300]= 1272139887;
assign addr[29301]= 1013581418;
assign addr[29302]= 734482665;
assign addr[29303]= 440499581;
assign addr[29304]= 137589750;
assign addr[29305]= -168108346;
assign addr[29306]= -470399716;
assign addr[29307]= -763158411;
assign addr[29308]= -1040451659;
assign addr[29309]= -1296660098;
assign addr[29310]= -1526591649;
assign addr[29311]= -1725586737;
assign addr[29312]= -1889612716;
assign addr[29313]= -2015345591;
assign addr[29314]= -2100237377;
assign addr[29315]= -2142567738;
assign addr[29316]= -2141478848;
assign addr[29317]= -2096992772;
assign addr[29318]= -2010011024;
assign addr[29319]= -1882296293;
assign addr[29320]= -1716436725;
assign addr[29321]= -1515793473;
assign addr[29322]= -1284432584;
assign addr[29323]= -1027042599;
assign addr[29324]= -748839539;
assign addr[29325]= -455461206;
assign addr[29326]= -152852926;
assign addr[29327]= 152852926;
assign addr[29328]= 455461206;
assign addr[29329]= 748839539;
assign addr[29330]= 1027042599;
assign addr[29331]= 1284432584;
assign addr[29332]= 1515793473;
assign addr[29333]= 1716436725;
assign addr[29334]= 1882296293;
assign addr[29335]= 2010011024;
assign addr[29336]= 2096992772;
assign addr[29337]= 2141478848;
assign addr[29338]= 2142567738;
assign addr[29339]= 2100237377;
assign addr[29340]= 2015345591;
assign addr[29341]= 1889612716;
assign addr[29342]= 1725586737;
assign addr[29343]= 1526591649;
assign addr[29344]= 1296660098;
assign addr[29345]= 1040451659;
assign addr[29346]= 763158411;
assign addr[29347]= 470399716;
assign addr[29348]= 168108346;
assign addr[29349]= -137589750;
assign addr[29350]= -440499581;
assign addr[29351]= -734482665;
assign addr[29352]= -1013581418;
assign addr[29353]= -1272139887;
assign addr[29354]= -1504918373;
assign addr[29355]= -1707199606;
assign addr[29356]= -1874884346;
assign addr[29357]= -2004574453;
assign addr[29358]= -2093641749;
assign addr[29359]= -2140281282;
assign addr[29360]= -2143547897;
assign addr[29361]= -2103375398;
assign addr[29362]= -2020577882;
assign addr[29363]= -1896833245;
assign addr[29364]= -1734649179;
assign addr[29365]= -1537312353;
assign addr[29366]= -1308821808;
assign addr[29367]= -1053807919;
assign addr[29368]= -777438554;
assign addr[29369]= -485314355;
assign addr[29370]= -183355234;
assign addr[29371]= 122319591;
assign addr[29372]= 425515602;
assign addr[29373]= 720088517;
assign addr[29374]= 1000068799;
assign addr[29375]= 1259782632;
assign addr[29376]= 1493966902;
assign addr[29377]= 1697875851;
assign addr[29378]= 1867377253;
assign addr[29379]= 1999036154;
assign addr[29380]= 2090184478;
assign addr[29381]= 2138975100;
assign addr[29382]= 2144419275;
assign addr[29383]= 2106406677;
assign addr[29384]= 2025707632;
assign addr[29385]= 1903957513;
assign addr[29386]= 1743623590;
assign addr[29387]= 1547955041;
assign addr[29388]= 1320917099;
assign addr[29389]= 1067110699;
assign addr[29390]= 791679244;
assign addr[29391]= 500204365;
assign addr[29392]= 198592817;
assign addr[29393]= -107043224;
assign addr[29394]= -410510029;
assign addr[29395]= -705657826;
assign addr[29396]= -986505429;
assign addr[29397]= -1247361445;
assign addr[29398]= -1482939614;
assign addr[29399]= -1688465931;
assign addr[29400]= -1859775393;
assign addr[29401]= -1993396407;
assign addr[29402]= -2086621133;
assign addr[29403]= -2137560369;
assign addr[29404]= -2145181827;
assign addr[29405]= -2109331059;
assign addr[29406]= -2030734582;
assign addr[29407]= -1910985158;
assign addr[29408]= -1752509516;
assign addr[29409]= -1558519173;
assign addr[29410]= -1332945355;
assign addr[29411]= -1080359326;
assign addr[29412]= -805879757;
assign addr[29413]= -515068990;
assign addr[29414]= -213820322;
assign addr[29415]= 91761426;
assign addr[29416]= 395483624;
assign addr[29417]= 691191324;
assign addr[29418]= 972891995;
assign addr[29419]= 1234876957;
assign addr[29420]= 1471837070;
assign addr[29421]= 1678970324;
assign addr[29422]= 1852079154;
assign addr[29423]= 1987655498;
assign addr[29424]= 2082951896;
assign addr[29425]= 2136037160;
assign addr[29426]= 2145835515;
assign addr[29427]= 2112148396;
assign addr[29428]= 2035658475;
assign addr[29429]= 1917915825;
assign addr[29430]= 1761306505;
assign addr[29431]= 1569004214;
assign addr[29432]= 1344905966;
assign addr[29433]= 1093553126;
assign addr[29434]= 820039373;
assign addr[29435]= 529907477;
assign addr[29436]= 229036977;
assign addr[29437]= -76474970;
assign addr[29438]= -380437148;
assign addr[29439]= -676689746;
assign addr[29440]= -959229189;
assign addr[29441]= -1222329801;
assign addr[29442]= -1460659832;
assign addr[29443]= -1669389513;
assign addr[29444]= -1844288924;
assign addr[29445]= -1981813720;
assign addr[29446]= -2079176953;
assign addr[29447]= -2134405552;
assign addr[29448]= -2146380306;
assign addr[29449]= -2114858546;
assign addr[29450]= -2040479063;
assign addr[29451]= -1924749160;
assign addr[29452]= -1770014111;
assign addr[29453]= -1579409630;
assign addr[29454]= -1356798326;
assign addr[29455]= -1106691431;
assign addr[29456]= -834157373;
assign addr[29457]= -544719071;
assign addr[29458]= -244242007;
assign addr[29459]= 61184634;
assign addr[29460]= 365371365;
assign addr[29461]= 662153826;
assign addr[29462]= 945517704;
assign addr[29463]= 1209720613;
assign addr[29464]= 1449408469;
assign addr[29465]= 1659723983;
assign addr[29466]= 1836405100;
assign addr[29467]= 1975871368;
assign addr[29468]= 2075296495;
assign addr[29469]= 2132665626;
assign addr[29470]= 2146816171;
assign addr[29471]= 2117461370;
assign addr[29472]= 2045196100;
assign addr[29473]= 1931484818;
assign addr[29474]= 1778631892;
assign addr[29475]= 1589734894;
assign addr[29476]= 1368621831;
assign addr[29477]= 1119773573;
assign addr[29478]= 848233042;
assign addr[29479]= 559503022;
assign addr[29480]= 259434643;
assign addr[29481]= -45891193;
assign addr[29482]= -350287041;
assign addr[29483]= -647584304;
assign addr[29484]= -931758235;
assign addr[29485]= -1197050035;
assign addr[29486]= -1438083551;
assign addr[29487]= -1649974225;
assign addr[29488]= -1828428082;
assign addr[29489]= -1969828744;
assign addr[29490]= -2071310720;
assign addr[29491]= -2130817471;
assign addr[29492]= -2147143090;
assign addr[29493]= -2119956737;
assign addr[29494]= -2049809346;
assign addr[29495]= -1938122457;
assign addr[29496]= -1787159411;
assign addr[29497]= -1599979481;
assign addr[29498]= -1380375881;
assign addr[29499]= -1132798888;
assign addr[29500]= -862265664;
assign addr[29501]= -574258580;
assign addr[29502]= -274614114;
assign addr[29503]= 30595422;
assign addr[29504]= 335184940;
assign addr[29505]= 632981917;
assign addr[29506]= 917951481;
assign addr[29507]= 1184318708;
assign addr[29508]= 1426685652;
assign addr[29509]= 1640140734;
assign addr[29510]= 1820358275;
assign addr[29511]= 1963686155;
assign addr[29512]= 2067219829;
assign addr[29513]= 2128861181;
assign addr[29514]= 2147361045;
assign addr[29515]= 2122344521;
assign addr[29516]= 2054318569;
assign addr[29517]= 1944661739;
assign addr[29518]= 1795596234;
assign addr[29519]= 1610142873;
assign addr[29520]= 1392059879;
assign addr[29521]= 1145766716;
assign addr[29522]= 876254528;
assign addr[29523]= 588984994;
assign addr[29524]= 289779648;
assign addr[29525]= -15298099;
assign addr[29526]= -320065829;
assign addr[29527]= -618347408;
assign addr[29528]= -904098143;
assign addr[29529]= -1171527280;
assign addr[29530]= -1415215352;
assign addr[29531]= -1630224009;
assign addr[29532]= -1812196087;
assign addr[29533]= -1957443913;
assign addr[29534]= -2063024031;
assign addr[29535]= -2126796855;
assign addr[29536]= -2147470025;
assign addr[29537]= -2124624598;
assign addr[29538]= -2058723538;
assign addr[29539]= -1951102334;
assign addr[29540]= -1803941934;
assign addr[29541]= -1620224553;
assign addr[29542]= -1403673233;
assign addr[29543]= -1158676398;
assign addr[29544]= -890198924;
assign addr[29545]= -603681519;
assign addr[29546]= -304930476;
assign addr[29547]= 0;
assign addr[29548]= 304930476;
assign addr[29549]= 603681519;
assign addr[29550]= 890198924;
assign addr[29551]= 1158676398;
assign addr[29552]= 1403673233;
assign addr[29553]= 1620224553;
assign addr[29554]= 1803941934;
assign addr[29555]= 1951102334;
assign addr[29556]= 2058723538;
assign addr[29557]= 2124624598;
assign addr[29558]= 2147470025;
assign addr[29559]= 2126796855;
assign addr[29560]= 2063024031;
assign addr[29561]= 1957443913;
assign addr[29562]= 1812196087;
assign addr[29563]= 1630224009;
assign addr[29564]= 1415215352;
assign addr[29565]= 1171527280;
assign addr[29566]= 904098143;
assign addr[29567]= 618347408;
assign addr[29568]= 320065829;
assign addr[29569]= 15298099;
assign addr[29570]= -289779648;
assign addr[29571]= -588984994;
assign addr[29572]= -876254528;
assign addr[29573]= -1145766716;
assign addr[29574]= -1392059879;
assign addr[29575]= -1610142873;
assign addr[29576]= -1795596234;
assign addr[29577]= -1944661739;
assign addr[29578]= -2054318569;
assign addr[29579]= -2122344521;
assign addr[29580]= -2147361045;
assign addr[29581]= -2128861181;
assign addr[29582]= -2067219829;
assign addr[29583]= -1963686155;
assign addr[29584]= -1820358275;
assign addr[29585]= -1640140734;
assign addr[29586]= -1426685652;
assign addr[29587]= -1184318708;
assign addr[29588]= -917951481;
assign addr[29589]= -632981917;
assign addr[29590]= -335184940;
assign addr[29591]= -30595422;
assign addr[29592]= 274614114;
assign addr[29593]= 574258580;
assign addr[29594]= 862265664;
assign addr[29595]= 1132798888;
assign addr[29596]= 1380375881;
assign addr[29597]= 1599979481;
assign addr[29598]= 1787159411;
assign addr[29599]= 1938122457;
assign addr[29600]= 2049809346;
assign addr[29601]= 2119956737;
assign addr[29602]= 2147143090;
assign addr[29603]= 2130817471;
assign addr[29604]= 2071310720;
assign addr[29605]= 1969828744;
assign addr[29606]= 1828428082;
assign addr[29607]= 1649974225;
assign addr[29608]= 1438083551;
assign addr[29609]= 1197050035;
assign addr[29610]= 931758235;
assign addr[29611]= 647584304;
assign addr[29612]= 350287041;
assign addr[29613]= 45891193;
assign addr[29614]= -259434643;
assign addr[29615]= -559503022;
assign addr[29616]= -848233042;
assign addr[29617]= -1119773573;
assign addr[29618]= -1368621831;
assign addr[29619]= -1589734894;
assign addr[29620]= -1778631892;
assign addr[29621]= -1931484818;
assign addr[29622]= -2045196100;
assign addr[29623]= -2117461370;
assign addr[29624]= -2146816171;
assign addr[29625]= -2132665626;
assign addr[29626]= -2075296495;
assign addr[29627]= -1975871368;
assign addr[29628]= -1836405100;
assign addr[29629]= -1659723983;
assign addr[29630]= -1449408469;
assign addr[29631]= -1209720613;
assign addr[29632]= -945517704;
assign addr[29633]= -662153826;
assign addr[29634]= -365371365;
assign addr[29635]= -61184634;
assign addr[29636]= 244242007;
assign addr[29637]= 544719071;
assign addr[29638]= 834157373;
assign addr[29639]= 1106691431;
assign addr[29640]= 1356798326;
assign addr[29641]= 1579409630;
assign addr[29642]= 1770014111;
assign addr[29643]= 1924749160;
assign addr[29644]= 2040479063;
assign addr[29645]= 2114858546;
assign addr[29646]= 2146380306;
assign addr[29647]= 2134405552;
assign addr[29648]= 2079176953;
assign addr[29649]= 1981813720;
assign addr[29650]= 1844288924;
assign addr[29651]= 1669389513;
assign addr[29652]= 1460659832;
assign addr[29653]= 1222329801;
assign addr[29654]= 959229189;
assign addr[29655]= 676689746;
assign addr[29656]= 380437148;
assign addr[29657]= 76474970;
assign addr[29658]= -229036977;
assign addr[29659]= -529907477;
assign addr[29660]= -820039373;
assign addr[29661]= -1093553126;
assign addr[29662]= -1344905966;
assign addr[29663]= -1569004214;
assign addr[29664]= -1761306505;
assign addr[29665]= -1917915825;
assign addr[29666]= -2035658475;
assign addr[29667]= -2112148396;
assign addr[29668]= -2145835515;
assign addr[29669]= -2136037160;
assign addr[29670]= -2082951896;
assign addr[29671]= -1987655498;
assign addr[29672]= -1852079154;
assign addr[29673]= -1678970324;
assign addr[29674]= -1471837070;
assign addr[29675]= -1234876957;
assign addr[29676]= -972891995;
assign addr[29677]= -691191324;
assign addr[29678]= -395483624;
assign addr[29679]= -91761426;
assign addr[29680]= 213820322;
assign addr[29681]= 515068990;
assign addr[29682]= 805879757;
assign addr[29683]= 1080359326;
assign addr[29684]= 1332945355;
assign addr[29685]= 1558519173;
assign addr[29686]= 1752509516;
assign addr[29687]= 1910985158;
assign addr[29688]= 2030734582;
assign addr[29689]= 2109331059;
assign addr[29690]= 2145181827;
assign addr[29691]= 2137560369;
assign addr[29692]= 2086621133;
assign addr[29693]= 1993396407;
assign addr[29694]= 1859775393;
assign addr[29695]= 1688465931;
assign addr[29696]= 1482939614;
assign addr[29697]= 1247361445;
assign addr[29698]= 986505429;
assign addr[29699]= 705657826;
assign addr[29700]= 410510029;
assign addr[29701]= 107043224;
assign addr[29702]= -198592817;
assign addr[29703]= -500204365;
assign addr[29704]= -791679244;
assign addr[29705]= -1067110699;
assign addr[29706]= -1320917099;
assign addr[29707]= -1547955041;
assign addr[29708]= -1743623590;
assign addr[29709]= -1903957513;
assign addr[29710]= -2025707632;
assign addr[29711]= -2106406677;
assign addr[29712]= -2144419275;
assign addr[29713]= -2138975100;
assign addr[29714]= -2090184478;
assign addr[29715]= -1999036154;
assign addr[29716]= -1867377253;
assign addr[29717]= -1697875851;
assign addr[29718]= -1493966902;
assign addr[29719]= -1259782632;
assign addr[29720]= -1000068799;
assign addr[29721]= -720088517;
assign addr[29722]= -425515602;
assign addr[29723]= -122319591;
assign addr[29724]= 183355234;
assign addr[29725]= 485314355;
assign addr[29726]= 777438554;
assign addr[29727]= 1053807919;
assign addr[29728]= 1308821808;
assign addr[29729]= 1537312353;
assign addr[29730]= 1734649179;
assign addr[29731]= 1896833245;
assign addr[29732]= 2020577882;
assign addr[29733]= 2103375398;
assign addr[29734]= 2143547897;
assign addr[29735]= 2140281282;
assign addr[29736]= 2093641749;
assign addr[29737]= 2004574453;
assign addr[29738]= 1874884346;
assign addr[29739]= 1707199606;
assign addr[29740]= 1504918373;
assign addr[29741]= 1272139887;
assign addr[29742]= 1013581418;
assign addr[29743]= 734482665;
assign addr[29744]= 440499581;
assign addr[29745]= 137589750;
assign addr[29746]= -168108346;
assign addr[29747]= -470399716;
assign addr[29748]= -763158411;
assign addr[29749]= -1040451659;
assign addr[29750]= -1296660098;
assign addr[29751]= -1526591649;
assign addr[29752]= -1725586737;
assign addr[29753]= -1889612716;
assign addr[29754]= -2015345591;
assign addr[29755]= -2100237377;
assign addr[29756]= -2142567738;
assign addr[29757]= -2141478848;
assign addr[29758]= -2096992772;
assign addr[29759]= -2010011024;
assign addr[29760]= -1882296293;
assign addr[29761]= -1716436725;
assign addr[29762]= -1515793473;
assign addr[29763]= -1284432584;
assign addr[29764]= -1027042599;
assign addr[29765]= -748839539;
assign addr[29766]= -455461206;
assign addr[29767]= -152852926;
assign addr[29768]= 152852926;
assign addr[29769]= 455461206;
assign addr[29770]= 748839539;
assign addr[29771]= 1027042599;
assign addr[29772]= 1284432584;
assign addr[29773]= 1515793473;
assign addr[29774]= 1716436725;
assign addr[29775]= 1882296293;
assign addr[29776]= 2010011024;
assign addr[29777]= 2096992772;
assign addr[29778]= 2141478848;
assign addr[29779]= 2142567738;
assign addr[29780]= 2100237377;
assign addr[29781]= 2015345591;
assign addr[29782]= 1889612716;
assign addr[29783]= 1725586737;
assign addr[29784]= 1526591649;
assign addr[29785]= 1296660098;
assign addr[29786]= 1040451659;
assign addr[29787]= 763158411;
assign addr[29788]= 470399716;
assign addr[29789]= 168108346;
assign addr[29790]= -137589750;
assign addr[29791]= -440499581;
assign addr[29792]= -734482665;
assign addr[29793]= -1013581418;
assign addr[29794]= -1272139887;
assign addr[29795]= -1504918373;
assign addr[29796]= -1707199606;
assign addr[29797]= -1874884346;
assign addr[29798]= -2004574453;
assign addr[29799]= -2093641749;
assign addr[29800]= -2140281282;
assign addr[29801]= -2143547897;
assign addr[29802]= -2103375398;
assign addr[29803]= -2020577882;
assign addr[29804]= -1896833245;
assign addr[29805]= -1734649179;
assign addr[29806]= -1537312353;
assign addr[29807]= -1308821808;
assign addr[29808]= -1053807919;
assign addr[29809]= -777438554;
assign addr[29810]= -485314355;
assign addr[29811]= -183355234;
assign addr[29812]= 122319591;
assign addr[29813]= 425515602;
assign addr[29814]= 720088517;
assign addr[29815]= 1000068799;
assign addr[29816]= 1259782632;
assign addr[29817]= 1493966902;
assign addr[29818]= 1697875851;
assign addr[29819]= 1867377253;
assign addr[29820]= 1999036154;
assign addr[29821]= 2090184478;
assign addr[29822]= 2138975100;
assign addr[29823]= 2144419275;
assign addr[29824]= 2106406677;
assign addr[29825]= 2025707632;
assign addr[29826]= 1903957513;
assign addr[29827]= 1743623590;
assign addr[29828]= 1547955041;
assign addr[29829]= 1320917099;
assign addr[29830]= 1067110699;
assign addr[29831]= 791679244;
assign addr[29832]= 500204365;
assign addr[29833]= 198592817;
assign addr[29834]= -107043224;
assign addr[29835]= -410510029;
assign addr[29836]= -705657826;
assign addr[29837]= -986505429;
assign addr[29838]= -1247361445;
assign addr[29839]= -1482939614;
assign addr[29840]= -1688465931;
assign addr[29841]= -1859775393;
assign addr[29842]= -1993396407;
assign addr[29843]= -2086621133;
assign addr[29844]= -2137560369;
assign addr[29845]= -2145181827;
assign addr[29846]= -2109331059;
assign addr[29847]= -2030734582;
assign addr[29848]= -1910985158;
assign addr[29849]= -1752509516;
assign addr[29850]= -1558519173;
assign addr[29851]= -1332945355;
assign addr[29852]= -1080359326;
assign addr[29853]= -805879757;
assign addr[29854]= -515068990;
assign addr[29855]= -213820322;
assign addr[29856]= 91761426;
assign addr[29857]= 395483624;
assign addr[29858]= 691191324;
assign addr[29859]= 972891995;
assign addr[29860]= 1234876957;
assign addr[29861]= 1471837070;
assign addr[29862]= 1678970324;
assign addr[29863]= 1852079154;
assign addr[29864]= 1987655498;
assign addr[29865]= 2082951896;
assign addr[29866]= 2136037160;
assign addr[29867]= 2145835515;
assign addr[29868]= 2112148396;
assign addr[29869]= 2035658475;
assign addr[29870]= 1917915825;
assign addr[29871]= 1761306505;
assign addr[29872]= 1569004214;
assign addr[29873]= 1344905966;
assign addr[29874]= 1093553126;
assign addr[29875]= 820039373;
assign addr[29876]= 529907477;
assign addr[29877]= 229036977;
assign addr[29878]= -76474970;
assign addr[29879]= -380437148;
assign addr[29880]= -676689746;
assign addr[29881]= -959229189;
assign addr[29882]= -1222329801;
assign addr[29883]= -1460659832;
assign addr[29884]= -1669389513;
assign addr[29885]= -1844288924;
assign addr[29886]= -1981813720;
assign addr[29887]= -2079176953;
assign addr[29888]= -2134405552;
assign addr[29889]= -2146380306;
assign addr[29890]= -2114858546;
assign addr[29891]= -2040479063;
assign addr[29892]= -1924749160;
assign addr[29893]= -1770014111;
assign addr[29894]= -1579409630;
assign addr[29895]= -1356798326;
assign addr[29896]= -1106691431;
assign addr[29897]= -834157373;
assign addr[29898]= -544719071;
assign addr[29899]= -244242007;
assign addr[29900]= 61184634;
assign addr[29901]= 365371365;
assign addr[29902]= 662153826;
assign addr[29903]= 945517704;
assign addr[29904]= 1209720613;
assign addr[29905]= 1449408469;
assign addr[29906]= 1659723983;
assign addr[29907]= 1836405100;
assign addr[29908]= 1975871368;
assign addr[29909]= 2075296495;
assign addr[29910]= 2132665626;
assign addr[29911]= 2146816171;
assign addr[29912]= 2117461370;
assign addr[29913]= 2045196100;
assign addr[29914]= 1931484818;
assign addr[29915]= 1778631892;
assign addr[29916]= 1589734894;
assign addr[29917]= 1368621831;
assign addr[29918]= 1119773573;
assign addr[29919]= 848233042;
assign addr[29920]= 559503022;
assign addr[29921]= 259434643;
assign addr[29922]= -45891193;
assign addr[29923]= -350287041;
assign addr[29924]= -647584304;
assign addr[29925]= -931758235;
assign addr[29926]= -1197050035;
assign addr[29927]= -1438083551;
assign addr[29928]= -1649974225;
assign addr[29929]= -1828428082;
assign addr[29930]= -1969828744;
assign addr[29931]= -2071310720;
assign addr[29932]= -2130817471;
assign addr[29933]= -2147143090;
assign addr[29934]= -2119956737;
assign addr[29935]= -2049809346;
assign addr[29936]= -1938122457;
assign addr[29937]= -1787159411;
assign addr[29938]= -1599979481;
assign addr[29939]= -1380375881;
assign addr[29940]= -1132798888;
assign addr[29941]= -862265664;
assign addr[29942]= -574258580;
assign addr[29943]= -274614114;
assign addr[29944]= 30595422;
assign addr[29945]= 335184940;
assign addr[29946]= 632981917;
assign addr[29947]= 917951481;
assign addr[29948]= 1184318708;
assign addr[29949]= 1426685652;
assign addr[29950]= 1640140734;
assign addr[29951]= 1820358275;
assign addr[29952]= 1963686155;
assign addr[29953]= 2067219829;
assign addr[29954]= 2128861181;
assign addr[29955]= 2147361045;
assign addr[29956]= 2122344521;
assign addr[29957]= 2054318569;
assign addr[29958]= 1944661739;
assign addr[29959]= 1795596234;
assign addr[29960]= 1610142873;
assign addr[29961]= 1392059879;
assign addr[29962]= 1145766716;
assign addr[29963]= 876254528;
assign addr[29964]= 588984994;
assign addr[29965]= 289779648;
assign addr[29966]= -15298099;
assign addr[29967]= -320065829;
assign addr[29968]= -618347408;
assign addr[29969]= -904098143;
assign addr[29970]= -1171527280;
assign addr[29971]= -1415215352;
assign addr[29972]= -1630224009;
assign addr[29973]= -1812196087;
assign addr[29974]= -1957443913;
assign addr[29975]= -2063024031;
assign addr[29976]= -2126796855;
assign addr[29977]= -2147470025;
assign addr[29978]= -2124624598;
assign addr[29979]= -2058723538;
assign addr[29980]= -1951102334;
assign addr[29981]= -1803941934;
assign addr[29982]= -1620224553;
assign addr[29983]= -1403673233;
assign addr[29984]= -1158676398;
assign addr[29985]= -890198924;
assign addr[29986]= -603681519;
assign addr[29987]= -304930476;
assign addr[29988]= 0;
assign addr[29989]= 304930476;
assign addr[29990]= 603681519;
assign addr[29991]= 890198924;
assign addr[29992]= 1158676398;
assign addr[29993]= 1403673233;
assign addr[29994]= 1620224553;
assign addr[29995]= 1803941934;
assign addr[29996]= 1951102334;
assign addr[29997]= 2058723538;
assign addr[29998]= 2124624598;
assign addr[29999]= 2147470025;
assign addr[30000]= 2126796855;
assign addr[30001]= 2063024031;
assign addr[30002]= 1957443913;
assign addr[30003]= 1812196087;
assign addr[30004]= 1630224009;
assign addr[30005]= 1415215352;
assign addr[30006]= 1171527280;
assign addr[30007]= 904098143;
assign addr[30008]= 618347408;
assign addr[30009]= 320065829;
assign addr[30010]= 15298099;
assign addr[30011]= -289779648;
assign addr[30012]= -588984994;
assign addr[30013]= -876254528;
assign addr[30014]= -1145766716;
assign addr[30015]= -1392059879;
assign addr[30016]= -1610142873;
assign addr[30017]= -1795596234;
assign addr[30018]= -1944661739;
assign addr[30019]= -2054318569;
assign addr[30020]= -2122344521;
assign addr[30021]= -2147361045;
assign addr[30022]= -2128861181;
assign addr[30023]= -2067219829;
assign addr[30024]= -1963686155;
assign addr[30025]= -1820358275;
assign addr[30026]= -1640140734;
assign addr[30027]= -1426685652;
assign addr[30028]= -1184318708;
assign addr[30029]= -917951481;
assign addr[30030]= -632981917;
assign addr[30031]= -335184940;
assign addr[30032]= -30595422;
assign addr[30033]= 274614114;
assign addr[30034]= 574258580;
assign addr[30035]= 862265664;
assign addr[30036]= 1132798888;
assign addr[30037]= 1380375881;
assign addr[30038]= 1599979481;
assign addr[30039]= 1787159411;
assign addr[30040]= 1938122457;
assign addr[30041]= 2049809346;
assign addr[30042]= 2119956737;
assign addr[30043]= 2147143090;
assign addr[30044]= 2130817471;
assign addr[30045]= 2071310720;
assign addr[30046]= 1969828744;
assign addr[30047]= 1828428082;
assign addr[30048]= 1649974225;
assign addr[30049]= 1438083551;
assign addr[30050]= 1197050035;
assign addr[30051]= 931758235;
assign addr[30052]= 647584304;
assign addr[30053]= 350287041;
assign addr[30054]= 45891193;
assign addr[30055]= -259434643;
assign addr[30056]= -559503022;
assign addr[30057]= -848233042;
assign addr[30058]= -1119773573;
assign addr[30059]= -1368621831;
assign addr[30060]= -1589734894;
assign addr[30061]= -1778631892;
assign addr[30062]= -1931484818;
assign addr[30063]= -2045196100;
assign addr[30064]= -2117461370;
assign addr[30065]= -2146816171;
assign addr[30066]= -2132665626;
assign addr[30067]= -2075296495;
assign addr[30068]= -1975871368;
assign addr[30069]= -1836405100;
assign addr[30070]= -1659723983;
assign addr[30071]= -1449408469;
assign addr[30072]= -1209720613;
assign addr[30073]= -945517704;
assign addr[30074]= -662153826;
assign addr[30075]= -365371365;
assign addr[30076]= -61184634;
assign addr[30077]= 244242007;
assign addr[30078]= 544719071;
assign addr[30079]= 834157373;
assign addr[30080]= 1106691431;
assign addr[30081]= 1356798326;
assign addr[30082]= 1579409630;
assign addr[30083]= 1770014111;
assign addr[30084]= 1924749160;
assign addr[30085]= 2040479063;
assign addr[30086]= 2114858546;
assign addr[30087]= 2146380306;
assign addr[30088]= 2134405552;
assign addr[30089]= 2079176953;
assign addr[30090]= 1981813720;
assign addr[30091]= 1844288924;
assign addr[30092]= 1669389513;
assign addr[30093]= 1460659832;
assign addr[30094]= 1222329801;
assign addr[30095]= 959229189;
assign addr[30096]= 676689746;
assign addr[30097]= 380437148;
assign addr[30098]= 76474970;
assign addr[30099]= -229036977;
assign addr[30100]= -529907477;
assign addr[30101]= -820039373;
assign addr[30102]= -1093553126;
assign addr[30103]= -1344905966;
assign addr[30104]= -1569004214;
assign addr[30105]= -1761306505;
assign addr[30106]= -1917915825;
assign addr[30107]= -2035658475;
assign addr[30108]= -2112148396;
assign addr[30109]= -2145835515;
assign addr[30110]= -2136037160;
assign addr[30111]= -2082951896;
assign addr[30112]= -1987655498;
assign addr[30113]= -1852079154;
assign addr[30114]= -1678970324;
assign addr[30115]= -1471837070;
assign addr[30116]= -1234876957;
assign addr[30117]= -972891995;
assign addr[30118]= -691191324;
assign addr[30119]= -395483624;
assign addr[30120]= -91761426;
assign addr[30121]= 213820322;
assign addr[30122]= 515068990;
assign addr[30123]= 805879757;
assign addr[30124]= 1080359326;
assign addr[30125]= 1332945355;
assign addr[30126]= 1558519173;
assign addr[30127]= 1752509516;
assign addr[30128]= 1910985158;
assign addr[30129]= 2030734582;
assign addr[30130]= 2109331059;
assign addr[30131]= 2145181827;
assign addr[30132]= 2137560369;
assign addr[30133]= 2086621133;
assign addr[30134]= 1993396407;
assign addr[30135]= 1859775393;
assign addr[30136]= 1688465931;
assign addr[30137]= 1482939614;
assign addr[30138]= 1247361445;
assign addr[30139]= 986505429;
assign addr[30140]= 705657826;
assign addr[30141]= 410510029;
assign addr[30142]= 107043224;
assign addr[30143]= -198592817;
assign addr[30144]= -500204365;
assign addr[30145]= -791679244;
assign addr[30146]= -1067110699;
assign addr[30147]= -1320917099;
assign addr[30148]= -1547955041;
assign addr[30149]= -1743623590;
assign addr[30150]= -1903957513;
assign addr[30151]= -2025707632;
assign addr[30152]= -2106406677;
assign addr[30153]= -2144419275;
assign addr[30154]= -2138975100;
assign addr[30155]= -2090184478;
assign addr[30156]= -1999036154;
assign addr[30157]= -1867377253;
assign addr[30158]= -1697875851;
assign addr[30159]= -1493966902;
assign addr[30160]= -1259782632;
assign addr[30161]= -1000068799;
assign addr[30162]= -720088517;
assign addr[30163]= -425515602;
assign addr[30164]= -122319591;
assign addr[30165]= 183355234;
assign addr[30166]= 485314355;
assign addr[30167]= 777438554;
assign addr[30168]= 1053807919;
assign addr[30169]= 1308821808;
assign addr[30170]= 1537312353;
assign addr[30171]= 1734649179;
assign addr[30172]= 1896833245;
assign addr[30173]= 2020577882;
assign addr[30174]= 2103375398;
assign addr[30175]= 2143547897;
assign addr[30176]= 2140281282;
assign addr[30177]= 2093641749;
assign addr[30178]= 2004574453;
assign addr[30179]= 1874884346;
assign addr[30180]= 1707199606;
assign addr[30181]= 1504918373;
assign addr[30182]= 1272139887;
assign addr[30183]= 1013581418;
assign addr[30184]= 734482665;
assign addr[30185]= 440499581;
assign addr[30186]= 137589750;
assign addr[30187]= -168108346;
assign addr[30188]= -470399716;
assign addr[30189]= -763158411;
assign addr[30190]= -1040451659;
assign addr[30191]= -1296660098;
assign addr[30192]= -1526591649;
assign addr[30193]= -1725586737;
assign addr[30194]= -1889612716;
assign addr[30195]= -2015345591;
assign addr[30196]= -2100237377;
assign addr[30197]= -2142567738;
assign addr[30198]= -2141478848;
assign addr[30199]= -2096992772;
assign addr[30200]= -2010011024;
assign addr[30201]= -1882296293;
assign addr[30202]= -1716436725;
assign addr[30203]= -1515793473;
assign addr[30204]= -1284432584;
assign addr[30205]= -1027042599;
assign addr[30206]= -748839539;
assign addr[30207]= -455461206;
assign addr[30208]= -152852926;
assign addr[30209]= 152852926;
assign addr[30210]= 455461206;
assign addr[30211]= 748839539;
assign addr[30212]= 1027042599;
assign addr[30213]= 1284432584;
assign addr[30214]= 1515793473;
assign addr[30215]= 1716436725;
assign addr[30216]= 1882296293;
assign addr[30217]= 2010011024;
assign addr[30218]= 2096992772;
assign addr[30219]= 2141478848;
assign addr[30220]= 2142567738;
assign addr[30221]= 2100237377;
assign addr[30222]= 2015345591;
assign addr[30223]= 1889612716;
assign addr[30224]= 1725586737;
assign addr[30225]= 1526591649;
assign addr[30226]= 1296660098;
assign addr[30227]= 1040451659;
assign addr[30228]= 763158411;
assign addr[30229]= 470399716;
assign addr[30230]= 168108346;
assign addr[30231]= -137589750;
assign addr[30232]= -440499581;
assign addr[30233]= -734482665;
assign addr[30234]= -1013581418;
assign addr[30235]= -1272139887;
assign addr[30236]= -1504918373;
assign addr[30237]= -1707199606;
assign addr[30238]= -1874884346;
assign addr[30239]= -2004574453;
assign addr[30240]= -2093641749;
assign addr[30241]= -2140281282;
assign addr[30242]= -2143547897;
assign addr[30243]= -2103375398;
assign addr[30244]= -2020577882;
assign addr[30245]= -1896833245;
assign addr[30246]= -1734649179;
assign addr[30247]= -1537312353;
assign addr[30248]= -1308821808;
assign addr[30249]= -1053807919;
assign addr[30250]= -777438554;
assign addr[30251]= -485314355;
assign addr[30252]= -183355234;
assign addr[30253]= 122319591;
assign addr[30254]= 425515602;
assign addr[30255]= 720088517;
assign addr[30256]= 1000068799;
assign addr[30257]= 1259782632;
assign addr[30258]= 1493966902;
assign addr[30259]= 1697875851;
assign addr[30260]= 1867377253;
assign addr[30261]= 1999036154;
assign addr[30262]= 2090184478;
assign addr[30263]= 2138975100;
assign addr[30264]= 2144419275;
assign addr[30265]= 2106406677;
assign addr[30266]= 2025707632;
assign addr[30267]= 1903957513;
assign addr[30268]= 1743623590;
assign addr[30269]= 1547955041;
assign addr[30270]= 1320917099;
assign addr[30271]= 1067110699;
assign addr[30272]= 791679244;
assign addr[30273]= 500204365;
assign addr[30274]= 198592817;
assign addr[30275]= -107043224;
assign addr[30276]= -410510029;
assign addr[30277]= -705657826;
assign addr[30278]= -986505429;
assign addr[30279]= -1247361445;
assign addr[30280]= -1482939614;
assign addr[30281]= -1688465931;
assign addr[30282]= -1859775393;
assign addr[30283]= -1993396407;
assign addr[30284]= -2086621133;
assign addr[30285]= -2137560369;
assign addr[30286]= -2145181827;
assign addr[30287]= -2109331059;
assign addr[30288]= -2030734582;
assign addr[30289]= -1910985158;
assign addr[30290]= -1752509516;
assign addr[30291]= -1558519173;
assign addr[30292]= -1332945355;
assign addr[30293]= -1080359326;
assign addr[30294]= -805879757;
assign addr[30295]= -515068990;
assign addr[30296]= -213820322;
assign addr[30297]= 91761426;
assign addr[30298]= 395483624;
assign addr[30299]= 691191324;
assign addr[30300]= 972891995;
assign addr[30301]= 1234876957;
assign addr[30302]= 1471837070;
assign addr[30303]= 1678970324;
assign addr[30304]= 1852079154;
assign addr[30305]= 1987655498;
assign addr[30306]= 2082951896;
assign addr[30307]= 2136037160;
assign addr[30308]= 2145835515;
assign addr[30309]= 2112148396;
assign addr[30310]= 2035658475;
assign addr[30311]= 1917915825;
assign addr[30312]= 1761306505;
assign addr[30313]= 1569004214;
assign addr[30314]= 1344905966;
assign addr[30315]= 1093553126;
assign addr[30316]= 820039373;
assign addr[30317]= 529907477;
assign addr[30318]= 229036977;
assign addr[30319]= -76474970;
assign addr[30320]= -380437148;
assign addr[30321]= -676689746;
assign addr[30322]= -959229189;
assign addr[30323]= -1222329801;
assign addr[30324]= -1460659832;
assign addr[30325]= -1669389513;
assign addr[30326]= -1844288924;
assign addr[30327]= -1981813720;
assign addr[30328]= -2079176953;
assign addr[30329]= -2134405552;
assign addr[30330]= -2146380306;
assign addr[30331]= -2114858546;
assign addr[30332]= -2040479063;
assign addr[30333]= -1924749160;
assign addr[30334]= -1770014111;
assign addr[30335]= -1579409630;
assign addr[30336]= -1356798326;
assign addr[30337]= -1106691431;
assign addr[30338]= -834157373;
assign addr[30339]= -544719071;
assign addr[30340]= -244242007;
assign addr[30341]= 61184634;
assign addr[30342]= 365371365;
assign addr[30343]= 662153826;
assign addr[30344]= 945517704;
assign addr[30345]= 1209720613;
assign addr[30346]= 1449408469;
assign addr[30347]= 1659723983;
assign addr[30348]= 1836405100;
assign addr[30349]= 1975871368;
assign addr[30350]= 2075296495;
assign addr[30351]= 2132665626;
assign addr[30352]= 2146816171;
assign addr[30353]= 2117461370;
assign addr[30354]= 2045196100;
assign addr[30355]= 1931484818;
assign addr[30356]= 1778631892;
assign addr[30357]= 1589734894;
assign addr[30358]= 1368621831;
assign addr[30359]= 1119773573;
assign addr[30360]= 848233042;
assign addr[30361]= 559503022;
assign addr[30362]= 259434643;
assign addr[30363]= -45891193;
assign addr[30364]= -350287041;
assign addr[30365]= -647584304;
assign addr[30366]= -931758235;
assign addr[30367]= -1197050035;
assign addr[30368]= -1438083551;
assign addr[30369]= -1649974225;
assign addr[30370]= -1828428082;
assign addr[30371]= -1969828744;
assign addr[30372]= -2071310720;
assign addr[30373]= -2130817471;
assign addr[30374]= -2147143090;
assign addr[30375]= -2119956737;
assign addr[30376]= -2049809346;
assign addr[30377]= -1938122457;
assign addr[30378]= -1787159411;
assign addr[30379]= -1599979481;
assign addr[30380]= -1380375881;
assign addr[30381]= -1132798888;
assign addr[30382]= -862265664;
assign addr[30383]= -574258580;
assign addr[30384]= -274614114;
assign addr[30385]= 30595422;
assign addr[30386]= 335184940;
assign addr[30387]= 632981917;
assign addr[30388]= 917951481;
assign addr[30389]= 1184318708;
assign addr[30390]= 1426685652;
assign addr[30391]= 1640140734;
assign addr[30392]= 1820358275;
assign addr[30393]= 1963686155;
assign addr[30394]= 2067219829;
assign addr[30395]= 2128861181;
assign addr[30396]= 2147361045;
assign addr[30397]= 2122344521;
assign addr[30398]= 2054318569;
assign addr[30399]= 1944661739;
assign addr[30400]= 1795596234;
assign addr[30401]= 1610142873;
assign addr[30402]= 1392059879;
assign addr[30403]= 1145766716;
assign addr[30404]= 876254528;
assign addr[30405]= 588984994;
assign addr[30406]= 289779648;
assign addr[30407]= -15298099;
assign addr[30408]= -320065829;
assign addr[30409]= -618347408;
assign addr[30410]= -904098143;
assign addr[30411]= -1171527280;
assign addr[30412]= -1415215352;
assign addr[30413]= -1630224009;
assign addr[30414]= -1812196087;
assign addr[30415]= -1957443913;
assign addr[30416]= -2063024031;
assign addr[30417]= -2126796855;
assign addr[30418]= -2147470025;
assign addr[30419]= -2124624598;
assign addr[30420]= -2058723538;
assign addr[30421]= -1951102334;
assign addr[30422]= -1803941934;
assign addr[30423]= -1620224553;
assign addr[30424]= -1403673233;
assign addr[30425]= -1158676398;
assign addr[30426]= -890198924;
assign addr[30427]= -603681519;
assign addr[30428]= -304930476;
assign addr[30429]= 0;
assign addr[30430]= 304930476;
assign addr[30431]= 603681519;
assign addr[30432]= 890198924;
assign addr[30433]= 1158676398;
assign addr[30434]= 1403673233;
assign addr[30435]= 1620224553;
assign addr[30436]= 1803941934;
assign addr[30437]= 1951102334;
assign addr[30438]= 2058723538;
assign addr[30439]= 2124624598;
assign addr[30440]= 2147470025;
assign addr[30441]= 2126796855;
assign addr[30442]= 2063024031;
assign addr[30443]= 1957443913;
assign addr[30444]= 1812196087;
assign addr[30445]= 1630224009;
assign addr[30446]= 1415215352;
assign addr[30447]= 1171527280;
assign addr[30448]= 904098143;
assign addr[30449]= 618347408;
assign addr[30450]= 320065829;
assign addr[30451]= 15298099;
assign addr[30452]= -289779648;
assign addr[30453]= -588984994;
assign addr[30454]= -876254528;
assign addr[30455]= -1145766716;
assign addr[30456]= -1392059879;
assign addr[30457]= -1610142873;
assign addr[30458]= -1795596234;
assign addr[30459]= -1944661739;
assign addr[30460]= -2054318569;
assign addr[30461]= -2122344521;
assign addr[30462]= -2147361045;
assign addr[30463]= -2128861181;
assign addr[30464]= -2067219829;
assign addr[30465]= -1963686155;
assign addr[30466]= -1820358275;
assign addr[30467]= -1640140734;
assign addr[30468]= -1426685652;
assign addr[30469]= -1184318708;
assign addr[30470]= -917951481;
assign addr[30471]= -632981917;
assign addr[30472]= -335184940;
assign addr[30473]= -30595422;
assign addr[30474]= 274614114;
assign addr[30475]= 574258580;
assign addr[30476]= 862265664;
assign addr[30477]= 1132798888;
assign addr[30478]= 1380375881;
assign addr[30479]= 1599979481;
assign addr[30480]= 1787159411;
assign addr[30481]= 1938122457;
assign addr[30482]= 2049809346;
assign addr[30483]= 2119956737;
assign addr[30484]= 2147143090;
assign addr[30485]= 2130817471;
assign addr[30486]= 2071310720;
assign addr[30487]= 1969828744;
assign addr[30488]= 1828428082;
assign addr[30489]= 1649974225;
assign addr[30490]= 1438083551;
assign addr[30491]= 1197050035;
assign addr[30492]= 931758235;
assign addr[30493]= 647584304;
assign addr[30494]= 350287041;
assign addr[30495]= 45891193;
assign addr[30496]= -259434643;
assign addr[30497]= -559503022;
assign addr[30498]= -848233042;
assign addr[30499]= -1119773573;
assign addr[30500]= -1368621831;
assign addr[30501]= -1589734894;
assign addr[30502]= -1778631892;
assign addr[30503]= -1931484818;
assign addr[30504]= -2045196100;
assign addr[30505]= -2117461370;
assign addr[30506]= -2146816171;
assign addr[30507]= -2132665626;
assign addr[30508]= -2075296495;
assign addr[30509]= -1975871368;
assign addr[30510]= -1836405100;
assign addr[30511]= -1659723983;
assign addr[30512]= -1449408469;
assign addr[30513]= -1209720613;
assign addr[30514]= -945517704;
assign addr[30515]= -662153826;
assign addr[30516]= -365371365;
assign addr[30517]= -61184634;
assign addr[30518]= 244242007;
assign addr[30519]= 544719071;
assign addr[30520]= 834157373;
assign addr[30521]= 1106691431;
assign addr[30522]= 1356798326;
assign addr[30523]= 1579409630;
assign addr[30524]= 1770014111;
assign addr[30525]= 1924749160;
assign addr[30526]= 2040479063;
assign addr[30527]= 2114858546;
assign addr[30528]= 2146380306;
assign addr[30529]= 2134405552;
assign addr[30530]= 2079176953;
assign addr[30531]= 1981813720;
assign addr[30532]= 1844288924;
assign addr[30533]= 1669389513;
assign addr[30534]= 1460659832;
assign addr[30535]= 1222329801;
assign addr[30536]= 959229189;
assign addr[30537]= 676689746;
assign addr[30538]= 380437148;
assign addr[30539]= 76474970;
assign addr[30540]= -229036977;
assign addr[30541]= -529907477;
assign addr[30542]= -820039373;
assign addr[30543]= -1093553126;
assign addr[30544]= -1344905966;
assign addr[30545]= -1569004214;
assign addr[30546]= -1761306505;
assign addr[30547]= -1917915825;
assign addr[30548]= -2035658475;
assign addr[30549]= -2112148396;
assign addr[30550]= -2145835515;
assign addr[30551]= -2136037160;
assign addr[30552]= -2082951896;
assign addr[30553]= -1987655498;
assign addr[30554]= -1852079154;
assign addr[30555]= -1678970324;
assign addr[30556]= -1471837070;
assign addr[30557]= -1234876957;
assign addr[30558]= -972891995;
assign addr[30559]= -691191324;
assign addr[30560]= -395483624;
assign addr[30561]= -91761426;
assign addr[30562]= 213820322;
assign addr[30563]= 515068990;
assign addr[30564]= 805879757;
assign addr[30565]= 1080359326;
assign addr[30566]= 1332945355;
assign addr[30567]= 1558519173;
assign addr[30568]= 1752509516;
assign addr[30569]= 1910985158;
assign addr[30570]= 2030734582;
assign addr[30571]= 2109331059;
assign addr[30572]= 2145181827;
assign addr[30573]= 2137560369;
assign addr[30574]= 2086621133;
assign addr[30575]= 1993396407;
assign addr[30576]= 1859775393;
assign addr[30577]= 1688465931;
assign addr[30578]= 1482939614;
assign addr[30579]= 1247361445;
assign addr[30580]= 986505429;
assign addr[30581]= 705657826;
assign addr[30582]= 410510029;
assign addr[30583]= 107043224;
assign addr[30584]= -198592817;
assign addr[30585]= -500204365;
assign addr[30586]= -791679244;
assign addr[30587]= -1067110699;
assign addr[30588]= -1320917099;
assign addr[30589]= -1547955041;
assign addr[30590]= -1743623590;
assign addr[30591]= -1903957513;
assign addr[30592]= -2025707632;
assign addr[30593]= -2106406677;
assign addr[30594]= -2144419275;
assign addr[30595]= -2138975100;
assign addr[30596]= -2090184478;
assign addr[30597]= -1999036154;
assign addr[30598]= -1867377253;
assign addr[30599]= -1697875851;
assign addr[30600]= -1493966902;
assign addr[30601]= -1259782632;
assign addr[30602]= -1000068799;
assign addr[30603]= -720088517;
assign addr[30604]= -425515602;
assign addr[30605]= -122319591;
assign addr[30606]= 183355234;
assign addr[30607]= 485314355;
assign addr[30608]= 777438554;
assign addr[30609]= 1053807919;
assign addr[30610]= 1308821808;
assign addr[30611]= 1537312353;
assign addr[30612]= 1734649179;
assign addr[30613]= 1896833245;
assign addr[30614]= 2020577882;
assign addr[30615]= 2103375398;
assign addr[30616]= 2143547897;
assign addr[30617]= 2140281282;
assign addr[30618]= 2093641749;
assign addr[30619]= 2004574453;
assign addr[30620]= 1874884346;
assign addr[30621]= 1707199606;
assign addr[30622]= 1504918373;
assign addr[30623]= 1272139887;
assign addr[30624]= 1013581418;
assign addr[30625]= 734482665;
assign addr[30626]= 440499581;
assign addr[30627]= 137589750;
assign addr[30628]= -168108346;
assign addr[30629]= -470399716;
assign addr[30630]= -763158411;
assign addr[30631]= -1040451659;
assign addr[30632]= -1296660098;
assign addr[30633]= -1526591649;
assign addr[30634]= -1725586737;
assign addr[30635]= -1889612716;
assign addr[30636]= -2015345591;
assign addr[30637]= -2100237377;
assign addr[30638]= -2142567738;
assign addr[30639]= -2141478848;
assign addr[30640]= -2096992772;
assign addr[30641]= -2010011024;
assign addr[30642]= -1882296293;
assign addr[30643]= -1716436725;
assign addr[30644]= -1515793473;
assign addr[30645]= -1284432584;
assign addr[30646]= -1027042599;
assign addr[30647]= -748839539;
assign addr[30648]= -455461206;
assign addr[30649]= -152852926;
assign addr[30650]= 152852926;
assign addr[30651]= 455461206;
assign addr[30652]= 748839539;
assign addr[30653]= 1027042599;
assign addr[30654]= 1284432584;
assign addr[30655]= 1515793473;
assign addr[30656]= 1716436725;
assign addr[30657]= 1882296293;
assign addr[30658]= 2010011024;
assign addr[30659]= 2096992772;
assign addr[30660]= 2141478848;
assign addr[30661]= 2142567738;
assign addr[30662]= 2100237377;
assign addr[30663]= 2015345591;
assign addr[30664]= 1889612716;
assign addr[30665]= 1725586737;
assign addr[30666]= 1526591649;
assign addr[30667]= 1296660098;
assign addr[30668]= 1040451659;
assign addr[30669]= 763158411;
assign addr[30670]= 470399716;
assign addr[30671]= 168108346;
assign addr[30672]= -137589750;
assign addr[30673]= -440499581;
assign addr[30674]= -734482665;
assign addr[30675]= -1013581418;
assign addr[30676]= -1272139887;
assign addr[30677]= -1504918373;
assign addr[30678]= -1707199606;
assign addr[30679]= -1874884346;
assign addr[30680]= -2004574453;
assign addr[30681]= -2093641749;
assign addr[30682]= -2140281282;
assign addr[30683]= -2143547897;
assign addr[30684]= -2103375398;
assign addr[30685]= -2020577882;
assign addr[30686]= -1896833245;
assign addr[30687]= -1734649179;
assign addr[30688]= -1537312353;
assign addr[30689]= -1308821808;
assign addr[30690]= -1053807919;
assign addr[30691]= -777438554;
assign addr[30692]= -485314355;
assign addr[30693]= -183355234;
assign addr[30694]= 122319591;
assign addr[30695]= 425515602;
assign addr[30696]= 720088517;
assign addr[30697]= 1000068799;
assign addr[30698]= 1259782632;
assign addr[30699]= 1493966902;
assign addr[30700]= 1697875851;
assign addr[30701]= 1867377253;
assign addr[30702]= 1999036154;
assign addr[30703]= 2090184478;
assign addr[30704]= 2138975100;
assign addr[30705]= 2144419275;
assign addr[30706]= 2106406677;
assign addr[30707]= 2025707632;
assign addr[30708]= 1903957513;
assign addr[30709]= 1743623590;
assign addr[30710]= 1547955041;
assign addr[30711]= 1320917099;
assign addr[30712]= 1067110699;
assign addr[30713]= 791679244;
assign addr[30714]= 500204365;
assign addr[30715]= 198592817;
assign addr[30716]= -107043224;
assign addr[30717]= -410510029;
assign addr[30718]= -705657826;
assign addr[30719]= -986505429;
assign addr[30720]= -1247361445;
assign addr[30721]= -1482939614;
assign addr[30722]= -1688465931;
assign addr[30723]= -1859775393;
assign addr[30724]= -1993396407;
assign addr[30725]= -2086621133;
assign addr[30726]= -2137560369;
assign addr[30727]= -2145181827;
assign addr[30728]= -2109331059;
assign addr[30729]= -2030734582;
assign addr[30730]= -1910985158;
assign addr[30731]= -1752509516;
assign addr[30732]= -1558519173;
assign addr[30733]= -1332945355;
assign addr[30734]= -1080359326;
assign addr[30735]= -805879757;
assign addr[30736]= -515068990;
assign addr[30737]= -213820322;
assign addr[30738]= 91761426;
assign addr[30739]= 395483624;
assign addr[30740]= 691191324;
assign addr[30741]= 972891995;
assign addr[30742]= 1234876957;
assign addr[30743]= 1471837070;
assign addr[30744]= 1678970324;
assign addr[30745]= 1852079154;
assign addr[30746]= 1987655498;
assign addr[30747]= 2082951896;
assign addr[30748]= 2136037160;
assign addr[30749]= 2145835515;
assign addr[30750]= 2112148396;
assign addr[30751]= 2035658475;
assign addr[30752]= 1917915825;
assign addr[30753]= 1761306505;
assign addr[30754]= 1569004214;
assign addr[30755]= 1344905966;
assign addr[30756]= 1093553126;
assign addr[30757]= 820039373;
assign addr[30758]= 529907477;
assign addr[30759]= 229036977;
assign addr[30760]= -76474970;
assign addr[30761]= -380437148;
assign addr[30762]= -676689746;
assign addr[30763]= -959229189;
assign addr[30764]= -1222329801;
assign addr[30765]= -1460659832;
assign addr[30766]= -1669389513;
assign addr[30767]= -1844288924;
assign addr[30768]= -1981813720;
assign addr[30769]= -2079176953;
assign addr[30770]= -2134405552;
assign addr[30771]= -2146380306;
assign addr[30772]= -2114858546;
assign addr[30773]= -2040479063;
assign addr[30774]= -1924749160;
assign addr[30775]= -1770014111;
assign addr[30776]= -1579409630;
assign addr[30777]= -1356798326;
assign addr[30778]= -1106691431;
assign addr[30779]= -834157373;
assign addr[30780]= -544719071;
assign addr[30781]= -244242007;
assign addr[30782]= 61184634;
assign addr[30783]= 365371365;
assign addr[30784]= 662153826;
assign addr[30785]= 945517704;
assign addr[30786]= 1209720613;
assign addr[30787]= 1449408469;
assign addr[30788]= 1659723983;
assign addr[30789]= 1836405100;
assign addr[30790]= 1975871368;
assign addr[30791]= 2075296495;
assign addr[30792]= 2132665626;
assign addr[30793]= 2146816171;
assign addr[30794]= 2117461370;
assign addr[30795]= 2045196100;
assign addr[30796]= 1931484818;
assign addr[30797]= 1778631892;
assign addr[30798]= 1589734894;
assign addr[30799]= 1368621831;
assign addr[30800]= 1119773573;
assign addr[30801]= 848233042;
assign addr[30802]= 559503022;
assign addr[30803]= 259434643;
assign addr[30804]= -45891193;
assign addr[30805]= -350287041;
assign addr[30806]= -647584304;
assign addr[30807]= -931758235;
assign addr[30808]= -1197050035;
assign addr[30809]= -1438083551;
assign addr[30810]= -1649974225;
assign addr[30811]= -1828428082;
assign addr[30812]= -1969828744;
assign addr[30813]= -2071310720;
assign addr[30814]= -2130817471;
assign addr[30815]= -2147143090;
assign addr[30816]= -2119956737;
assign addr[30817]= -2049809346;
assign addr[30818]= -1938122457;
assign addr[30819]= -1787159411;
assign addr[30820]= -1599979481;
assign addr[30821]= -1380375881;
assign addr[30822]= -1132798888;
assign addr[30823]= -862265664;
assign addr[30824]= -574258580;
assign addr[30825]= -274614114;
assign addr[30826]= 30595422;
assign addr[30827]= 335184940;
assign addr[30828]= 632981917;
assign addr[30829]= 917951481;
assign addr[30830]= 1184318708;
assign addr[30831]= 1426685652;
assign addr[30832]= 1640140734;
assign addr[30833]= 1820358275;
assign addr[30834]= 1963686155;
assign addr[30835]= 2067219829;
assign addr[30836]= 2128861181;
assign addr[30837]= 2147361045;
assign addr[30838]= 2122344521;
assign addr[30839]= 2054318569;
assign addr[30840]= 1944661739;
assign addr[30841]= 1795596234;
assign addr[30842]= 1610142873;
assign addr[30843]= 1392059879;
assign addr[30844]= 1145766716;
assign addr[30845]= 876254528;
assign addr[30846]= 588984994;
assign addr[30847]= 289779648;
assign addr[30848]= -15298099;
assign addr[30849]= -320065829;
assign addr[30850]= -618347408;
assign addr[30851]= -904098143;
assign addr[30852]= -1171527280;
assign addr[30853]= -1415215352;
assign addr[30854]= -1630224009;
assign addr[30855]= -1812196087;
assign addr[30856]= -1957443913;
assign addr[30857]= -2063024031;
assign addr[30858]= -2126796855;
assign addr[30859]= -2147470025;
assign addr[30860]= -2124624598;
assign addr[30861]= -2058723538;
assign addr[30862]= -1951102334;
assign addr[30863]= -1803941934;
assign addr[30864]= -1620224553;
assign addr[30865]= -1403673233;
assign addr[30866]= -1158676398;
assign addr[30867]= -890198924;
assign addr[30868]= -603681519;
assign addr[30869]= -304930476;
assign addr[30870]= 0;
assign addr[30871]= 304930476;
assign addr[30872]= 603681519;
assign addr[30873]= 890198924;
assign addr[30874]= 1158676398;
assign addr[30875]= 1403673233;
assign addr[30876]= 1620224553;
assign addr[30877]= 1803941934;
assign addr[30878]= 1951102334;
assign addr[30879]= 2058723538;
assign addr[30880]= 2124624598;
assign addr[30881]= 2147470025;
assign addr[30882]= 2126796855;
assign addr[30883]= 2063024031;
assign addr[30884]= 1957443913;
assign addr[30885]= 1812196087;
assign addr[30886]= 1630224009;
assign addr[30887]= 1415215352;
assign addr[30888]= 1171527280;
assign addr[30889]= 904098143;
assign addr[30890]= 618347408;
assign addr[30891]= 320065829;
assign addr[30892]= 15298099;
assign addr[30893]= -289779648;
assign addr[30894]= -588984994;
assign addr[30895]= -876254528;
assign addr[30896]= -1145766716;
assign addr[30897]= -1392059879;
assign addr[30898]= -1610142873;
assign addr[30899]= -1795596234;
assign addr[30900]= -1944661739;
assign addr[30901]= -2054318569;
assign addr[30902]= -2122344521;
assign addr[30903]= -2147361045;
assign addr[30904]= -2128861181;
assign addr[30905]= -2067219829;
assign addr[30906]= -1963686155;
assign addr[30907]= -1820358275;
assign addr[30908]= -1640140734;
assign addr[30909]= -1426685652;
assign addr[30910]= -1184318708;
assign addr[30911]= -917951481;
assign addr[30912]= -632981917;
assign addr[30913]= -335184940;
assign addr[30914]= -30595422;
assign addr[30915]= 274614114;
assign addr[30916]= 574258580;
assign addr[30917]= 862265664;
assign addr[30918]= 1132798888;
assign addr[30919]= 1380375881;
assign addr[30920]= 1599979481;
assign addr[30921]= 1787159411;
assign addr[30922]= 1938122457;
assign addr[30923]= 2049809346;
assign addr[30924]= 2119956737;
assign addr[30925]= 2147143090;
assign addr[30926]= 2130817471;
assign addr[30927]= 2071310720;
assign addr[30928]= 1969828744;
assign addr[30929]= 1828428082;
assign addr[30930]= 1649974225;
assign addr[30931]= 1438083551;
assign addr[30932]= 1197050035;
assign addr[30933]= 931758235;
assign addr[30934]= 647584304;
assign addr[30935]= 350287041;
assign addr[30936]= 45891193;
assign addr[30937]= -259434643;
assign addr[30938]= -559503022;
assign addr[30939]= -848233042;
assign addr[30940]= -1119773573;
assign addr[30941]= -1368621831;
assign addr[30942]= -1589734894;
assign addr[30943]= -1778631892;
assign addr[30944]= -1931484818;
assign addr[30945]= -2045196100;
assign addr[30946]= -2117461370;
assign addr[30947]= -2146816171;
assign addr[30948]= -2132665626;
assign addr[30949]= -2075296495;
assign addr[30950]= -1975871368;
assign addr[30951]= -1836405100;
assign addr[30952]= -1659723983;
assign addr[30953]= -1449408469;
assign addr[30954]= -1209720613;
assign addr[30955]= -945517704;
assign addr[30956]= -662153826;
assign addr[30957]= -365371365;
assign addr[30958]= -61184634;
assign addr[30959]= 244242007;
assign addr[30960]= 544719071;
assign addr[30961]= 834157373;
assign addr[30962]= 1106691431;
assign addr[30963]= 1356798326;
assign addr[30964]= 1579409630;
assign addr[30965]= 1770014111;
assign addr[30966]= 1924749160;
assign addr[30967]= 2040479063;
assign addr[30968]= 2114858546;
assign addr[30969]= 2146380306;
assign addr[30970]= 2134405552;
assign addr[30971]= 2079176953;
assign addr[30972]= 1981813720;
assign addr[30973]= 1844288924;
assign addr[30974]= 1669389513;
assign addr[30975]= 1460659832;
assign addr[30976]= 1222329801;
assign addr[30977]= 959229189;
assign addr[30978]= 676689746;
assign addr[30979]= 380437148;
assign addr[30980]= 76474970;
assign addr[30981]= -229036977;
assign addr[30982]= -529907477;
assign addr[30983]= -820039373;
assign addr[30984]= -1093553126;
assign addr[30985]= -1344905966;
assign addr[30986]= -1569004214;
assign addr[30987]= -1761306505;
assign addr[30988]= -1917915825;
assign addr[30989]= -2035658475;
assign addr[30990]= -2112148396;
assign addr[30991]= -2145835515;
assign addr[30992]= -2136037160;
assign addr[30993]= -2082951896;
assign addr[30994]= -1987655498;
assign addr[30995]= -1852079154;
assign addr[30996]= -1678970324;
assign addr[30997]= -1471837070;
assign addr[30998]= -1234876957;
assign addr[30999]= -972891995;
assign addr[31000]= -691191324;
assign addr[31001]= -395483624;
assign addr[31002]= -91761426;
assign addr[31003]= 213820322;
assign addr[31004]= 515068990;
assign addr[31005]= 805879757;
assign addr[31006]= 1080359326;
assign addr[31007]= 1332945355;
assign addr[31008]= 1558519173;
assign addr[31009]= 1752509516;
assign addr[31010]= 1910985158;
assign addr[31011]= 2030734582;
assign addr[31012]= 2109331059;
assign addr[31013]= 2145181827;
assign addr[31014]= 2137560369;
assign addr[31015]= 2086621133;
assign addr[31016]= 1993396407;
assign addr[31017]= 1859775393;
assign addr[31018]= 1688465931;
assign addr[31019]= 1482939614;
assign addr[31020]= 1247361445;
assign addr[31021]= 986505429;
assign addr[31022]= 705657826;
assign addr[31023]= 410510029;
assign addr[31024]= 107043224;
assign addr[31025]= -198592817;
assign addr[31026]= -500204365;
assign addr[31027]= -791679244;
assign addr[31028]= -1067110699;
assign addr[31029]= -1320917099;
assign addr[31030]= -1547955041;
assign addr[31031]= -1743623590;
assign addr[31032]= -1903957513;
assign addr[31033]= -2025707632;
assign addr[31034]= -2106406677;
assign addr[31035]= -2144419275;
assign addr[31036]= -2138975100;
assign addr[31037]= -2090184478;
assign addr[31038]= -1999036154;
assign addr[31039]= -1867377253;
assign addr[31040]= -1697875851;
assign addr[31041]= -1493966902;
assign addr[31042]= -1259782632;
assign addr[31043]= -1000068799;
assign addr[31044]= -720088517;
assign addr[31045]= -425515602;
assign addr[31046]= -122319591;
assign addr[31047]= 183355234;
assign addr[31048]= 485314355;
assign addr[31049]= 777438554;
assign addr[31050]= 1053807919;
assign addr[31051]= 1308821808;
assign addr[31052]= 1537312353;
assign addr[31053]= 1734649179;
assign addr[31054]= 1896833245;
assign addr[31055]= 2020577882;
assign addr[31056]= 2103375398;
assign addr[31057]= 2143547897;
assign addr[31058]= 2140281282;
assign addr[31059]= 2093641749;
assign addr[31060]= 2004574453;
assign addr[31061]= 1874884346;
assign addr[31062]= 1707199606;
assign addr[31063]= 1504918373;
assign addr[31064]= 1272139887;
assign addr[31065]= 1013581418;
assign addr[31066]= 734482665;
assign addr[31067]= 440499581;
assign addr[31068]= 137589750;
assign addr[31069]= -168108346;
assign addr[31070]= -470399716;
assign addr[31071]= -763158411;
assign addr[31072]= -1040451659;
assign addr[31073]= -1296660098;
assign addr[31074]= -1526591649;
assign addr[31075]= -1725586737;
assign addr[31076]= -1889612716;
assign addr[31077]= -2015345591;
assign addr[31078]= -2100237377;
assign addr[31079]= -2142567738;
assign addr[31080]= -2141478848;
assign addr[31081]= -2096992772;
assign addr[31082]= -2010011024;
assign addr[31083]= -1882296293;
assign addr[31084]= -1716436725;
assign addr[31085]= -1515793473;
assign addr[31086]= -1284432584;
assign addr[31087]= -1027042599;
assign addr[31088]= -748839539;
assign addr[31089]= -455461206;
assign addr[31090]= -152852926;
assign addr[31091]= 152852926;
assign addr[31092]= 455461206;
assign addr[31093]= 748839539;
assign addr[31094]= 1027042599;
assign addr[31095]= 1284432584;
assign addr[31096]= 1515793473;
assign addr[31097]= 1716436725;
assign addr[31098]= 1882296293;
assign addr[31099]= 2010011024;
assign addr[31100]= 2096992772;
assign addr[31101]= 2141478848;
assign addr[31102]= 2142567738;
assign addr[31103]= 2100237377;
assign addr[31104]= 2015345591;
assign addr[31105]= 1889612716;
assign addr[31106]= 1725586737;
assign addr[31107]= 1526591649;
assign addr[31108]= 1296660098;
assign addr[31109]= 1040451659;
assign addr[31110]= 763158411;
assign addr[31111]= 470399716;
assign addr[31112]= 168108346;
assign addr[31113]= -137589750;
assign addr[31114]= -440499581;
assign addr[31115]= -734482665;
assign addr[31116]= -1013581418;
assign addr[31117]= -1272139887;
assign addr[31118]= -1504918373;
assign addr[31119]= -1707199606;
assign addr[31120]= -1874884346;
assign addr[31121]= -2004574453;
assign addr[31122]= -2093641749;
assign addr[31123]= -2140281282;
assign addr[31124]= -2143547897;
assign addr[31125]= -2103375398;
assign addr[31126]= -2020577882;
assign addr[31127]= -1896833245;
assign addr[31128]= -1734649179;
assign addr[31129]= -1537312353;
assign addr[31130]= -1308821808;
assign addr[31131]= -1053807919;
assign addr[31132]= -777438554;
assign addr[31133]= -485314355;
assign addr[31134]= -183355234;
assign addr[31135]= 122319591;
assign addr[31136]= 425515602;
assign addr[31137]= 720088517;
assign addr[31138]= 1000068799;
assign addr[31139]= 1259782632;
assign addr[31140]= 1493966902;
assign addr[31141]= 1697875851;
assign addr[31142]= 1867377253;
assign addr[31143]= 1999036154;
assign addr[31144]= 2090184478;
assign addr[31145]= 2138975100;
assign addr[31146]= 2144419275;
assign addr[31147]= 2106406677;
assign addr[31148]= 2025707632;
assign addr[31149]= 1903957513;
assign addr[31150]= 1743623590;
assign addr[31151]= 1547955041;
assign addr[31152]= 1320917099;
assign addr[31153]= 1067110699;
assign addr[31154]= 791679244;
assign addr[31155]= 500204365;
assign addr[31156]= 198592817;
assign addr[31157]= -107043224;
assign addr[31158]= -410510029;
assign addr[31159]= -705657826;
assign addr[31160]= -986505429;
assign addr[31161]= -1247361445;
assign addr[31162]= -1482939614;
assign addr[31163]= -1688465931;
assign addr[31164]= -1859775393;
assign addr[31165]= -1993396407;
assign addr[31166]= -2086621133;
assign addr[31167]= -2137560369;
assign addr[31168]= -2145181827;
assign addr[31169]= -2109331059;
assign addr[31170]= -2030734582;
assign addr[31171]= -1910985158;
assign addr[31172]= -1752509516;
assign addr[31173]= -1558519173;
assign addr[31174]= -1332945355;
assign addr[31175]= -1080359326;
assign addr[31176]= -805879757;
assign addr[31177]= -515068990;
assign addr[31178]= -213820322;
assign addr[31179]= 91761426;
assign addr[31180]= 395483624;
assign addr[31181]= 691191324;
assign addr[31182]= 972891995;
assign addr[31183]= 1234876957;
assign addr[31184]= 1471837070;
assign addr[31185]= 1678970324;
assign addr[31186]= 1852079154;
assign addr[31187]= 1987655498;
assign addr[31188]= 2082951896;
assign addr[31189]= 2136037160;
assign addr[31190]= 2145835515;
assign addr[31191]= 2112148396;
assign addr[31192]= 2035658475;
assign addr[31193]= 1917915825;
assign addr[31194]= 1761306505;
assign addr[31195]= 1569004214;
assign addr[31196]= 1344905966;
assign addr[31197]= 1093553126;
assign addr[31198]= 820039373;
assign addr[31199]= 529907477;
assign addr[31200]= 229036977;
assign addr[31201]= -76474970;
assign addr[31202]= -380437148;
assign addr[31203]= -676689746;
assign addr[31204]= -959229189;
assign addr[31205]= -1222329801;
assign addr[31206]= -1460659832;
assign addr[31207]= -1669389513;
assign addr[31208]= -1844288924;
assign addr[31209]= -1981813720;
assign addr[31210]= -2079176953;
assign addr[31211]= -2134405552;
assign addr[31212]= -2146380306;
assign addr[31213]= -2114858546;
assign addr[31214]= -2040479063;
assign addr[31215]= -1924749160;
assign addr[31216]= -1770014111;
assign addr[31217]= -1579409630;
assign addr[31218]= -1356798326;
assign addr[31219]= -1106691431;
assign addr[31220]= -834157373;
assign addr[31221]= -544719071;
assign addr[31222]= -244242007;
assign addr[31223]= 61184634;
assign addr[31224]= 365371365;
assign addr[31225]= 662153826;
assign addr[31226]= 945517704;
assign addr[31227]= 1209720613;
assign addr[31228]= 1449408469;
assign addr[31229]= 1659723983;
assign addr[31230]= 1836405100;
assign addr[31231]= 1975871368;
assign addr[31232]= 2075296495;
assign addr[31233]= 2132665626;
assign addr[31234]= 2146816171;
assign addr[31235]= 2117461370;
assign addr[31236]= 2045196100;
assign addr[31237]= 1931484818;
assign addr[31238]= 1778631892;
assign addr[31239]= 1589734894;
assign addr[31240]= 1368621831;
assign addr[31241]= 1119773573;
assign addr[31242]= 848233042;
assign addr[31243]= 559503022;
assign addr[31244]= 259434643;
assign addr[31245]= -45891193;
assign addr[31246]= -350287041;
assign addr[31247]= -647584304;
assign addr[31248]= -931758235;
assign addr[31249]= -1197050035;
assign addr[31250]= -1438083551;
assign addr[31251]= -1649974225;
assign addr[31252]= -1828428082;
assign addr[31253]= -1969828744;
assign addr[31254]= -2071310720;
assign addr[31255]= -2130817471;
assign addr[31256]= -2147143090;
assign addr[31257]= -2119956737;
assign addr[31258]= -2049809346;
assign addr[31259]= -1938122457;
assign addr[31260]= -1787159411;
assign addr[31261]= -1599979481;
assign addr[31262]= -1380375881;
assign addr[31263]= -1132798888;
assign addr[31264]= -862265664;
assign addr[31265]= -574258580;
assign addr[31266]= -274614114;
assign addr[31267]= 30595422;
assign addr[31268]= 335184940;
assign addr[31269]= 632981917;
assign addr[31270]= 917951481;
assign addr[31271]= 1184318708;
assign addr[31272]= 1426685652;
assign addr[31273]= 1640140734;
assign addr[31274]= 1820358275;
assign addr[31275]= 1963686155;
assign addr[31276]= 2067219829;
assign addr[31277]= 2128861181;
assign addr[31278]= 2147361045;
assign addr[31279]= 2122344521;
assign addr[31280]= 2054318569;
assign addr[31281]= 1944661739;
assign addr[31282]= 1795596234;
assign addr[31283]= 1610142873;
assign addr[31284]= 1392059879;
assign addr[31285]= 1145766716;
assign addr[31286]= 876254528;
assign addr[31287]= 588984994;
assign addr[31288]= 289779648;
assign addr[31289]= -15298099;
assign addr[31290]= -320065829;
assign addr[31291]= -618347408;
assign addr[31292]= -904098143;
assign addr[31293]= -1171527280;
assign addr[31294]= -1415215352;
assign addr[31295]= -1630224009;
assign addr[31296]= -1812196087;
assign addr[31297]= -1957443913;
assign addr[31298]= -2063024031;
assign addr[31299]= -2126796855;
assign addr[31300]= -2147470025;
assign addr[31301]= -2124624598;
assign addr[31302]= -2058723538;
assign addr[31303]= -1951102334;
assign addr[31304]= -1803941934;
assign addr[31305]= -1620224553;
assign addr[31306]= -1403673233;
assign addr[31307]= -1158676398;
assign addr[31308]= -890198924;
assign addr[31309]= -603681519;
assign addr[31310]= -304930476;
assign addr[31311]= 0;
assign addr[31312]= 304930476;
assign addr[31313]= 603681519;
assign addr[31314]= 890198924;
assign addr[31315]= 1158676398;
assign addr[31316]= 1403673233;
assign addr[31317]= 1620224553;
assign addr[31318]= 1803941934;
assign addr[31319]= 1951102334;
assign addr[31320]= 2058723538;
assign addr[31321]= 2124624598;
assign addr[31322]= 2147470025;
assign addr[31323]= 2126796855;
assign addr[31324]= 2063024031;
assign addr[31325]= 1957443913;
assign addr[31326]= 1812196087;
assign addr[31327]= 1630224009;
assign addr[31328]= 1415215352;
assign addr[31329]= 1171527280;
assign addr[31330]= 904098143;
assign addr[31331]= 618347408;
assign addr[31332]= 320065829;
assign addr[31333]= 15298099;
assign addr[31334]= -289779648;
assign addr[31335]= -588984994;
assign addr[31336]= -876254528;
assign addr[31337]= -1145766716;
assign addr[31338]= -1392059879;
assign addr[31339]= -1610142873;
assign addr[31340]= -1795596234;
assign addr[31341]= -1944661739;
assign addr[31342]= -2054318569;
assign addr[31343]= -2122344521;
assign addr[31344]= -2147361045;
assign addr[31345]= -2128861181;
assign addr[31346]= -2067219829;
assign addr[31347]= -1963686155;
assign addr[31348]= -1820358275;
assign addr[31349]= -1640140734;
assign addr[31350]= -1426685652;
assign addr[31351]= -1184318708;
assign addr[31352]= -917951481;
assign addr[31353]= -632981917;
assign addr[31354]= -335184940;
assign addr[31355]= -30595422;
assign addr[31356]= 274614114;
assign addr[31357]= 574258580;
assign addr[31358]= 862265664;
assign addr[31359]= 1132798888;
assign addr[31360]= 1380375881;
assign addr[31361]= 1599979481;
assign addr[31362]= 1787159411;
assign addr[31363]= 1938122457;
assign addr[31364]= 2049809346;
assign addr[31365]= 2119956737;
assign addr[31366]= 2147143090;
assign addr[31367]= 2130817471;
assign addr[31368]= 2071310720;
assign addr[31369]= 1969828744;
assign addr[31370]= 1828428082;
assign addr[31371]= 1649974225;
assign addr[31372]= 1438083551;
assign addr[31373]= 1197050035;
assign addr[31374]= 931758235;
assign addr[31375]= 647584304;
assign addr[31376]= 350287041;
assign addr[31377]= 45891193;
assign addr[31378]= -259434643;
assign addr[31379]= -559503022;
assign addr[31380]= -848233042;
assign addr[31381]= -1119773573;
assign addr[31382]= -1368621831;
assign addr[31383]= -1589734894;
assign addr[31384]= -1778631892;
assign addr[31385]= -1931484818;
assign addr[31386]= -2045196100;
assign addr[31387]= -2117461370;
assign addr[31388]= -2146816171;
assign addr[31389]= -2132665626;
assign addr[31390]= -2075296495;
assign addr[31391]= -1975871368;
assign addr[31392]= -1836405100;
assign addr[31393]= -1659723983;
assign addr[31394]= -1449408469;
assign addr[31395]= -1209720613;
assign addr[31396]= -945517704;
assign addr[31397]= -662153826;
assign addr[31398]= -365371365;
assign addr[31399]= -61184634;
assign addr[31400]= 244242007;
assign addr[31401]= 544719071;
assign addr[31402]= 834157373;
assign addr[31403]= 1106691431;
assign addr[31404]= 1356798326;
assign addr[31405]= 1579409630;
assign addr[31406]= 1770014111;
assign addr[31407]= 1924749160;
assign addr[31408]= 2040479063;
assign addr[31409]= 2114858546;
assign addr[31410]= 2146380306;
assign addr[31411]= 2134405552;
assign addr[31412]= 2079176953;
assign addr[31413]= 1981813720;
assign addr[31414]= 1844288924;
assign addr[31415]= 1669389513;
assign addr[31416]= 1460659832;
assign addr[31417]= 1222329801;
assign addr[31418]= 959229189;
assign addr[31419]= 676689746;
assign addr[31420]= 380437148;
assign addr[31421]= 76474970;
assign addr[31422]= -229036977;
assign addr[31423]= -529907477;
assign addr[31424]= -820039373;
assign addr[31425]= -1093553126;
assign addr[31426]= -1344905966;
assign addr[31427]= -1569004214;
assign addr[31428]= -1761306505;
assign addr[31429]= -1917915825;
assign addr[31430]= -2035658475;
assign addr[31431]= -2112148396;
assign addr[31432]= -2145835515;
assign addr[31433]= -2136037160;
assign addr[31434]= -2082951896;
assign addr[31435]= -1987655498;
assign addr[31436]= -1852079154;
assign addr[31437]= -1678970324;
assign addr[31438]= -1471837070;
assign addr[31439]= -1234876957;
assign addr[31440]= -972891995;
assign addr[31441]= -691191324;
assign addr[31442]= -395483624;
assign addr[31443]= -91761426;
assign addr[31444]= 213820322;
assign addr[31445]= 515068990;
assign addr[31446]= 805879757;
assign addr[31447]= 1080359326;
assign addr[31448]= 1332945355;
assign addr[31449]= 1558519173;
assign addr[31450]= 1752509516;
assign addr[31451]= 1910985158;
assign addr[31452]= 2030734582;
assign addr[31453]= 2109331059;
assign addr[31454]= 2145181827;
assign addr[31455]= 2137560369;
assign addr[31456]= 2086621133;
assign addr[31457]= 1993396407;
assign addr[31458]= 1859775393;
assign addr[31459]= 1688465931;
assign addr[31460]= 1482939614;
assign addr[31461]= 1247361445;
assign addr[31462]= 986505429;
assign addr[31463]= 705657826;
assign addr[31464]= 410510029;
assign addr[31465]= 107043224;
assign addr[31466]= -198592817;
assign addr[31467]= -500204365;
assign addr[31468]= -791679244;
assign addr[31469]= -1067110699;
assign addr[31470]= -1320917099;
assign addr[31471]= -1547955041;
assign addr[31472]= -1743623590;
assign addr[31473]= -1903957513;
assign addr[31474]= -2025707632;
assign addr[31475]= -2106406677;
assign addr[31476]= -2144419275;
assign addr[31477]= -2138975100;
assign addr[31478]= -2090184478;
assign addr[31479]= -1999036154;
assign addr[31480]= -1867377253;
assign addr[31481]= -1697875851;
assign addr[31482]= -1493966902;
assign addr[31483]= -1259782632;
assign addr[31484]= -1000068799;
assign addr[31485]= -720088517;
assign addr[31486]= -425515602;
assign addr[31487]= -122319591;
assign addr[31488]= 183355234;
assign addr[31489]= 485314355;
assign addr[31490]= 777438554;
assign addr[31491]= 1053807919;
assign addr[31492]= 1308821808;
assign addr[31493]= 1537312353;
assign addr[31494]= 1734649179;
assign addr[31495]= 1896833245;
assign addr[31496]= 2020577882;
assign addr[31497]= 2103375398;
assign addr[31498]= 2143547897;
assign addr[31499]= 2140281282;
assign addr[31500]= 2093641749;
assign addr[31501]= 2004574453;
assign addr[31502]= 1874884346;
assign addr[31503]= 1707199606;
assign addr[31504]= 1504918373;
assign addr[31505]= 1272139887;
assign addr[31506]= 1013581418;
assign addr[31507]= 734482665;
assign addr[31508]= 440499581;
assign addr[31509]= 137589750;
assign addr[31510]= -168108346;
assign addr[31511]= -470399716;
assign addr[31512]= -763158411;
assign addr[31513]= -1040451659;
assign addr[31514]= -1296660098;
assign addr[31515]= -1526591649;
assign addr[31516]= -1725586737;
assign addr[31517]= -1889612716;
assign addr[31518]= -2015345591;
assign addr[31519]= -2100237377;
assign addr[31520]= -2142567738;
assign addr[31521]= -2141478848;
assign addr[31522]= -2096992772;
assign addr[31523]= -2010011024;
assign addr[31524]= -1882296293;
assign addr[31525]= -1716436725;
assign addr[31526]= -1515793473;
assign addr[31527]= -1284432584;
assign addr[31528]= -1027042599;
assign addr[31529]= -748839539;
assign addr[31530]= -455461206;
assign addr[31531]= -152852926;
assign addr[31532]= 152852926;
assign addr[31533]= 455461206;
assign addr[31534]= 748839539;
assign addr[31535]= 1027042599;
assign addr[31536]= 1284432584;
assign addr[31537]= 1515793473;
assign addr[31538]= 1716436725;
assign addr[31539]= 1882296293;
assign addr[31540]= 2010011024;
assign addr[31541]= 2096992772;
assign addr[31542]= 2141478848;
assign addr[31543]= 2142567738;
assign addr[31544]= 2100237377;
assign addr[31545]= 2015345591;
assign addr[31546]= 1889612716;
assign addr[31547]= 1725586737;
assign addr[31548]= 1526591649;
assign addr[31549]= 1296660098;
assign addr[31550]= 1040451659;
assign addr[31551]= 763158411;
assign addr[31552]= 470399716;
assign addr[31553]= 168108346;
assign addr[31554]= -137589750;
assign addr[31555]= -440499581;
assign addr[31556]= -734482665;
assign addr[31557]= -1013581418;
assign addr[31558]= -1272139887;
assign addr[31559]= -1504918373;
assign addr[31560]= -1707199606;
assign addr[31561]= -1874884346;
assign addr[31562]= -2004574453;
assign addr[31563]= -2093641749;
assign addr[31564]= -2140281282;
assign addr[31565]= -2143547897;
assign addr[31566]= -2103375398;
assign addr[31567]= -2020577882;
assign addr[31568]= -1896833245;
assign addr[31569]= -1734649179;
assign addr[31570]= -1537312353;
assign addr[31571]= -1308821808;
assign addr[31572]= -1053807919;
assign addr[31573]= -777438554;
assign addr[31574]= -485314355;
assign addr[31575]= -183355234;
assign addr[31576]= 122319591;
assign addr[31577]= 425515602;
assign addr[31578]= 720088517;
assign addr[31579]= 1000068799;
assign addr[31580]= 1259782632;
assign addr[31581]= 1493966902;
assign addr[31582]= 1697875851;
assign addr[31583]= 1867377253;
assign addr[31584]= 1999036154;
assign addr[31585]= 2090184478;
assign addr[31586]= 2138975100;
assign addr[31587]= 2144419275;
assign addr[31588]= 2106406677;
assign addr[31589]= 2025707632;
assign addr[31590]= 1903957513;
assign addr[31591]= 1743623590;
assign addr[31592]= 1547955041;
assign addr[31593]= 1320917099;
assign addr[31594]= 1067110699;
assign addr[31595]= 791679244;
assign addr[31596]= 500204365;
assign addr[31597]= 198592817;
assign addr[31598]= -107043224;
assign addr[31599]= -410510029;
assign addr[31600]= -705657826;
assign addr[31601]= -986505429;
assign addr[31602]= -1247361445;
assign addr[31603]= -1482939614;
assign addr[31604]= -1688465931;
assign addr[31605]= -1859775393;
assign addr[31606]= -1993396407;
assign addr[31607]= -2086621133;
assign addr[31608]= -2137560369;
assign addr[31609]= -2145181827;
assign addr[31610]= -2109331059;
assign addr[31611]= -2030734582;
assign addr[31612]= -1910985158;
assign addr[31613]= -1752509516;
assign addr[31614]= -1558519173;
assign addr[31615]= -1332945355;
assign addr[31616]= -1080359326;
assign addr[31617]= -805879757;
assign addr[31618]= -515068990;
assign addr[31619]= -213820322;
assign addr[31620]= 91761426;
assign addr[31621]= 395483624;
assign addr[31622]= 691191324;
assign addr[31623]= 972891995;
assign addr[31624]= 1234876957;
assign addr[31625]= 1471837070;
assign addr[31626]= 1678970324;
assign addr[31627]= 1852079154;
assign addr[31628]= 1987655498;
assign addr[31629]= 2082951896;
assign addr[31630]= 2136037160;
assign addr[31631]= 2145835515;
assign addr[31632]= 2112148396;
assign addr[31633]= 2035658475;
assign addr[31634]= 1917915825;
assign addr[31635]= 1761306505;
assign addr[31636]= 1569004214;
assign addr[31637]= 1344905966;
assign addr[31638]= 1093553126;
assign addr[31639]= 820039373;
assign addr[31640]= 529907477;
assign addr[31641]= 229036977;
assign addr[31642]= -76474970;
assign addr[31643]= -380437148;
assign addr[31644]= -676689746;
assign addr[31645]= -959229189;
assign addr[31646]= -1222329801;
assign addr[31647]= -1460659832;
assign addr[31648]= -1669389513;
assign addr[31649]= -1844288924;
assign addr[31650]= -1981813720;
assign addr[31651]= -2079176953;
assign addr[31652]= -2134405552;
assign addr[31653]= -2146380306;
assign addr[31654]= -2114858546;
assign addr[31655]= -2040479063;
assign addr[31656]= -1924749160;
assign addr[31657]= -1770014111;
assign addr[31658]= -1579409630;
assign addr[31659]= -1356798326;
assign addr[31660]= -1106691431;
assign addr[31661]= -834157373;
assign addr[31662]= -544719071;
assign addr[31663]= -244242007;
assign addr[31664]= 61184634;
assign addr[31665]= 365371365;
assign addr[31666]= 662153826;
assign addr[31667]= 945517704;
assign addr[31668]= 1209720613;
assign addr[31669]= 1449408469;
assign addr[31670]= 1659723983;
assign addr[31671]= 1836405100;
assign addr[31672]= 1975871368;
assign addr[31673]= 2075296495;
assign addr[31674]= 2132665626;
assign addr[31675]= 2146816171;
assign addr[31676]= 2117461370;
assign addr[31677]= 2045196100;
assign addr[31678]= 1931484818;
assign addr[31679]= 1778631892;
assign addr[31680]= 1589734894;
assign addr[31681]= 1368621831;
assign addr[31682]= 1119773573;
assign addr[31683]= 848233042;
assign addr[31684]= 559503022;
assign addr[31685]= 259434643;
assign addr[31686]= -45891193;
assign addr[31687]= -350287041;
assign addr[31688]= -647584304;
assign addr[31689]= -931758235;
assign addr[31690]= -1197050035;
assign addr[31691]= -1438083551;
assign addr[31692]= -1649974225;
assign addr[31693]= -1828428082;
assign addr[31694]= -1969828744;
assign addr[31695]= -2071310720;
assign addr[31696]= -2130817471;
assign addr[31697]= -2147143090;
assign addr[31698]= -2119956737;
assign addr[31699]= -2049809346;
assign addr[31700]= -1938122457;
assign addr[31701]= -1787159411;
assign addr[31702]= -1599979481;
assign addr[31703]= -1380375881;
assign addr[31704]= -1132798888;
assign addr[31705]= -862265664;
assign addr[31706]= -574258580;
assign addr[31707]= -274614114;
assign addr[31708]= 30595422;
assign addr[31709]= 335184940;
assign addr[31710]= 632981917;
assign addr[31711]= 917951481;
assign addr[31712]= 1184318708;
assign addr[31713]= 1426685652;
assign addr[31714]= 1640140734;
assign addr[31715]= 1820358275;
assign addr[31716]= 1963686155;
assign addr[31717]= 2067219829;
assign addr[31718]= 2128861181;
assign addr[31719]= 2147361045;
assign addr[31720]= 2122344521;
assign addr[31721]= 2054318569;
assign addr[31722]= 1944661739;
assign addr[31723]= 1795596234;
assign addr[31724]= 1610142873;
assign addr[31725]= 1392059879;
assign addr[31726]= 1145766716;
assign addr[31727]= 876254528;
assign addr[31728]= 588984994;
assign addr[31729]= 289779648;
assign addr[31730]= -15298099;
assign addr[31731]= -320065829;
assign addr[31732]= -618347408;
assign addr[31733]= -904098143;
assign addr[31734]= -1171527280;
assign addr[31735]= -1415215352;
assign addr[31736]= -1630224009;
assign addr[31737]= -1812196087;
assign addr[31738]= -1957443913;
assign addr[31739]= -2063024031;
assign addr[31740]= -2126796855;
assign addr[31741]= -2147470025;
assign addr[31742]= -2124624598;
assign addr[31743]= -2058723538;
assign addr[31744]= -1951102334;
assign addr[31745]= -1803941934;
assign addr[31746]= -1620224553;
assign addr[31747]= -1403673233;
assign addr[31748]= -1158676398;
assign addr[31749]= -890198924;
assign addr[31750]= -603681519;
assign addr[31751]= -304930476;
assign addr[31752]= 0;
assign addr[31753]= 304930476;
assign addr[31754]= 603681519;
assign addr[31755]= 890198924;
assign addr[31756]= 1158676398;
assign addr[31757]= 1403673233;
assign addr[31758]= 1620224553;
assign addr[31759]= 1803941934;
assign addr[31760]= 1951102334;
assign addr[31761]= 2058723538;
assign addr[31762]= 2124624598;
assign addr[31763]= 2147470025;
assign addr[31764]= 2126796855;
assign addr[31765]= 2063024031;
assign addr[31766]= 1957443913;
assign addr[31767]= 1812196087;
assign addr[31768]= 1630224009;
assign addr[31769]= 1415215352;
assign addr[31770]= 1171527280;
assign addr[31771]= 904098143;
assign addr[31772]= 618347408;
assign addr[31773]= 320065829;
assign addr[31774]= 15298099;
assign addr[31775]= -289779648;
assign addr[31776]= -588984994;
assign addr[31777]= -876254528;
assign addr[31778]= -1145766716;
assign addr[31779]= -1392059879;
assign addr[31780]= -1610142873;
assign addr[31781]= -1795596234;
assign addr[31782]= -1944661739;
assign addr[31783]= -2054318569;
assign addr[31784]= -2122344521;
assign addr[31785]= -2147361045;
assign addr[31786]= -2128861181;
assign addr[31787]= -2067219829;
assign addr[31788]= -1963686155;
assign addr[31789]= -1820358275;
assign addr[31790]= -1640140734;
assign addr[31791]= -1426685652;
assign addr[31792]= -1184318708;
assign addr[31793]= -917951481;
assign addr[31794]= -632981917;
assign addr[31795]= -335184940;
assign addr[31796]= -30595422;
assign addr[31797]= 274614114;
assign addr[31798]= 574258580;
assign addr[31799]= 862265664;
assign addr[31800]= 1132798888;
assign addr[31801]= 1380375881;
assign addr[31802]= 1599979481;
assign addr[31803]= 1787159411;
assign addr[31804]= 1938122457;
assign addr[31805]= 2049809346;
assign addr[31806]= 2119956737;
assign addr[31807]= 2147143090;
assign addr[31808]= 2130817471;
assign addr[31809]= 2071310720;
assign addr[31810]= 1969828744;
assign addr[31811]= 1828428082;
assign addr[31812]= 1649974225;
assign addr[31813]= 1438083551;
assign addr[31814]= 1197050035;
assign addr[31815]= 931758235;
assign addr[31816]= 647584304;
assign addr[31817]= 350287041;
assign addr[31818]= 45891193;
assign addr[31819]= -259434643;
assign addr[31820]= -559503022;
assign addr[31821]= -848233042;
assign addr[31822]= -1119773573;
assign addr[31823]= -1368621831;
assign addr[31824]= -1589734894;
assign addr[31825]= -1778631892;
assign addr[31826]= -1931484818;
assign addr[31827]= -2045196100;
assign addr[31828]= -2117461370;
assign addr[31829]= -2146816171;
assign addr[31830]= -2132665626;
assign addr[31831]= -2075296495;
assign addr[31832]= -1975871368;
assign addr[31833]= -1836405100;
assign addr[31834]= -1659723983;
assign addr[31835]= -1449408469;
assign addr[31836]= -1209720613;
assign addr[31837]= -945517704;
assign addr[31838]= -662153826;
assign addr[31839]= -365371365;
assign addr[31840]= -61184634;
assign addr[31841]= 244242007;
assign addr[31842]= 544719071;
assign addr[31843]= 834157373;
assign addr[31844]= 1106691431;
assign addr[31845]= 1356798326;
assign addr[31846]= 1579409630;
assign addr[31847]= 1770014111;
assign addr[31848]= 1924749160;
assign addr[31849]= 2040479063;
assign addr[31850]= 2114858546;
assign addr[31851]= 2146380306;
assign addr[31852]= 2134405552;
assign addr[31853]= 2079176953;
assign addr[31854]= 1981813720;
assign addr[31855]= 1844288924;
assign addr[31856]= 1669389513;
assign addr[31857]= 1460659832;
assign addr[31858]= 1222329801;
assign addr[31859]= 959229189;
assign addr[31860]= 676689746;
assign addr[31861]= 380437148;
assign addr[31862]= 76474970;
assign addr[31863]= -229036977;
assign addr[31864]= -529907477;
assign addr[31865]= -820039373;
assign addr[31866]= -1093553126;
assign addr[31867]= -1344905966;
assign addr[31868]= -1569004214;
assign addr[31869]= -1761306505;
assign addr[31870]= -1917915825;
assign addr[31871]= -2035658475;
assign addr[31872]= -2112148396;
assign addr[31873]= -2145835515;
assign addr[31874]= -2136037160;
assign addr[31875]= -2082951896;
assign addr[31876]= -1987655498;
assign addr[31877]= -1852079154;
assign addr[31878]= -1678970324;
assign addr[31879]= -1471837070;
assign addr[31880]= -1234876957;
assign addr[31881]= -972891995;
assign addr[31882]= -691191324;
assign addr[31883]= -395483624;
assign addr[31884]= -91761426;
assign addr[31885]= 213820322;
assign addr[31886]= 515068990;
assign addr[31887]= 805879757;
assign addr[31888]= 1080359326;
assign addr[31889]= 1332945355;
assign addr[31890]= 1558519173;
assign addr[31891]= 1752509516;
assign addr[31892]= 1910985158;
assign addr[31893]= 2030734582;
assign addr[31894]= 2109331059;
assign addr[31895]= 2145181827;
assign addr[31896]= 2137560369;
assign addr[31897]= 2086621133;
assign addr[31898]= 1993396407;
assign addr[31899]= 1859775393;
assign addr[31900]= 1688465931;
assign addr[31901]= 1482939614;
assign addr[31902]= 1247361445;
assign addr[31903]= 986505429;
assign addr[31904]= 705657826;
assign addr[31905]= 410510029;
assign addr[31906]= 107043224;
assign addr[31907]= -198592817;
assign addr[31908]= -500204365;
assign addr[31909]= -791679244;
assign addr[31910]= -1067110699;
assign addr[31911]= -1320917099;
assign addr[31912]= -1547955041;
assign addr[31913]= -1743623590;
assign addr[31914]= -1903957513;
assign addr[31915]= -2025707632;
assign addr[31916]= -2106406677;
assign addr[31917]= -2144419275;
assign addr[31918]= -2138975100;
assign addr[31919]= -2090184478;
assign addr[31920]= -1999036154;
assign addr[31921]= -1867377253;
assign addr[31922]= -1697875851;
assign addr[31923]= -1493966902;
assign addr[31924]= -1259782632;
assign addr[31925]= -1000068799;
assign addr[31926]= -720088517;
assign addr[31927]= -425515602;
assign addr[31928]= -122319591;
assign addr[31929]= 183355234;
assign addr[31930]= 485314355;
assign addr[31931]= 777438554;
assign addr[31932]= 1053807919;
assign addr[31933]= 1308821808;
assign addr[31934]= 1537312353;
assign addr[31935]= 1734649179;
assign addr[31936]= 1896833245;
assign addr[31937]= 2020577882;
assign addr[31938]= 2103375398;
assign addr[31939]= 2143547897;
assign addr[31940]= 2140281282;
assign addr[31941]= 2093641749;
assign addr[31942]= 2004574453;
assign addr[31943]= 1874884346;
assign addr[31944]= 1707199606;
assign addr[31945]= 1504918373;
assign addr[31946]= 1272139887;
assign addr[31947]= 1013581418;
assign addr[31948]= 734482665;
assign addr[31949]= 440499581;
assign addr[31950]= 137589750;
assign addr[31951]= -168108346;
assign addr[31952]= -470399716;
assign addr[31953]= -763158411;
assign addr[31954]= -1040451659;
assign addr[31955]= -1296660098;
assign addr[31956]= -1526591649;
assign addr[31957]= -1725586737;
assign addr[31958]= -1889612716;
assign addr[31959]= -2015345591;
assign addr[31960]= -2100237377;
assign addr[31961]= -2142567738;
assign addr[31962]= -2141478848;
assign addr[31963]= -2096992772;
assign addr[31964]= -2010011024;
assign addr[31965]= -1882296293;
assign addr[31966]= -1716436725;
assign addr[31967]= -1515793473;
assign addr[31968]= -1284432584;
assign addr[31969]= -1027042599;
assign addr[31970]= -748839539;
assign addr[31971]= -455461206;
assign addr[31972]= -152852926;
assign addr[31973]= 152852926;
assign addr[31974]= 455461206;
assign addr[31975]= 748839539;
assign addr[31976]= 1027042599;
assign addr[31977]= 1284432584;
assign addr[31978]= 1515793473;
assign addr[31979]= 1716436725;
assign addr[31980]= 1882296293;
assign addr[31981]= 2010011024;
assign addr[31982]= 2096992772;
assign addr[31983]= 2141478848;
assign addr[31984]= 2142567738;
assign addr[31985]= 2100237377;
assign addr[31986]= 2015345591;
assign addr[31987]= 1889612716;
assign addr[31988]= 1725586737;
assign addr[31989]= 1526591649;
assign addr[31990]= 1296660098;
assign addr[31991]= 1040451659;
assign addr[31992]= 763158411;
assign addr[31993]= 470399716;
assign addr[31994]= 168108346;
assign addr[31995]= -137589750;
assign addr[31996]= -440499581;
assign addr[31997]= -734482665;
assign addr[31998]= -1013581418;
assign addr[31999]= -1272139887;
assign addr[32000]= -1504918373;
assign addr[32001]= -1707199606;
assign addr[32002]= -1874884346;
assign addr[32003]= -2004574453;
assign addr[32004]= -2093641749;
assign addr[32005]= -2140281282;
assign addr[32006]= -2143547897;
assign addr[32007]= -2103375398;
assign addr[32008]= -2020577882;
assign addr[32009]= -1896833245;
assign addr[32010]= -1734649179;
assign addr[32011]= -1537312353;
assign addr[32012]= -1308821808;
assign addr[32013]= -1053807919;
assign addr[32014]= -777438554;
assign addr[32015]= -485314355;
assign addr[32016]= -183355234;
assign addr[32017]= 122319591;
assign addr[32018]= 425515602;
assign addr[32019]= 720088517;
assign addr[32020]= 1000068799;
assign addr[32021]= 1259782632;
assign addr[32022]= 1493966902;
assign addr[32023]= 1697875851;
assign addr[32024]= 1867377253;
assign addr[32025]= 1999036154;
assign addr[32026]= 2090184478;
assign addr[32027]= 2138975100;
assign addr[32028]= 2144419275;
assign addr[32029]= 2106406677;
assign addr[32030]= 2025707632;
assign addr[32031]= 1903957513;
assign addr[32032]= 1743623590;
assign addr[32033]= 1547955041;
assign addr[32034]= 1320917099;
assign addr[32035]= 1067110699;
assign addr[32036]= 791679244;
assign addr[32037]= 500204365;
assign addr[32038]= 198592817;
assign addr[32039]= -107043224;
assign addr[32040]= -410510029;
assign addr[32041]= -705657826;
assign addr[32042]= -986505429;
assign addr[32043]= -1247361445;
assign addr[32044]= -1482939614;
assign addr[32045]= -1688465931;
assign addr[32046]= -1859775393;
assign addr[32047]= -1993396407;
assign addr[32048]= -2086621133;
assign addr[32049]= -2137560369;
assign addr[32050]= -2145181827;
assign addr[32051]= -2109331059;
assign addr[32052]= -2030734582;
assign addr[32053]= -1910985158;
assign addr[32054]= -1752509516;
assign addr[32055]= -1558519173;
assign addr[32056]= -1332945355;
assign addr[32057]= -1080359326;
assign addr[32058]= -805879757;
assign addr[32059]= -515068990;
assign addr[32060]= -213820322;
assign addr[32061]= 91761426;
assign addr[32062]= 395483624;
assign addr[32063]= 691191324;
assign addr[32064]= 972891995;
assign addr[32065]= 1234876957;
assign addr[32066]= 1471837070;
assign addr[32067]= 1678970324;
assign addr[32068]= 1852079154;
assign addr[32069]= 1987655498;
assign addr[32070]= 2082951896;
assign addr[32071]= 2136037160;
assign addr[32072]= 2145835515;
assign addr[32073]= 2112148396;
assign addr[32074]= 2035658475;
assign addr[32075]= 1917915825;
assign addr[32076]= 1761306505;
assign addr[32077]= 1569004214;
assign addr[32078]= 1344905966;
assign addr[32079]= 1093553126;
assign addr[32080]= 820039373;
assign addr[32081]= 529907477;
assign addr[32082]= 229036977;
assign addr[32083]= -76474970;
assign addr[32084]= -380437148;
assign addr[32085]= -676689746;
assign addr[32086]= -959229189;
assign addr[32087]= -1222329801;
assign addr[32088]= -1460659832;
assign addr[32089]= -1669389513;
assign addr[32090]= -1844288924;
assign addr[32091]= -1981813720;
assign addr[32092]= -2079176953;
assign addr[32093]= -2134405552;
assign addr[32094]= -2146380306;
assign addr[32095]= -2114858546;
assign addr[32096]= -2040479063;
assign addr[32097]= -1924749160;
assign addr[32098]= -1770014111;
assign addr[32099]= -1579409630;
assign addr[32100]= -1356798326;
assign addr[32101]= -1106691431;
assign addr[32102]= -834157373;
assign addr[32103]= -544719071;
assign addr[32104]= -244242007;
assign addr[32105]= 61184634;
assign addr[32106]= 365371365;
assign addr[32107]= 662153826;
assign addr[32108]= 945517704;
assign addr[32109]= 1209720613;
assign addr[32110]= 1449408469;
assign addr[32111]= 1659723983;
assign addr[32112]= 1836405100;
assign addr[32113]= 1975871368;
assign addr[32114]= 2075296495;
assign addr[32115]= 2132665626;
assign addr[32116]= 2146816171;
assign addr[32117]= 2117461370;
assign addr[32118]= 2045196100;
assign addr[32119]= 1931484818;
assign addr[32120]= 1778631892;
assign addr[32121]= 1589734894;
assign addr[32122]= 1368621831;
assign addr[32123]= 1119773573;
assign addr[32124]= 848233042;
assign addr[32125]= 559503022;
assign addr[32126]= 259434643;
assign addr[32127]= -45891193;
assign addr[32128]= -350287041;
assign addr[32129]= -647584304;
assign addr[32130]= -931758235;
assign addr[32131]= -1197050035;
assign addr[32132]= -1438083551;
assign addr[32133]= -1649974225;
assign addr[32134]= -1828428082;
assign addr[32135]= -1969828744;
assign addr[32136]= -2071310720;
assign addr[32137]= -2130817471;
assign addr[32138]= -2147143090;
assign addr[32139]= -2119956737;
assign addr[32140]= -2049809346;
assign addr[32141]= -1938122457;
assign addr[32142]= -1787159411;
assign addr[32143]= -1599979481;
assign addr[32144]= -1380375881;
assign addr[32145]= -1132798888;
assign addr[32146]= -862265664;
assign addr[32147]= -574258580;
assign addr[32148]= -274614114;
assign addr[32149]= 30595422;
assign addr[32150]= 335184940;
assign addr[32151]= 632981917;
assign addr[32152]= 917951481;
assign addr[32153]= 1184318708;
assign addr[32154]= 1426685652;
assign addr[32155]= 1640140734;
assign addr[32156]= 1820358275;
assign addr[32157]= 1963686155;
assign addr[32158]= 2067219829;
assign addr[32159]= 2128861181;
assign addr[32160]= 2147361045;
assign addr[32161]= 2122344521;
assign addr[32162]= 2054318569;
assign addr[32163]= 1944661739;
assign addr[32164]= 1795596234;
assign addr[32165]= 1610142873;
assign addr[32166]= 1392059879;
assign addr[32167]= 1145766716;
assign addr[32168]= 876254528;
assign addr[32169]= 588984994;
assign addr[32170]= 289779648;
assign addr[32171]= -15298099;
assign addr[32172]= -320065829;
assign addr[32173]= -618347408;
assign addr[32174]= -904098143;
assign addr[32175]= -1171527280;
assign addr[32176]= -1415215352;
assign addr[32177]= -1630224009;
assign addr[32178]= -1812196087;
assign addr[32179]= -1957443913;
assign addr[32180]= -2063024031;
assign addr[32181]= -2126796855;
assign addr[32182]= -2147470025;
assign addr[32183]= -2124624598;
assign addr[32184]= -2058723538;
assign addr[32185]= -1951102334;
assign addr[32186]= -1803941934;
assign addr[32187]= -1620224553;
assign addr[32188]= -1403673233;
assign addr[32189]= -1158676398;
assign addr[32190]= -890198924;
assign addr[32191]= -603681519;
assign addr[32192]= -304930476;
assign addr[32193]= 0;
assign addr[32194]= 304930476;
assign addr[32195]= 603681519;
assign addr[32196]= 890198924;
assign addr[32197]= 1158676398;
assign addr[32198]= 1403673233;
assign addr[32199]= 1620224553;
assign addr[32200]= 1803941934;
assign addr[32201]= 1951102334;
assign addr[32202]= 2058723538;
assign addr[32203]= 2124624598;
assign addr[32204]= 2147470025;
assign addr[32205]= 2126796855;
assign addr[32206]= 2063024031;
assign addr[32207]= 1957443913;
assign addr[32208]= 1812196087;
assign addr[32209]= 1630224009;
assign addr[32210]= 1415215352;
assign addr[32211]= 1171527280;
assign addr[32212]= 904098143;
assign addr[32213]= 618347408;
assign addr[32214]= 320065829;
assign addr[32215]= 15298099;
assign addr[32216]= -289779648;
assign addr[32217]= -588984994;
assign addr[32218]= -876254528;
assign addr[32219]= -1145766716;
assign addr[32220]= -1392059879;
assign addr[32221]= -1610142873;
assign addr[32222]= -1795596234;
assign addr[32223]= -1944661739;
assign addr[32224]= -2054318569;
assign addr[32225]= -2122344521;
assign addr[32226]= -2147361045;
assign addr[32227]= -2128861181;
assign addr[32228]= -2067219829;
assign addr[32229]= -1963686155;
assign addr[32230]= -1820358275;
assign addr[32231]= -1640140734;
assign addr[32232]= -1426685652;
assign addr[32233]= -1184318708;
assign addr[32234]= -917951481;
assign addr[32235]= -632981917;
assign addr[32236]= -335184940;
assign addr[32237]= -30595422;
assign addr[32238]= 274614114;
assign addr[32239]= 574258580;
assign addr[32240]= 862265664;
assign addr[32241]= 1132798888;
assign addr[32242]= 1380375881;
assign addr[32243]= 1599979481;
assign addr[32244]= 1787159411;
assign addr[32245]= 1938122457;
assign addr[32246]= 2049809346;
assign addr[32247]= 2119956737;
assign addr[32248]= 2147143090;
assign addr[32249]= 2130817471;
assign addr[32250]= 2071310720;
assign addr[32251]= 1969828744;
assign addr[32252]= 1828428082;
assign addr[32253]= 1649974225;
assign addr[32254]= 1438083551;
assign addr[32255]= 1197050035;
assign addr[32256]= 931758235;
assign addr[32257]= 647584304;
assign addr[32258]= 350287041;
assign addr[32259]= 45891193;
assign addr[32260]= -259434643;
assign addr[32261]= -559503022;
assign addr[32262]= -848233042;
assign addr[32263]= -1119773573;
assign addr[32264]= -1368621831;
assign addr[32265]= -1589734894;
assign addr[32266]= -1778631892;
assign addr[32267]= -1931484818;
assign addr[32268]= -2045196100;
assign addr[32269]= -2117461370;
assign addr[32270]= -2146816171;
assign addr[32271]= -2132665626;
assign addr[32272]= -2075296495;
assign addr[32273]= -1975871368;
assign addr[32274]= -1836405100;
assign addr[32275]= -1659723983;
assign addr[32276]= -1449408469;
assign addr[32277]= -1209720613;
assign addr[32278]= -945517704;
assign addr[32279]= -662153826;
assign addr[32280]= -365371365;
assign addr[32281]= -61184634;
assign addr[32282]= 244242007;
assign addr[32283]= 544719071;
assign addr[32284]= 834157373;
assign addr[32285]= 1106691431;
assign addr[32286]= 1356798326;
assign addr[32287]= 1579409630;
assign addr[32288]= 1770014111;
assign addr[32289]= 1924749160;
assign addr[32290]= 2040479063;
assign addr[32291]= 2114858546;
assign addr[32292]= 2146380306;
assign addr[32293]= 2134405552;
assign addr[32294]= 2079176953;
assign addr[32295]= 1981813720;
assign addr[32296]= 1844288924;
assign addr[32297]= 1669389513;
assign addr[32298]= 1460659832;
assign addr[32299]= 1222329801;
assign addr[32300]= 959229189;
assign addr[32301]= 676689746;
assign addr[32302]= 380437148;
assign addr[32303]= 76474970;
assign addr[32304]= -229036977;
assign addr[32305]= -529907477;
assign addr[32306]= -820039373;
assign addr[32307]= -1093553126;
assign addr[32308]= -1344905966;
assign addr[32309]= -1569004214;
assign addr[32310]= -1761306505;
assign addr[32311]= -1917915825;
assign addr[32312]= -2035658475;
assign addr[32313]= -2112148396;
assign addr[32314]= -2145835515;
assign addr[32315]= -2136037160;
assign addr[32316]= -2082951896;
assign addr[32317]= -1987655498;
assign addr[32318]= -1852079154;
assign addr[32319]= -1678970324;
assign addr[32320]= -1471837070;
assign addr[32321]= -1234876957;
assign addr[32322]= -972891995;
assign addr[32323]= -691191324;
assign addr[32324]= -395483624;
assign addr[32325]= -91761426;
assign addr[32326]= 213820322;
assign addr[32327]= 515068990;
assign addr[32328]= 805879757;
assign addr[32329]= 1080359326;
assign addr[32330]= 1332945355;
assign addr[32331]= 1558519173;
assign addr[32332]= 1752509516;
assign addr[32333]= 1910985158;
assign addr[32334]= 2030734582;
assign addr[32335]= 2109331059;
assign addr[32336]= 2145181827;
assign addr[32337]= 2137560369;
assign addr[32338]= 2086621133;
assign addr[32339]= 1993396407;
assign addr[32340]= 1859775393;
assign addr[32341]= 1688465931;
assign addr[32342]= 1482939614;
assign addr[32343]= 1247361445;
assign addr[32344]= 986505429;
assign addr[32345]= 705657826;
assign addr[32346]= 410510029;
assign addr[32347]= 107043224;
assign addr[32348]= -198592817;
assign addr[32349]= -500204365;
assign addr[32350]= -791679244;
assign addr[32351]= -1067110699;
assign addr[32352]= -1320917099;
assign addr[32353]= -1547955041;
assign addr[32354]= -1743623590;
assign addr[32355]= -1903957513;
assign addr[32356]= -2025707632;
assign addr[32357]= -2106406677;
assign addr[32358]= -2144419275;
assign addr[32359]= -2138975100;
assign addr[32360]= -2090184478;
assign addr[32361]= -1999036154;
assign addr[32362]= -1867377253;
assign addr[32363]= -1697875851;
assign addr[32364]= -1493966902;
assign addr[32365]= -1259782632;
assign addr[32366]= -1000068799;
assign addr[32367]= -720088517;
assign addr[32368]= -425515602;
assign addr[32369]= -122319591;
assign addr[32370]= 183355234;
assign addr[32371]= 485314355;
assign addr[32372]= 777438554;
assign addr[32373]= 1053807919;
assign addr[32374]= 1308821808;
assign addr[32375]= 1537312353;
assign addr[32376]= 1734649179;
assign addr[32377]= 1896833245;
assign addr[32378]= 2020577882;
assign addr[32379]= 2103375398;
assign addr[32380]= 2143547897;
assign addr[32381]= 2140281282;
assign addr[32382]= 2093641749;
assign addr[32383]= 2004574453;
assign addr[32384]= 1874884346;
assign addr[32385]= 1707199606;
assign addr[32386]= 1504918373;
assign addr[32387]= 1272139887;
assign addr[32388]= 1013581418;
assign addr[32389]= 734482665;
assign addr[32390]= 440499581;
assign addr[32391]= 137589750;
assign addr[32392]= -168108346;
assign addr[32393]= -470399716;
assign addr[32394]= -763158411;
assign addr[32395]= -1040451659;
assign addr[32396]= -1296660098;
assign addr[32397]= -1526591649;
assign addr[32398]= -1725586737;
assign addr[32399]= -1889612716;
assign addr[32400]= -2015345591;
assign addr[32401]= -2100237377;
assign addr[32402]= -2142567738;
assign addr[32403]= -2141478848;
assign addr[32404]= -2096992772;
assign addr[32405]= -2010011024;
assign addr[32406]= -1882296293;
assign addr[32407]= -1716436725;
assign addr[32408]= -1515793473;
assign addr[32409]= -1284432584;
assign addr[32410]= -1027042599;
assign addr[32411]= -748839539;
assign addr[32412]= -455461206;
assign addr[32413]= -152852926;
assign addr[32414]= 152852926;
assign addr[32415]= 455461206;
assign addr[32416]= 748839539;
assign addr[32417]= 1027042599;
assign addr[32418]= 1284432584;
assign addr[32419]= 1515793473;
assign addr[32420]= 1716436725;
assign addr[32421]= 1882296293;
assign addr[32422]= 2010011024;
assign addr[32423]= 2096992772;
assign addr[32424]= 2141478848;
assign addr[32425]= 2142567738;
assign addr[32426]= 2100237377;
assign addr[32427]= 2015345591;
assign addr[32428]= 1889612716;
assign addr[32429]= 1725586737;
assign addr[32430]= 1526591649;
assign addr[32431]= 1296660098;
assign addr[32432]= 1040451659;
assign addr[32433]= 763158411;
assign addr[32434]= 470399716;
assign addr[32435]= 168108346;
assign addr[32436]= -137589750;
assign addr[32437]= -440499581;
assign addr[32438]= -734482665;
assign addr[32439]= -1013581418;
assign addr[32440]= -1272139887;
assign addr[32441]= -1504918373;
assign addr[32442]= -1707199606;
assign addr[32443]= -1874884346;
assign addr[32444]= -2004574453;
assign addr[32445]= -2093641749;
assign addr[32446]= -2140281282;
assign addr[32447]= -2143547897;
assign addr[32448]= -2103375398;
assign addr[32449]= -2020577882;
assign addr[32450]= -1896833245;
assign addr[32451]= -1734649179;
assign addr[32452]= -1537312353;
assign addr[32453]= -1308821808;
assign addr[32454]= -1053807919;
assign addr[32455]= -777438554;
assign addr[32456]= -485314355;
assign addr[32457]= -183355234;
assign addr[32458]= 122319591;
assign addr[32459]= 425515602;
assign addr[32460]= 720088517;
assign addr[32461]= 1000068799;
assign addr[32462]= 1259782632;
assign addr[32463]= 1493966902;
assign addr[32464]= 1697875851;
assign addr[32465]= 1867377253;
assign addr[32466]= 1999036154;
assign addr[32467]= 2090184478;
assign addr[32468]= 2138975100;
assign addr[32469]= 2144419275;
assign addr[32470]= 2106406677;
assign addr[32471]= 2025707632;
assign addr[32472]= 1903957513;
assign addr[32473]= 1743623590;
assign addr[32474]= 1547955041;
assign addr[32475]= 1320917099;
assign addr[32476]= 1067110699;
assign addr[32477]= 791679244;
assign addr[32478]= 500204365;
assign addr[32479]= 198592817;
assign addr[32480]= -107043224;
assign addr[32481]= -410510029;
assign addr[32482]= -705657826;
assign addr[32483]= -986505429;
assign addr[32484]= -1247361445;
assign addr[32485]= -1482939614;
assign addr[32486]= -1688465931;
assign addr[32487]= -1859775393;
assign addr[32488]= -1993396407;
assign addr[32489]= -2086621133;
assign addr[32490]= -2137560369;
assign addr[32491]= -2145181827;
assign addr[32492]= -2109331059;
assign addr[32493]= -2030734582;
assign addr[32494]= -1910985158;
assign addr[32495]= -1752509516;
assign addr[32496]= -1558519173;
assign addr[32497]= -1332945355;
assign addr[32498]= -1080359326;
assign addr[32499]= -805879757;
assign addr[32500]= -515068990;
assign addr[32501]= -213820322;
assign addr[32502]= 91761426;
assign addr[32503]= 395483624;
assign addr[32504]= 691191324;
assign addr[32505]= 972891995;
assign addr[32506]= 1234876957;
assign addr[32507]= 1471837070;
assign addr[32508]= 1678970324;
assign addr[32509]= 1852079154;
assign addr[32510]= 1987655498;
assign addr[32511]= 2082951896;
assign addr[32512]= 2136037160;
assign addr[32513]= 2145835515;
assign addr[32514]= 2112148396;
assign addr[32515]= 2035658475;
assign addr[32516]= 1917915825;
assign addr[32517]= 1761306505;
assign addr[32518]= 1569004214;
assign addr[32519]= 1344905966;
assign addr[32520]= 1093553126;
assign addr[32521]= 820039373;
assign addr[32522]= 529907477;
assign addr[32523]= 229036977;
assign addr[32524]= -76474970;
assign addr[32525]= -380437148;
assign addr[32526]= -676689746;
assign addr[32527]= -959229189;
assign addr[32528]= -1222329801;
assign addr[32529]= -1460659832;
assign addr[32530]= -1669389513;
assign addr[32531]= -1844288924;
assign addr[32532]= -1981813720;
assign addr[32533]= -2079176953;
assign addr[32534]= -2134405552;
assign addr[32535]= -2146380306;
assign addr[32536]= -2114858546;
assign addr[32537]= -2040479063;
assign addr[32538]= -1924749160;
assign addr[32539]= -1770014111;
assign addr[32540]= -1579409630;
assign addr[32541]= -1356798326;
assign addr[32542]= -1106691431;
assign addr[32543]= -834157373;
assign addr[32544]= -544719071;
assign addr[32545]= -244242007;
assign addr[32546]= 61184634;
assign addr[32547]= 365371365;
assign addr[32548]= 662153826;
assign addr[32549]= 945517704;
assign addr[32550]= 1209720613;
assign addr[32551]= 1449408469;
assign addr[32552]= 1659723983;
assign addr[32553]= 1836405100;
assign addr[32554]= 1975871368;
assign addr[32555]= 2075296495;
assign addr[32556]= 2132665626;
assign addr[32557]= 2146816171;
assign addr[32558]= 2117461370;
assign addr[32559]= 2045196100;
assign addr[32560]= 1931484818;
assign addr[32561]= 1778631892;
assign addr[32562]= 1589734894;
assign addr[32563]= 1368621831;
assign addr[32564]= 1119773573;
assign addr[32565]= 848233042;
assign addr[32566]= 559503022;
assign addr[32567]= 259434643;
assign addr[32568]= -45891193;
assign addr[32569]= -350287041;
assign addr[32570]= -647584304;
assign addr[32571]= -931758235;
assign addr[32572]= -1197050035;
assign addr[32573]= -1438083551;
assign addr[32574]= -1649974225;
assign addr[32575]= -1828428082;
assign addr[32576]= -1969828744;
assign addr[32577]= -2071310720;
assign addr[32578]= -2130817471;
assign addr[32579]= -2147143090;
assign addr[32580]= -2119956737;
assign addr[32581]= -2049809346;
assign addr[32582]= -1938122457;
assign addr[32583]= -1787159411;
assign addr[32584]= -1599979481;
assign addr[32585]= -1380375881;
assign addr[32586]= -1132798888;
assign addr[32587]= -862265664;
assign addr[32588]= -574258580;
assign addr[32589]= -274614114;
assign addr[32590]= 30595422;
assign addr[32591]= 335184940;
assign addr[32592]= 632981917;
assign addr[32593]= 917951481;
assign addr[32594]= 1184318708;
assign addr[32595]= 1426685652;
assign addr[32596]= 1640140734;
assign addr[32597]= 1820358275;
assign addr[32598]= 1963686155;
assign addr[32599]= 2067219829;
assign addr[32600]= 2128861181;
assign addr[32601]= 2147361045;
assign addr[32602]= 2122344521;
assign addr[32603]= 2054318569;
assign addr[32604]= 1944661739;
assign addr[32605]= 1795596234;
assign addr[32606]= 1610142873;
assign addr[32607]= 1392059879;
assign addr[32608]= 1145766716;
assign addr[32609]= 876254528;
assign addr[32610]= 588984994;
assign addr[32611]= 289779648;
assign addr[32612]= -15298099;
assign addr[32613]= -320065829;
assign addr[32614]= -618347408;
assign addr[32615]= -904098143;
assign addr[32616]= -1171527280;
assign addr[32617]= -1415215352;
assign addr[32618]= -1630224009;
assign addr[32619]= -1812196087;
assign addr[32620]= -1957443913;
assign addr[32621]= -2063024031;
assign addr[32622]= -2126796855;
assign addr[32623]= -2147470025;
assign addr[32624]= -2124624598;
assign addr[32625]= -2058723538;
assign addr[32626]= -1951102334;
assign addr[32627]= -1803941934;
assign addr[32628]= -1620224553;
assign addr[32629]= -1403673233;
assign addr[32630]= -1158676398;
assign addr[32631]= -890198924;
assign addr[32632]= -603681519;
assign addr[32633]= -304930476;
assign addr[32634]= 0;
assign addr[32635]= 304930476;
assign addr[32636]= 603681519;
assign addr[32637]= 890198924;
assign addr[32638]= 1158676398;
assign addr[32639]= 1403673233;
assign addr[32640]= 1620224553;
assign addr[32641]= 1803941934;
assign addr[32642]= 1951102334;
assign addr[32643]= 2058723538;
assign addr[32644]= 2124624598;
assign addr[32645]= 2147470025;
assign addr[32646]= 2126796855;
assign addr[32647]= 2063024031;
assign addr[32648]= 1957443913;
assign addr[32649]= 1812196087;
assign addr[32650]= 1630224009;
assign addr[32651]= 1415215352;
assign addr[32652]= 1171527280;
assign addr[32653]= 904098143;
assign addr[32654]= 618347408;
assign addr[32655]= 320065829;
assign addr[32656]= 15298099;
assign addr[32657]= -289779648;
assign addr[32658]= -588984994;
assign addr[32659]= -876254528;
assign addr[32660]= -1145766716;
assign addr[32661]= -1392059879;
assign addr[32662]= -1610142873;
assign addr[32663]= -1795596234;
assign addr[32664]= -1944661739;
assign addr[32665]= -2054318569;
assign addr[32666]= -2122344521;
assign addr[32667]= -2147361045;
assign addr[32668]= -2128861181;
assign addr[32669]= -2067219829;
assign addr[32670]= -1963686155;
assign addr[32671]= -1820358275;
assign addr[32672]= -1640140734;
assign addr[32673]= -1426685652;
assign addr[32674]= -1184318708;
assign addr[32675]= -917951481;
assign addr[32676]= -632981917;
assign addr[32677]= -335184940;
assign addr[32678]= -30595422;
assign addr[32679]= 274614114;
assign addr[32680]= 574258580;
assign addr[32681]= 862265664;
assign addr[32682]= 1132798888;
assign addr[32683]= 1380375881;
assign addr[32684]= 1599979481;
assign addr[32685]= 1787159411;
assign addr[32686]= 1938122457;
assign addr[32687]= 2049809346;
assign addr[32688]= 2119956737;
assign addr[32689]= 2147143090;
assign addr[32690]= 2130817471;
assign addr[32691]= 2071310720;
assign addr[32692]= 1969828744;
assign addr[32693]= 1828428082;
assign addr[32694]= 1649974225;
assign addr[32695]= 1438083551;
assign addr[32696]= 1197050035;
assign addr[32697]= 931758235;
assign addr[32698]= 647584304;
assign addr[32699]= 350287041;
assign addr[32700]= 45891193;
assign addr[32701]= -259434643;
assign addr[32702]= -559503022;
assign addr[32703]= -848233042;
assign addr[32704]= -1119773573;
assign addr[32705]= -1368621831;
assign addr[32706]= -1589734894;
assign addr[32707]= -1778631892;
assign addr[32708]= -1931484818;
assign addr[32709]= -2045196100;
assign addr[32710]= -2117461370;
assign addr[32711]= -2146816171;
assign addr[32712]= -2132665626;
assign addr[32713]= -2075296495;
assign addr[32714]= -1975871368;
assign addr[32715]= -1836405100;
assign addr[32716]= -1659723983;
assign addr[32717]= -1449408469;
assign addr[32718]= -1209720613;
assign addr[32719]= -945517704;
assign addr[32720]= -662153826;
assign addr[32721]= -365371365;
assign addr[32722]= -61184634;
assign addr[32723]= 244242007;
assign addr[32724]= 544719071;
assign addr[32725]= 834157373;
assign addr[32726]= 1106691431;
assign addr[32727]= 1356798326;
assign addr[32728]= 1579409630;
assign addr[32729]= 1770014111;
assign addr[32730]= 1924749160;
assign addr[32731]= 2040479063;
assign addr[32732]= 2114858546;
assign addr[32733]= 2146380306;
assign addr[32734]= 2134405552;
assign addr[32735]= 2079176953;
assign addr[32736]= 1981813720;
assign addr[32737]= 1844288924;
assign addr[32738]= 1669389513;
assign addr[32739]= 1460659832;
assign addr[32740]= 1222329801;
assign addr[32741]= 959229189;
assign addr[32742]= 676689746;
assign addr[32743]= 380437148;
assign addr[32744]= 76474970;
assign addr[32745]= -229036977;
assign addr[32746]= -529907477;
assign addr[32747]= -820039373;
assign addr[32748]= -1093553126;
assign addr[32749]= -1344905966;
assign addr[32750]= -1569004214;
assign addr[32751]= -1761306505;
assign addr[32752]= -1917915825;
assign addr[32753]= -2035658475;
assign addr[32754]= -2112148396;
assign addr[32755]= -2145835515;
assign addr[32756]= -2136037160;
assign addr[32757]= -2082951896;
assign addr[32758]= -1987655498;
assign addr[32759]= -1852079154;
assign addr[32760]= -1678970324;
assign addr[32761]= -1471837070;
assign addr[32762]= -1234876957;
assign addr[32763]= -972891995;
assign addr[32764]= -691191324;
assign addr[32765]= -395483624;
assign addr[32766]= -91761426;
assign addr[32767]= 213820322;
assign addr[32768]= 515068990;
assign addr[32769]= 805879757;
assign addr[32770]= 1080359326;
assign addr[32771]= 1332945355;
assign addr[32772]= 1558519173;
assign addr[32773]= 1752509516;
assign addr[32774]= 1910985158;
assign addr[32775]= 2030734582;
assign addr[32776]= 2109331059;
assign addr[32777]= 2145181827;
assign addr[32778]= 2137560369;
assign addr[32779]= 2086621133;
assign addr[32780]= 1993396407;
assign addr[32781]= 1859775393;
assign addr[32782]= 1688465931;
assign addr[32783]= 1482939614;
assign addr[32784]= 1247361445;
assign addr[32785]= 986505429;
assign addr[32786]= 705657826;
assign addr[32787]= 410510029;
assign addr[32788]= 107043224;
assign addr[32789]= -198592817;
assign addr[32790]= -500204365;
assign addr[32791]= -791679244;
assign addr[32792]= -1067110699;
assign addr[32793]= -1320917099;
assign addr[32794]= -1547955041;
assign addr[32795]= -1743623590;
assign addr[32796]= -1903957513;
assign addr[32797]= -2025707632;
assign addr[32798]= -2106406677;
assign addr[32799]= -2144419275;
assign addr[32800]= -2138975100;
assign addr[32801]= -2090184478;
assign addr[32802]= -1999036154;
assign addr[32803]= -1867377253;
assign addr[32804]= -1697875851;
assign addr[32805]= -1493966902;
assign addr[32806]= -1259782632;
assign addr[32807]= -1000068799;
assign addr[32808]= -720088517;
assign addr[32809]= -425515602;
assign addr[32810]= -122319591;
assign addr[32811]= 183355234;
assign addr[32812]= 485314355;
assign addr[32813]= 777438554;
assign addr[32814]= 1053807919;
assign addr[32815]= 1308821808;
assign addr[32816]= 1537312353;
assign addr[32817]= 1734649179;
assign addr[32818]= 1896833245;
assign addr[32819]= 2020577882;
assign addr[32820]= 2103375398;
assign addr[32821]= 2143547897;
assign addr[32822]= 2140281282;
assign addr[32823]= 2093641749;
assign addr[32824]= 2004574453;
assign addr[32825]= 1874884346;
assign addr[32826]= 1707199606;
assign addr[32827]= 1504918373;
assign addr[32828]= 1272139887;
assign addr[32829]= 1013581418;
assign addr[32830]= 734482665;
assign addr[32831]= 440499581;
assign addr[32832]= 137589750;
assign addr[32833]= -168108346;
assign addr[32834]= -470399716;
assign addr[32835]= -763158411;
assign addr[32836]= -1040451659;
assign addr[32837]= -1296660098;
assign addr[32838]= -1526591649;
assign addr[32839]= -1725586737;
assign addr[32840]= -1889612716;
assign addr[32841]= -2015345591;
assign addr[32842]= -2100237377;
assign addr[32843]= -2142567738;
assign addr[32844]= -2141478848;
assign addr[32845]= -2096992772;
assign addr[32846]= -2010011024;
assign addr[32847]= -1882296293;
assign addr[32848]= -1716436725;
assign addr[32849]= -1515793473;
assign addr[32850]= -1284432584;
assign addr[32851]= -1027042599;
assign addr[32852]= -748839539;
assign addr[32853]= -455461206;
assign addr[32854]= -152852926;
assign addr[32855]= 152852926;
assign addr[32856]= 455461206;
assign addr[32857]= 748839539;
assign addr[32858]= 1027042599;
assign addr[32859]= 1284432584;
assign addr[32860]= 1515793473;
assign addr[32861]= 1716436725;
assign addr[32862]= 1882296293;
assign addr[32863]= 2010011024;
assign addr[32864]= 2096992772;
assign addr[32865]= 2141478848;
assign addr[32866]= 2142567738;
assign addr[32867]= 2100237377;
assign addr[32868]= 2015345591;
assign addr[32869]= 1889612716;
assign addr[32870]= 1725586737;
assign addr[32871]= 1526591649;
assign addr[32872]= 1296660098;
assign addr[32873]= 1040451659;
assign addr[32874]= 763158411;
assign addr[32875]= 470399716;
assign addr[32876]= 168108346;
assign addr[32877]= -137589750;
assign addr[32878]= -440499581;
assign addr[32879]= -734482665;
assign addr[32880]= -1013581418;
assign addr[32881]= -1272139887;
assign addr[32882]= -1504918373;
assign addr[32883]= -1707199606;
assign addr[32884]= -1874884346;
assign addr[32885]= -2004574453;
assign addr[32886]= -2093641749;
assign addr[32887]= -2140281282;
assign addr[32888]= -2143547897;
assign addr[32889]= -2103375398;
assign addr[32890]= -2020577882;
assign addr[32891]= -1896833245;
assign addr[32892]= -1734649179;
assign addr[32893]= -1537312353;
assign addr[32894]= -1308821808;
assign addr[32895]= -1053807919;
assign addr[32896]= -777438554;
assign addr[32897]= -485314355;
assign addr[32898]= -183355234;
assign addr[32899]= 122319591;
assign addr[32900]= 425515602;
assign addr[32901]= 720088517;
assign addr[32902]= 1000068799;
assign addr[32903]= 1259782632;
assign addr[32904]= 1493966902;
assign addr[32905]= 1697875851;
assign addr[32906]= 1867377253;
assign addr[32907]= 1999036154;
assign addr[32908]= 2090184478;
assign addr[32909]= 2138975100;
assign addr[32910]= 2144419275;
assign addr[32911]= 2106406677;
assign addr[32912]= 2025707632;
assign addr[32913]= 1903957513;
assign addr[32914]= 1743623590;
assign addr[32915]= 1547955041;
assign addr[32916]= 1320917099;
assign addr[32917]= 1067110699;
assign addr[32918]= 791679244;
assign addr[32919]= 500204365;
assign addr[32920]= 198592817;
assign addr[32921]= -107043224;
assign addr[32922]= -410510029;
assign addr[32923]= -705657826;
assign addr[32924]= -986505429;
assign addr[32925]= -1247361445;
assign addr[32926]= -1482939614;
assign addr[32927]= -1688465931;
assign addr[32928]= -1859775393;
assign addr[32929]= -1993396407;
assign addr[32930]= -2086621133;
assign addr[32931]= -2137560369;
assign addr[32932]= -2145181827;
assign addr[32933]= -2109331059;
assign addr[32934]= -2030734582;
assign addr[32935]= -1910985158;
assign addr[32936]= -1752509516;
assign addr[32937]= -1558519173;
assign addr[32938]= -1332945355;
assign addr[32939]= -1080359326;
assign addr[32940]= -805879757;
assign addr[32941]= -515068990;
assign addr[32942]= -213820322;
assign addr[32943]= 91761426;
assign addr[32944]= 395483624;
assign addr[32945]= 691191324;
assign addr[32946]= 972891995;
assign addr[32947]= 1234876957;
assign addr[32948]= 1471837070;
assign addr[32949]= 1678970324;
assign addr[32950]= 1852079154;
assign addr[32951]= 1987655498;
assign addr[32952]= 2082951896;
assign addr[32953]= 2136037160;
assign addr[32954]= 2145835515;
assign addr[32955]= 2112148396;
assign addr[32956]= 2035658475;
assign addr[32957]= 1917915825;
assign addr[32958]= 1761306505;
assign addr[32959]= 1569004214;
assign addr[32960]= 1344905966;
assign addr[32961]= 1093553126;
assign addr[32962]= 820039373;
assign addr[32963]= 529907477;
assign addr[32964]= 229036977;
assign addr[32965]= -76474970;
assign addr[32966]= -380437148;
assign addr[32967]= -676689746;
assign addr[32968]= -959229189;
assign addr[32969]= -1222329801;
assign addr[32970]= -1460659832;
assign addr[32971]= -1669389513;
assign addr[32972]= -1844288924;
assign addr[32973]= -1981813720;
assign addr[32974]= -2079176953;
assign addr[32975]= -2134405552;
assign addr[32976]= -2146380306;
assign addr[32977]= -2114858546;
assign addr[32978]= -2040479063;
assign addr[32979]= -1924749160;
assign addr[32980]= -1770014111;
assign addr[32981]= -1579409630;
assign addr[32982]= -1356798326;
assign addr[32983]= -1106691431;
assign addr[32984]= -834157373;
assign addr[32985]= -544719071;
assign addr[32986]= -244242007;
assign addr[32987]= 61184634;
assign addr[32988]= 365371365;
assign addr[32989]= 662153826;
assign addr[32990]= 945517704;
assign addr[32991]= 1209720613;
assign addr[32992]= 1449408469;
assign addr[32993]= 1659723983;
assign addr[32994]= 1836405100;
assign addr[32995]= 1975871368;
assign addr[32996]= 2075296495;
assign addr[32997]= 2132665626;
assign addr[32998]= 2146816171;
assign addr[32999]= 2117461370;
assign addr[33000]= 2045196100;
assign addr[33001]= 1931484818;
assign addr[33002]= 1778631892;
assign addr[33003]= 1589734894;
assign addr[33004]= 1368621831;
assign addr[33005]= 1119773573;
assign addr[33006]= 848233042;
assign addr[33007]= 559503022;
assign addr[33008]= 259434643;
assign addr[33009]= -45891193;
assign addr[33010]= -350287041;
assign addr[33011]= -647584304;
assign addr[33012]= -931758235;
assign addr[33013]= -1197050035;
assign addr[33014]= -1438083551;
assign addr[33015]= -1649974225;
assign addr[33016]= -1828428082;
assign addr[33017]= -1969828744;
assign addr[33018]= -2071310720;
assign addr[33019]= -2130817471;
assign addr[33020]= -2147143090;
assign addr[33021]= -2119956737;
assign addr[33022]= -2049809346;
assign addr[33023]= -1938122457;
assign addr[33024]= -1787159411;
assign addr[33025]= -1599979481;
assign addr[33026]= -1380375881;
assign addr[33027]= -1132798888;
assign addr[33028]= -862265664;
assign addr[33029]= -574258580;
assign addr[33030]= -274614114;
assign addr[33031]= 30595422;
assign addr[33032]= 335184940;
assign addr[33033]= 632981917;
assign addr[33034]= 917951481;
assign addr[33035]= 1184318708;
assign addr[33036]= 1426685652;
assign addr[33037]= 1640140734;
assign addr[33038]= 1820358275;
assign addr[33039]= 1963686155;
assign addr[33040]= 2067219829;
assign addr[33041]= 2128861181;
assign addr[33042]= 2147361045;
assign addr[33043]= 2122344521;
assign addr[33044]= 2054318569;
assign addr[33045]= 1944661739;
assign addr[33046]= 1795596234;
assign addr[33047]= 1610142873;
assign addr[33048]= 1392059879;
assign addr[33049]= 1145766716;
assign addr[33050]= 876254528;
assign addr[33051]= 588984994;
assign addr[33052]= 289779648;
assign addr[33053]= -15298099;
assign addr[33054]= -320065829;
assign addr[33055]= -618347408;
assign addr[33056]= -904098143;
assign addr[33057]= -1171527280;
assign addr[33058]= -1415215352;
assign addr[33059]= -1630224009;
assign addr[33060]= -1812196087;
assign addr[33061]= -1957443913;
assign addr[33062]= -2063024031;
assign addr[33063]= -2126796855;
assign addr[33064]= -2147470025;
assign addr[33065]= -2124624598;
assign addr[33066]= -2058723538;
assign addr[33067]= -1951102334;
assign addr[33068]= -1803941934;
assign addr[33069]= -1620224553;
assign addr[33070]= -1403673233;
assign addr[33071]= -1158676398;
assign addr[33072]= -890198924;
assign addr[33073]= -603681519;
assign addr[33074]= -304930476;
assign addr[33075]= 0;
assign addr[33076]= 304930476;
assign addr[33077]= 603681519;
assign addr[33078]= 890198924;
assign addr[33079]= 1158676398;
assign addr[33080]= 1403673233;
assign addr[33081]= 1620224553;
assign addr[33082]= 1803941934;
assign addr[33083]= 1951102334;
assign addr[33084]= 2058723538;
assign addr[33085]= 2124624598;
assign addr[33086]= 2147470025;
assign addr[33087]= 2126796855;
assign addr[33088]= 2063024031;
assign addr[33089]= 1957443913;
assign addr[33090]= 1812196087;
assign addr[33091]= 1630224009;
assign addr[33092]= 1415215352;
assign addr[33093]= 1171527280;
assign addr[33094]= 904098143;
assign addr[33095]= 618347408;
assign addr[33096]= 320065829;
assign addr[33097]= 15298099;
assign addr[33098]= -289779648;
assign addr[33099]= -588984994;
assign addr[33100]= -876254528;
assign addr[33101]= -1145766716;
assign addr[33102]= -1392059879;
assign addr[33103]= -1610142873;
assign addr[33104]= -1795596234;
assign addr[33105]= -1944661739;
assign addr[33106]= -2054318569;
assign addr[33107]= -2122344521;
assign addr[33108]= -2147361045;
assign addr[33109]= -2128861181;
assign addr[33110]= -2067219829;
assign addr[33111]= -1963686155;
assign addr[33112]= -1820358275;
assign addr[33113]= -1640140734;
assign addr[33114]= -1426685652;
assign addr[33115]= -1184318708;
assign addr[33116]= -917951481;
assign addr[33117]= -632981917;
assign addr[33118]= -335184940;
assign addr[33119]= -30595422;
assign addr[33120]= 274614114;
assign addr[33121]= 574258580;
assign addr[33122]= 862265664;
assign addr[33123]= 1132798888;
assign addr[33124]= 1380375881;
assign addr[33125]= 1599979481;
assign addr[33126]= 1787159411;
assign addr[33127]= 1938122457;
assign addr[33128]= 2049809346;
assign addr[33129]= 2119956737;
assign addr[33130]= 2147143090;
assign addr[33131]= 2130817471;
assign addr[33132]= 2071310720;
assign addr[33133]= 1969828744;
assign addr[33134]= 1828428082;
assign addr[33135]= 1649974225;
assign addr[33136]= 1438083551;
assign addr[33137]= 1197050035;
assign addr[33138]= 931758235;
assign addr[33139]= 647584304;
assign addr[33140]= 350287041;
assign addr[33141]= 45891193;
assign addr[33142]= -259434643;
assign addr[33143]= -559503022;
assign addr[33144]= -848233042;
assign addr[33145]= -1119773573;
assign addr[33146]= -1368621831;
assign addr[33147]= -1589734894;
assign addr[33148]= -1778631892;
assign addr[33149]= -1931484818;
assign addr[33150]= -2045196100;
assign addr[33151]= -2117461370;
assign addr[33152]= -2146816171;
assign addr[33153]= -2132665626;
assign addr[33154]= -2075296495;
assign addr[33155]= -1975871368;
assign addr[33156]= -1836405100;
assign addr[33157]= -1659723983;
assign addr[33158]= -1449408469;
assign addr[33159]= -1209720613;
assign addr[33160]= -945517704;
assign addr[33161]= -662153826;
assign addr[33162]= -365371365;
assign addr[33163]= -61184634;
assign addr[33164]= 244242007;
assign addr[33165]= 544719071;
assign addr[33166]= 834157373;
assign addr[33167]= 1106691431;
assign addr[33168]= 1356798326;
assign addr[33169]= 1579409630;
assign addr[33170]= 1770014111;
assign addr[33171]= 1924749160;
assign addr[33172]= 2040479063;
assign addr[33173]= 2114858546;
assign addr[33174]= 2146380306;
assign addr[33175]= 2134405552;
assign addr[33176]= 2079176953;
assign addr[33177]= 1981813720;
assign addr[33178]= 1844288924;
assign addr[33179]= 1669389513;
assign addr[33180]= 1460659832;
assign addr[33181]= 1222329801;
assign addr[33182]= 959229189;
assign addr[33183]= 676689746;
assign addr[33184]= 380437148;
assign addr[33185]= 76474970;
assign addr[33186]= -229036977;
assign addr[33187]= -529907477;
assign addr[33188]= -820039373;
assign addr[33189]= -1093553126;
assign addr[33190]= -1344905966;
assign addr[33191]= -1569004214;
assign addr[33192]= -1761306505;
assign addr[33193]= -1917915825;
assign addr[33194]= -2035658475;
assign addr[33195]= -2112148396;
assign addr[33196]= -2145835515;
assign addr[33197]= -2136037160;
assign addr[33198]= -2082951896;
assign addr[33199]= -1987655498;
assign addr[33200]= -1852079154;
assign addr[33201]= -1678970324;
assign addr[33202]= -1471837070;
assign addr[33203]= -1234876957;
assign addr[33204]= -972891995;
assign addr[33205]= -691191324;
assign addr[33206]= -395483624;
assign addr[33207]= -91761426;
assign addr[33208]= 213820322;
assign addr[33209]= 515068990;
assign addr[33210]= 805879757;
assign addr[33211]= 1080359326;
assign addr[33212]= 1332945355;
assign addr[33213]= 1558519173;
assign addr[33214]= 1752509516;
assign addr[33215]= 1910985158;
assign addr[33216]= 2030734582;
assign addr[33217]= 2109331059;
assign addr[33218]= 2145181827;
assign addr[33219]= 2137560369;
assign addr[33220]= 2086621133;
assign addr[33221]= 1993396407;
assign addr[33222]= 1859775393;
assign addr[33223]= 1688465931;
assign addr[33224]= 1482939614;
assign addr[33225]= 1247361445;
assign addr[33226]= 986505429;
assign addr[33227]= 705657826;
assign addr[33228]= 410510029;
assign addr[33229]= 107043224;
assign addr[33230]= -198592817;
assign addr[33231]= -500204365;
assign addr[33232]= -791679244;
assign addr[33233]= -1067110699;
assign addr[33234]= -1320917099;
assign addr[33235]= -1547955041;
assign addr[33236]= -1743623590;
assign addr[33237]= -1903957513;
assign addr[33238]= -2025707632;
assign addr[33239]= -2106406677;
assign addr[33240]= -2144419275;
assign addr[33241]= -2138975100;
assign addr[33242]= -2090184478;
assign addr[33243]= -1999036154;
assign addr[33244]= -1867377253;
assign addr[33245]= -1697875851;
assign addr[33246]= -1493966902;
assign addr[33247]= -1259782632;
assign addr[33248]= -1000068799;
assign addr[33249]= -720088517;
assign addr[33250]= -425515602;
assign addr[33251]= -122319591;
assign addr[33252]= 183355234;
assign addr[33253]= 485314355;
assign addr[33254]= 777438554;
assign addr[33255]= 1053807919;
assign addr[33256]= 1308821808;
assign addr[33257]= 1537312353;
assign addr[33258]= 1734649179;
assign addr[33259]= 1896833245;
assign addr[33260]= 2020577882;
assign addr[33261]= 2103375398;
assign addr[33262]= 2143547897;
assign addr[33263]= 2140281282;
assign addr[33264]= 2093641749;
assign addr[33265]= 2004574453;
assign addr[33266]= 1874884346;
assign addr[33267]= 1707199606;
assign addr[33268]= 1504918373;
assign addr[33269]= 1272139887;
assign addr[33270]= 1013581418;
assign addr[33271]= 734482665;
assign addr[33272]= 440499581;
assign addr[33273]= 137589750;
assign addr[33274]= -168108346;
assign addr[33275]= -470399716;
assign addr[33276]= -763158411;
assign addr[33277]= -1040451659;
assign addr[33278]= -1296660098;
assign addr[33279]= -1526591649;
assign addr[33280]= -1725586737;
assign addr[33281]= -1889612716;
assign addr[33282]= -2015345591;
assign addr[33283]= -2100237377;
assign addr[33284]= -2142567738;
assign addr[33285]= -2141478848;
assign addr[33286]= -2096992772;
assign addr[33287]= -2010011024;
assign addr[33288]= -1882296293;
assign addr[33289]= -1716436725;
assign addr[33290]= -1515793473;
assign addr[33291]= -1284432584;
assign addr[33292]= -1027042599;
assign addr[33293]= -748839539;
assign addr[33294]= -455461206;
assign addr[33295]= -152852926;
assign addr[33296]= 152852926;
assign addr[33297]= 455461206;
assign addr[33298]= 748839539;
assign addr[33299]= 1027042599;
assign addr[33300]= 1284432584;
assign addr[33301]= 1515793473;
assign addr[33302]= 1716436725;
assign addr[33303]= 1882296293;
assign addr[33304]= 2010011024;
assign addr[33305]= 2096992772;
assign addr[33306]= 2141478848;
assign addr[33307]= 2142567738;
assign addr[33308]= 2100237377;
assign addr[33309]= 2015345591;
assign addr[33310]= 1889612716;
assign addr[33311]= 1725586737;
assign addr[33312]= 1526591649;
assign addr[33313]= 1296660098;
assign addr[33314]= 1040451659;
assign addr[33315]= 763158411;
assign addr[33316]= 470399716;
assign addr[33317]= 168108346;
assign addr[33318]= -137589750;
assign addr[33319]= -440499581;
assign addr[33320]= -734482665;
assign addr[33321]= -1013581418;
assign addr[33322]= -1272139887;
assign addr[33323]= -1504918373;
assign addr[33324]= -1707199606;
assign addr[33325]= -1874884346;
assign addr[33326]= -2004574453;
assign addr[33327]= -2093641749;
assign addr[33328]= -2140281282;
assign addr[33329]= -2143547897;
assign addr[33330]= -2103375398;
assign addr[33331]= -2020577882;
assign addr[33332]= -1896833245;
assign addr[33333]= -1734649179;
assign addr[33334]= -1537312353;
assign addr[33335]= -1308821808;
assign addr[33336]= -1053807919;
assign addr[33337]= -777438554;
assign addr[33338]= -485314355;
assign addr[33339]= -183355234;
assign addr[33340]= 122319591;
assign addr[33341]= 425515602;
assign addr[33342]= 720088517;
assign addr[33343]= 1000068799;
assign addr[33344]= 1259782632;
assign addr[33345]= 1493966902;
assign addr[33346]= 1697875851;
assign addr[33347]= 1867377253;
assign addr[33348]= 1999036154;
assign addr[33349]= 2090184478;
assign addr[33350]= 2138975100;
assign addr[33351]= 2144419275;
assign addr[33352]= 2106406677;
assign addr[33353]= 2025707632;
assign addr[33354]= 1903957513;
assign addr[33355]= 1743623590;
assign addr[33356]= 1547955041;
assign addr[33357]= 1320917099;
assign addr[33358]= 1067110699;
assign addr[33359]= 791679244;
assign addr[33360]= 500204365;
assign addr[33361]= 198592817;
assign addr[33362]= -107043224;
assign addr[33363]= -410510029;
assign addr[33364]= -705657826;
assign addr[33365]= -986505429;
assign addr[33366]= -1247361445;
assign addr[33367]= -1482939614;
assign addr[33368]= -1688465931;
assign addr[33369]= -1859775393;
assign addr[33370]= -1993396407;
assign addr[33371]= -2086621133;
assign addr[33372]= -2137560369;
assign addr[33373]= -2145181827;
assign addr[33374]= -2109331059;
assign addr[33375]= -2030734582;
assign addr[33376]= -1910985158;
assign addr[33377]= -1752509516;
assign addr[33378]= -1558519173;
assign addr[33379]= -1332945355;
assign addr[33380]= -1080359326;
assign addr[33381]= -805879757;
assign addr[33382]= -515068990;
assign addr[33383]= -213820322;
assign addr[33384]= 91761426;
assign addr[33385]= 395483624;
assign addr[33386]= 691191324;
assign addr[33387]= 972891995;
assign addr[33388]= 1234876957;
assign addr[33389]= 1471837070;
assign addr[33390]= 1678970324;
assign addr[33391]= 1852079154;
assign addr[33392]= 1987655498;
assign addr[33393]= 2082951896;
assign addr[33394]= 2136037160;
assign addr[33395]= 2145835515;
assign addr[33396]= 2112148396;
assign addr[33397]= 2035658475;
assign addr[33398]= 1917915825;
assign addr[33399]= 1761306505;
assign addr[33400]= 1569004214;
assign addr[33401]= 1344905966;
assign addr[33402]= 1093553126;
assign addr[33403]= 820039373;
assign addr[33404]= 529907477;
assign addr[33405]= 229036977;
assign addr[33406]= -76474970;
assign addr[33407]= -380437148;
assign addr[33408]= -676689746;
assign addr[33409]= -959229189;
assign addr[33410]= -1222329801;
assign addr[33411]= -1460659832;
assign addr[33412]= -1669389513;
assign addr[33413]= -1844288924;
assign addr[33414]= -1981813720;
assign addr[33415]= -2079176953;
assign addr[33416]= -2134405552;
assign addr[33417]= -2146380306;
assign addr[33418]= -2114858546;
assign addr[33419]= -2040479063;
assign addr[33420]= -1924749160;
assign addr[33421]= -1770014111;
assign addr[33422]= -1579409630;
assign addr[33423]= -1356798326;
assign addr[33424]= -1106691431;
assign addr[33425]= -834157373;
assign addr[33426]= -544719071;
assign addr[33427]= -244242007;
assign addr[33428]= 61184634;
assign addr[33429]= 365371365;
assign addr[33430]= 662153826;
assign addr[33431]= 945517704;
assign addr[33432]= 1209720613;
assign addr[33433]= 1449408469;
assign addr[33434]= 1659723983;
assign addr[33435]= 1836405100;
assign addr[33436]= 1975871368;
assign addr[33437]= 2075296495;
assign addr[33438]= 2132665626;
assign addr[33439]= 2146816171;
assign addr[33440]= 2117461370;
assign addr[33441]= 2045196100;
assign addr[33442]= 1931484818;
assign addr[33443]= 1778631892;
assign addr[33444]= 1589734894;
assign addr[33445]= 1368621831;
assign addr[33446]= 1119773573;
assign addr[33447]= 848233042;
assign addr[33448]= 559503022;
assign addr[33449]= 259434643;
assign addr[33450]= -45891193;
assign addr[33451]= -350287041;
assign addr[33452]= -647584304;
assign addr[33453]= -931758235;
assign addr[33454]= -1197050035;
assign addr[33455]= -1438083551;
assign addr[33456]= -1649974225;
assign addr[33457]= -1828428082;
assign addr[33458]= -1969828744;
assign addr[33459]= -2071310720;
assign addr[33460]= -2130817471;
assign addr[33461]= -2147143090;
assign addr[33462]= -2119956737;
assign addr[33463]= -2049809346;
assign addr[33464]= -1938122457;
assign addr[33465]= -1787159411;
assign addr[33466]= -1599979481;
assign addr[33467]= -1380375881;
assign addr[33468]= -1132798888;
assign addr[33469]= -862265664;
assign addr[33470]= -574258580;
assign addr[33471]= -274614114;
assign addr[33472]= 30595422;
assign addr[33473]= 335184940;
assign addr[33474]= 632981917;
assign addr[33475]= 917951481;
assign addr[33476]= 1184318708;
assign addr[33477]= 1426685652;
assign addr[33478]= 1640140734;
assign addr[33479]= 1820358275;
assign addr[33480]= 1963686155;
assign addr[33481]= 2067219829;
assign addr[33482]= 2128861181;
assign addr[33483]= 2147361045;
assign addr[33484]= 2122344521;
assign addr[33485]= 2054318569;
assign addr[33486]= 1944661739;
assign addr[33487]= 1795596234;
assign addr[33488]= 1610142873;
assign addr[33489]= 1392059879;
assign addr[33490]= 1145766716;
assign addr[33491]= 876254528;
assign addr[33492]= 588984994;
assign addr[33493]= 289779648;
assign addr[33494]= -15298099;
assign addr[33495]= -320065829;
assign addr[33496]= -618347408;
assign addr[33497]= -904098143;
assign addr[33498]= -1171527280;
assign addr[33499]= -1415215352;
assign addr[33500]= -1630224009;
assign addr[33501]= -1812196087;
assign addr[33502]= -1957443913;
assign addr[33503]= -2063024031;
assign addr[33504]= -2126796855;
assign addr[33505]= -2147470025;
assign addr[33506]= -2124624598;
assign addr[33507]= -2058723538;
assign addr[33508]= -1951102334;
assign addr[33509]= -1803941934;
assign addr[33510]= -1620224553;
assign addr[33511]= -1403673233;
assign addr[33512]= -1158676398;
assign addr[33513]= -890198924;
assign addr[33514]= -603681519;
assign addr[33515]= -304930476;
assign addr[33516]= 0;
assign addr[33517]= 304930476;
assign addr[33518]= 603681519;
assign addr[33519]= 890198924;
assign addr[33520]= 1158676398;
assign addr[33521]= 1403673233;
assign addr[33522]= 1620224553;
assign addr[33523]= 1803941934;
assign addr[33524]= 1951102334;
assign addr[33525]= 2058723538;
assign addr[33526]= 2124624598;
assign addr[33527]= 2147470025;
assign addr[33528]= 2126796855;
assign addr[33529]= 2063024031;
assign addr[33530]= 1957443913;
assign addr[33531]= 1812196087;
assign addr[33532]= 1630224009;
assign addr[33533]= 1415215352;
assign addr[33534]= 1171527280;
assign addr[33535]= 904098143;
assign addr[33536]= 618347408;
assign addr[33537]= 320065829;
assign addr[33538]= 15298099;
assign addr[33539]= -289779648;
assign addr[33540]= -588984994;
assign addr[33541]= -876254528;
assign addr[33542]= -1145766716;
assign addr[33543]= -1392059879;
assign addr[33544]= -1610142873;
assign addr[33545]= -1795596234;
assign addr[33546]= -1944661739;
assign addr[33547]= -2054318569;
assign addr[33548]= -2122344521;
assign addr[33549]= -2147361045;
assign addr[33550]= -2128861181;
assign addr[33551]= -2067219829;
assign addr[33552]= -1963686155;
assign addr[33553]= -1820358275;
assign addr[33554]= -1640140734;
assign addr[33555]= -1426685652;
assign addr[33556]= -1184318708;
assign addr[33557]= -917951481;
assign addr[33558]= -632981917;
assign addr[33559]= -335184940;
assign addr[33560]= -30595422;
assign addr[33561]= 274614114;
assign addr[33562]= 574258580;
assign addr[33563]= 862265664;
assign addr[33564]= 1132798888;
assign addr[33565]= 1380375881;
assign addr[33566]= 1599979481;
assign addr[33567]= 1787159411;
assign addr[33568]= 1938122457;
assign addr[33569]= 2049809346;
assign addr[33570]= 2119956737;
assign addr[33571]= 2147143090;
assign addr[33572]= 2130817471;
assign addr[33573]= 2071310720;
assign addr[33574]= 1969828744;
assign addr[33575]= 1828428082;
assign addr[33576]= 1649974225;
assign addr[33577]= 1438083551;
assign addr[33578]= 1197050035;
assign addr[33579]= 931758235;
assign addr[33580]= 647584304;
assign addr[33581]= 350287041;
assign addr[33582]= 45891193;
assign addr[33583]= -259434643;
assign addr[33584]= -559503022;
assign addr[33585]= -848233042;
assign addr[33586]= -1119773573;
assign addr[33587]= -1368621831;
assign addr[33588]= -1589734894;
assign addr[33589]= -1778631892;
assign addr[33590]= -1931484818;
assign addr[33591]= -2045196100;
assign addr[33592]= -2117461370;
assign addr[33593]= -2146816171;
assign addr[33594]= -2132665626;
assign addr[33595]= -2075296495;
assign addr[33596]= -1975871368;
assign addr[33597]= -1836405100;
assign addr[33598]= -1659723983;
assign addr[33599]= -1449408469;
assign addr[33600]= -1209720613;
assign addr[33601]= -945517704;
assign addr[33602]= -662153826;
assign addr[33603]= -365371365;
assign addr[33604]= -61184634;
assign addr[33605]= 244242007;
assign addr[33606]= 544719071;
assign addr[33607]= 834157373;
assign addr[33608]= 1106691431;
assign addr[33609]= 1356798326;
assign addr[33610]= 1579409630;
assign addr[33611]= 1770014111;
assign addr[33612]= 1924749160;
assign addr[33613]= 2040479063;
assign addr[33614]= 2114858546;
assign addr[33615]= 2146380306;
assign addr[33616]= 2134405552;
assign addr[33617]= 2079176953;
assign addr[33618]= 1981813720;
assign addr[33619]= 1844288924;
assign addr[33620]= 1669389513;
assign addr[33621]= 1460659832;
assign addr[33622]= 1222329801;
assign addr[33623]= 959229189;
assign addr[33624]= 676689746;
assign addr[33625]= 380437148;
assign addr[33626]= 76474970;
assign addr[33627]= -229036977;
assign addr[33628]= -529907477;
assign addr[33629]= -820039373;
assign addr[33630]= -1093553126;
assign addr[33631]= -1344905966;
assign addr[33632]= -1569004214;
assign addr[33633]= -1761306505;
assign addr[33634]= -1917915825;
assign addr[33635]= -2035658475;
assign addr[33636]= -2112148396;
assign addr[33637]= -2145835515;
assign addr[33638]= -2136037160;
assign addr[33639]= -2082951896;
assign addr[33640]= -1987655498;
assign addr[33641]= -1852079154;
assign addr[33642]= -1678970324;
assign addr[33643]= -1471837070;
assign addr[33644]= -1234876957;
assign addr[33645]= -972891995;
assign addr[33646]= -691191324;
assign addr[33647]= -395483624;
assign addr[33648]= -91761426;
assign addr[33649]= 213820322;
assign addr[33650]= 515068990;
assign addr[33651]= 805879757;
assign addr[33652]= 1080359326;
assign addr[33653]= 1332945355;
assign addr[33654]= 1558519173;
assign addr[33655]= 1752509516;
assign addr[33656]= 1910985158;
assign addr[33657]= 2030734582;
assign addr[33658]= 2109331059;
assign addr[33659]= 2145181827;
assign addr[33660]= 2137560369;
assign addr[33661]= 2086621133;
assign addr[33662]= 1993396407;
assign addr[33663]= 1859775393;
assign addr[33664]= 1688465931;
assign addr[33665]= 1482939614;
assign addr[33666]= 1247361445;
assign addr[33667]= 986505429;
assign addr[33668]= 705657826;
assign addr[33669]= 410510029;
assign addr[33670]= 107043224;
assign addr[33671]= -198592817;
assign addr[33672]= -500204365;
assign addr[33673]= -791679244;
assign addr[33674]= -1067110699;
assign addr[33675]= -1320917099;
assign addr[33676]= -1547955041;
assign addr[33677]= -1743623590;
assign addr[33678]= -1903957513;
assign addr[33679]= -2025707632;
assign addr[33680]= -2106406677;
assign addr[33681]= -2144419275;
assign addr[33682]= -2138975100;
assign addr[33683]= -2090184478;
assign addr[33684]= -1999036154;
assign addr[33685]= -1867377253;
assign addr[33686]= -1697875851;
assign addr[33687]= -1493966902;
assign addr[33688]= -1259782632;
assign addr[33689]= -1000068799;
assign addr[33690]= -720088517;
assign addr[33691]= -425515602;
assign addr[33692]= -122319591;
assign addr[33693]= 183355234;
assign addr[33694]= 485314355;
assign addr[33695]= 777438554;
assign addr[33696]= 1053807919;
assign addr[33697]= 1308821808;
assign addr[33698]= 1537312353;
assign addr[33699]= 1734649179;
assign addr[33700]= 1896833245;
assign addr[33701]= 2020577882;
assign addr[33702]= 2103375398;
assign addr[33703]= 2143547897;
assign addr[33704]= 2140281282;
assign addr[33705]= 2093641749;
assign addr[33706]= 2004574453;
assign addr[33707]= 1874884346;
assign addr[33708]= 1707199606;
assign addr[33709]= 1504918373;
assign addr[33710]= 1272139887;
assign addr[33711]= 1013581418;
assign addr[33712]= 734482665;
assign addr[33713]= 440499581;
assign addr[33714]= 137589750;
assign addr[33715]= -168108346;
assign addr[33716]= -470399716;
assign addr[33717]= -763158411;
assign addr[33718]= -1040451659;
assign addr[33719]= -1296660098;
assign addr[33720]= -1526591649;
assign addr[33721]= -1725586737;
assign addr[33722]= -1889612716;
assign addr[33723]= -2015345591;
assign addr[33724]= -2100237377;
assign addr[33725]= -2142567738;
assign addr[33726]= -2141478848;
assign addr[33727]= -2096992772;
assign addr[33728]= -2010011024;
assign addr[33729]= -1882296293;
assign addr[33730]= -1716436725;
assign addr[33731]= -1515793473;
assign addr[33732]= -1284432584;
assign addr[33733]= -1027042599;
assign addr[33734]= -748839539;
assign addr[33735]= -455461206;
assign addr[33736]= -152852926;
assign addr[33737]= 152852926;
assign addr[33738]= 455461206;
assign addr[33739]= 748839539;
assign addr[33740]= 1027042599;
assign addr[33741]= 1284432584;
assign addr[33742]= 1515793473;
assign addr[33743]= 1716436725;
assign addr[33744]= 1882296293;
assign addr[33745]= 2010011024;
assign addr[33746]= 2096992772;
assign addr[33747]= 2141478848;
assign addr[33748]= 2142567738;
assign addr[33749]= 2100237377;
assign addr[33750]= 2015345591;
assign addr[33751]= 1889612716;
assign addr[33752]= 1725586737;
assign addr[33753]= 1526591649;
assign addr[33754]= 1296660098;
assign addr[33755]= 1040451659;
assign addr[33756]= 763158411;
assign addr[33757]= 470399716;
assign addr[33758]= 168108346;
assign addr[33759]= -137589750;
assign addr[33760]= -440499581;
assign addr[33761]= -734482665;
assign addr[33762]= -1013581418;
assign addr[33763]= -1272139887;
assign addr[33764]= -1504918373;
assign addr[33765]= -1707199606;
assign addr[33766]= -1874884346;
assign addr[33767]= -2004574453;
assign addr[33768]= -2093641749;
assign addr[33769]= -2140281282;
assign addr[33770]= -2143547897;
assign addr[33771]= -2103375398;
assign addr[33772]= -2020577882;
assign addr[33773]= -1896833245;
assign addr[33774]= -1734649179;
assign addr[33775]= -1537312353;
assign addr[33776]= -1308821808;
assign addr[33777]= -1053807919;
assign addr[33778]= -777438554;
assign addr[33779]= -485314355;
assign addr[33780]= -183355234;
assign addr[33781]= 122319591;
assign addr[33782]= 425515602;
assign addr[33783]= 720088517;
assign addr[33784]= 1000068799;
assign addr[33785]= 1259782632;
assign addr[33786]= 1493966902;
assign addr[33787]= 1697875851;
assign addr[33788]= 1867377253;
assign addr[33789]= 1999036154;
assign addr[33790]= 2090184478;
assign addr[33791]= 2138975100;
assign addr[33792]= 2144419275;
assign addr[33793]= 2106406677;
assign addr[33794]= 2025707632;
assign addr[33795]= 1903957513;
assign addr[33796]= 1743623590;
assign addr[33797]= 1547955041;
assign addr[33798]= 1320917099;
assign addr[33799]= 1067110699;
assign addr[33800]= 791679244;
assign addr[33801]= 500204365;
assign addr[33802]= 198592817;
assign addr[33803]= -107043224;
assign addr[33804]= -410510029;
assign addr[33805]= -705657826;
assign addr[33806]= -986505429;
assign addr[33807]= -1247361445;
assign addr[33808]= -1482939614;
assign addr[33809]= -1688465931;
assign addr[33810]= -1859775393;
assign addr[33811]= -1993396407;
assign addr[33812]= -2086621133;
assign addr[33813]= -2137560369;
assign addr[33814]= -2145181827;
assign addr[33815]= -2109331059;
assign addr[33816]= -2030734582;
assign addr[33817]= -1910985158;
assign addr[33818]= -1752509516;
assign addr[33819]= -1558519173;
assign addr[33820]= -1332945355;
assign addr[33821]= -1080359326;
assign addr[33822]= -805879757;
assign addr[33823]= -515068990;
assign addr[33824]= -213820322;
assign addr[33825]= 91761426;
assign addr[33826]= 395483624;
assign addr[33827]= 691191324;
assign addr[33828]= 972891995;
assign addr[33829]= 1234876957;
assign addr[33830]= 1471837070;
assign addr[33831]= 1678970324;
assign addr[33832]= 1852079154;
assign addr[33833]= 1987655498;
assign addr[33834]= 2082951896;
assign addr[33835]= 2136037160;
assign addr[33836]= 2145835515;
assign addr[33837]= 2112148396;
assign addr[33838]= 2035658475;
assign addr[33839]= 1917915825;
assign addr[33840]= 1761306505;
assign addr[33841]= 1569004214;
assign addr[33842]= 1344905966;
assign addr[33843]= 1093553126;
assign addr[33844]= 820039373;
assign addr[33845]= 529907477;
assign addr[33846]= 229036977;
assign addr[33847]= -76474970;
assign addr[33848]= -380437148;
assign addr[33849]= -676689746;
assign addr[33850]= -959229189;
assign addr[33851]= -1222329801;
assign addr[33852]= -1460659832;
assign addr[33853]= -1669389513;
assign addr[33854]= -1844288924;
assign addr[33855]= -1981813720;
assign addr[33856]= -2079176953;
assign addr[33857]= -2134405552;
assign addr[33858]= -2146380306;
assign addr[33859]= -2114858546;
assign addr[33860]= -2040479063;
assign addr[33861]= -1924749160;
assign addr[33862]= -1770014111;
assign addr[33863]= -1579409630;
assign addr[33864]= -1356798326;
assign addr[33865]= -1106691431;
assign addr[33866]= -834157373;
assign addr[33867]= -544719071;
assign addr[33868]= -244242007;
assign addr[33869]= 61184634;
assign addr[33870]= 365371365;
assign addr[33871]= 662153826;
assign addr[33872]= 945517704;
assign addr[33873]= 1209720613;
assign addr[33874]= 1449408469;
assign addr[33875]= 1659723983;
assign addr[33876]= 1836405100;
assign addr[33877]= 1975871368;
assign addr[33878]= 2075296495;
assign addr[33879]= 2132665626;
assign addr[33880]= 2146816171;
assign addr[33881]= 2117461370;
assign addr[33882]= 2045196100;
assign addr[33883]= 1931484818;
assign addr[33884]= 1778631892;
assign addr[33885]= 1589734894;
assign addr[33886]= 1368621831;
assign addr[33887]= 1119773573;
assign addr[33888]= 848233042;
assign addr[33889]= 559503022;
assign addr[33890]= 259434643;
assign addr[33891]= -45891193;
assign addr[33892]= -350287041;
assign addr[33893]= -647584304;
assign addr[33894]= -931758235;
assign addr[33895]= -1197050035;
assign addr[33896]= -1438083551;
assign addr[33897]= -1649974225;
assign addr[33898]= -1828428082;
assign addr[33899]= -1969828744;
assign addr[33900]= -2071310720;
assign addr[33901]= -2130817471;
assign addr[33902]= -2147143090;
assign addr[33903]= -2119956737;
assign addr[33904]= -2049809346;
assign addr[33905]= -1938122457;
assign addr[33906]= -1787159411;
assign addr[33907]= -1599979481;
assign addr[33908]= -1380375881;
assign addr[33909]= -1132798888;
assign addr[33910]= -862265664;
assign addr[33911]= -574258580;
assign addr[33912]= -274614114;
assign addr[33913]= 30595422;
assign addr[33914]= 335184940;
assign addr[33915]= 632981917;
assign addr[33916]= 917951481;
assign addr[33917]= 1184318708;
assign addr[33918]= 1426685652;
assign addr[33919]= 1640140734;
assign addr[33920]= 1820358275;
assign addr[33921]= 1963686155;
assign addr[33922]= 2067219829;
assign addr[33923]= 2128861181;
assign addr[33924]= 2147361045;
assign addr[33925]= 2122344521;
assign addr[33926]= 2054318569;
assign addr[33927]= 1944661739;
assign addr[33928]= 1795596234;
assign addr[33929]= 1610142873;
assign addr[33930]= 1392059879;
assign addr[33931]= 1145766716;
assign addr[33932]= 876254528;
assign addr[33933]= 588984994;
assign addr[33934]= 289779648;
assign addr[33935]= -15298099;
assign addr[33936]= -320065829;
assign addr[33937]= -618347408;
assign addr[33938]= -904098143;
assign addr[33939]= -1171527280;
assign addr[33940]= -1415215352;
assign addr[33941]= -1630224009;
assign addr[33942]= -1812196087;
assign addr[33943]= -1957443913;
assign addr[33944]= -2063024031;
assign addr[33945]= -2126796855;
assign addr[33946]= -2147470025;
assign addr[33947]= -2124624598;
assign addr[33948]= -2058723538;
assign addr[33949]= -1951102334;
assign addr[33950]= -1803941934;
assign addr[33951]= -1620224553;
assign addr[33952]= -1403673233;
assign addr[33953]= -1158676398;
assign addr[33954]= -890198924;
assign addr[33955]= -603681519;
assign addr[33956]= -304930476;
assign addr[33957]= 0;
assign addr[33958]= 304930476;
assign addr[33959]= 603681519;
assign addr[33960]= 890198924;
assign addr[33961]= 1158676398;
assign addr[33962]= 1403673233;
assign addr[33963]= 1620224553;
assign addr[33964]= 1803941934;
assign addr[33965]= 1951102334;
assign addr[33966]= 2058723538;
assign addr[33967]= 2124624598;
assign addr[33968]= 2147470025;
assign addr[33969]= 2126796855;
assign addr[33970]= 2063024031;
assign addr[33971]= 1957443913;
assign addr[33972]= 1812196087;
assign addr[33973]= 1630224009;
assign addr[33974]= 1415215352;
assign addr[33975]= 1171527280;
assign addr[33976]= 904098143;
assign addr[33977]= 618347408;
assign addr[33978]= 320065829;
assign addr[33979]= 15298099;
assign addr[33980]= -289779648;
assign addr[33981]= -588984994;
assign addr[33982]= -876254528;
assign addr[33983]= -1145766716;
assign addr[33984]= -1392059879;
assign addr[33985]= -1610142873;
assign addr[33986]= -1795596234;
assign addr[33987]= -1944661739;
assign addr[33988]= -2054318569;
assign addr[33989]= -2122344521;
assign addr[33990]= -2147361045;
assign addr[33991]= -2128861181;
assign addr[33992]= -2067219829;
assign addr[33993]= -1963686155;
assign addr[33994]= -1820358275;
assign addr[33995]= -1640140734;
assign addr[33996]= -1426685652;
assign addr[33997]= -1184318708;
assign addr[33998]= -917951481;
assign addr[33999]= -632981917;
assign addr[34000]= -335184940;
assign addr[34001]= -30595422;
assign addr[34002]= 274614114;
assign addr[34003]= 574258580;
assign addr[34004]= 862265664;
assign addr[34005]= 1132798888;
assign addr[34006]= 1380375881;
assign addr[34007]= 1599979481;
assign addr[34008]= 1787159411;
assign addr[34009]= 1938122457;
assign addr[34010]= 2049809346;
assign addr[34011]= 2119956737;
assign addr[34012]= 2147143090;
assign addr[34013]= 2130817471;
assign addr[34014]= 2071310720;
assign addr[34015]= 1969828744;
assign addr[34016]= 1828428082;
assign addr[34017]= 1649974225;
assign addr[34018]= 1438083551;
assign addr[34019]= 1197050035;
assign addr[34020]= 931758235;
assign addr[34021]= 647584304;
assign addr[34022]= 350287041;
assign addr[34023]= 45891193;
assign addr[34024]= -259434643;
assign addr[34025]= -559503022;
assign addr[34026]= -848233042;
assign addr[34027]= -1119773573;
assign addr[34028]= -1368621831;
assign addr[34029]= -1589734894;
assign addr[34030]= -1778631892;
assign addr[34031]= -1931484818;
assign addr[34032]= -2045196100;
assign addr[34033]= -2117461370;
assign addr[34034]= -2146816171;
assign addr[34035]= -2132665626;
assign addr[34036]= -2075296495;
assign addr[34037]= -1975871368;
assign addr[34038]= -1836405100;
assign addr[34039]= -1659723983;
assign addr[34040]= -1449408469;
assign addr[34041]= -1209720613;
assign addr[34042]= -945517704;
assign addr[34043]= -662153826;
assign addr[34044]= -365371365;
assign addr[34045]= -61184634;
assign addr[34046]= 244242007;
assign addr[34047]= 544719071;
assign addr[34048]= 834157373;
assign addr[34049]= 1106691431;
assign addr[34050]= 1356798326;
assign addr[34051]= 1579409630;
assign addr[34052]= 1770014111;
assign addr[34053]= 1924749160;
assign addr[34054]= 2040479063;
assign addr[34055]= 2114858546;
assign addr[34056]= 2146380306;
assign addr[34057]= 2134405552;
assign addr[34058]= 2079176953;
assign addr[34059]= 1981813720;
assign addr[34060]= 1844288924;
assign addr[34061]= 1669389513;
assign addr[34062]= 1460659832;
assign addr[34063]= 1222329801;
assign addr[34064]= 959229189;
assign addr[34065]= 676689746;
assign addr[34066]= 380437148;
assign addr[34067]= 76474970;
assign addr[34068]= -229036977;
assign addr[34069]= -529907477;
assign addr[34070]= -820039373;
assign addr[34071]= -1093553126;
assign addr[34072]= -1344905966;
assign addr[34073]= -1569004214;
assign addr[34074]= -1761306505;
assign addr[34075]= -1917915825;
assign addr[34076]= -2035658475;
assign addr[34077]= -2112148396;
assign addr[34078]= -2145835515;
assign addr[34079]= -2136037160;
assign addr[34080]= -2082951896;
assign addr[34081]= -1987655498;
assign addr[34082]= -1852079154;
assign addr[34083]= -1678970324;
assign addr[34084]= -1471837070;
assign addr[34085]= -1234876957;
assign addr[34086]= -972891995;
assign addr[34087]= -691191324;
assign addr[34088]= -395483624;
assign addr[34089]= -91761426;
assign addr[34090]= 213820322;
assign addr[34091]= 515068990;
assign addr[34092]= 805879757;
assign addr[34093]= 1080359326;
assign addr[34094]= 1332945355;
assign addr[34095]= 1558519173;
assign addr[34096]= 1752509516;
assign addr[34097]= 1910985158;
assign addr[34098]= 2030734582;
assign addr[34099]= 2109331059;
assign addr[34100]= 2145181827;
assign addr[34101]= 2137560369;
assign addr[34102]= 2086621133;
assign addr[34103]= 1993396407;
assign addr[34104]= 1859775393;
assign addr[34105]= 1688465931;
assign addr[34106]= 1482939614;
assign addr[34107]= 1247361445;
assign addr[34108]= 986505429;
assign addr[34109]= 705657826;
assign addr[34110]= 410510029;
assign addr[34111]= 107043224;
assign addr[34112]= -198592817;
assign addr[34113]= -500204365;
assign addr[34114]= -791679244;
assign addr[34115]= -1067110699;
assign addr[34116]= -1320917099;
assign addr[34117]= -1547955041;
assign addr[34118]= -1743623590;
assign addr[34119]= -1903957513;
assign addr[34120]= -2025707632;
assign addr[34121]= -2106406677;
assign addr[34122]= -2144419275;
assign addr[34123]= -2138975100;
assign addr[34124]= -2090184478;
assign addr[34125]= -1999036154;
assign addr[34126]= -1867377253;
assign addr[34127]= -1697875851;
assign addr[34128]= -1493966902;
assign addr[34129]= -1259782632;
assign addr[34130]= -1000068799;
assign addr[34131]= -720088517;
assign addr[34132]= -425515602;
assign addr[34133]= -122319591;
assign addr[34134]= 183355234;
assign addr[34135]= 485314355;
assign addr[34136]= 777438554;
assign addr[34137]= 1053807919;
assign addr[34138]= 1308821808;
assign addr[34139]= 1537312353;
assign addr[34140]= 1734649179;
assign addr[34141]= 1896833245;
assign addr[34142]= 2020577882;
assign addr[34143]= 2103375398;
assign addr[34144]= 2143547897;
assign addr[34145]= 2140281282;
assign addr[34146]= 2093641749;
assign addr[34147]= 2004574453;
assign addr[34148]= 1874884346;
assign addr[34149]= 1707199606;
assign addr[34150]= 1504918373;
assign addr[34151]= 1272139887;
assign addr[34152]= 1013581418;
assign addr[34153]= 734482665;
assign addr[34154]= 440499581;
assign addr[34155]= 137589750;
assign addr[34156]= -168108346;
assign addr[34157]= -470399716;
assign addr[34158]= -763158411;
assign addr[34159]= -1040451659;
assign addr[34160]= -1296660098;
assign addr[34161]= -1526591649;
assign addr[34162]= -1725586737;
assign addr[34163]= -1889612716;
assign addr[34164]= -2015345591;
assign addr[34165]= -2100237377;
assign addr[34166]= -2142567738;
assign addr[34167]= -2141478848;
assign addr[34168]= -2096992772;
assign addr[34169]= -2010011024;
assign addr[34170]= -1882296293;
assign addr[34171]= -1716436725;
assign addr[34172]= -1515793473;
assign addr[34173]= -1284432584;
assign addr[34174]= -1027042599;
assign addr[34175]= -748839539;
assign addr[34176]= -455461206;
assign addr[34177]= -152852926;
assign addr[34178]= 152852926;
assign addr[34179]= 455461206;
assign addr[34180]= 748839539;
assign addr[34181]= 1027042599;
assign addr[34182]= 1284432584;
assign addr[34183]= 1515793473;
assign addr[34184]= 1716436725;
assign addr[34185]= 1882296293;
assign addr[34186]= 2010011024;
assign addr[34187]= 2096992772;
assign addr[34188]= 2141478848;
assign addr[34189]= 2142567738;
assign addr[34190]= 2100237377;
assign addr[34191]= 2015345591;
assign addr[34192]= 1889612716;
assign addr[34193]= 1725586737;
assign addr[34194]= 1526591649;
assign addr[34195]= 1296660098;
assign addr[34196]= 1040451659;
assign addr[34197]= 763158411;
assign addr[34198]= 470399716;
assign addr[34199]= 168108346;
assign addr[34200]= -137589750;
assign addr[34201]= -440499581;
assign addr[34202]= -734482665;
assign addr[34203]= -1013581418;
assign addr[34204]= -1272139887;
assign addr[34205]= -1504918373;
assign addr[34206]= -1707199606;
assign addr[34207]= -1874884346;
assign addr[34208]= -2004574453;
assign addr[34209]= -2093641749;
assign addr[34210]= -2140281282;
assign addr[34211]= -2143547897;
assign addr[34212]= -2103375398;
assign addr[34213]= -2020577882;
assign addr[34214]= -1896833245;
assign addr[34215]= -1734649179;
assign addr[34216]= -1537312353;
assign addr[34217]= -1308821808;
assign addr[34218]= -1053807919;
assign addr[34219]= -777438554;
assign addr[34220]= -485314355;
assign addr[34221]= -183355234;
assign addr[34222]= 122319591;
assign addr[34223]= 425515602;
assign addr[34224]= 720088517;
assign addr[34225]= 1000068799;
assign addr[34226]= 1259782632;
assign addr[34227]= 1493966902;
assign addr[34228]= 1697875851;
assign addr[34229]= 1867377253;
assign addr[34230]= 1999036154;
assign addr[34231]= 2090184478;
assign addr[34232]= 2138975100;
assign addr[34233]= 2144419275;
assign addr[34234]= 2106406677;
assign addr[34235]= 2025707632;
assign addr[34236]= 1903957513;
assign addr[34237]= 1743623590;
assign addr[34238]= 1547955041;
assign addr[34239]= 1320917099;
assign addr[34240]= 1067110699;
assign addr[34241]= 791679244;
assign addr[34242]= 500204365;
assign addr[34243]= 198592817;
assign addr[34244]= -107043224;
assign addr[34245]= -410510029;
assign addr[34246]= -705657826;
assign addr[34247]= -986505429;
assign addr[34248]= -1247361445;
assign addr[34249]= -1482939614;
assign addr[34250]= -1688465931;
assign addr[34251]= -1859775393;
assign addr[34252]= -1993396407;
assign addr[34253]= -2086621133;
assign addr[34254]= -2137560369;
assign addr[34255]= -2145181827;
assign addr[34256]= -2109331059;
assign addr[34257]= -2030734582;
assign addr[34258]= -1910985158;
assign addr[34259]= -1752509516;
assign addr[34260]= -1558519173;
assign addr[34261]= -1332945355;
assign addr[34262]= -1080359326;
assign addr[34263]= -805879757;
assign addr[34264]= -515068990;
assign addr[34265]= -213820322;
assign addr[34266]= 91761426;
assign addr[34267]= 395483624;
assign addr[34268]= 691191324;
assign addr[34269]= 972891995;
assign addr[34270]= 1234876957;
assign addr[34271]= 1471837070;
assign addr[34272]= 1678970324;
assign addr[34273]= 1852079154;
assign addr[34274]= 1987655498;
assign addr[34275]= 2082951896;
assign addr[34276]= 2136037160;
assign addr[34277]= 2145835515;
assign addr[34278]= 2112148396;
assign addr[34279]= 2035658475;
assign addr[34280]= 1917915825;
assign addr[34281]= 1761306505;
assign addr[34282]= 1569004214;
assign addr[34283]= 1344905966;
assign addr[34284]= 1093553126;
assign addr[34285]= 820039373;
assign addr[34286]= 529907477;
assign addr[34287]= 229036977;
assign addr[34288]= -76474970;
assign addr[34289]= -380437148;
assign addr[34290]= -676689746;
assign addr[34291]= -959229189;
assign addr[34292]= -1222329801;
assign addr[34293]= -1460659832;
assign addr[34294]= -1669389513;
assign addr[34295]= -1844288924;
assign addr[34296]= -1981813720;
assign addr[34297]= -2079176953;
assign addr[34298]= -2134405552;
assign addr[34299]= -2146380306;
assign addr[34300]= -2114858546;
assign addr[34301]= -2040479063;
assign addr[34302]= -1924749160;
assign addr[34303]= -1770014111;
assign addr[34304]= -1579409630;
assign addr[34305]= -1356798326;
assign addr[34306]= -1106691431;
assign addr[34307]= -834157373;
assign addr[34308]= -544719071;
assign addr[34309]= -244242007;
assign addr[34310]= 61184634;
assign addr[34311]= 365371365;
assign addr[34312]= 662153826;
assign addr[34313]= 945517704;
assign addr[34314]= 1209720613;
assign addr[34315]= 1449408469;
assign addr[34316]= 1659723983;
assign addr[34317]= 1836405100;
assign addr[34318]= 1975871368;
assign addr[34319]= 2075296495;
assign addr[34320]= 2132665626;
assign addr[34321]= 2146816171;
assign addr[34322]= 2117461370;
assign addr[34323]= 2045196100;
assign addr[34324]= 1931484818;
assign addr[34325]= 1778631892;
assign addr[34326]= 1589734894;
assign addr[34327]= 1368621831;
assign addr[34328]= 1119773573;
assign addr[34329]= 848233042;
assign addr[34330]= 559503022;
assign addr[34331]= 259434643;
assign addr[34332]= -45891193;
assign addr[34333]= -350287041;
assign addr[34334]= -647584304;
assign addr[34335]= -931758235;
assign addr[34336]= -1197050035;
assign addr[34337]= -1438083551;
assign addr[34338]= -1649974225;
assign addr[34339]= -1828428082;
assign addr[34340]= -1969828744;
assign addr[34341]= -2071310720;
assign addr[34342]= -2130817471;
assign addr[34343]= -2147143090;
assign addr[34344]= -2119956737;
assign addr[34345]= -2049809346;
assign addr[34346]= -1938122457;
assign addr[34347]= -1787159411;
assign addr[34348]= -1599979481;
assign addr[34349]= -1380375881;
assign addr[34350]= -1132798888;
assign addr[34351]= -862265664;
assign addr[34352]= -574258580;
assign addr[34353]= -274614114;
assign addr[34354]= 30595422;
assign addr[34355]= 335184940;
assign addr[34356]= 632981917;
assign addr[34357]= 917951481;
assign addr[34358]= 1184318708;
assign addr[34359]= 1426685652;
assign addr[34360]= 1640140734;
assign addr[34361]= 1820358275;
assign addr[34362]= 1963686155;
assign addr[34363]= 2067219829;
assign addr[34364]= 2128861181;
assign addr[34365]= 2147361045;
assign addr[34366]= 2122344521;
assign addr[34367]= 2054318569;
assign addr[34368]= 1944661739;
assign addr[34369]= 1795596234;
assign addr[34370]= 1610142873;
assign addr[34371]= 1392059879;
assign addr[34372]= 1145766716;
assign addr[34373]= 876254528;
assign addr[34374]= 588984994;
assign addr[34375]= 289779648;
assign addr[34376]= -15298099;
assign addr[34377]= -320065829;
assign addr[34378]= -618347408;
assign addr[34379]= -904098143;
assign addr[34380]= -1171527280;
assign addr[34381]= -1415215352;
assign addr[34382]= -1630224009;
assign addr[34383]= -1812196087;
assign addr[34384]= -1957443913;
assign addr[34385]= -2063024031;
assign addr[34386]= -2126796855;
assign addr[34387]= -2147470025;
assign addr[34388]= -2124624598;
assign addr[34389]= -2058723538;
assign addr[34390]= -1951102334;
assign addr[34391]= -1803941934;
assign addr[34392]= -1620224553;
assign addr[34393]= -1403673233;
assign addr[34394]= -1158676398;
assign addr[34395]= -890198924;
assign addr[34396]= -603681519;
assign addr[34397]= -304930476;
assign addr[34398]= 0;
assign addr[34399]= 304930476;
assign addr[34400]= 603681519;
assign addr[34401]= 890198924;
assign addr[34402]= 1158676398;
assign addr[34403]= 1403673233;
assign addr[34404]= 1620224553;
assign addr[34405]= 1803941934;
assign addr[34406]= 1951102334;
assign addr[34407]= 2058723538;
assign addr[34408]= 2124624598;
assign addr[34409]= 2147470025;
assign addr[34410]= 2126796855;
assign addr[34411]= 2063024031;
assign addr[34412]= 1957443913;
assign addr[34413]= 1812196087;
assign addr[34414]= 1630224009;
assign addr[34415]= 1415215352;
assign addr[34416]= 1171527280;
assign addr[34417]= 904098143;
assign addr[34418]= 618347408;
assign addr[34419]= 320065829;
assign addr[34420]= 15298099;
assign addr[34421]= -289779648;
assign addr[34422]= -588984994;
assign addr[34423]= -876254528;
assign addr[34424]= -1145766716;
assign addr[34425]= -1392059879;
assign addr[34426]= -1610142873;
assign addr[34427]= -1795596234;
assign addr[34428]= -1944661739;
assign addr[34429]= -2054318569;
assign addr[34430]= -2122344521;
assign addr[34431]= -2147361045;
assign addr[34432]= -2128861181;
assign addr[34433]= -2067219829;
assign addr[34434]= -1963686155;
assign addr[34435]= -1820358275;
assign addr[34436]= -1640140734;
assign addr[34437]= -1426685652;
assign addr[34438]= -1184318708;
assign addr[34439]= -917951481;
assign addr[34440]= -632981917;
assign addr[34441]= -335184940;
assign addr[34442]= -30595422;
assign addr[34443]= 274614114;
assign addr[34444]= 574258580;
assign addr[34445]= 862265664;
assign addr[34446]= 1132798888;
assign addr[34447]= 1380375881;
assign addr[34448]= 1599979481;
assign addr[34449]= 1787159411;
assign addr[34450]= 1938122457;
assign addr[34451]= 2049809346;
assign addr[34452]= 2119956737;
assign addr[34453]= 2147143090;
assign addr[34454]= 2130817471;
assign addr[34455]= 2071310720;
assign addr[34456]= 1969828744;
assign addr[34457]= 1828428082;
assign addr[34458]= 1649974225;
assign addr[34459]= 1438083551;
assign addr[34460]= 1197050035;
assign addr[34461]= 931758235;
assign addr[34462]= 647584304;
assign addr[34463]= 350287041;
assign addr[34464]= 45891193;
assign addr[34465]= -259434643;
assign addr[34466]= -559503022;
assign addr[34467]= -848233042;
assign addr[34468]= -1119773573;
assign addr[34469]= -1368621831;
assign addr[34470]= -1589734894;
assign addr[34471]= -1778631892;
assign addr[34472]= -1931484818;
assign addr[34473]= -2045196100;
assign addr[34474]= -2117461370;
assign addr[34475]= -2146816171;
assign addr[34476]= -2132665626;
assign addr[34477]= -2075296495;
assign addr[34478]= -1975871368;
assign addr[34479]= -1836405100;
assign addr[34480]= -1659723983;
assign addr[34481]= -1449408469;
assign addr[34482]= -1209720613;
assign addr[34483]= -945517704;
assign addr[34484]= -662153826;
assign addr[34485]= -365371365;
assign addr[34486]= -61184634;
assign addr[34487]= 244242007;
assign addr[34488]= 544719071;
assign addr[34489]= 834157373;
assign addr[34490]= 1106691431;
assign addr[34491]= 1356798326;
assign addr[34492]= 1579409630;
assign addr[34493]= 1770014111;
assign addr[34494]= 1924749160;
assign addr[34495]= 2040479063;
assign addr[34496]= 2114858546;
assign addr[34497]= 2146380306;
assign addr[34498]= 2134405552;
assign addr[34499]= 2079176953;
assign addr[34500]= 1981813720;
assign addr[34501]= 1844288924;
assign addr[34502]= 1669389513;
assign addr[34503]= 1460659832;
assign addr[34504]= 1222329801;
assign addr[34505]= 959229189;
assign addr[34506]= 676689746;
assign addr[34507]= 380437148;
assign addr[34508]= 76474970;
assign addr[34509]= -229036977;
assign addr[34510]= -529907477;
assign addr[34511]= -820039373;
assign addr[34512]= -1093553126;
assign addr[34513]= -1344905966;
assign addr[34514]= -1569004214;
assign addr[34515]= -1761306505;
assign addr[34516]= -1917915825;
assign addr[34517]= -2035658475;
assign addr[34518]= -2112148396;
assign addr[34519]= -2145835515;
assign addr[34520]= -2136037160;
assign addr[34521]= -2082951896;
assign addr[34522]= -1987655498;
assign addr[34523]= -1852079154;
assign addr[34524]= -1678970324;
assign addr[34525]= -1471837070;
assign addr[34526]= -1234876957;
assign addr[34527]= -972891995;
assign addr[34528]= -691191324;
assign addr[34529]= -395483624;
assign addr[34530]= -91761426;
assign addr[34531]= 213820322;
assign addr[34532]= 515068990;
assign addr[34533]= 805879757;
assign addr[34534]= 1080359326;
assign addr[34535]= 1332945355;
assign addr[34536]= 1558519173;
assign addr[34537]= 1752509516;
assign addr[34538]= 1910985158;
assign addr[34539]= 2030734582;
assign addr[34540]= 2109331059;
assign addr[34541]= 2145181827;
assign addr[34542]= 2137560369;
assign addr[34543]= 2086621133;
assign addr[34544]= 1993396407;
assign addr[34545]= 1859775393;
assign addr[34546]= 1688465931;
assign addr[34547]= 1482939614;
assign addr[34548]= 1247361445;
assign addr[34549]= 986505429;
assign addr[34550]= 705657826;
assign addr[34551]= 410510029;
assign addr[34552]= 107043224;
assign addr[34553]= -198592817;
assign addr[34554]= -500204365;
assign addr[34555]= -791679244;
assign addr[34556]= -1067110699;
assign addr[34557]= -1320917099;
assign addr[34558]= -1547955041;
assign addr[34559]= -1743623590;
assign addr[34560]= -1903957513;
assign addr[34561]= -2025707632;
assign addr[34562]= -2106406677;
assign addr[34563]= -2144419275;
assign addr[34564]= -2138975100;
assign addr[34565]= -2090184478;
assign addr[34566]= -1999036154;
assign addr[34567]= -1867377253;
assign addr[34568]= -1697875851;
assign addr[34569]= -1493966902;
assign addr[34570]= -1259782632;
assign addr[34571]= -1000068799;
assign addr[34572]= -720088517;
assign addr[34573]= -425515602;
assign addr[34574]= -122319591;
assign addr[34575]= 183355234;
assign addr[34576]= 485314355;
assign addr[34577]= 777438554;
assign addr[34578]= 1053807919;
assign addr[34579]= 1308821808;
assign addr[34580]= 1537312353;
assign addr[34581]= 1734649179;
assign addr[34582]= 1896833245;
assign addr[34583]= 2020577882;
assign addr[34584]= 2103375398;
assign addr[34585]= 2143547897;
assign addr[34586]= 2140281282;
assign addr[34587]= 2093641749;
assign addr[34588]= 2004574453;
assign addr[34589]= 1874884346;
assign addr[34590]= 1707199606;
assign addr[34591]= 1504918373;
assign addr[34592]= 1272139887;
assign addr[34593]= 1013581418;
assign addr[34594]= 734482665;
assign addr[34595]= 440499581;
assign addr[34596]= 137589750;
assign addr[34597]= -168108346;
assign addr[34598]= -470399716;
assign addr[34599]= -763158411;
assign addr[34600]= -1040451659;
assign addr[34601]= -1296660098;
assign addr[34602]= -1526591649;
assign addr[34603]= -1725586737;
assign addr[34604]= -1889612716;
assign addr[34605]= -2015345591;
assign addr[34606]= -2100237377;
assign addr[34607]= -2142567738;
assign addr[34608]= -2141478848;
assign addr[34609]= -2096992772;
assign addr[34610]= -2010011024;
assign addr[34611]= -1882296293;
assign addr[34612]= -1716436725;
assign addr[34613]= -1515793473;
assign addr[34614]= -1284432584;
assign addr[34615]= -1027042599;
assign addr[34616]= -748839539;
assign addr[34617]= -455461206;
assign addr[34618]= -152852926;
assign addr[34619]= 152852926;
assign addr[34620]= 455461206;
assign addr[34621]= 748839539;
assign addr[34622]= 1027042599;
assign addr[34623]= 1284432584;
assign addr[34624]= 1515793473;
assign addr[34625]= 1716436725;
assign addr[34626]= 1882296293;
assign addr[34627]= 2010011024;
assign addr[34628]= 2096992772;
assign addr[34629]= 2141478848;
assign addr[34630]= 2142567738;
assign addr[34631]= 2100237377;
assign addr[34632]= 2015345591;
assign addr[34633]= 1889612716;
assign addr[34634]= 1725586737;
assign addr[34635]= 1526591649;
assign addr[34636]= 1296660098;
assign addr[34637]= 1040451659;
assign addr[34638]= 763158411;
assign addr[34639]= 470399716;
assign addr[34640]= 168108346;
assign addr[34641]= -137589750;
assign addr[34642]= -440499581;
assign addr[34643]= -734482665;
assign addr[34644]= -1013581418;
assign addr[34645]= -1272139887;
assign addr[34646]= -1504918373;
assign addr[34647]= -1707199606;
assign addr[34648]= -1874884346;
assign addr[34649]= -2004574453;
assign addr[34650]= -2093641749;
assign addr[34651]= -2140281282;
assign addr[34652]= -2143547897;
assign addr[34653]= -2103375398;
assign addr[34654]= -2020577882;
assign addr[34655]= -1896833245;
assign addr[34656]= -1734649179;
assign addr[34657]= -1537312353;
assign addr[34658]= -1308821808;
assign addr[34659]= -1053807919;
assign addr[34660]= -777438554;
assign addr[34661]= -485314355;
assign addr[34662]= -183355234;
assign addr[34663]= 122319591;
assign addr[34664]= 425515602;
assign addr[34665]= 720088517;
assign addr[34666]= 1000068799;
assign addr[34667]= 1259782632;
assign addr[34668]= 1493966902;
assign addr[34669]= 1697875851;
assign addr[34670]= 1867377253;
assign addr[34671]= 1999036154;
assign addr[34672]= 2090184478;
assign addr[34673]= 2138975100;
assign addr[34674]= 2144419275;
assign addr[34675]= 2106406677;
assign addr[34676]= 2025707632;
assign addr[34677]= 1903957513;
assign addr[34678]= 1743623590;
assign addr[34679]= 1547955041;
assign addr[34680]= 1320917099;
assign addr[34681]= 1067110699;
assign addr[34682]= 791679244;
assign addr[34683]= 500204365;
assign addr[34684]= 198592817;
assign addr[34685]= -107043224;
assign addr[34686]= -410510029;
assign addr[34687]= -705657826;
assign addr[34688]= -986505429;
assign addr[34689]= -1247361445;
assign addr[34690]= -1482939614;
assign addr[34691]= -1688465931;
assign addr[34692]= -1859775393;
assign addr[34693]= -1993396407;
assign addr[34694]= -2086621133;
assign addr[34695]= -2137560369;
assign addr[34696]= -2145181827;
assign addr[34697]= -2109331059;
assign addr[34698]= -2030734582;
assign addr[34699]= -1910985158;
assign addr[34700]= -1752509516;
assign addr[34701]= -1558519173;
assign addr[34702]= -1332945355;
assign addr[34703]= -1080359326;
assign addr[34704]= -805879757;
assign addr[34705]= -515068990;
assign addr[34706]= -213820322;
assign addr[34707]= 91761426;
assign addr[34708]= 395483624;
assign addr[34709]= 691191324;
assign addr[34710]= 972891995;
assign addr[34711]= 1234876957;
assign addr[34712]= 1471837070;
assign addr[34713]= 1678970324;
assign addr[34714]= 1852079154;
assign addr[34715]= 1987655498;
assign addr[34716]= 2082951896;
assign addr[34717]= 2136037160;
assign addr[34718]= 2145835515;
assign addr[34719]= 2112148396;
assign addr[34720]= 2035658475;
assign addr[34721]= 1917915825;
assign addr[34722]= 1761306505;
assign addr[34723]= 1569004214;
assign addr[34724]= 1344905966;
assign addr[34725]= 1093553126;
assign addr[34726]= 820039373;
assign addr[34727]= 529907477;
assign addr[34728]= 229036977;
assign addr[34729]= -76474970;
assign addr[34730]= -380437148;
assign addr[34731]= -676689746;
assign addr[34732]= -959229189;
assign addr[34733]= -1222329801;
assign addr[34734]= -1460659832;
assign addr[34735]= -1669389513;
assign addr[34736]= -1844288924;
assign addr[34737]= -1981813720;
assign addr[34738]= -2079176953;
assign addr[34739]= -2134405552;
assign addr[34740]= -2146380306;
assign addr[34741]= -2114858546;
assign addr[34742]= -2040479063;
assign addr[34743]= -1924749160;
assign addr[34744]= -1770014111;
assign addr[34745]= -1579409630;
assign addr[34746]= -1356798326;
assign addr[34747]= -1106691431;
assign addr[34748]= -834157373;
assign addr[34749]= -544719071;
assign addr[34750]= -244242007;
assign addr[34751]= 61184634;
assign addr[34752]= 365371365;
assign addr[34753]= 662153826;
assign addr[34754]= 945517704;
assign addr[34755]= 1209720613;
assign addr[34756]= 1449408469;
assign addr[34757]= 1659723983;
assign addr[34758]= 1836405100;
assign addr[34759]= 1975871368;
assign addr[34760]= 2075296495;
assign addr[34761]= 2132665626;
assign addr[34762]= 2146816171;
assign addr[34763]= 2117461370;
assign addr[34764]= 2045196100;
assign addr[34765]= 1931484818;
assign addr[34766]= 1778631892;
assign addr[34767]= 1589734894;
assign addr[34768]= 1368621831;
assign addr[34769]= 1119773573;
assign addr[34770]= 848233042;
assign addr[34771]= 559503022;
assign addr[34772]= 259434643;
assign addr[34773]= -45891193;
assign addr[34774]= -350287041;
assign addr[34775]= -647584304;
assign addr[34776]= -931758235;
assign addr[34777]= -1197050035;
assign addr[34778]= -1438083551;
assign addr[34779]= -1649974225;
assign addr[34780]= -1828428082;
assign addr[34781]= -1969828744;
assign addr[34782]= -2071310720;
assign addr[34783]= -2130817471;
assign addr[34784]= -2147143090;
assign addr[34785]= -2119956737;
assign addr[34786]= -2049809346;
assign addr[34787]= -1938122457;
assign addr[34788]= -1787159411;
assign addr[34789]= -1599979481;
assign addr[34790]= -1380375881;
assign addr[34791]= -1132798888;
assign addr[34792]= -862265664;
assign addr[34793]= -574258580;
assign addr[34794]= -274614114;
assign addr[34795]= 30595422;
assign addr[34796]= 335184940;
assign addr[34797]= 632981917;
assign addr[34798]= 917951481;
assign addr[34799]= 1184318708;
assign addr[34800]= 1426685652;
assign addr[34801]= 1640140734;
assign addr[34802]= 1820358275;
assign addr[34803]= 1963686155;
assign addr[34804]= 2067219829;
assign addr[34805]= 2128861181;
assign addr[34806]= 2147361045;
assign addr[34807]= 2122344521;
assign addr[34808]= 2054318569;
assign addr[34809]= 1944661739;
assign addr[34810]= 1795596234;
assign addr[34811]= 1610142873;
assign addr[34812]= 1392059879;
assign addr[34813]= 1145766716;
assign addr[34814]= 876254528;
assign addr[34815]= 588984994;
assign addr[34816]= 289779648;
assign addr[34817]= -15298099;
assign addr[34818]= -320065829;
assign addr[34819]= -618347408;
assign addr[34820]= -904098143;
assign addr[34821]= -1171527280;
assign addr[34822]= -1415215352;
assign addr[34823]= -1630224009;
assign addr[34824]= -1812196087;
assign addr[34825]= -1957443913;
assign addr[34826]= -2063024031;
assign addr[34827]= -2126796855;
assign addr[34828]= -2147470025;
assign addr[34829]= -2124624598;
assign addr[34830]= -2058723538;
assign addr[34831]= -1951102334;
assign addr[34832]= -1803941934;
assign addr[34833]= -1620224553;
assign addr[34834]= -1403673233;
assign addr[34835]= -1158676398;
assign addr[34836]= -890198924;
assign addr[34837]= -603681519;
assign addr[34838]= -304930476;
assign addr[34839]= 0;
assign addr[34840]= 304930476;
assign addr[34841]= 603681519;
assign addr[34842]= 890198924;
assign addr[34843]= 1158676398;
assign addr[34844]= 1403673233;
assign addr[34845]= 1620224553;
assign addr[34846]= 1803941934;
assign addr[34847]= 1951102334;
assign addr[34848]= 2058723538;
assign addr[34849]= 2124624598;
assign addr[34850]= 2147470025;
assign addr[34851]= 2126796855;
assign addr[34852]= 2063024031;
assign addr[34853]= 1957443913;
assign addr[34854]= 1812196087;
assign addr[34855]= 1630224009;
assign addr[34856]= 1415215352;
assign addr[34857]= 1171527280;
assign addr[34858]= 904098143;
assign addr[34859]= 618347408;
assign addr[34860]= 320065829;
assign addr[34861]= 15298099;
assign addr[34862]= -289779648;
assign addr[34863]= -588984994;
assign addr[34864]= -876254528;
assign addr[34865]= -1145766716;
assign addr[34866]= -1392059879;
assign addr[34867]= -1610142873;
assign addr[34868]= -1795596234;
assign addr[34869]= -1944661739;
assign addr[34870]= -2054318569;
assign addr[34871]= -2122344521;
assign addr[34872]= -2147361045;
assign addr[34873]= -2128861181;
assign addr[34874]= -2067219829;
assign addr[34875]= -1963686155;
assign addr[34876]= -1820358275;
assign addr[34877]= -1640140734;
assign addr[34878]= -1426685652;
assign addr[34879]= -1184318708;
assign addr[34880]= -917951481;
assign addr[34881]= -632981917;
assign addr[34882]= -335184940;
assign addr[34883]= -30595422;
assign addr[34884]= 274614114;
assign addr[34885]= 574258580;
assign addr[34886]= 862265664;
assign addr[34887]= 1132798888;
assign addr[34888]= 1380375881;
assign addr[34889]= 1599979481;
assign addr[34890]= 1787159411;
assign addr[34891]= 1938122457;
assign addr[34892]= 2049809346;
assign addr[34893]= 2119956737;
assign addr[34894]= 2147143090;
assign addr[34895]= 2130817471;
assign addr[34896]= 2071310720;
assign addr[34897]= 1969828744;
assign addr[34898]= 1828428082;
assign addr[34899]= 1649974225;
assign addr[34900]= 1438083551;
assign addr[34901]= 1197050035;
assign addr[34902]= 931758235;
assign addr[34903]= 647584304;
assign addr[34904]= 350287041;
assign addr[34905]= 45891193;
assign addr[34906]= -259434643;
assign addr[34907]= -559503022;
assign addr[34908]= -848233042;
assign addr[34909]= -1119773573;
assign addr[34910]= -1368621831;
assign addr[34911]= -1589734894;
assign addr[34912]= -1778631892;
assign addr[34913]= -1931484818;
assign addr[34914]= -2045196100;
assign addr[34915]= -2117461370;
assign addr[34916]= -2146816171;
assign addr[34917]= -2132665626;
assign addr[34918]= -2075296495;
assign addr[34919]= -1975871368;
assign addr[34920]= -1836405100;
assign addr[34921]= -1659723983;
assign addr[34922]= -1449408469;
assign addr[34923]= -1209720613;
assign addr[34924]= -945517704;
assign addr[34925]= -662153826;
assign addr[34926]= -365371365;
assign addr[34927]= -61184634;
assign addr[34928]= 244242007;
assign addr[34929]= 544719071;
assign addr[34930]= 834157373;
assign addr[34931]= 1106691431;
assign addr[34932]= 1356798326;
assign addr[34933]= 1579409630;
assign addr[34934]= 1770014111;
assign addr[34935]= 1924749160;
assign addr[34936]= 2040479063;
assign addr[34937]= 2114858546;
assign addr[34938]= 2146380306;
assign addr[34939]= 2134405552;
assign addr[34940]= 2079176953;
assign addr[34941]= 1981813720;
assign addr[34942]= 1844288924;
assign addr[34943]= 1669389513;
assign addr[34944]= 1460659832;
assign addr[34945]= 1222329801;
assign addr[34946]= 959229189;
assign addr[34947]= 676689746;
assign addr[34948]= 380437148;
assign addr[34949]= 76474970;
assign addr[34950]= -229036977;
assign addr[34951]= -529907477;
assign addr[34952]= -820039373;
assign addr[34953]= -1093553126;
assign addr[34954]= -1344905966;
assign addr[34955]= -1569004214;
assign addr[34956]= -1761306505;
assign addr[34957]= -1917915825;
assign addr[34958]= -2035658475;
assign addr[34959]= -2112148396;
assign addr[34960]= -2145835515;
assign addr[34961]= -2136037160;
assign addr[34962]= -2082951896;
assign addr[34963]= -1987655498;
assign addr[34964]= -1852079154;
assign addr[34965]= -1678970324;
assign addr[34966]= -1471837070;
assign addr[34967]= -1234876957;
assign addr[34968]= -972891995;
assign addr[34969]= -691191324;
assign addr[34970]= -395483624;
assign addr[34971]= -91761426;
assign addr[34972]= 213820322;
assign addr[34973]= 515068990;
assign addr[34974]= 805879757;
assign addr[34975]= 1080359326;
assign addr[34976]= 1332945355;
assign addr[34977]= 1558519173;
assign addr[34978]= 1752509516;
assign addr[34979]= 1910985158;
assign addr[34980]= 2030734582;
assign addr[34981]= 2109331059;
assign addr[34982]= 2145181827;
assign addr[34983]= 2137560369;
assign addr[34984]= 2086621133;
assign addr[34985]= 1993396407;
assign addr[34986]= 1859775393;
assign addr[34987]= 1688465931;
assign addr[34988]= 1482939614;
assign addr[34989]= 1247361445;
assign addr[34990]= 986505429;
assign addr[34991]= 705657826;
assign addr[34992]= 410510029;
assign addr[34993]= 107043224;
assign addr[34994]= -198592817;
assign addr[34995]= -500204365;
assign addr[34996]= -791679244;
assign addr[34997]= -1067110699;
assign addr[34998]= -1320917099;
assign addr[34999]= -1547955041;
assign addr[35000]= -1743623590;
assign addr[35001]= -1903957513;
assign addr[35002]= -2025707632;
assign addr[35003]= -2106406677;
assign addr[35004]= -2144419275;
assign addr[35005]= -2138975100;
assign addr[35006]= -2090184478;
assign addr[35007]= -1999036154;
assign addr[35008]= -1867377253;
assign addr[35009]= -1697875851;
assign addr[35010]= -1493966902;
assign addr[35011]= -1259782632;
assign addr[35012]= -1000068799;
assign addr[35013]= -720088517;
assign addr[35014]= -425515602;
assign addr[35015]= -122319591;
assign addr[35016]= 183355234;
assign addr[35017]= 485314355;
assign addr[35018]= 777438554;
assign addr[35019]= 1053807919;
assign addr[35020]= 1308821808;
assign addr[35021]= 1537312353;
assign addr[35022]= 1734649179;
assign addr[35023]= 1896833245;
assign addr[35024]= 2020577882;
assign addr[35025]= 2103375398;
assign addr[35026]= 2143547897;
assign addr[35027]= 2140281282;
assign addr[35028]= 2093641749;
assign addr[35029]= 2004574453;
assign addr[35030]= 1874884346;
assign addr[35031]= 1707199606;
assign addr[35032]= 1504918373;
assign addr[35033]= 1272139887;
assign addr[35034]= 1013581418;
assign addr[35035]= 734482665;
assign addr[35036]= 440499581;
assign addr[35037]= 137589750;
assign addr[35038]= -168108346;
assign addr[35039]= -470399716;
assign addr[35040]= -763158411;
assign addr[35041]= -1040451659;
assign addr[35042]= -1296660098;
assign addr[35043]= -1526591649;
assign addr[35044]= -1725586737;
assign addr[35045]= -1889612716;
assign addr[35046]= -2015345591;
assign addr[35047]= -2100237377;
assign addr[35048]= -2142567738;
assign addr[35049]= -2141478848;
assign addr[35050]= -2096992772;
assign addr[35051]= -2010011024;
assign addr[35052]= -1882296293;
assign addr[35053]= -1716436725;
assign addr[35054]= -1515793473;
assign addr[35055]= -1284432584;
assign addr[35056]= -1027042599;
assign addr[35057]= -748839539;
assign addr[35058]= -455461206;
assign addr[35059]= -152852926;
assign addr[35060]= 152852926;
assign addr[35061]= 455461206;
assign addr[35062]= 748839539;
assign addr[35063]= 1027042599;
assign addr[35064]= 1284432584;
assign addr[35065]= 1515793473;
assign addr[35066]= 1716436725;
assign addr[35067]= 1882296293;
assign addr[35068]= 2010011024;
assign addr[35069]= 2096992772;
assign addr[35070]= 2141478848;
assign addr[35071]= 2142567738;
assign addr[35072]= 2100237377;
assign addr[35073]= 2015345591;
assign addr[35074]= 1889612716;
assign addr[35075]= 1725586737;
assign addr[35076]= 1526591649;
assign addr[35077]= 1296660098;
assign addr[35078]= 1040451659;
assign addr[35079]= 763158411;
assign addr[35080]= 470399716;
assign addr[35081]= 168108346;
assign addr[35082]= -137589750;
assign addr[35083]= -440499581;
assign addr[35084]= -734482665;
assign addr[35085]= -1013581418;
assign addr[35086]= -1272139887;
assign addr[35087]= -1504918373;
assign addr[35088]= -1707199606;
assign addr[35089]= -1874884346;
assign addr[35090]= -2004574453;
assign addr[35091]= -2093641749;
assign addr[35092]= -2140281282;
assign addr[35093]= -2143547897;
assign addr[35094]= -2103375398;
assign addr[35095]= -2020577882;
assign addr[35096]= -1896833245;
assign addr[35097]= -1734649179;
assign addr[35098]= -1537312353;
assign addr[35099]= -1308821808;
assign addr[35100]= -1053807919;
assign addr[35101]= -777438554;
assign addr[35102]= -485314355;
assign addr[35103]= -183355234;
assign addr[35104]= 122319591;
assign addr[35105]= 425515602;
assign addr[35106]= 720088517;
assign addr[35107]= 1000068799;
assign addr[35108]= 1259782632;
assign addr[35109]= 1493966902;
assign addr[35110]= 1697875851;
assign addr[35111]= 1867377253;
assign addr[35112]= 1999036154;
assign addr[35113]= 2090184478;
assign addr[35114]= 2138975100;
assign addr[35115]= 2144419275;
assign addr[35116]= 2106406677;
assign addr[35117]= 2025707632;
assign addr[35118]= 1903957513;
assign addr[35119]= 1743623590;
assign addr[35120]= 1547955041;
assign addr[35121]= 1320917099;
assign addr[35122]= 1067110699;
assign addr[35123]= 791679244;
assign addr[35124]= 500204365;
assign addr[35125]= 198592817;
assign addr[35126]= -107043224;
assign addr[35127]= -410510029;
assign addr[35128]= -705657826;
assign addr[35129]= -986505429;
assign addr[35130]= -1247361445;
assign addr[35131]= -1482939614;
assign addr[35132]= -1688465931;
assign addr[35133]= -1859775393;
assign addr[35134]= -1993396407;
assign addr[35135]= -2086621133;
assign addr[35136]= -2137560369;
assign addr[35137]= -2145181827;
assign addr[35138]= -2109331059;
assign addr[35139]= -2030734582;
assign addr[35140]= -1910985158;
assign addr[35141]= -1752509516;
assign addr[35142]= -1558519173;
assign addr[35143]= -1332945355;
assign addr[35144]= -1080359326;
assign addr[35145]= -805879757;
assign addr[35146]= -515068990;
assign addr[35147]= -213820322;
assign addr[35148]= 91761426;
assign addr[35149]= 395483624;
assign addr[35150]= 691191324;
assign addr[35151]= 972891995;
assign addr[35152]= 1234876957;
assign addr[35153]= 1471837070;
assign addr[35154]= 1678970324;
assign addr[35155]= 1852079154;
assign addr[35156]= 1987655498;
assign addr[35157]= 2082951896;
assign addr[35158]= 2136037160;
assign addr[35159]= 2145835515;
assign addr[35160]= 2112148396;
assign addr[35161]= 2035658475;
assign addr[35162]= 1917915825;
assign addr[35163]= 1761306505;
assign addr[35164]= 1569004214;
assign addr[35165]= 1344905966;
assign addr[35166]= 1093553126;
assign addr[35167]= 820039373;
assign addr[35168]= 529907477;
assign addr[35169]= 229036977;
assign addr[35170]= -76474970;
assign addr[35171]= -380437148;
assign addr[35172]= -676689746;
assign addr[35173]= -959229189;
assign addr[35174]= -1222329801;
assign addr[35175]= -1460659832;
assign addr[35176]= -1669389513;
assign addr[35177]= -1844288924;
assign addr[35178]= -1981813720;
assign addr[35179]= -2079176953;
assign addr[35180]= -2134405552;
assign addr[35181]= -2146380306;
assign addr[35182]= -2114858546;
assign addr[35183]= -2040479063;
assign addr[35184]= -1924749160;
assign addr[35185]= -1770014111;
assign addr[35186]= -1579409630;
assign addr[35187]= -1356798326;
assign addr[35188]= -1106691431;
assign addr[35189]= -834157373;
assign addr[35190]= -544719071;
assign addr[35191]= -244242007;
assign addr[35192]= 61184634;
assign addr[35193]= 365371365;
assign addr[35194]= 662153826;
assign addr[35195]= 945517704;
assign addr[35196]= 1209720613;
assign addr[35197]= 1449408469;
assign addr[35198]= 1659723983;
assign addr[35199]= 1836405100;
assign addr[35200]= 1975871368;
assign addr[35201]= 2075296495;
assign addr[35202]= 2132665626;
assign addr[35203]= 2146816171;
assign addr[35204]= 2117461370;
assign addr[35205]= 2045196100;
assign addr[35206]= 1931484818;
assign addr[35207]= 1778631892;
assign addr[35208]= 1589734894;
assign addr[35209]= 1368621831;
assign addr[35210]= 1119773573;
assign addr[35211]= 848233042;
assign addr[35212]= 559503022;
assign addr[35213]= 259434643;
assign addr[35214]= -45891193;
assign addr[35215]= -350287041;
assign addr[35216]= -647584304;
assign addr[35217]= -931758235;
assign addr[35218]= -1197050035;
assign addr[35219]= -1438083551;
assign addr[35220]= -1649974225;
assign addr[35221]= -1828428082;
assign addr[35222]= -1969828744;
assign addr[35223]= -2071310720;
assign addr[35224]= -2130817471;
assign addr[35225]= -2147143090;
assign addr[35226]= -2119956737;
assign addr[35227]= -2049809346;
assign addr[35228]= -1938122457;
assign addr[35229]= -1787159411;
assign addr[35230]= -1599979481;
assign addr[35231]= -1380375881;
assign addr[35232]= -1132798888;
assign addr[35233]= -862265664;
assign addr[35234]= -574258580;
assign addr[35235]= -274614114;
assign addr[35236]= 30595422;
assign addr[35237]= 335184940;
assign addr[35238]= 632981917;
assign addr[35239]= 917951481;
assign addr[35240]= 1184318708;
assign addr[35241]= 1426685652;
assign addr[35242]= 1640140734;
assign addr[35243]= 1820358275;
assign addr[35244]= 1963686155;
assign addr[35245]= 2067219829;
assign addr[35246]= 2128861181;
assign addr[35247]= 2147361045;
assign addr[35248]= 2122344521;
assign addr[35249]= 2054318569;
assign addr[35250]= 1944661739;
assign addr[35251]= 1795596234;
assign addr[35252]= 1610142873;
assign addr[35253]= 1392059879;
assign addr[35254]= 1145766716;
assign addr[35255]= 876254528;
assign addr[35256]= 588984994;
assign addr[35257]= 289779648;
assign addr[35258]= -15298099;
assign addr[35259]= -320065829;
assign addr[35260]= -618347408;
assign addr[35261]= -904098143;
assign addr[35262]= -1171527280;
assign addr[35263]= -1415215352;
assign addr[35264]= -1630224009;
assign addr[35265]= -1812196087;
assign addr[35266]= -1957443913;
assign addr[35267]= -2063024031;
assign addr[35268]= -2126796855;
assign addr[35269]= -2147470025;
assign addr[35270]= -2124624598;
assign addr[35271]= -2058723538;
assign addr[35272]= -1951102334;
assign addr[35273]= -1803941934;
assign addr[35274]= -1620224553;
assign addr[35275]= -1403673233;
assign addr[35276]= -1158676398;
assign addr[35277]= -890198924;
assign addr[35278]= -603681519;
assign addr[35279]= -304930476;
assign addr[35280]= 0;
assign addr[35281]= 304930476;
assign addr[35282]= 603681519;
assign addr[35283]= 890198924;
assign addr[35284]= 1158676398;
assign addr[35285]= 1403673233;
assign addr[35286]= 1620224553;
assign addr[35287]= 1803941934;
assign addr[35288]= 1951102334;
assign addr[35289]= 2058723538;
assign addr[35290]= 2124624598;
assign addr[35291]= 2147470025;
assign addr[35292]= 2126796855;
assign addr[35293]= 2063024031;
assign addr[35294]= 1957443913;
assign addr[35295]= 1812196087;
assign addr[35296]= 1630224009;
assign addr[35297]= 1415215352;
assign addr[35298]= 1171527280;
assign addr[35299]= 904098143;
assign addr[35300]= 618347408;
assign addr[35301]= 320065829;
assign addr[35302]= 15298099;
assign addr[35303]= -289779648;
assign addr[35304]= -588984994;
assign addr[35305]= -876254528;
assign addr[35306]= -1145766716;
assign addr[35307]= -1392059879;
assign addr[35308]= -1610142873;
assign addr[35309]= -1795596234;
assign addr[35310]= -1944661739;
assign addr[35311]= -2054318569;
assign addr[35312]= -2122344521;
assign addr[35313]= -2147361045;
assign addr[35314]= -2128861181;
assign addr[35315]= -2067219829;
assign addr[35316]= -1963686155;
assign addr[35317]= -1820358275;
assign addr[35318]= -1640140734;
assign addr[35319]= -1426685652;
assign addr[35320]= -1184318708;
assign addr[35321]= -917951481;
assign addr[35322]= -632981917;
assign addr[35323]= -335184940;
assign addr[35324]= -30595422;
assign addr[35325]= 274614114;
assign addr[35326]= 574258580;
assign addr[35327]= 862265664;
assign addr[35328]= 1132798888;
assign addr[35329]= 1380375881;
assign addr[35330]= 1599979481;
assign addr[35331]= 1787159411;
assign addr[35332]= 1938122457;
assign addr[35333]= 2049809346;
assign addr[35334]= 2119956737;
assign addr[35335]= 2147143090;
assign addr[35336]= 2130817471;
assign addr[35337]= 2071310720;
assign addr[35338]= 1969828744;
assign addr[35339]= 1828428082;
assign addr[35340]= 1649974225;
assign addr[35341]= 1438083551;
assign addr[35342]= 1197050035;
assign addr[35343]= 931758235;
assign addr[35344]= 647584304;
assign addr[35345]= 350287041;
assign addr[35346]= 45891193;
assign addr[35347]= -259434643;
assign addr[35348]= -559503022;
assign addr[35349]= -848233042;
assign addr[35350]= -1119773573;
assign addr[35351]= -1368621831;
assign addr[35352]= -1589734894;
assign addr[35353]= -1778631892;
assign addr[35354]= -1931484818;
assign addr[35355]= -2045196100;
assign addr[35356]= -2117461370;
assign addr[35357]= -2146816171;
assign addr[35358]= -2132665626;
assign addr[35359]= -2075296495;
assign addr[35360]= -1975871368;
assign addr[35361]= -1836405100;
assign addr[35362]= -1659723983;
assign addr[35363]= -1449408469;
assign addr[35364]= -1209720613;
assign addr[35365]= -945517704;
assign addr[35366]= -662153826;
assign addr[35367]= -365371365;
assign addr[35368]= -61184634;
assign addr[35369]= 244242007;
assign addr[35370]= 544719071;
assign addr[35371]= 834157373;
assign addr[35372]= 1106691431;
assign addr[35373]= 1356798326;
assign addr[35374]= 1579409630;
assign addr[35375]= 1770014111;
assign addr[35376]= 1924749160;
assign addr[35377]= 2040479063;
assign addr[35378]= 2114858546;
assign addr[35379]= 2146380306;
assign addr[35380]= 2134405552;
assign addr[35381]= 2079176953;
assign addr[35382]= 1981813720;
assign addr[35383]= 1844288924;
assign addr[35384]= 1669389513;
assign addr[35385]= 1460659832;
assign addr[35386]= 1222329801;
assign addr[35387]= 959229189;
assign addr[35388]= 676689746;
assign addr[35389]= 380437148;
assign addr[35390]= 76474970;
assign addr[35391]= -229036977;
assign addr[35392]= -529907477;
assign addr[35393]= -820039373;
assign addr[35394]= -1093553126;
assign addr[35395]= -1344905966;
assign addr[35396]= -1569004214;
assign addr[35397]= -1761306505;
assign addr[35398]= -1917915825;
assign addr[35399]= -2035658475;
assign addr[35400]= -2112148396;
assign addr[35401]= -2145835515;
assign addr[35402]= -2136037160;
assign addr[35403]= -2082951896;
assign addr[35404]= -1987655498;
assign addr[35405]= -1852079154;
assign addr[35406]= -1678970324;
assign addr[35407]= -1471837070;
assign addr[35408]= -1234876957;
assign addr[35409]= -972891995;
assign addr[35410]= -691191324;
assign addr[35411]= -395483624;
assign addr[35412]= -91761426;
assign addr[35413]= 213820322;
assign addr[35414]= 515068990;
assign addr[35415]= 805879757;
assign addr[35416]= 1080359326;
assign addr[35417]= 1332945355;
assign addr[35418]= 1558519173;
assign addr[35419]= 1752509516;
assign addr[35420]= 1910985158;
assign addr[35421]= 2030734582;
assign addr[35422]= 2109331059;
assign addr[35423]= 2145181827;
assign addr[35424]= 2137560369;
assign addr[35425]= 2086621133;
assign addr[35426]= 1993396407;
assign addr[35427]= 1859775393;
assign addr[35428]= 1688465931;
assign addr[35429]= 1482939614;
assign addr[35430]= 1247361445;
assign addr[35431]= 986505429;
assign addr[35432]= 705657826;
assign addr[35433]= 410510029;
assign addr[35434]= 107043224;
assign addr[35435]= -198592817;
assign addr[35436]= -500204365;
assign addr[35437]= -791679244;
assign addr[35438]= -1067110699;
assign addr[35439]= -1320917099;
assign addr[35440]= -1547955041;
assign addr[35441]= -1743623590;
assign addr[35442]= -1903957513;
assign addr[35443]= -2025707632;
assign addr[35444]= -2106406677;
assign addr[35445]= -2144419275;
assign addr[35446]= -2138975100;
assign addr[35447]= -2090184478;
assign addr[35448]= -1999036154;
assign addr[35449]= -1867377253;
assign addr[35450]= -1697875851;
assign addr[35451]= -1493966902;
assign addr[35452]= -1259782632;
assign addr[35453]= -1000068799;
assign addr[35454]= -720088517;
assign addr[35455]= -425515602;
assign addr[35456]= -122319591;
assign addr[35457]= 183355234;
assign addr[35458]= 485314355;
assign addr[35459]= 777438554;
assign addr[35460]= 1053807919;
assign addr[35461]= 1308821808;
assign addr[35462]= 1537312353;
assign addr[35463]= 1734649179;
assign addr[35464]= 1896833245;
assign addr[35465]= 2020577882;
assign addr[35466]= 2103375398;
assign addr[35467]= 2143547897;
assign addr[35468]= 2140281282;
assign addr[35469]= 2093641749;
assign addr[35470]= 2004574453;
assign addr[35471]= 1874884346;
assign addr[35472]= 1707199606;
assign addr[35473]= 1504918373;
assign addr[35474]= 1272139887;
assign addr[35475]= 1013581418;
assign addr[35476]= 734482665;
assign addr[35477]= 440499581;
assign addr[35478]= 137589750;
assign addr[35479]= -168108346;
assign addr[35480]= -470399716;
assign addr[35481]= -763158411;
assign addr[35482]= -1040451659;
assign addr[35483]= -1296660098;
assign addr[35484]= -1526591649;
assign addr[35485]= -1725586737;
assign addr[35486]= -1889612716;
assign addr[35487]= -2015345591;
assign addr[35488]= -2100237377;
assign addr[35489]= -2142567738;
assign addr[35490]= -2141478848;
assign addr[35491]= -2096992772;
assign addr[35492]= -2010011024;
assign addr[35493]= -1882296293;
assign addr[35494]= -1716436725;
assign addr[35495]= -1515793473;
assign addr[35496]= -1284432584;
assign addr[35497]= -1027042599;
assign addr[35498]= -748839539;
assign addr[35499]= -455461206;
assign addr[35500]= -152852926;
assign addr[35501]= 152852926;
assign addr[35502]= 455461206;
assign addr[35503]= 748839539;
assign addr[35504]= 1027042599;
assign addr[35505]= 1284432584;
assign addr[35506]= 1515793473;
assign addr[35507]= 1716436725;
assign addr[35508]= 1882296293;
assign addr[35509]= 2010011024;
assign addr[35510]= 2096992772;
assign addr[35511]= 2141478848;
assign addr[35512]= 2142567738;
assign addr[35513]= 2100237377;
assign addr[35514]= 2015345591;
assign addr[35515]= 1889612716;
assign addr[35516]= 1725586737;
assign addr[35517]= 1526591649;
assign addr[35518]= 1296660098;
assign addr[35519]= 1040451659;
assign addr[35520]= 763158411;
assign addr[35521]= 470399716;
assign addr[35522]= 168108346;
assign addr[35523]= -137589750;
assign addr[35524]= -440499581;
assign addr[35525]= -734482665;
assign addr[35526]= -1013581418;
assign addr[35527]= -1272139887;
assign addr[35528]= -1504918373;
assign addr[35529]= -1707199606;
assign addr[35530]= -1874884346;
assign addr[35531]= -2004574453;
assign addr[35532]= -2093641749;
assign addr[35533]= -2140281282;
assign addr[35534]= -2143547897;
assign addr[35535]= -2103375398;
assign addr[35536]= -2020577882;
assign addr[35537]= -1896833245;
assign addr[35538]= -1734649179;
assign addr[35539]= -1537312353;
assign addr[35540]= -1308821808;
assign addr[35541]= -1053807919;
assign addr[35542]= -777438554;
assign addr[35543]= -485314355;
assign addr[35544]= -183355234;
assign addr[35545]= 122319591;
assign addr[35546]= 425515602;
assign addr[35547]= 720088517;
assign addr[35548]= 1000068799;
assign addr[35549]= 1259782632;
assign addr[35550]= 1493966902;
assign addr[35551]= 1697875851;
assign addr[35552]= 1867377253;
assign addr[35553]= 1999036154;
assign addr[35554]= 2090184478;
assign addr[35555]= 2138975100;
assign addr[35556]= 2144419275;
assign addr[35557]= 2106406677;
assign addr[35558]= 2025707632;
assign addr[35559]= 1903957513;
assign addr[35560]= 1743623590;
assign addr[35561]= 1547955041;
assign addr[35562]= 1320917099;
assign addr[35563]= 1067110699;
assign addr[35564]= 791679244;
assign addr[35565]= 500204365;
assign addr[35566]= 198592817;
assign addr[35567]= -107043224;
assign addr[35568]= -410510029;
assign addr[35569]= -705657826;
assign addr[35570]= -986505429;
assign addr[35571]= -1247361445;
assign addr[35572]= -1482939614;
assign addr[35573]= -1688465931;
assign addr[35574]= -1859775393;
assign addr[35575]= -1993396407;
assign addr[35576]= -2086621133;
assign addr[35577]= -2137560369;
assign addr[35578]= -2145181827;
assign addr[35579]= -2109331059;
assign addr[35580]= -2030734582;
assign addr[35581]= -1910985158;
assign addr[35582]= -1752509516;
assign addr[35583]= -1558519173;
assign addr[35584]= -1332945355;
assign addr[35585]= -1080359326;
assign addr[35586]= -805879757;
assign addr[35587]= -515068990;
assign addr[35588]= -213820322;
assign addr[35589]= 91761426;
assign addr[35590]= 395483624;
assign addr[35591]= 691191324;
assign addr[35592]= 972891995;
assign addr[35593]= 1234876957;
assign addr[35594]= 1471837070;
assign addr[35595]= 1678970324;
assign addr[35596]= 1852079154;
assign addr[35597]= 1987655498;
assign addr[35598]= 2082951896;
assign addr[35599]= 2136037160;
assign addr[35600]= 2145835515;
assign addr[35601]= 2112148396;
assign addr[35602]= 2035658475;
assign addr[35603]= 1917915825;
assign addr[35604]= 1761306505;
assign addr[35605]= 1569004214;
assign addr[35606]= 1344905966;
assign addr[35607]= 1093553126;
assign addr[35608]= 820039373;
assign addr[35609]= 529907477;
assign addr[35610]= 229036977;
assign addr[35611]= -76474970;
assign addr[35612]= -380437148;
assign addr[35613]= -676689746;
assign addr[35614]= -959229189;
assign addr[35615]= -1222329801;
assign addr[35616]= -1460659832;
assign addr[35617]= -1669389513;
assign addr[35618]= -1844288924;
assign addr[35619]= -1981813720;
assign addr[35620]= -2079176953;
assign addr[35621]= -2134405552;
assign addr[35622]= -2146380306;
assign addr[35623]= -2114858546;
assign addr[35624]= -2040479063;
assign addr[35625]= -1924749160;
assign addr[35626]= -1770014111;
assign addr[35627]= -1579409630;
assign addr[35628]= -1356798326;
assign addr[35629]= -1106691431;
assign addr[35630]= -834157373;
assign addr[35631]= -544719071;
assign addr[35632]= -244242007;
assign addr[35633]= 61184634;
assign addr[35634]= 365371365;
assign addr[35635]= 662153826;
assign addr[35636]= 945517704;
assign addr[35637]= 1209720613;
assign addr[35638]= 1449408469;
assign addr[35639]= 1659723983;
assign addr[35640]= 1836405100;
assign addr[35641]= 1975871368;
assign addr[35642]= 2075296495;
assign addr[35643]= 2132665626;
assign addr[35644]= 2146816171;
assign addr[35645]= 2117461370;
assign addr[35646]= 2045196100;
assign addr[35647]= 1931484818;
assign addr[35648]= 1778631892;
assign addr[35649]= 1589734894;
assign addr[35650]= 1368621831;
assign addr[35651]= 1119773573;
assign addr[35652]= 848233042;
assign addr[35653]= 559503022;
assign addr[35654]= 259434643;
assign addr[35655]= -45891193;
assign addr[35656]= -350287041;
assign addr[35657]= -647584304;
assign addr[35658]= -931758235;
assign addr[35659]= -1197050035;
assign addr[35660]= -1438083551;
assign addr[35661]= -1649974225;
assign addr[35662]= -1828428082;
assign addr[35663]= -1969828744;
assign addr[35664]= -2071310720;
assign addr[35665]= -2130817471;
assign addr[35666]= -2147143090;
assign addr[35667]= -2119956737;
assign addr[35668]= -2049809346;
assign addr[35669]= -1938122457;
assign addr[35670]= -1787159411;
assign addr[35671]= -1599979481;
assign addr[35672]= -1380375881;
assign addr[35673]= -1132798888;
assign addr[35674]= -862265664;
assign addr[35675]= -574258580;
assign addr[35676]= -274614114;
assign addr[35677]= 30595422;
assign addr[35678]= 335184940;
assign addr[35679]= 632981917;
assign addr[35680]= 917951481;
assign addr[35681]= 1184318708;
assign addr[35682]= 1426685652;
assign addr[35683]= 1640140734;
assign addr[35684]= 1820358275;
assign addr[35685]= 1963686155;
assign addr[35686]= 2067219829;
assign addr[35687]= 2128861181;
assign addr[35688]= 2147361045;
assign addr[35689]= 2122344521;
assign addr[35690]= 2054318569;
assign addr[35691]= 1944661739;
assign addr[35692]= 1795596234;
assign addr[35693]= 1610142873;
assign addr[35694]= 1392059879;
assign addr[35695]= 1145766716;
assign addr[35696]= 876254528;
assign addr[35697]= 588984994;
assign addr[35698]= 289779648;
assign addr[35699]= -15298099;
assign addr[35700]= -320065829;
assign addr[35701]= -618347408;
assign addr[35702]= -904098143;
assign addr[35703]= -1171527280;
assign addr[35704]= -1415215352;
assign addr[35705]= -1630224009;
assign addr[35706]= -1812196087;
assign addr[35707]= -1957443913;
assign addr[35708]= -2063024031;
assign addr[35709]= -2126796855;
assign addr[35710]= -2147470025;
assign addr[35711]= -2124624598;
assign addr[35712]= -2058723538;
assign addr[35713]= -1951102334;
assign addr[35714]= -1803941934;
assign addr[35715]= -1620224553;
assign addr[35716]= -1403673233;
assign addr[35717]= -1158676398;
assign addr[35718]= -890198924;
assign addr[35719]= -603681519;
assign addr[35720]= -304930476;
assign addr[35721]= 0;
assign addr[35722]= 304930476;
assign addr[35723]= 603681519;
assign addr[35724]= 890198924;
assign addr[35725]= 1158676398;
assign addr[35726]= 1403673233;
assign addr[35727]= 1620224553;
assign addr[35728]= 1803941934;
assign addr[35729]= 1951102334;
assign addr[35730]= 2058723538;
assign addr[35731]= 2124624598;
assign addr[35732]= 2147470025;
assign addr[35733]= 2126796855;
assign addr[35734]= 2063024031;
assign addr[35735]= 1957443913;
assign addr[35736]= 1812196087;
assign addr[35737]= 1630224009;
assign addr[35738]= 1415215352;
assign addr[35739]= 1171527280;
assign addr[35740]= 904098143;
assign addr[35741]= 618347408;
assign addr[35742]= 320065829;
assign addr[35743]= 15298099;
assign addr[35744]= -289779648;
assign addr[35745]= -588984994;
assign addr[35746]= -876254528;
assign addr[35747]= -1145766716;
assign addr[35748]= -1392059879;
assign addr[35749]= -1610142873;
assign addr[35750]= -1795596234;
assign addr[35751]= -1944661739;
assign addr[35752]= -2054318569;
assign addr[35753]= -2122344521;
assign addr[35754]= -2147361045;
assign addr[35755]= -2128861181;
assign addr[35756]= -2067219829;
assign addr[35757]= -1963686155;
assign addr[35758]= -1820358275;
assign addr[35759]= -1640140734;
assign addr[35760]= -1426685652;
assign addr[35761]= -1184318708;
assign addr[35762]= -917951481;
assign addr[35763]= -632981917;
assign addr[35764]= -335184940;
assign addr[35765]= -30595422;
assign addr[35766]= 274614114;
assign addr[35767]= 574258580;
assign addr[35768]= 862265664;
assign addr[35769]= 1132798888;
assign addr[35770]= 1380375881;
assign addr[35771]= 1599979481;
assign addr[35772]= 1787159411;
assign addr[35773]= 1938122457;
assign addr[35774]= 2049809346;
assign addr[35775]= 2119956737;
assign addr[35776]= 2147143090;
assign addr[35777]= 2130817471;
assign addr[35778]= 2071310720;
assign addr[35779]= 1969828744;
assign addr[35780]= 1828428082;
assign addr[35781]= 1649974225;
assign addr[35782]= 1438083551;
assign addr[35783]= 1197050035;
assign addr[35784]= 931758235;
assign addr[35785]= 647584304;
assign addr[35786]= 350287041;
assign addr[35787]= 45891193;
assign addr[35788]= -259434643;
assign addr[35789]= -559503022;
assign addr[35790]= -848233042;
assign addr[35791]= -1119773573;
assign addr[35792]= -1368621831;
assign addr[35793]= -1589734894;
assign addr[35794]= -1778631892;
assign addr[35795]= -1931484818;
assign addr[35796]= -2045196100;
assign addr[35797]= -2117461370;
assign addr[35798]= -2146816171;
assign addr[35799]= -2132665626;
assign addr[35800]= -2075296495;
assign addr[35801]= -1975871368;
assign addr[35802]= -1836405100;
assign addr[35803]= -1659723983;
assign addr[35804]= -1449408469;
assign addr[35805]= -1209720613;
assign addr[35806]= -945517704;
assign addr[35807]= -662153826;
assign addr[35808]= -365371365;
assign addr[35809]= -61184634;
assign addr[35810]= 244242007;
assign addr[35811]= 544719071;
assign addr[35812]= 834157373;
assign addr[35813]= 1106691431;
assign addr[35814]= 1356798326;
assign addr[35815]= 1579409630;
assign addr[35816]= 1770014111;
assign addr[35817]= 1924749160;
assign addr[35818]= 2040479063;
assign addr[35819]= 2114858546;
assign addr[35820]= 2146380306;
assign addr[35821]= 2134405552;
assign addr[35822]= 2079176953;
assign addr[35823]= 1981813720;
assign addr[35824]= 1844288924;
assign addr[35825]= 1669389513;
assign addr[35826]= 1460659832;
assign addr[35827]= 1222329801;
assign addr[35828]= 959229189;
assign addr[35829]= 676689746;
assign addr[35830]= 380437148;
assign addr[35831]= 76474970;
assign addr[35832]= -229036977;
assign addr[35833]= -529907477;
assign addr[35834]= -820039373;
assign addr[35835]= -1093553126;
assign addr[35836]= -1344905966;
assign addr[35837]= -1569004214;
assign addr[35838]= -1761306505;
assign addr[35839]= -1917915825;
assign addr[35840]= -2035658475;
assign addr[35841]= -2112148396;
assign addr[35842]= -2145835515;
assign addr[35843]= -2136037160;
assign addr[35844]= -2082951896;
assign addr[35845]= -1987655498;
assign addr[35846]= -1852079154;
assign addr[35847]= -1678970324;
assign addr[35848]= -1471837070;
assign addr[35849]= -1234876957;
assign addr[35850]= -972891995;
assign addr[35851]= -691191324;
assign addr[35852]= -395483624;
assign addr[35853]= -91761426;
assign addr[35854]= 213820322;
assign addr[35855]= 515068990;
assign addr[35856]= 805879757;
assign addr[35857]= 1080359326;
assign addr[35858]= 1332945355;
assign addr[35859]= 1558519173;
assign addr[35860]= 1752509516;
assign addr[35861]= 1910985158;
assign addr[35862]= 2030734582;
assign addr[35863]= 2109331059;
assign addr[35864]= 2145181827;
assign addr[35865]= 2137560369;
assign addr[35866]= 2086621133;
assign addr[35867]= 1993396407;
assign addr[35868]= 1859775393;
assign addr[35869]= 1688465931;
assign addr[35870]= 1482939614;
assign addr[35871]= 1247361445;
assign addr[35872]= 986505429;
assign addr[35873]= 705657826;
assign addr[35874]= 410510029;
assign addr[35875]= 107043224;
assign addr[35876]= -198592817;
assign addr[35877]= -500204365;
assign addr[35878]= -791679244;
assign addr[35879]= -1067110699;
assign addr[35880]= -1320917099;
assign addr[35881]= -1547955041;
assign addr[35882]= -1743623590;
assign addr[35883]= -1903957513;
assign addr[35884]= -2025707632;
assign addr[35885]= -2106406677;
assign addr[35886]= -2144419275;
assign addr[35887]= -2138975100;
assign addr[35888]= -2090184478;
assign addr[35889]= -1999036154;
assign addr[35890]= -1867377253;
assign addr[35891]= -1697875851;
assign addr[35892]= -1493966902;
assign addr[35893]= -1259782632;
assign addr[35894]= -1000068799;
assign addr[35895]= -720088517;
assign addr[35896]= -425515602;
assign addr[35897]= -122319591;
assign addr[35898]= 183355234;
assign addr[35899]= 485314355;
assign addr[35900]= 777438554;
assign addr[35901]= 1053807919;
assign addr[35902]= 1308821808;
assign addr[35903]= 1537312353;
assign addr[35904]= 1734649179;
assign addr[35905]= 1896833245;
assign addr[35906]= 2020577882;
assign addr[35907]= 2103375398;
assign addr[35908]= 2143547897;
assign addr[35909]= 2140281282;
assign addr[35910]= 2093641749;
assign addr[35911]= 2004574453;
assign addr[35912]= 1874884346;
assign addr[35913]= 1707199606;
assign addr[35914]= 1504918373;
assign addr[35915]= 1272139887;
assign addr[35916]= 1013581418;
assign addr[35917]= 734482665;
assign addr[35918]= 440499581;
assign addr[35919]= 137589750;
assign addr[35920]= -168108346;
assign addr[35921]= -470399716;
assign addr[35922]= -763158411;
assign addr[35923]= -1040451659;
assign addr[35924]= -1296660098;
assign addr[35925]= -1526591649;
assign addr[35926]= -1725586737;
assign addr[35927]= -1889612716;
assign addr[35928]= -2015345591;
assign addr[35929]= -2100237377;
assign addr[35930]= -2142567738;
assign addr[35931]= -2141478848;
assign addr[35932]= -2096992772;
assign addr[35933]= -2010011024;
assign addr[35934]= -1882296293;
assign addr[35935]= -1716436725;
assign addr[35936]= -1515793473;
assign addr[35937]= -1284432584;
assign addr[35938]= -1027042599;
assign addr[35939]= -748839539;
assign addr[35940]= -455461206;
assign addr[35941]= -152852926;
assign addr[35942]= 152852926;
assign addr[35943]= 455461206;
assign addr[35944]= 748839539;
assign addr[35945]= 1027042599;
assign addr[35946]= 1284432584;
assign addr[35947]= 1515793473;
assign addr[35948]= 1716436725;
assign addr[35949]= 1882296293;
assign addr[35950]= 2010011024;
assign addr[35951]= 2096992772;
assign addr[35952]= 2141478848;
assign addr[35953]= 2142567738;
assign addr[35954]= 2100237377;
assign addr[35955]= 2015345591;
assign addr[35956]= 1889612716;
assign addr[35957]= 1725586737;
assign addr[35958]= 1526591649;
assign addr[35959]= 1296660098;
assign addr[35960]= 1040451659;
assign addr[35961]= 763158411;
assign addr[35962]= 470399716;
assign addr[35963]= 168108346;
assign addr[35964]= -137589750;
assign addr[35965]= -440499581;
assign addr[35966]= -734482665;
assign addr[35967]= -1013581418;
assign addr[35968]= -1272139887;
assign addr[35969]= -1504918373;
assign addr[35970]= -1707199606;
assign addr[35971]= -1874884346;
assign addr[35972]= -2004574453;
assign addr[35973]= -2093641749;
assign addr[35974]= -2140281282;
assign addr[35975]= -2143547897;
assign addr[35976]= -2103375398;
assign addr[35977]= -2020577882;
assign addr[35978]= -1896833245;
assign addr[35979]= -1734649179;
assign addr[35980]= -1537312353;
assign addr[35981]= -1308821808;
assign addr[35982]= -1053807919;
assign addr[35983]= -777438554;
assign addr[35984]= -485314355;
assign addr[35985]= -183355234;
assign addr[35986]= 122319591;
assign addr[35987]= 425515602;
assign addr[35988]= 720088517;
assign addr[35989]= 1000068799;
assign addr[35990]= 1259782632;
assign addr[35991]= 1493966902;
assign addr[35992]= 1697875851;
assign addr[35993]= 1867377253;
assign addr[35994]= 1999036154;
assign addr[35995]= 2090184478;
assign addr[35996]= 2138975100;
assign addr[35997]= 2144419275;
assign addr[35998]= 2106406677;
assign addr[35999]= 2025707632;
assign addr[36000]= 1903957513;
assign addr[36001]= 1743623590;
assign addr[36002]= 1547955041;
assign addr[36003]= 1320917099;
assign addr[36004]= 1067110699;
assign addr[36005]= 791679244;
assign addr[36006]= 500204365;
assign addr[36007]= 198592817;
assign addr[36008]= -107043224;
assign addr[36009]= -410510029;
assign addr[36010]= -705657826;
assign addr[36011]= -986505429;
assign addr[36012]= -1247361445;
assign addr[36013]= -1482939614;
assign addr[36014]= -1688465931;
assign addr[36015]= -1859775393;
assign addr[36016]= -1993396407;
assign addr[36017]= -2086621133;
assign addr[36018]= -2137560369;
assign addr[36019]= -2145181827;
assign addr[36020]= -2109331059;
assign addr[36021]= -2030734582;
assign addr[36022]= -1910985158;
assign addr[36023]= -1752509516;
assign addr[36024]= -1558519173;
assign addr[36025]= -1332945355;
assign addr[36026]= -1080359326;
assign addr[36027]= -805879757;
assign addr[36028]= -515068990;
assign addr[36029]= -213820322;
assign addr[36030]= 91761426;
assign addr[36031]= 395483624;
assign addr[36032]= 691191324;
assign addr[36033]= 972891995;
assign addr[36034]= 1234876957;
assign addr[36035]= 1471837070;
assign addr[36036]= 1678970324;
assign addr[36037]= 1852079154;
assign addr[36038]= 1987655498;
assign addr[36039]= 2082951896;
assign addr[36040]= 2136037160;
assign addr[36041]= 2145835515;
assign addr[36042]= 2112148396;
assign addr[36043]= 2035658475;
assign addr[36044]= 1917915825;
assign addr[36045]= 1761306505;
assign addr[36046]= 1569004214;
assign addr[36047]= 1344905966;
assign addr[36048]= 1093553126;
assign addr[36049]= 820039373;
assign addr[36050]= 529907477;
assign addr[36051]= 229036977;
assign addr[36052]= -76474970;
assign addr[36053]= -380437148;
assign addr[36054]= -676689746;
assign addr[36055]= -959229189;
assign addr[36056]= -1222329801;
assign addr[36057]= -1460659832;
assign addr[36058]= -1669389513;
assign addr[36059]= -1844288924;
assign addr[36060]= -1981813720;
assign addr[36061]= -2079176953;
assign addr[36062]= -2134405552;
assign addr[36063]= -2146380306;
assign addr[36064]= -2114858546;
assign addr[36065]= -2040479063;
assign addr[36066]= -1924749160;
assign addr[36067]= -1770014111;
assign addr[36068]= -1579409630;
assign addr[36069]= -1356798326;
assign addr[36070]= -1106691431;
assign addr[36071]= -834157373;
assign addr[36072]= -544719071;
assign addr[36073]= -244242007;
assign addr[36074]= 61184634;
assign addr[36075]= 365371365;
assign addr[36076]= 662153826;
assign addr[36077]= 945517704;
assign addr[36078]= 1209720613;
assign addr[36079]= 1449408469;
assign addr[36080]= 1659723983;
assign addr[36081]= 1836405100;
assign addr[36082]= 1975871368;
assign addr[36083]= 2075296495;
assign addr[36084]= 2132665626;
assign addr[36085]= 2146816171;
assign addr[36086]= 2117461370;
assign addr[36087]= 2045196100;
assign addr[36088]= 1931484818;
assign addr[36089]= 1778631892;
assign addr[36090]= 1589734894;
assign addr[36091]= 1368621831;
assign addr[36092]= 1119773573;
assign addr[36093]= 848233042;
assign addr[36094]= 559503022;
assign addr[36095]= 259434643;
assign addr[36096]= -45891193;
assign addr[36097]= -350287041;
assign addr[36098]= -647584304;
assign addr[36099]= -931758235;
assign addr[36100]= -1197050035;
assign addr[36101]= -1438083551;
assign addr[36102]= -1649974225;
assign addr[36103]= -1828428082;
assign addr[36104]= -1969828744;
assign addr[36105]= -2071310720;
assign addr[36106]= -2130817471;
assign addr[36107]= -2147143090;
assign addr[36108]= -2119956737;
assign addr[36109]= -2049809346;
assign addr[36110]= -1938122457;
assign addr[36111]= -1787159411;
assign addr[36112]= -1599979481;
assign addr[36113]= -1380375881;
assign addr[36114]= -1132798888;
assign addr[36115]= -862265664;
assign addr[36116]= -574258580;
assign addr[36117]= -274614114;
assign addr[36118]= 30595422;
assign addr[36119]= 335184940;
assign addr[36120]= 632981917;
assign addr[36121]= 917951481;
assign addr[36122]= 1184318708;
assign addr[36123]= 1426685652;
assign addr[36124]= 1640140734;
assign addr[36125]= 1820358275;
assign addr[36126]= 1963686155;
assign addr[36127]= 2067219829;
assign addr[36128]= 2128861181;
assign addr[36129]= 2147361045;
assign addr[36130]= 2122344521;
assign addr[36131]= 2054318569;
assign addr[36132]= 1944661739;
assign addr[36133]= 1795596234;
assign addr[36134]= 1610142873;
assign addr[36135]= 1392059879;
assign addr[36136]= 1145766716;
assign addr[36137]= 876254528;
assign addr[36138]= 588984994;
assign addr[36139]= 289779648;
assign addr[36140]= -15298099;
assign addr[36141]= -320065829;
assign addr[36142]= -618347408;
assign addr[36143]= -904098143;
assign addr[36144]= -1171527280;
assign addr[36145]= -1415215352;
assign addr[36146]= -1630224009;
assign addr[36147]= -1812196087;
assign addr[36148]= -1957443913;
assign addr[36149]= -2063024031;
assign addr[36150]= -2126796855;
assign addr[36151]= -2147470025;
assign addr[36152]= -2124624598;
assign addr[36153]= -2058723538;
assign addr[36154]= -1951102334;
assign addr[36155]= -1803941934;
assign addr[36156]= -1620224553;
assign addr[36157]= -1403673233;
assign addr[36158]= -1158676398;
assign addr[36159]= -890198924;
assign addr[36160]= -603681519;
assign addr[36161]= -304930476;
assign addr[36162]= 0;
assign addr[36163]= 304930476;
assign addr[36164]= 603681519;
assign addr[36165]= 890198924;
assign addr[36166]= 1158676398;
assign addr[36167]= 1403673233;
assign addr[36168]= 1620224553;
assign addr[36169]= 1803941934;
assign addr[36170]= 1951102334;
assign addr[36171]= 2058723538;
assign addr[36172]= 2124624598;
assign addr[36173]= 2147470025;
assign addr[36174]= 2126796855;
assign addr[36175]= 2063024031;
assign addr[36176]= 1957443913;
assign addr[36177]= 1812196087;
assign addr[36178]= 1630224009;
assign addr[36179]= 1415215352;
assign addr[36180]= 1171527280;
assign addr[36181]= 904098143;
assign addr[36182]= 618347408;
assign addr[36183]= 320065829;
assign addr[36184]= 15298099;
assign addr[36185]= -289779648;
assign addr[36186]= -588984994;
assign addr[36187]= -876254528;
assign addr[36188]= -1145766716;
assign addr[36189]= -1392059879;
assign addr[36190]= -1610142873;
assign addr[36191]= -1795596234;
assign addr[36192]= -1944661739;
assign addr[36193]= -2054318569;
assign addr[36194]= -2122344521;
assign addr[36195]= -2147361045;
assign addr[36196]= -2128861181;
assign addr[36197]= -2067219829;
assign addr[36198]= -1963686155;
assign addr[36199]= -1820358275;
assign addr[36200]= -1640140734;
assign addr[36201]= -1426685652;
assign addr[36202]= -1184318708;
assign addr[36203]= -917951481;
assign addr[36204]= -632981917;
assign addr[36205]= -335184940;
assign addr[36206]= -30595422;
assign addr[36207]= 274614114;
assign addr[36208]= 574258580;
assign addr[36209]= 862265664;
assign addr[36210]= 1132798888;
assign addr[36211]= 1380375881;
assign addr[36212]= 1599979481;
assign addr[36213]= 1787159411;
assign addr[36214]= 1938122457;
assign addr[36215]= 2049809346;
assign addr[36216]= 2119956737;
assign addr[36217]= 2147143090;
assign addr[36218]= 2130817471;
assign addr[36219]= 2071310720;
assign addr[36220]= 1969828744;
assign addr[36221]= 1828428082;
assign addr[36222]= 1649974225;
assign addr[36223]= 1438083551;
assign addr[36224]= 1197050035;
assign addr[36225]= 931758235;
assign addr[36226]= 647584304;
assign addr[36227]= 350287041;
assign addr[36228]= 45891193;
assign addr[36229]= -259434643;
assign addr[36230]= -559503022;
assign addr[36231]= -848233042;
assign addr[36232]= -1119773573;
assign addr[36233]= -1368621831;
assign addr[36234]= -1589734894;
assign addr[36235]= -1778631892;
assign addr[36236]= -1931484818;
assign addr[36237]= -2045196100;
assign addr[36238]= -2117461370;
assign addr[36239]= -2146816171;
assign addr[36240]= -2132665626;
assign addr[36241]= -2075296495;
assign addr[36242]= -1975871368;
assign addr[36243]= -1836405100;
assign addr[36244]= -1659723983;
assign addr[36245]= -1449408469;
assign addr[36246]= -1209720613;
assign addr[36247]= -945517704;
assign addr[36248]= -662153826;
assign addr[36249]= -365371365;
assign addr[36250]= -61184634;
assign addr[36251]= 244242007;
assign addr[36252]= 544719071;
assign addr[36253]= 834157373;
assign addr[36254]= 1106691431;
assign addr[36255]= 1356798326;
assign addr[36256]= 1579409630;
assign addr[36257]= 1770014111;
assign addr[36258]= 1924749160;
assign addr[36259]= 2040479063;
assign addr[36260]= 2114858546;
assign addr[36261]= 2146380306;
assign addr[36262]= 2134405552;
assign addr[36263]= 2079176953;
assign addr[36264]= 1981813720;
assign addr[36265]= 1844288924;
assign addr[36266]= 1669389513;
assign addr[36267]= 1460659832;
assign addr[36268]= 1222329801;
assign addr[36269]= 959229189;
assign addr[36270]= 676689746;
assign addr[36271]= 380437148;
assign addr[36272]= 76474970;
assign addr[36273]= -229036977;
assign addr[36274]= -529907477;
assign addr[36275]= -820039373;
assign addr[36276]= -1093553126;
assign addr[36277]= -1344905966;
assign addr[36278]= -1569004214;
assign addr[36279]= -1761306505;
assign addr[36280]= -1917915825;
assign addr[36281]= -2035658475;
assign addr[36282]= -2112148396;
assign addr[36283]= -2145835515;
assign addr[36284]= -2136037160;
assign addr[36285]= -2082951896;
assign addr[36286]= -1987655498;
assign addr[36287]= -1852079154;
assign addr[36288]= -1678970324;
assign addr[36289]= -1471837070;
assign addr[36290]= -1234876957;
assign addr[36291]= -972891995;
assign addr[36292]= -691191324;
assign addr[36293]= -395483624;
assign addr[36294]= -91761426;
assign addr[36295]= 213820322;
assign addr[36296]= 515068990;
assign addr[36297]= 805879757;
assign addr[36298]= 1080359326;
assign addr[36299]= 1332945355;
assign addr[36300]= 1558519173;
assign addr[36301]= 1752509516;
assign addr[36302]= 1910985158;
assign addr[36303]= 2030734582;
assign addr[36304]= 2109331059;
assign addr[36305]= 2145181827;
assign addr[36306]= 2137560369;
assign addr[36307]= 2086621133;
assign addr[36308]= 1993396407;
assign addr[36309]= 1859775393;
assign addr[36310]= 1688465931;
assign addr[36311]= 1482939614;
assign addr[36312]= 1247361445;
assign addr[36313]= 986505429;
assign addr[36314]= 705657826;
assign addr[36315]= 410510029;
assign addr[36316]= 107043224;
assign addr[36317]= -198592817;
assign addr[36318]= -500204365;
assign addr[36319]= -791679244;
assign addr[36320]= -1067110699;
assign addr[36321]= -1320917099;
assign addr[36322]= -1547955041;
assign addr[36323]= -1743623590;
assign addr[36324]= -1903957513;
assign addr[36325]= -2025707632;
assign addr[36326]= -2106406677;
assign addr[36327]= -2144419275;
assign addr[36328]= -2138975100;
assign addr[36329]= -2090184478;
assign addr[36330]= -1999036154;
assign addr[36331]= -1867377253;
assign addr[36332]= -1697875851;
assign addr[36333]= -1493966902;
assign addr[36334]= -1259782632;
assign addr[36335]= -1000068799;
assign addr[36336]= -720088517;
assign addr[36337]= -425515602;
assign addr[36338]= -122319591;
assign addr[36339]= 183355234;
assign addr[36340]= 485314355;
assign addr[36341]= 777438554;
assign addr[36342]= 1053807919;
assign addr[36343]= 1308821808;
assign addr[36344]= 1537312353;
assign addr[36345]= 1734649179;
assign addr[36346]= 1896833245;
assign addr[36347]= 2020577882;
assign addr[36348]= 2103375398;
assign addr[36349]= 2143547897;
assign addr[36350]= 2140281282;
assign addr[36351]= 2093641749;
assign addr[36352]= 2004574453;
assign addr[36353]= 1874884346;
assign addr[36354]= 1707199606;
assign addr[36355]= 1504918373;
assign addr[36356]= 1272139887;
assign addr[36357]= 1013581418;
assign addr[36358]= 734482665;
assign addr[36359]= 440499581;
assign addr[36360]= 137589750;
assign addr[36361]= -168108346;
assign addr[36362]= -470399716;
assign addr[36363]= -763158411;
assign addr[36364]= -1040451659;
assign addr[36365]= -1296660098;
assign addr[36366]= -1526591649;
assign addr[36367]= -1725586737;
assign addr[36368]= -1889612716;
assign addr[36369]= -2015345591;
assign addr[36370]= -2100237377;
assign addr[36371]= -2142567738;
assign addr[36372]= -2141478848;
assign addr[36373]= -2096992772;
assign addr[36374]= -2010011024;
assign addr[36375]= -1882296293;
assign addr[36376]= -1716436725;
assign addr[36377]= -1515793473;
assign addr[36378]= -1284432584;
assign addr[36379]= -1027042599;
assign addr[36380]= -748839539;
assign addr[36381]= -455461206;
assign addr[36382]= -152852926;
assign addr[36383]= 152852926;
assign addr[36384]= 455461206;
assign addr[36385]= 748839539;
assign addr[36386]= 1027042599;
assign addr[36387]= 1284432584;
assign addr[36388]= 1515793473;
assign addr[36389]= 1716436725;
assign addr[36390]= 1882296293;
assign addr[36391]= 2010011024;
assign addr[36392]= 2096992772;
assign addr[36393]= 2141478848;
assign addr[36394]= 2142567738;
assign addr[36395]= 2100237377;
assign addr[36396]= 2015345591;
assign addr[36397]= 1889612716;
assign addr[36398]= 1725586737;
assign addr[36399]= 1526591649;
assign addr[36400]= 1296660098;
assign addr[36401]= 1040451659;
assign addr[36402]= 763158411;
assign addr[36403]= 470399716;
assign addr[36404]= 168108346;
assign addr[36405]= -137589750;
assign addr[36406]= -440499581;
assign addr[36407]= -734482665;
assign addr[36408]= -1013581418;
assign addr[36409]= -1272139887;
assign addr[36410]= -1504918373;
assign addr[36411]= -1707199606;
assign addr[36412]= -1874884346;
assign addr[36413]= -2004574453;
assign addr[36414]= -2093641749;
assign addr[36415]= -2140281282;
assign addr[36416]= -2143547897;
assign addr[36417]= -2103375398;
assign addr[36418]= -2020577882;
assign addr[36419]= -1896833245;
assign addr[36420]= -1734649179;
assign addr[36421]= -1537312353;
assign addr[36422]= -1308821808;
assign addr[36423]= -1053807919;
assign addr[36424]= -777438554;
assign addr[36425]= -485314355;
assign addr[36426]= -183355234;
assign addr[36427]= 122319591;
assign addr[36428]= 425515602;
assign addr[36429]= 720088517;
assign addr[36430]= 1000068799;
assign addr[36431]= 1259782632;
assign addr[36432]= 1493966902;
assign addr[36433]= 1697875851;
assign addr[36434]= 1867377253;
assign addr[36435]= 1999036154;
assign addr[36436]= 2090184478;
assign addr[36437]= 2138975100;
assign addr[36438]= 2144419275;
assign addr[36439]= 2106406677;
assign addr[36440]= 2025707632;
assign addr[36441]= 1903957513;
assign addr[36442]= 1743623590;
assign addr[36443]= 1547955041;
assign addr[36444]= 1320917099;
assign addr[36445]= 1067110699;
assign addr[36446]= 791679244;
assign addr[36447]= 500204365;
assign addr[36448]= 198592817;
assign addr[36449]= -107043224;
assign addr[36450]= -410510029;
assign addr[36451]= -705657826;
assign addr[36452]= -986505429;
assign addr[36453]= -1247361445;
assign addr[36454]= -1482939614;
assign addr[36455]= -1688465931;
assign addr[36456]= -1859775393;
assign addr[36457]= -1993396407;
assign addr[36458]= -2086621133;
assign addr[36459]= -2137560369;
assign addr[36460]= -2145181827;
assign addr[36461]= -2109331059;
assign addr[36462]= -2030734582;
assign addr[36463]= -1910985158;
assign addr[36464]= -1752509516;
assign addr[36465]= -1558519173;
assign addr[36466]= -1332945355;
assign addr[36467]= -1080359326;
assign addr[36468]= -805879757;
assign addr[36469]= -515068990;
assign addr[36470]= -213820322;
assign addr[36471]= 91761426;
assign addr[36472]= 395483624;
assign addr[36473]= 691191324;
assign addr[36474]= 972891995;
assign addr[36475]= 1234876957;
assign addr[36476]= 1471837070;
assign addr[36477]= 1678970324;
assign addr[36478]= 1852079154;
assign addr[36479]= 1987655498;
assign addr[36480]= 2082951896;
assign addr[36481]= 2136037160;
assign addr[36482]= 2145835515;
assign addr[36483]= 2112148396;
assign addr[36484]= 2035658475;
assign addr[36485]= 1917915825;
assign addr[36486]= 1761306505;
assign addr[36487]= 1569004214;
assign addr[36488]= 1344905966;
assign addr[36489]= 1093553126;
assign addr[36490]= 820039373;
assign addr[36491]= 529907477;
assign addr[36492]= 229036977;
assign addr[36493]= -76474970;
assign addr[36494]= -380437148;
assign addr[36495]= -676689746;
assign addr[36496]= -959229189;
assign addr[36497]= -1222329801;
assign addr[36498]= -1460659832;
assign addr[36499]= -1669389513;
assign addr[36500]= -1844288924;
assign addr[36501]= -1981813720;
assign addr[36502]= -2079176953;
assign addr[36503]= -2134405552;
assign addr[36504]= -2146380306;
assign addr[36505]= -2114858546;
assign addr[36506]= -2040479063;
assign addr[36507]= -1924749160;
assign addr[36508]= -1770014111;
assign addr[36509]= -1579409630;
assign addr[36510]= -1356798326;
assign addr[36511]= -1106691431;
assign addr[36512]= -834157373;
assign addr[36513]= -544719071;
assign addr[36514]= -244242007;
assign addr[36515]= 61184634;
assign addr[36516]= 365371365;
assign addr[36517]= 662153826;
assign addr[36518]= 945517704;
assign addr[36519]= 1209720613;
assign addr[36520]= 1449408469;
assign addr[36521]= 1659723983;
assign addr[36522]= 1836405100;
assign addr[36523]= 1975871368;
assign addr[36524]= 2075296495;
assign addr[36525]= 2132665626;
assign addr[36526]= 2146816171;
assign addr[36527]= 2117461370;
assign addr[36528]= 2045196100;
assign addr[36529]= 1931484818;
assign addr[36530]= 1778631892;
assign addr[36531]= 1589734894;
assign addr[36532]= 1368621831;
assign addr[36533]= 1119773573;
assign addr[36534]= 848233042;
assign addr[36535]= 559503022;
assign addr[36536]= 259434643;
assign addr[36537]= -45891193;
assign addr[36538]= -350287041;
assign addr[36539]= -647584304;
assign addr[36540]= -931758235;
assign addr[36541]= -1197050035;
assign addr[36542]= -1438083551;
assign addr[36543]= -1649974225;
assign addr[36544]= -1828428082;
assign addr[36545]= -1969828744;
assign addr[36546]= -2071310720;
assign addr[36547]= -2130817471;
assign addr[36548]= -2147143090;
assign addr[36549]= -2119956737;
assign addr[36550]= -2049809346;
assign addr[36551]= -1938122457;
assign addr[36552]= -1787159411;
assign addr[36553]= -1599979481;
assign addr[36554]= -1380375881;
assign addr[36555]= -1132798888;
assign addr[36556]= -862265664;
assign addr[36557]= -574258580;
assign addr[36558]= -274614114;
assign addr[36559]= 30595422;
assign addr[36560]= 335184940;
assign addr[36561]= 632981917;
assign addr[36562]= 917951481;
assign addr[36563]= 1184318708;
assign addr[36564]= 1426685652;
assign addr[36565]= 1640140734;
assign addr[36566]= 1820358275;
assign addr[36567]= 1963686155;
assign addr[36568]= 2067219829;
assign addr[36569]= 2128861181;
assign addr[36570]= 2147361045;
assign addr[36571]= 2122344521;
assign addr[36572]= 2054318569;
assign addr[36573]= 1944661739;
assign addr[36574]= 1795596234;
assign addr[36575]= 1610142873;
assign addr[36576]= 1392059879;
assign addr[36577]= 1145766716;
assign addr[36578]= 876254528;
assign addr[36579]= 588984994;
assign addr[36580]= 289779648;
assign addr[36581]= -15298099;
assign addr[36582]= -320065829;
assign addr[36583]= -618347408;
assign addr[36584]= -904098143;
assign addr[36585]= -1171527280;
assign addr[36586]= -1415215352;
assign addr[36587]= -1630224009;
assign addr[36588]= -1812196087;
assign addr[36589]= -1957443913;
assign addr[36590]= -2063024031;
assign addr[36591]= -2126796855;
assign addr[36592]= -2147470025;
assign addr[36593]= -2124624598;
assign addr[36594]= -2058723538;
assign addr[36595]= -1951102334;
assign addr[36596]= -1803941934;
assign addr[36597]= -1620224553;
assign addr[36598]= -1403673233;
assign addr[36599]= -1158676398;
assign addr[36600]= -890198924;
assign addr[36601]= -603681519;
assign addr[36602]= -304930476;
assign addr[36603]= 0;
assign addr[36604]= 304930476;
assign addr[36605]= 603681519;
assign addr[36606]= 890198924;
assign addr[36607]= 1158676398;
assign addr[36608]= 1403673233;
assign addr[36609]= 1620224553;
assign addr[36610]= 1803941934;
assign addr[36611]= 1951102334;
assign addr[36612]= 2058723538;
assign addr[36613]= 2124624598;
assign addr[36614]= 2147470025;
assign addr[36615]= 2126796855;
assign addr[36616]= 2063024031;
assign addr[36617]= 1957443913;
assign addr[36618]= 1812196087;
assign addr[36619]= 1630224009;
assign addr[36620]= 1415215352;
assign addr[36621]= 1171527280;
assign addr[36622]= 904098143;
assign addr[36623]= 618347408;
assign addr[36624]= 320065829;
assign addr[36625]= 15298099;
assign addr[36626]= -289779648;
assign addr[36627]= -588984994;
assign addr[36628]= -876254528;
assign addr[36629]= -1145766716;
assign addr[36630]= -1392059879;
assign addr[36631]= -1610142873;
assign addr[36632]= -1795596234;
assign addr[36633]= -1944661739;
assign addr[36634]= -2054318569;
assign addr[36635]= -2122344521;
assign addr[36636]= -2147361045;
assign addr[36637]= -2128861181;
assign addr[36638]= -2067219829;
assign addr[36639]= -1963686155;
assign addr[36640]= -1820358275;
assign addr[36641]= -1640140734;
assign addr[36642]= -1426685652;
assign addr[36643]= -1184318708;
assign addr[36644]= -917951481;
assign addr[36645]= -632981917;
assign addr[36646]= -335184940;
assign addr[36647]= -30595422;
assign addr[36648]= 274614114;
assign addr[36649]= 574258580;
assign addr[36650]= 862265664;
assign addr[36651]= 1132798888;
assign addr[36652]= 1380375881;
assign addr[36653]= 1599979481;
assign addr[36654]= 1787159411;
assign addr[36655]= 1938122457;
assign addr[36656]= 2049809346;
assign addr[36657]= 2119956737;
assign addr[36658]= 2147143090;
assign addr[36659]= 2130817471;
assign addr[36660]= 2071310720;
assign addr[36661]= 1969828744;
assign addr[36662]= 1828428082;
assign addr[36663]= 1649974225;
assign addr[36664]= 1438083551;
assign addr[36665]= 1197050035;
assign addr[36666]= 931758235;
assign addr[36667]= 647584304;
assign addr[36668]= 350287041;
assign addr[36669]= 45891193;
assign addr[36670]= -259434643;
assign addr[36671]= -559503022;
assign addr[36672]= -848233042;
assign addr[36673]= -1119773573;
assign addr[36674]= -1368621831;
assign addr[36675]= -1589734894;
assign addr[36676]= -1778631892;
assign addr[36677]= -1931484818;
assign addr[36678]= -2045196100;
assign addr[36679]= -2117461370;
assign addr[36680]= -2146816171;
assign addr[36681]= -2132665626;
assign addr[36682]= -2075296495;
assign addr[36683]= -1975871368;
assign addr[36684]= -1836405100;
assign addr[36685]= -1659723983;
assign addr[36686]= -1449408469;
assign addr[36687]= -1209720613;
assign addr[36688]= -945517704;
assign addr[36689]= -662153826;
assign addr[36690]= -365371365;
assign addr[36691]= -61184634;
assign addr[36692]= 244242007;
assign addr[36693]= 544719071;
assign addr[36694]= 834157373;
assign addr[36695]= 1106691431;
assign addr[36696]= 1356798326;
assign addr[36697]= 1579409630;
assign addr[36698]= 1770014111;
assign addr[36699]= 1924749160;
assign addr[36700]= 2040479063;
assign addr[36701]= 2114858546;
assign addr[36702]= 2146380306;
assign addr[36703]= 2134405552;
assign addr[36704]= 2079176953;
assign addr[36705]= 1981813720;
assign addr[36706]= 1844288924;
assign addr[36707]= 1669389513;
assign addr[36708]= 1460659832;
assign addr[36709]= 1222329801;
assign addr[36710]= 959229189;
assign addr[36711]= 676689746;
assign addr[36712]= 380437148;
assign addr[36713]= 76474970;
assign addr[36714]= -229036977;
assign addr[36715]= -529907477;
assign addr[36716]= -820039373;
assign addr[36717]= -1093553126;
assign addr[36718]= -1344905966;
assign addr[36719]= -1569004214;
assign addr[36720]= -1761306505;
assign addr[36721]= -1917915825;
assign addr[36722]= -2035658475;
assign addr[36723]= -2112148396;
assign addr[36724]= -2145835515;
assign addr[36725]= -2136037160;
assign addr[36726]= -2082951896;
assign addr[36727]= -1987655498;
assign addr[36728]= -1852079154;
assign addr[36729]= -1678970324;
assign addr[36730]= -1471837070;
assign addr[36731]= -1234876957;
assign addr[36732]= -972891995;
assign addr[36733]= -691191324;
assign addr[36734]= -395483624;
assign addr[36735]= -91761426;
assign addr[36736]= 213820322;
assign addr[36737]= 515068990;
assign addr[36738]= 805879757;
assign addr[36739]= 1080359326;
assign addr[36740]= 1332945355;
assign addr[36741]= 1558519173;
assign addr[36742]= 1752509516;
assign addr[36743]= 1910985158;
assign addr[36744]= 2030734582;
assign addr[36745]= 2109331059;
assign addr[36746]= 2145181827;
assign addr[36747]= 2137560369;
assign addr[36748]= 2086621133;
assign addr[36749]= 1993396407;
assign addr[36750]= 1859775393;
assign addr[36751]= 1688465931;
assign addr[36752]= 1482939614;
assign addr[36753]= 1247361445;
assign addr[36754]= 986505429;
assign addr[36755]= 705657826;
assign addr[36756]= 410510029;
assign addr[36757]= 107043224;
assign addr[36758]= -198592817;
assign addr[36759]= -500204365;
assign addr[36760]= -791679244;
assign addr[36761]= -1067110699;
assign addr[36762]= -1320917099;
assign addr[36763]= -1547955041;
assign addr[36764]= -1743623590;
assign addr[36765]= -1903957513;
assign addr[36766]= -2025707632;
assign addr[36767]= -2106406677;
assign addr[36768]= -2144419275;
assign addr[36769]= -2138975100;
assign addr[36770]= -2090184478;
assign addr[36771]= -1999036154;
assign addr[36772]= -1867377253;
assign addr[36773]= -1697875851;
assign addr[36774]= -1493966902;
assign addr[36775]= -1259782632;
assign addr[36776]= -1000068799;
assign addr[36777]= -720088517;
assign addr[36778]= -425515602;
assign addr[36779]= -122319591;
assign addr[36780]= 183355234;
assign addr[36781]= 485314355;
assign addr[36782]= 777438554;
assign addr[36783]= 1053807919;
assign addr[36784]= 1308821808;
assign addr[36785]= 1537312353;
assign addr[36786]= 1734649179;
assign addr[36787]= 1896833245;
assign addr[36788]= 2020577882;
assign addr[36789]= 2103375398;
assign addr[36790]= 2143547897;
assign addr[36791]= 2140281282;
assign addr[36792]= 2093641749;
assign addr[36793]= 2004574453;
assign addr[36794]= 1874884346;
assign addr[36795]= 1707199606;
assign addr[36796]= 1504918373;
assign addr[36797]= 1272139887;
assign addr[36798]= 1013581418;
assign addr[36799]= 734482665;
assign addr[36800]= 440499581;
assign addr[36801]= 137589750;
assign addr[36802]= -168108346;
assign addr[36803]= -470399716;
assign addr[36804]= -763158411;
assign addr[36805]= -1040451659;
assign addr[36806]= -1296660098;
assign addr[36807]= -1526591649;
assign addr[36808]= -1725586737;
assign addr[36809]= -1889612716;
assign addr[36810]= -2015345591;
assign addr[36811]= -2100237377;
assign addr[36812]= -2142567738;
assign addr[36813]= -2141478848;
assign addr[36814]= -2096992772;
assign addr[36815]= -2010011024;
assign addr[36816]= -1882296293;
assign addr[36817]= -1716436725;
assign addr[36818]= -1515793473;
assign addr[36819]= -1284432584;
assign addr[36820]= -1027042599;
assign addr[36821]= -748839539;
assign addr[36822]= -455461206;
assign addr[36823]= -152852926;
assign addr[36824]= 152852926;
assign addr[36825]= 455461206;
assign addr[36826]= 748839539;
assign addr[36827]= 1027042599;
assign addr[36828]= 1284432584;
assign addr[36829]= 1515793473;
assign addr[36830]= 1716436725;
assign addr[36831]= 1882296293;
assign addr[36832]= 2010011024;
assign addr[36833]= 2096992772;
assign addr[36834]= 2141478848;
assign addr[36835]= 2142567738;
assign addr[36836]= 2100237377;
assign addr[36837]= 2015345591;
assign addr[36838]= 1889612716;
assign addr[36839]= 1725586737;
assign addr[36840]= 1526591649;
assign addr[36841]= 1296660098;
assign addr[36842]= 1040451659;
assign addr[36843]= 763158411;
assign addr[36844]= 470399716;
assign addr[36845]= 168108346;
assign addr[36846]= -137589750;
assign addr[36847]= -440499581;
assign addr[36848]= -734482665;
assign addr[36849]= -1013581418;
assign addr[36850]= -1272139887;
assign addr[36851]= -1504918373;
assign addr[36852]= -1707199606;
assign addr[36853]= -1874884346;
assign addr[36854]= -2004574453;
assign addr[36855]= -2093641749;
assign addr[36856]= -2140281282;
assign addr[36857]= -2143547897;
assign addr[36858]= -2103375398;
assign addr[36859]= -2020577882;
assign addr[36860]= -1896833245;
assign addr[36861]= -1734649179;
assign addr[36862]= -1537312353;
assign addr[36863]= -1308821808;
assign addr[36864]= -1053807919;
assign addr[36865]= -777438554;
assign addr[36866]= -485314355;
assign addr[36867]= -183355234;
assign addr[36868]= 122319591;
assign addr[36869]= 425515602;
assign addr[36870]= 720088517;
assign addr[36871]= 1000068799;
assign addr[36872]= 1259782632;
assign addr[36873]= 1493966902;
assign addr[36874]= 1697875851;
assign addr[36875]= 1867377253;
assign addr[36876]= 1999036154;
assign addr[36877]= 2090184478;
assign addr[36878]= 2138975100;
assign addr[36879]= 2144419275;
assign addr[36880]= 2106406677;
assign addr[36881]= 2025707632;
assign addr[36882]= 1903957513;
assign addr[36883]= 1743623590;
assign addr[36884]= 1547955041;
assign addr[36885]= 1320917099;
assign addr[36886]= 1067110699;
assign addr[36887]= 791679244;
assign addr[36888]= 500204365;
assign addr[36889]= 198592817;
assign addr[36890]= -107043224;
assign addr[36891]= -410510029;
assign addr[36892]= -705657826;
assign addr[36893]= -986505429;
assign addr[36894]= -1247361445;
assign addr[36895]= -1482939614;
assign addr[36896]= -1688465931;
assign addr[36897]= -1859775393;
assign addr[36898]= -1993396407;
assign addr[36899]= -2086621133;
assign addr[36900]= -2137560369;
assign addr[36901]= -2145181827;
assign addr[36902]= -2109331059;
assign addr[36903]= -2030734582;
assign addr[36904]= -1910985158;
assign addr[36905]= -1752509516;
assign addr[36906]= -1558519173;
assign addr[36907]= -1332945355;
assign addr[36908]= -1080359326;
assign addr[36909]= -805879757;
assign addr[36910]= -515068990;
assign addr[36911]= -213820322;
assign addr[36912]= 91761426;
assign addr[36913]= 395483624;
assign addr[36914]= 691191324;
assign addr[36915]= 972891995;
assign addr[36916]= 1234876957;
assign addr[36917]= 1471837070;
assign addr[36918]= 1678970324;
assign addr[36919]= 1852079154;
assign addr[36920]= 1987655498;
assign addr[36921]= 2082951896;
assign addr[36922]= 2136037160;
assign addr[36923]= 2145835515;
assign addr[36924]= 2112148396;
assign addr[36925]= 2035658475;
assign addr[36926]= 1917915825;
assign addr[36927]= 1761306505;
assign addr[36928]= 1569004214;
assign addr[36929]= 1344905966;
assign addr[36930]= 1093553126;
assign addr[36931]= 820039373;
assign addr[36932]= 529907477;
assign addr[36933]= 229036977;
assign addr[36934]= -76474970;
assign addr[36935]= -380437148;
assign addr[36936]= -676689746;
assign addr[36937]= -959229189;
assign addr[36938]= -1222329801;
assign addr[36939]= -1460659832;
assign addr[36940]= -1669389513;
assign addr[36941]= -1844288924;
assign addr[36942]= -1981813720;
assign addr[36943]= -2079176953;
assign addr[36944]= -2134405552;
assign addr[36945]= -2146380306;
assign addr[36946]= -2114858546;
assign addr[36947]= -2040479063;
assign addr[36948]= -1924749160;
assign addr[36949]= -1770014111;
assign addr[36950]= -1579409630;
assign addr[36951]= -1356798326;
assign addr[36952]= -1106691431;
assign addr[36953]= -834157373;
assign addr[36954]= -544719071;
assign addr[36955]= -244242007;
assign addr[36956]= 61184634;
assign addr[36957]= 365371365;
assign addr[36958]= 662153826;
assign addr[36959]= 945517704;
assign addr[36960]= 1209720613;
assign addr[36961]= 1449408469;
assign addr[36962]= 1659723983;
assign addr[36963]= 1836405100;
assign addr[36964]= 1975871368;
assign addr[36965]= 2075296495;
assign addr[36966]= 2132665626;
assign addr[36967]= 2146816171;
assign addr[36968]= 2117461370;
assign addr[36969]= 2045196100;
assign addr[36970]= 1931484818;
assign addr[36971]= 1778631892;
assign addr[36972]= 1589734894;
assign addr[36973]= 1368621831;
assign addr[36974]= 1119773573;
assign addr[36975]= 848233042;
assign addr[36976]= 559503022;
assign addr[36977]= 259434643;
assign addr[36978]= -45891193;
assign addr[36979]= -350287041;
assign addr[36980]= -647584304;
assign addr[36981]= -931758235;
assign addr[36982]= -1197050035;
assign addr[36983]= -1438083551;
assign addr[36984]= -1649974225;
assign addr[36985]= -1828428082;
assign addr[36986]= -1969828744;
assign addr[36987]= -2071310720;
assign addr[36988]= -2130817471;
assign addr[36989]= -2147143090;
assign addr[36990]= -2119956737;
assign addr[36991]= -2049809346;
assign addr[36992]= -1938122457;
assign addr[36993]= -1787159411;
assign addr[36994]= -1599979481;
assign addr[36995]= -1380375881;
assign addr[36996]= -1132798888;
assign addr[36997]= -862265664;
assign addr[36998]= -574258580;
assign addr[36999]= -274614114;
assign addr[37000]= 30595422;
assign addr[37001]= 335184940;
assign addr[37002]= 632981917;
assign addr[37003]= 917951481;
assign addr[37004]= 1184318708;
assign addr[37005]= 1426685652;
assign addr[37006]= 1640140734;
assign addr[37007]= 1820358275;
assign addr[37008]= 1963686155;
assign addr[37009]= 2067219829;
assign addr[37010]= 2128861181;
assign addr[37011]= 2147361045;
assign addr[37012]= 2122344521;
assign addr[37013]= 2054318569;
assign addr[37014]= 1944661739;
assign addr[37015]= 1795596234;
assign addr[37016]= 1610142873;
assign addr[37017]= 1392059879;
assign addr[37018]= 1145766716;
assign addr[37019]= 876254528;
assign addr[37020]= 588984994;
assign addr[37021]= 289779648;
assign addr[37022]= -15298099;
assign addr[37023]= -320065829;
assign addr[37024]= -618347408;
assign addr[37025]= -904098143;
assign addr[37026]= -1171527280;
assign addr[37027]= -1415215352;
assign addr[37028]= -1630224009;
assign addr[37029]= -1812196087;
assign addr[37030]= -1957443913;
assign addr[37031]= -2063024031;
assign addr[37032]= -2126796855;
assign addr[37033]= -2147470025;
assign addr[37034]= -2124624598;
assign addr[37035]= -2058723538;
assign addr[37036]= -1951102334;
assign addr[37037]= -1803941934;
assign addr[37038]= -1620224553;
assign addr[37039]= -1403673233;
assign addr[37040]= -1158676398;
assign addr[37041]= -890198924;
assign addr[37042]= -603681519;
assign addr[37043]= -304930476;
assign addr[37044]= 0;
assign addr[37045]= 304930476;
assign addr[37046]= 603681519;
assign addr[37047]= 890198924;
assign addr[37048]= 1158676398;
assign addr[37049]= 1403673233;
assign addr[37050]= 1620224553;
assign addr[37051]= 1803941934;
assign addr[37052]= 1951102334;
assign addr[37053]= 2058723538;
assign addr[37054]= 2124624598;
assign addr[37055]= 2147470025;
assign addr[37056]= 2126796855;
assign addr[37057]= 2063024031;
assign addr[37058]= 1957443913;
assign addr[37059]= 1812196087;
assign addr[37060]= 1630224009;
assign addr[37061]= 1415215352;
assign addr[37062]= 1171527280;
assign addr[37063]= 904098143;
assign addr[37064]= 618347408;
assign addr[37065]= 320065829;
assign addr[37066]= 15298099;
assign addr[37067]= -289779648;
assign addr[37068]= -588984994;
assign addr[37069]= -876254528;
assign addr[37070]= -1145766716;
assign addr[37071]= -1392059879;
assign addr[37072]= -1610142873;
assign addr[37073]= -1795596234;
assign addr[37074]= -1944661739;
assign addr[37075]= -2054318569;
assign addr[37076]= -2122344521;
assign addr[37077]= -2147361045;
assign addr[37078]= -2128861181;
assign addr[37079]= -2067219829;
assign addr[37080]= -1963686155;
assign addr[37081]= -1820358275;
assign addr[37082]= -1640140734;
assign addr[37083]= -1426685652;
assign addr[37084]= -1184318708;
assign addr[37085]= -917951481;
assign addr[37086]= -632981917;
assign addr[37087]= -335184940;
assign addr[37088]= -30595422;
assign addr[37089]= 274614114;
assign addr[37090]= 574258580;
assign addr[37091]= 862265664;
assign addr[37092]= 1132798888;
assign addr[37093]= 1380375881;
assign addr[37094]= 1599979481;
assign addr[37095]= 1787159411;
assign addr[37096]= 1938122457;
assign addr[37097]= 2049809346;
assign addr[37098]= 2119956737;
assign addr[37099]= 2147143090;
assign addr[37100]= 2130817471;
assign addr[37101]= 2071310720;
assign addr[37102]= 1969828744;
assign addr[37103]= 1828428082;
assign addr[37104]= 1649974225;
assign addr[37105]= 1438083551;
assign addr[37106]= 1197050035;
assign addr[37107]= 931758235;
assign addr[37108]= 647584304;
assign addr[37109]= 350287041;
assign addr[37110]= 45891193;
assign addr[37111]= -259434643;
assign addr[37112]= -559503022;
assign addr[37113]= -848233042;
assign addr[37114]= -1119773573;
assign addr[37115]= -1368621831;
assign addr[37116]= -1589734894;
assign addr[37117]= -1778631892;
assign addr[37118]= -1931484818;
assign addr[37119]= -2045196100;
assign addr[37120]= -2117461370;
assign addr[37121]= -2146816171;
assign addr[37122]= -2132665626;
assign addr[37123]= -2075296495;
assign addr[37124]= -1975871368;
assign addr[37125]= -1836405100;
assign addr[37126]= -1659723983;
assign addr[37127]= -1449408469;
assign addr[37128]= -1209720613;
assign addr[37129]= -945517704;
assign addr[37130]= -662153826;
assign addr[37131]= -365371365;
assign addr[37132]= -61184634;
assign addr[37133]= 244242007;
assign addr[37134]= 544719071;
assign addr[37135]= 834157373;
assign addr[37136]= 1106691431;
assign addr[37137]= 1356798326;
assign addr[37138]= 1579409630;
assign addr[37139]= 1770014111;
assign addr[37140]= 1924749160;
assign addr[37141]= 2040479063;
assign addr[37142]= 2114858546;
assign addr[37143]= 2146380306;
assign addr[37144]= 2134405552;
assign addr[37145]= 2079176953;
assign addr[37146]= 1981813720;
assign addr[37147]= 1844288924;
assign addr[37148]= 1669389513;
assign addr[37149]= 1460659832;
assign addr[37150]= 1222329801;
assign addr[37151]= 959229189;
assign addr[37152]= 676689746;
assign addr[37153]= 380437148;
assign addr[37154]= 76474970;
assign addr[37155]= -229036977;
assign addr[37156]= -529907477;
assign addr[37157]= -820039373;
assign addr[37158]= -1093553126;
assign addr[37159]= -1344905966;
assign addr[37160]= -1569004214;
assign addr[37161]= -1761306505;
assign addr[37162]= -1917915825;
assign addr[37163]= -2035658475;
assign addr[37164]= -2112148396;
assign addr[37165]= -2145835515;
assign addr[37166]= -2136037160;
assign addr[37167]= -2082951896;
assign addr[37168]= -1987655498;
assign addr[37169]= -1852079154;
assign addr[37170]= -1678970324;
assign addr[37171]= -1471837070;
assign addr[37172]= -1234876957;
assign addr[37173]= -972891995;
assign addr[37174]= -691191324;
assign addr[37175]= -395483624;
assign addr[37176]= -91761426;
assign addr[37177]= 213820322;
assign addr[37178]= 515068990;
assign addr[37179]= 805879757;
assign addr[37180]= 1080359326;
assign addr[37181]= 1332945355;
assign addr[37182]= 1558519173;
assign addr[37183]= 1752509516;
assign addr[37184]= 1910985158;
assign addr[37185]= 2030734582;
assign addr[37186]= 2109331059;
assign addr[37187]= 2145181827;
assign addr[37188]= 2137560369;
assign addr[37189]= 2086621133;
assign addr[37190]= 1993396407;
assign addr[37191]= 1859775393;
assign addr[37192]= 1688465931;
assign addr[37193]= 1482939614;
assign addr[37194]= 1247361445;
assign addr[37195]= 986505429;
assign addr[37196]= 705657826;
assign addr[37197]= 410510029;
assign addr[37198]= 107043224;
assign addr[37199]= -198592817;
assign addr[37200]= -500204365;
assign addr[37201]= -791679244;
assign addr[37202]= -1067110699;
assign addr[37203]= -1320917099;
assign addr[37204]= -1547955041;
assign addr[37205]= -1743623590;
assign addr[37206]= -1903957513;
assign addr[37207]= -2025707632;
assign addr[37208]= -2106406677;
assign addr[37209]= -2144419275;
assign addr[37210]= -2138975100;
assign addr[37211]= -2090184478;
assign addr[37212]= -1999036154;
assign addr[37213]= -1867377253;
assign addr[37214]= -1697875851;
assign addr[37215]= -1493966902;
assign addr[37216]= -1259782632;
assign addr[37217]= -1000068799;
assign addr[37218]= -720088517;
assign addr[37219]= -425515602;
assign addr[37220]= -122319591;
assign addr[37221]= 183355234;
assign addr[37222]= 485314355;
assign addr[37223]= 777438554;
assign addr[37224]= 1053807919;
assign addr[37225]= 1308821808;
assign addr[37226]= 1537312353;
assign addr[37227]= 1734649179;
assign addr[37228]= 1896833245;
assign addr[37229]= 2020577882;
assign addr[37230]= 2103375398;
assign addr[37231]= 2143547897;
assign addr[37232]= 2140281282;
assign addr[37233]= 2093641749;
assign addr[37234]= 2004574453;
assign addr[37235]= 1874884346;
assign addr[37236]= 1707199606;
assign addr[37237]= 1504918373;
assign addr[37238]= 1272139887;
assign addr[37239]= 1013581418;
assign addr[37240]= 734482665;
assign addr[37241]= 440499581;
assign addr[37242]= 137589750;
assign addr[37243]= -168108346;
assign addr[37244]= -470399716;
assign addr[37245]= -763158411;
assign addr[37246]= -1040451659;
assign addr[37247]= -1296660098;
assign addr[37248]= -1526591649;
assign addr[37249]= -1725586737;
assign addr[37250]= -1889612716;
assign addr[37251]= -2015345591;
assign addr[37252]= -2100237377;
assign addr[37253]= -2142567738;
assign addr[37254]= -2141478848;
assign addr[37255]= -2096992772;
assign addr[37256]= -2010011024;
assign addr[37257]= -1882296293;
assign addr[37258]= -1716436725;
assign addr[37259]= -1515793473;
assign addr[37260]= -1284432584;
assign addr[37261]= -1027042599;
assign addr[37262]= -748839539;
assign addr[37263]= -455461206;
assign addr[37264]= -152852926;
assign addr[37265]= 152852926;
assign addr[37266]= 455461206;
assign addr[37267]= 748839539;
assign addr[37268]= 1027042599;
assign addr[37269]= 1284432584;
assign addr[37270]= 1515793473;
assign addr[37271]= 1716436725;
assign addr[37272]= 1882296293;
assign addr[37273]= 2010011024;
assign addr[37274]= 2096992772;
assign addr[37275]= 2141478848;
assign addr[37276]= 2142567738;
assign addr[37277]= 2100237377;
assign addr[37278]= 2015345591;
assign addr[37279]= 1889612716;
assign addr[37280]= 1725586737;
assign addr[37281]= 1526591649;
assign addr[37282]= 1296660098;
assign addr[37283]= 1040451659;
assign addr[37284]= 763158411;
assign addr[37285]= 470399716;
assign addr[37286]= 168108346;
assign addr[37287]= -137589750;
assign addr[37288]= -440499581;
assign addr[37289]= -734482665;
assign addr[37290]= -1013581418;
assign addr[37291]= -1272139887;
assign addr[37292]= -1504918373;
assign addr[37293]= -1707199606;
assign addr[37294]= -1874884346;
assign addr[37295]= -2004574453;
assign addr[37296]= -2093641749;
assign addr[37297]= -2140281282;
assign addr[37298]= -2143547897;
assign addr[37299]= -2103375398;
assign addr[37300]= -2020577882;
assign addr[37301]= -1896833245;
assign addr[37302]= -1734649179;
assign addr[37303]= -1537312353;
assign addr[37304]= -1308821808;
assign addr[37305]= -1053807919;
assign addr[37306]= -777438554;
assign addr[37307]= -485314355;
assign addr[37308]= -183355234;
assign addr[37309]= 122319591;
assign addr[37310]= 425515602;
assign addr[37311]= 720088517;
assign addr[37312]= 1000068799;
assign addr[37313]= 1259782632;
assign addr[37314]= 1493966902;
assign addr[37315]= 1697875851;
assign addr[37316]= 1867377253;
assign addr[37317]= 1999036154;
assign addr[37318]= 2090184478;
assign addr[37319]= 2138975100;
assign addr[37320]= 2144419275;
assign addr[37321]= 2106406677;
assign addr[37322]= 2025707632;
assign addr[37323]= 1903957513;
assign addr[37324]= 1743623590;
assign addr[37325]= 1547955041;
assign addr[37326]= 1320917099;
assign addr[37327]= 1067110699;
assign addr[37328]= 791679244;
assign addr[37329]= 500204365;
assign addr[37330]= 198592817;
assign addr[37331]= -107043224;
assign addr[37332]= -410510029;
assign addr[37333]= -705657826;
assign addr[37334]= -986505429;
assign addr[37335]= -1247361445;
assign addr[37336]= -1482939614;
assign addr[37337]= -1688465931;
assign addr[37338]= -1859775393;
assign addr[37339]= -1993396407;
assign addr[37340]= -2086621133;
assign addr[37341]= -2137560369;
assign addr[37342]= -2145181827;
assign addr[37343]= -2109331059;
assign addr[37344]= -2030734582;
assign addr[37345]= -1910985158;
assign addr[37346]= -1752509516;
assign addr[37347]= -1558519173;
assign addr[37348]= -1332945355;
assign addr[37349]= -1080359326;
assign addr[37350]= -805879757;
assign addr[37351]= -515068990;
assign addr[37352]= -213820322;
assign addr[37353]= 91761426;
assign addr[37354]= 395483624;
assign addr[37355]= 691191324;
assign addr[37356]= 972891995;
assign addr[37357]= 1234876957;
assign addr[37358]= 1471837070;
assign addr[37359]= 1678970324;
assign addr[37360]= 1852079154;
assign addr[37361]= 1987655498;
assign addr[37362]= 2082951896;
assign addr[37363]= 2136037160;
assign addr[37364]= 2145835515;
assign addr[37365]= 2112148396;
assign addr[37366]= 2035658475;
assign addr[37367]= 1917915825;
assign addr[37368]= 1761306505;
assign addr[37369]= 1569004214;
assign addr[37370]= 1344905966;
assign addr[37371]= 1093553126;
assign addr[37372]= 820039373;
assign addr[37373]= 529907477;
assign addr[37374]= 229036977;
assign addr[37375]= -76474970;
assign addr[37376]= -380437148;
assign addr[37377]= -676689746;
assign addr[37378]= -959229189;
assign addr[37379]= -1222329801;
assign addr[37380]= -1460659832;
assign addr[37381]= -1669389513;
assign addr[37382]= -1844288924;
assign addr[37383]= -1981813720;
assign addr[37384]= -2079176953;
assign addr[37385]= -2134405552;
assign addr[37386]= -2146380306;
assign addr[37387]= -2114858546;
assign addr[37388]= -2040479063;
assign addr[37389]= -1924749160;
assign addr[37390]= -1770014111;
assign addr[37391]= -1579409630;
assign addr[37392]= -1356798326;
assign addr[37393]= -1106691431;
assign addr[37394]= -834157373;
assign addr[37395]= -544719071;
assign addr[37396]= -244242007;
assign addr[37397]= 61184634;
assign addr[37398]= 365371365;
assign addr[37399]= 662153826;
assign addr[37400]= 945517704;
assign addr[37401]= 1209720613;
assign addr[37402]= 1449408469;
assign addr[37403]= 1659723983;
assign addr[37404]= 1836405100;
assign addr[37405]= 1975871368;
assign addr[37406]= 2075296495;
assign addr[37407]= 2132665626;
assign addr[37408]= 2146816171;
assign addr[37409]= 2117461370;
assign addr[37410]= 2045196100;
assign addr[37411]= 1931484818;
assign addr[37412]= 1778631892;
assign addr[37413]= 1589734894;
assign addr[37414]= 1368621831;
assign addr[37415]= 1119773573;
assign addr[37416]= 848233042;
assign addr[37417]= 559503022;
assign addr[37418]= 259434643;
assign addr[37419]= -45891193;
assign addr[37420]= -350287041;
assign addr[37421]= -647584304;
assign addr[37422]= -931758235;
assign addr[37423]= -1197050035;
assign addr[37424]= -1438083551;
assign addr[37425]= -1649974225;
assign addr[37426]= -1828428082;
assign addr[37427]= -1969828744;
assign addr[37428]= -2071310720;
assign addr[37429]= -2130817471;
assign addr[37430]= -2147143090;
assign addr[37431]= -2119956737;
assign addr[37432]= -2049809346;
assign addr[37433]= -1938122457;
assign addr[37434]= -1787159411;
assign addr[37435]= -1599979481;
assign addr[37436]= -1380375881;
assign addr[37437]= -1132798888;
assign addr[37438]= -862265664;
assign addr[37439]= -574258580;
assign addr[37440]= -274614114;
assign addr[37441]= 30595422;
assign addr[37442]= 335184940;
assign addr[37443]= 632981917;
assign addr[37444]= 917951481;
assign addr[37445]= 1184318708;
assign addr[37446]= 1426685652;
assign addr[37447]= 1640140734;
assign addr[37448]= 1820358275;
assign addr[37449]= 1963686155;
assign addr[37450]= 2067219829;
assign addr[37451]= 2128861181;
assign addr[37452]= 2147361045;
assign addr[37453]= 2122344521;
assign addr[37454]= 2054318569;
assign addr[37455]= 1944661739;
assign addr[37456]= 1795596234;
assign addr[37457]= 1610142873;
assign addr[37458]= 1392059879;
assign addr[37459]= 1145766716;
assign addr[37460]= 876254528;
assign addr[37461]= 588984994;
assign addr[37462]= 289779648;
assign addr[37463]= -15298099;
assign addr[37464]= -320065829;
assign addr[37465]= -618347408;
assign addr[37466]= -904098143;
assign addr[37467]= -1171527280;
assign addr[37468]= -1415215352;
assign addr[37469]= -1630224009;
assign addr[37470]= -1812196087;
assign addr[37471]= -1957443913;
assign addr[37472]= -2063024031;
assign addr[37473]= -2126796855;
assign addr[37474]= -2147470025;
assign addr[37475]= -2124624598;
assign addr[37476]= -2058723538;
assign addr[37477]= -1951102334;
assign addr[37478]= -1803941934;
assign addr[37479]= -1620224553;
assign addr[37480]= -1403673233;
assign addr[37481]= -1158676398;
assign addr[37482]= -890198924;
assign addr[37483]= -603681519;
assign addr[37484]= -304930476;
assign addr[37485]= 0;
assign addr[37486]= 304930476;
assign addr[37487]= 603681519;
assign addr[37488]= 890198924;
assign addr[37489]= 1158676398;
assign addr[37490]= 1403673233;
assign addr[37491]= 1620224553;
assign addr[37492]= 1803941934;
assign addr[37493]= 1951102334;
assign addr[37494]= 2058723538;
assign addr[37495]= 2124624598;
assign addr[37496]= 2147470025;
assign addr[37497]= 2126796855;
assign addr[37498]= 2063024031;
assign addr[37499]= 1957443913;
assign addr[37500]= 1812196087;
assign addr[37501]= 1630224009;
assign addr[37502]= 1415215352;
assign addr[37503]= 1171527280;
assign addr[37504]= 904098143;
assign addr[37505]= 618347408;
assign addr[37506]= 320065829;
assign addr[37507]= 15298099;
assign addr[37508]= -289779648;
assign addr[37509]= -588984994;
assign addr[37510]= -876254528;
assign addr[37511]= -1145766716;
assign addr[37512]= -1392059879;
assign addr[37513]= -1610142873;
assign addr[37514]= -1795596234;
assign addr[37515]= -1944661739;
assign addr[37516]= -2054318569;
assign addr[37517]= -2122344521;
assign addr[37518]= -2147361045;
assign addr[37519]= -2128861181;
assign addr[37520]= -2067219829;
assign addr[37521]= -1963686155;
assign addr[37522]= -1820358275;
assign addr[37523]= -1640140734;
assign addr[37524]= -1426685652;
assign addr[37525]= -1184318708;
assign addr[37526]= -917951481;
assign addr[37527]= -632981917;
assign addr[37528]= -335184940;
assign addr[37529]= -30595422;
assign addr[37530]= 274614114;
assign addr[37531]= 574258580;
assign addr[37532]= 862265664;
assign addr[37533]= 1132798888;
assign addr[37534]= 1380375881;
assign addr[37535]= 1599979481;
assign addr[37536]= 1787159411;
assign addr[37537]= 1938122457;
assign addr[37538]= 2049809346;
assign addr[37539]= 2119956737;
assign addr[37540]= 2147143090;
assign addr[37541]= 2130817471;
assign addr[37542]= 2071310720;
assign addr[37543]= 1969828744;
assign addr[37544]= 1828428082;
assign addr[37545]= 1649974225;
assign addr[37546]= 1438083551;
assign addr[37547]= 1197050035;
assign addr[37548]= 931758235;
assign addr[37549]= 647584304;
assign addr[37550]= 350287041;
assign addr[37551]= 45891193;
assign addr[37552]= -259434643;
assign addr[37553]= -559503022;
assign addr[37554]= -848233042;
assign addr[37555]= -1119773573;
assign addr[37556]= -1368621831;
assign addr[37557]= -1589734894;
assign addr[37558]= -1778631892;
assign addr[37559]= -1931484818;
assign addr[37560]= -2045196100;
assign addr[37561]= -2117461370;
assign addr[37562]= -2146816171;
assign addr[37563]= -2132665626;
assign addr[37564]= -2075296495;
assign addr[37565]= -1975871368;
assign addr[37566]= -1836405100;
assign addr[37567]= -1659723983;
assign addr[37568]= -1449408469;
assign addr[37569]= -1209720613;
assign addr[37570]= -945517704;
assign addr[37571]= -662153826;
assign addr[37572]= -365371365;
assign addr[37573]= -61184634;
assign addr[37574]= 244242007;
assign addr[37575]= 544719071;
assign addr[37576]= 834157373;
assign addr[37577]= 1106691431;
assign addr[37578]= 1356798326;
assign addr[37579]= 1579409630;
assign addr[37580]= 1770014111;
assign addr[37581]= 1924749160;
assign addr[37582]= 2040479063;
assign addr[37583]= 2114858546;
assign addr[37584]= 2146380306;
assign addr[37585]= 2134405552;
assign addr[37586]= 2079176953;
assign addr[37587]= 1981813720;
assign addr[37588]= 1844288924;
assign addr[37589]= 1669389513;
assign addr[37590]= 1460659832;
assign addr[37591]= 1222329801;
assign addr[37592]= 959229189;
assign addr[37593]= 676689746;
assign addr[37594]= 380437148;
assign addr[37595]= 76474970;
assign addr[37596]= -229036977;
assign addr[37597]= -529907477;
assign addr[37598]= -820039373;
assign addr[37599]= -1093553126;
assign addr[37600]= -1344905966;
assign addr[37601]= -1569004214;
assign addr[37602]= -1761306505;
assign addr[37603]= -1917915825;
assign addr[37604]= -2035658475;
assign addr[37605]= -2112148396;
assign addr[37606]= -2145835515;
assign addr[37607]= -2136037160;
assign addr[37608]= -2082951896;
assign addr[37609]= -1987655498;
assign addr[37610]= -1852079154;
assign addr[37611]= -1678970324;
assign addr[37612]= -1471837070;
assign addr[37613]= -1234876957;
assign addr[37614]= -972891995;
assign addr[37615]= -691191324;
assign addr[37616]= -395483624;
assign addr[37617]= -91761426;
assign addr[37618]= 213820322;
assign addr[37619]= 515068990;
assign addr[37620]= 805879757;
assign addr[37621]= 1080359326;
assign addr[37622]= 1332945355;
assign addr[37623]= 1558519173;
assign addr[37624]= 1752509516;
assign addr[37625]= 1910985158;
assign addr[37626]= 2030734582;
assign addr[37627]= 2109331059;
assign addr[37628]= 2145181827;
assign addr[37629]= 2137560369;
assign addr[37630]= 2086621133;
assign addr[37631]= 1993396407;
assign addr[37632]= 1859775393;
assign addr[37633]= 1688465931;
assign addr[37634]= 1482939614;
assign addr[37635]= 1247361445;
assign addr[37636]= 986505429;
assign addr[37637]= 705657826;
assign addr[37638]= 410510029;
assign addr[37639]= 107043224;
assign addr[37640]= -198592817;
assign addr[37641]= -500204365;
assign addr[37642]= -791679244;
assign addr[37643]= -1067110699;
assign addr[37644]= -1320917099;
assign addr[37645]= -1547955041;
assign addr[37646]= -1743623590;
assign addr[37647]= -1903957513;
assign addr[37648]= -2025707632;
assign addr[37649]= -2106406677;
assign addr[37650]= -2144419275;
assign addr[37651]= -2138975100;
assign addr[37652]= -2090184478;
assign addr[37653]= -1999036154;
assign addr[37654]= -1867377253;
assign addr[37655]= -1697875851;
assign addr[37656]= -1493966902;
assign addr[37657]= -1259782632;
assign addr[37658]= -1000068799;
assign addr[37659]= -720088517;
assign addr[37660]= -425515602;
assign addr[37661]= -122319591;
assign addr[37662]= 183355234;
assign addr[37663]= 485314355;
assign addr[37664]= 777438554;
assign addr[37665]= 1053807919;
assign addr[37666]= 1308821808;
assign addr[37667]= 1537312353;
assign addr[37668]= 1734649179;
assign addr[37669]= 1896833245;
assign addr[37670]= 2020577882;
assign addr[37671]= 2103375398;
assign addr[37672]= 2143547897;
assign addr[37673]= 2140281282;
assign addr[37674]= 2093641749;
assign addr[37675]= 2004574453;
assign addr[37676]= 1874884346;
assign addr[37677]= 1707199606;
assign addr[37678]= 1504918373;
assign addr[37679]= 1272139887;
assign addr[37680]= 1013581418;
assign addr[37681]= 734482665;
assign addr[37682]= 440499581;
assign addr[37683]= 137589750;
assign addr[37684]= -168108346;
assign addr[37685]= -470399716;
assign addr[37686]= -763158411;
assign addr[37687]= -1040451659;
assign addr[37688]= -1296660098;
assign addr[37689]= -1526591649;
assign addr[37690]= -1725586737;
assign addr[37691]= -1889612716;
assign addr[37692]= -2015345591;
assign addr[37693]= -2100237377;
assign addr[37694]= -2142567738;
assign addr[37695]= -2141478848;
assign addr[37696]= -2096992772;
assign addr[37697]= -2010011024;
assign addr[37698]= -1882296293;
assign addr[37699]= -1716436725;
assign addr[37700]= -1515793473;
assign addr[37701]= -1284432584;
assign addr[37702]= -1027042599;
assign addr[37703]= -748839539;
assign addr[37704]= -455461206;
assign addr[37705]= -152852926;
assign addr[37706]= 152852926;
assign addr[37707]= 455461206;
assign addr[37708]= 748839539;
assign addr[37709]= 1027042599;
assign addr[37710]= 1284432584;
assign addr[37711]= 1515793473;
assign addr[37712]= 1716436725;
assign addr[37713]= 1882296293;
assign addr[37714]= 2010011024;
assign addr[37715]= 2096992772;
assign addr[37716]= 2141478848;
assign addr[37717]= 2142567738;
assign addr[37718]= 2100237377;
assign addr[37719]= 2015345591;
assign addr[37720]= 1889612716;
assign addr[37721]= 1725586737;
assign addr[37722]= 1526591649;
assign addr[37723]= 1296660098;
assign addr[37724]= 1040451659;
assign addr[37725]= 763158411;
assign addr[37726]= 470399716;
assign addr[37727]= 168108346;
assign addr[37728]= -137589750;
assign addr[37729]= -440499581;
assign addr[37730]= -734482665;
assign addr[37731]= -1013581418;
assign addr[37732]= -1272139887;
assign addr[37733]= -1504918373;
assign addr[37734]= -1707199606;
assign addr[37735]= -1874884346;
assign addr[37736]= -2004574453;
assign addr[37737]= -2093641749;
assign addr[37738]= -2140281282;
assign addr[37739]= -2143547897;
assign addr[37740]= -2103375398;
assign addr[37741]= -2020577882;
assign addr[37742]= -1896833245;
assign addr[37743]= -1734649179;
assign addr[37744]= -1537312353;
assign addr[37745]= -1308821808;
assign addr[37746]= -1053807919;
assign addr[37747]= -777438554;
assign addr[37748]= -485314355;
assign addr[37749]= -183355234;
assign addr[37750]= 122319591;
assign addr[37751]= 425515602;
assign addr[37752]= 720088517;
assign addr[37753]= 1000068799;
assign addr[37754]= 1259782632;
assign addr[37755]= 1493966902;
assign addr[37756]= 1697875851;
assign addr[37757]= 1867377253;
assign addr[37758]= 1999036154;
assign addr[37759]= 2090184478;
assign addr[37760]= 2138975100;
assign addr[37761]= 2144419275;
assign addr[37762]= 2106406677;
assign addr[37763]= 2025707632;
assign addr[37764]= 1903957513;
assign addr[37765]= 1743623590;
assign addr[37766]= 1547955041;
assign addr[37767]= 1320917099;
assign addr[37768]= 1067110699;
assign addr[37769]= 791679244;
assign addr[37770]= 500204365;
assign addr[37771]= 198592817;
assign addr[37772]= -107043224;
assign addr[37773]= -410510029;
assign addr[37774]= -705657826;
assign addr[37775]= -986505429;
assign addr[37776]= -1247361445;
assign addr[37777]= -1482939614;
assign addr[37778]= -1688465931;
assign addr[37779]= -1859775393;
assign addr[37780]= -1993396407;
assign addr[37781]= -2086621133;
assign addr[37782]= -2137560369;
assign addr[37783]= -2145181827;
assign addr[37784]= -2109331059;
assign addr[37785]= -2030734582;
assign addr[37786]= -1910985158;
assign addr[37787]= -1752509516;
assign addr[37788]= -1558519173;
assign addr[37789]= -1332945355;
assign addr[37790]= -1080359326;
assign addr[37791]= -805879757;
assign addr[37792]= -515068990;
assign addr[37793]= -213820322;
assign addr[37794]= 91761426;
assign addr[37795]= 395483624;
assign addr[37796]= 691191324;
assign addr[37797]= 972891995;
assign addr[37798]= 1234876957;
assign addr[37799]= 1471837070;
assign addr[37800]= 1678970324;
assign addr[37801]= 1852079154;
assign addr[37802]= 1987655498;
assign addr[37803]= 2082951896;
assign addr[37804]= 2136037160;
assign addr[37805]= 2145835515;
assign addr[37806]= 2112148396;
assign addr[37807]= 2035658475;
assign addr[37808]= 1917915825;
assign addr[37809]= 1761306505;
assign addr[37810]= 1569004214;
assign addr[37811]= 1344905966;
assign addr[37812]= 1093553126;
assign addr[37813]= 820039373;
assign addr[37814]= 529907477;
assign addr[37815]= 229036977;
assign addr[37816]= -76474970;
assign addr[37817]= -380437148;
assign addr[37818]= -676689746;
assign addr[37819]= -959229189;
assign addr[37820]= -1222329801;
assign addr[37821]= -1460659832;
assign addr[37822]= -1669389513;
assign addr[37823]= -1844288924;
assign addr[37824]= -1981813720;
assign addr[37825]= -2079176953;
assign addr[37826]= -2134405552;
assign addr[37827]= -2146380306;
assign addr[37828]= -2114858546;
assign addr[37829]= -2040479063;
assign addr[37830]= -1924749160;
assign addr[37831]= -1770014111;
assign addr[37832]= -1579409630;
assign addr[37833]= -1356798326;
assign addr[37834]= -1106691431;
assign addr[37835]= -834157373;
assign addr[37836]= -544719071;
assign addr[37837]= -244242007;
assign addr[37838]= 61184634;
assign addr[37839]= 365371365;
assign addr[37840]= 662153826;
assign addr[37841]= 945517704;
assign addr[37842]= 1209720613;
assign addr[37843]= 1449408469;
assign addr[37844]= 1659723983;
assign addr[37845]= 1836405100;
assign addr[37846]= 1975871368;
assign addr[37847]= 2075296495;
assign addr[37848]= 2132665626;
assign addr[37849]= 2146816171;
assign addr[37850]= 2117461370;
assign addr[37851]= 2045196100;
assign addr[37852]= 1931484818;
assign addr[37853]= 1778631892;
assign addr[37854]= 1589734894;
assign addr[37855]= 1368621831;
assign addr[37856]= 1119773573;
assign addr[37857]= 848233042;
assign addr[37858]= 559503022;
assign addr[37859]= 259434643;
assign addr[37860]= -45891193;
assign addr[37861]= -350287041;
assign addr[37862]= -647584304;
assign addr[37863]= -931758235;
assign addr[37864]= -1197050035;
assign addr[37865]= -1438083551;
assign addr[37866]= -1649974225;
assign addr[37867]= -1828428082;
assign addr[37868]= -1969828744;
assign addr[37869]= -2071310720;
assign addr[37870]= -2130817471;
assign addr[37871]= -2147143090;
assign addr[37872]= -2119956737;
assign addr[37873]= -2049809346;
assign addr[37874]= -1938122457;
assign addr[37875]= -1787159411;
assign addr[37876]= -1599979481;
assign addr[37877]= -1380375881;
assign addr[37878]= -1132798888;
assign addr[37879]= -862265664;
assign addr[37880]= -574258580;
assign addr[37881]= -274614114;
assign addr[37882]= 30595422;
assign addr[37883]= 335184940;
assign addr[37884]= 632981917;
assign addr[37885]= 917951481;
assign addr[37886]= 1184318708;
assign addr[37887]= 1426685652;
assign addr[37888]= 1640140734;
assign addr[37889]= 1820358275;
assign addr[37890]= 1963686155;
assign addr[37891]= 2067219829;
assign addr[37892]= 2128861181;
assign addr[37893]= 2147361045;
assign addr[37894]= 2122344521;
assign addr[37895]= 2054318569;
assign addr[37896]= 1944661739;
assign addr[37897]= 1795596234;
assign addr[37898]= 1610142873;
assign addr[37899]= 1392059879;
assign addr[37900]= 1145766716;
assign addr[37901]= 876254528;
assign addr[37902]= 588984994;
assign addr[37903]= 289779648;
assign addr[37904]= -15298099;
assign addr[37905]= -320065829;
assign addr[37906]= -618347408;
assign addr[37907]= -904098143;
assign addr[37908]= -1171527280;
assign addr[37909]= -1415215352;
assign addr[37910]= -1630224009;
assign addr[37911]= -1812196087;
assign addr[37912]= -1957443913;
assign addr[37913]= -2063024031;
assign addr[37914]= -2126796855;
assign addr[37915]= -2147470025;
assign addr[37916]= -2124624598;
assign addr[37917]= -2058723538;
assign addr[37918]= -1951102334;
assign addr[37919]= -1803941934;
assign addr[37920]= -1620224553;
assign addr[37921]= -1403673233;
assign addr[37922]= -1158676398;
assign addr[37923]= -890198924;
assign addr[37924]= -603681519;
assign addr[37925]= -304930476;
assign addr[37926]= 0;
assign addr[37927]= 304930476;
assign addr[37928]= 603681519;
assign addr[37929]= 890198924;
assign addr[37930]= 1158676398;
assign addr[37931]= 1403673233;
assign addr[37932]= 1620224553;
assign addr[37933]= 1803941934;
assign addr[37934]= 1951102334;
assign addr[37935]= 2058723538;
assign addr[37936]= 2124624598;
assign addr[37937]= 2147470025;
assign addr[37938]= 2126796855;
assign addr[37939]= 2063024031;
assign addr[37940]= 1957443913;
assign addr[37941]= 1812196087;
assign addr[37942]= 1630224009;
assign addr[37943]= 1415215352;
assign addr[37944]= 1171527280;
assign addr[37945]= 904098143;
assign addr[37946]= 618347408;
assign addr[37947]= 320065829;
assign addr[37948]= 15298099;
assign addr[37949]= -289779648;
assign addr[37950]= -588984994;
assign addr[37951]= -876254528;
assign addr[37952]= -1145766716;
assign addr[37953]= -1392059879;
assign addr[37954]= -1610142873;
assign addr[37955]= -1795596234;
assign addr[37956]= -1944661739;
assign addr[37957]= -2054318569;
assign addr[37958]= -2122344521;
assign addr[37959]= -2147361045;
assign addr[37960]= -2128861181;
assign addr[37961]= -2067219829;
assign addr[37962]= -1963686155;
assign addr[37963]= -1820358275;
assign addr[37964]= -1640140734;
assign addr[37965]= -1426685652;
assign addr[37966]= -1184318708;
assign addr[37967]= -917951481;
assign addr[37968]= -632981917;
assign addr[37969]= -335184940;
assign addr[37970]= -30595422;
assign addr[37971]= 274614114;
assign addr[37972]= 574258580;
assign addr[37973]= 862265664;
assign addr[37974]= 1132798888;
assign addr[37975]= 1380375881;
assign addr[37976]= 1599979481;
assign addr[37977]= 1787159411;
assign addr[37978]= 1938122457;
assign addr[37979]= 2049809346;
assign addr[37980]= 2119956737;
assign addr[37981]= 2147143090;
assign addr[37982]= 2130817471;
assign addr[37983]= 2071310720;
assign addr[37984]= 1969828744;
assign addr[37985]= 1828428082;
assign addr[37986]= 1649974225;
assign addr[37987]= 1438083551;
assign addr[37988]= 1197050035;
assign addr[37989]= 931758235;
assign addr[37990]= 647584304;
assign addr[37991]= 350287041;
assign addr[37992]= 45891193;
assign addr[37993]= -259434643;
assign addr[37994]= -559503022;
assign addr[37995]= -848233042;
assign addr[37996]= -1119773573;
assign addr[37997]= -1368621831;
assign addr[37998]= -1589734894;
assign addr[37999]= -1778631892;
assign addr[38000]= -1931484818;
assign addr[38001]= -2045196100;
assign addr[38002]= -2117461370;
assign addr[38003]= -2146816171;
assign addr[38004]= -2132665626;
assign addr[38005]= -2075296495;
assign addr[38006]= -1975871368;
assign addr[38007]= -1836405100;
assign addr[38008]= -1659723983;
assign addr[38009]= -1449408469;
assign addr[38010]= -1209720613;
assign addr[38011]= -945517704;
assign addr[38012]= -662153826;
assign addr[38013]= -365371365;
assign addr[38014]= -61184634;
assign addr[38015]= 244242007;
assign addr[38016]= 544719071;
assign addr[38017]= 834157373;
assign addr[38018]= 1106691431;
assign addr[38019]= 1356798326;
assign addr[38020]= 1579409630;
assign addr[38021]= 1770014111;
assign addr[38022]= 1924749160;
assign addr[38023]= 2040479063;
assign addr[38024]= 2114858546;
assign addr[38025]= 2146380306;
assign addr[38026]= 2134405552;
assign addr[38027]= 2079176953;
assign addr[38028]= 1981813720;
assign addr[38029]= 1844288924;
assign addr[38030]= 1669389513;
assign addr[38031]= 1460659832;
assign addr[38032]= 1222329801;
assign addr[38033]= 959229189;
assign addr[38034]= 676689746;
assign addr[38035]= 380437148;
assign addr[38036]= 76474970;
assign addr[38037]= -229036977;
assign addr[38038]= -529907477;
assign addr[38039]= -820039373;
assign addr[38040]= -1093553126;
assign addr[38041]= -1344905966;
assign addr[38042]= -1569004214;
assign addr[38043]= -1761306505;
assign addr[38044]= -1917915825;
assign addr[38045]= -2035658475;
assign addr[38046]= -2112148396;
assign addr[38047]= -2145835515;
assign addr[38048]= -2136037160;
assign addr[38049]= -2082951896;
assign addr[38050]= -1987655498;
assign addr[38051]= -1852079154;
assign addr[38052]= -1678970324;
assign addr[38053]= -1471837070;
assign addr[38054]= -1234876957;
assign addr[38055]= -972891995;
assign addr[38056]= -691191324;
assign addr[38057]= -395483624;
assign addr[38058]= -91761426;
assign addr[38059]= 213820322;
assign addr[38060]= 515068990;
assign addr[38061]= 805879757;
assign addr[38062]= 1080359326;
assign addr[38063]= 1332945355;
assign addr[38064]= 1558519173;
assign addr[38065]= 1752509516;
assign addr[38066]= 1910985158;
assign addr[38067]= 2030734582;
assign addr[38068]= 2109331059;
assign addr[38069]= 2145181827;
assign addr[38070]= 2137560369;
assign addr[38071]= 2086621133;
assign addr[38072]= 1993396407;
assign addr[38073]= 1859775393;
assign addr[38074]= 1688465931;
assign addr[38075]= 1482939614;
assign addr[38076]= 1247361445;
assign addr[38077]= 986505429;
assign addr[38078]= 705657826;
assign addr[38079]= 410510029;
assign addr[38080]= 107043224;
assign addr[38081]= -198592817;
assign addr[38082]= -500204365;
assign addr[38083]= -791679244;
assign addr[38084]= -1067110699;
assign addr[38085]= -1320917099;
assign addr[38086]= -1547955041;
assign addr[38087]= -1743623590;
assign addr[38088]= -1903957513;
assign addr[38089]= -2025707632;
assign addr[38090]= -2106406677;
assign addr[38091]= -2144419275;
assign addr[38092]= -2138975100;
assign addr[38093]= -2090184478;
assign addr[38094]= -1999036154;
assign addr[38095]= -1867377253;
assign addr[38096]= -1697875851;
assign addr[38097]= -1493966902;
assign addr[38098]= -1259782632;
assign addr[38099]= -1000068799;
assign addr[38100]= -720088517;
assign addr[38101]= -425515602;
assign addr[38102]= -122319591;
assign addr[38103]= 183355234;
assign addr[38104]= 485314355;
assign addr[38105]= 777438554;
assign addr[38106]= 1053807919;
assign addr[38107]= 1308821808;
assign addr[38108]= 1537312353;
assign addr[38109]= 1734649179;
assign addr[38110]= 1896833245;
assign addr[38111]= 2020577882;
assign addr[38112]= 2103375398;
assign addr[38113]= 2143547897;
assign addr[38114]= 2140281282;
assign addr[38115]= 2093641749;
assign addr[38116]= 2004574453;
assign addr[38117]= 1874884346;
assign addr[38118]= 1707199606;
assign addr[38119]= 1504918373;
assign addr[38120]= 1272139887;
assign addr[38121]= 1013581418;
assign addr[38122]= 734482665;
assign addr[38123]= 440499581;
assign addr[38124]= 137589750;
assign addr[38125]= -168108346;
assign addr[38126]= -470399716;
assign addr[38127]= -763158411;
assign addr[38128]= -1040451659;
assign addr[38129]= -1296660098;
assign addr[38130]= -1526591649;
assign addr[38131]= -1725586737;
assign addr[38132]= -1889612716;
assign addr[38133]= -2015345591;
assign addr[38134]= -2100237377;
assign addr[38135]= -2142567738;
assign addr[38136]= -2141478848;
assign addr[38137]= -2096992772;
assign addr[38138]= -2010011024;
assign addr[38139]= -1882296293;
assign addr[38140]= -1716436725;
assign addr[38141]= -1515793473;
assign addr[38142]= -1284432584;
assign addr[38143]= -1027042599;
assign addr[38144]= -748839539;
assign addr[38145]= -455461206;
assign addr[38146]= -152852926;
assign addr[38147]= 152852926;
assign addr[38148]= 455461206;
assign addr[38149]= 748839539;
assign addr[38150]= 1027042599;
assign addr[38151]= 1284432584;
assign addr[38152]= 1515793473;
assign addr[38153]= 1716436725;
assign addr[38154]= 1882296293;
assign addr[38155]= 2010011024;
assign addr[38156]= 2096992772;
assign addr[38157]= 2141478848;
assign addr[38158]= 2142567738;
assign addr[38159]= 2100237377;
assign addr[38160]= 2015345591;
assign addr[38161]= 1889612716;
assign addr[38162]= 1725586737;
assign addr[38163]= 1526591649;
assign addr[38164]= 1296660098;
assign addr[38165]= 1040451659;
assign addr[38166]= 763158411;
assign addr[38167]= 470399716;
assign addr[38168]= 168108346;
assign addr[38169]= -137589750;
assign addr[38170]= -440499581;
assign addr[38171]= -734482665;
assign addr[38172]= -1013581418;
assign addr[38173]= -1272139887;
assign addr[38174]= -1504918373;
assign addr[38175]= -1707199606;
assign addr[38176]= -1874884346;
assign addr[38177]= -2004574453;
assign addr[38178]= -2093641749;
assign addr[38179]= -2140281282;
assign addr[38180]= -2143547897;
assign addr[38181]= -2103375398;
assign addr[38182]= -2020577882;
assign addr[38183]= -1896833245;
assign addr[38184]= -1734649179;
assign addr[38185]= -1537312353;
assign addr[38186]= -1308821808;
assign addr[38187]= -1053807919;
assign addr[38188]= -777438554;
assign addr[38189]= -485314355;
assign addr[38190]= -183355234;
assign addr[38191]= 122319591;
assign addr[38192]= 425515602;
assign addr[38193]= 720088517;
assign addr[38194]= 1000068799;
assign addr[38195]= 1259782632;
assign addr[38196]= 1493966902;
assign addr[38197]= 1697875851;
assign addr[38198]= 1867377253;
assign addr[38199]= 1999036154;
assign addr[38200]= 2090184478;
assign addr[38201]= 2138975100;
assign addr[38202]= 2144419275;
assign addr[38203]= 2106406677;
assign addr[38204]= 2025707632;
assign addr[38205]= 1903957513;
assign addr[38206]= 1743623590;
assign addr[38207]= 1547955041;
assign addr[38208]= 1320917099;
assign addr[38209]= 1067110699;
assign addr[38210]= 791679244;
assign addr[38211]= 500204365;
assign addr[38212]= 198592817;
assign addr[38213]= -107043224;
assign addr[38214]= -410510029;
assign addr[38215]= -705657826;
assign addr[38216]= -986505429;
assign addr[38217]= -1247361445;
assign addr[38218]= -1482939614;
assign addr[38219]= -1688465931;
assign addr[38220]= -1859775393;
assign addr[38221]= -1993396407;
assign addr[38222]= -2086621133;
assign addr[38223]= -2137560369;
assign addr[38224]= -2145181827;
assign addr[38225]= -2109331059;
assign addr[38226]= -2030734582;
assign addr[38227]= -1910985158;
assign addr[38228]= -1752509516;
assign addr[38229]= -1558519173;
assign addr[38230]= -1332945355;
assign addr[38231]= -1080359326;
assign addr[38232]= -805879757;
assign addr[38233]= -515068990;
assign addr[38234]= -213820322;
assign addr[38235]= 91761426;
assign addr[38236]= 395483624;
assign addr[38237]= 691191324;
assign addr[38238]= 972891995;
assign addr[38239]= 1234876957;
assign addr[38240]= 1471837070;
assign addr[38241]= 1678970324;
assign addr[38242]= 1852079154;
assign addr[38243]= 1987655498;
assign addr[38244]= 2082951896;
assign addr[38245]= 2136037160;
assign addr[38246]= 2145835515;
assign addr[38247]= 2112148396;
assign addr[38248]= 2035658475;
assign addr[38249]= 1917915825;
assign addr[38250]= 1761306505;
assign addr[38251]= 1569004214;
assign addr[38252]= 1344905966;
assign addr[38253]= 1093553126;
assign addr[38254]= 820039373;
assign addr[38255]= 529907477;
assign addr[38256]= 229036977;
assign addr[38257]= -76474970;
assign addr[38258]= -380437148;
assign addr[38259]= -676689746;
assign addr[38260]= -959229189;
assign addr[38261]= -1222329801;
assign addr[38262]= -1460659832;
assign addr[38263]= -1669389513;
assign addr[38264]= -1844288924;
assign addr[38265]= -1981813720;
assign addr[38266]= -2079176953;
assign addr[38267]= -2134405552;
assign addr[38268]= -2146380306;
assign addr[38269]= -2114858546;
assign addr[38270]= -2040479063;
assign addr[38271]= -1924749160;
assign addr[38272]= -1770014111;
assign addr[38273]= -1579409630;
assign addr[38274]= -1356798326;
assign addr[38275]= -1106691431;
assign addr[38276]= -834157373;
assign addr[38277]= -544719071;
assign addr[38278]= -244242007;
assign addr[38279]= 61184634;
assign addr[38280]= 365371365;
assign addr[38281]= 662153826;
assign addr[38282]= 945517704;
assign addr[38283]= 1209720613;
assign addr[38284]= 1449408469;
assign addr[38285]= 1659723983;
assign addr[38286]= 1836405100;
assign addr[38287]= 1975871368;
assign addr[38288]= 2075296495;
assign addr[38289]= 2132665626;
assign addr[38290]= 2146816171;
assign addr[38291]= 2117461370;
assign addr[38292]= 2045196100;
assign addr[38293]= 1931484818;
assign addr[38294]= 1778631892;
assign addr[38295]= 1589734894;
assign addr[38296]= 1368621831;
assign addr[38297]= 1119773573;
assign addr[38298]= 848233042;
assign addr[38299]= 559503022;
assign addr[38300]= 259434643;
assign addr[38301]= -45891193;
assign addr[38302]= -350287041;
assign addr[38303]= -647584304;
assign addr[38304]= -931758235;
assign addr[38305]= -1197050035;
assign addr[38306]= -1438083551;
assign addr[38307]= -1649974225;
assign addr[38308]= -1828428082;
assign addr[38309]= -1969828744;
assign addr[38310]= -2071310720;
assign addr[38311]= -2130817471;
assign addr[38312]= -2147143090;
assign addr[38313]= -2119956737;
assign addr[38314]= -2049809346;
assign addr[38315]= -1938122457;
assign addr[38316]= -1787159411;
assign addr[38317]= -1599979481;
assign addr[38318]= -1380375881;
assign addr[38319]= -1132798888;
assign addr[38320]= -862265664;
assign addr[38321]= -574258580;
assign addr[38322]= -274614114;
assign addr[38323]= 30595422;
assign addr[38324]= 335184940;
assign addr[38325]= 632981917;
assign addr[38326]= 917951481;
assign addr[38327]= 1184318708;
assign addr[38328]= 1426685652;
assign addr[38329]= 1640140734;
assign addr[38330]= 1820358275;
assign addr[38331]= 1963686155;
assign addr[38332]= 2067219829;
assign addr[38333]= 2128861181;
assign addr[38334]= 2147361045;
assign addr[38335]= 2122344521;
assign addr[38336]= 2054318569;
assign addr[38337]= 1944661739;
assign addr[38338]= 1795596234;
assign addr[38339]= 1610142873;
assign addr[38340]= 1392059879;
assign addr[38341]= 1145766716;
assign addr[38342]= 876254528;
assign addr[38343]= 588984994;
assign addr[38344]= 289779648;
assign addr[38345]= -15298099;
assign addr[38346]= -320065829;
assign addr[38347]= -618347408;
assign addr[38348]= -904098143;
assign addr[38349]= -1171527280;
assign addr[38350]= -1415215352;
assign addr[38351]= -1630224009;
assign addr[38352]= -1812196087;
assign addr[38353]= -1957443913;
assign addr[38354]= -2063024031;
assign addr[38355]= -2126796855;
assign addr[38356]= -2147470025;
assign addr[38357]= -2124624598;
assign addr[38358]= -2058723538;
assign addr[38359]= -1951102334;
assign addr[38360]= -1803941934;
assign addr[38361]= -1620224553;
assign addr[38362]= -1403673233;
assign addr[38363]= -1158676398;
assign addr[38364]= -890198924;
assign addr[38365]= -603681519;
assign addr[38366]= -304930476;
assign addr[38367]= 0;
assign addr[38368]= 304930476;
assign addr[38369]= 603681519;
assign addr[38370]= 890198924;
assign addr[38371]= 1158676398;
assign addr[38372]= 1403673233;
assign addr[38373]= 1620224553;
assign addr[38374]= 1803941934;
assign addr[38375]= 1951102334;
assign addr[38376]= 2058723538;
assign addr[38377]= 2124624598;
assign addr[38378]= 2147470025;
assign addr[38379]= 2126796855;
assign addr[38380]= 2063024031;
assign addr[38381]= 1957443913;
assign addr[38382]= 1812196087;
assign addr[38383]= 1630224009;
assign addr[38384]= 1415215352;
assign addr[38385]= 1171527280;
assign addr[38386]= 904098143;
assign addr[38387]= 618347408;
assign addr[38388]= 320065829;
assign addr[38389]= 15298099;
assign addr[38390]= -289779648;
assign addr[38391]= -588984994;
assign addr[38392]= -876254528;
assign addr[38393]= -1145766716;
assign addr[38394]= -1392059879;
assign addr[38395]= -1610142873;
assign addr[38396]= -1795596234;
assign addr[38397]= -1944661739;
assign addr[38398]= -2054318569;
assign addr[38399]= -2122344521;
assign addr[38400]= -2147361045;
assign addr[38401]= -2128861181;
assign addr[38402]= -2067219829;
assign addr[38403]= -1963686155;
assign addr[38404]= -1820358275;
assign addr[38405]= -1640140734;
assign addr[38406]= -1426685652;
assign addr[38407]= -1184318708;
assign addr[38408]= -917951481;
assign addr[38409]= -632981917;
assign addr[38410]= -335184940;
assign addr[38411]= -30595422;
assign addr[38412]= 274614114;
assign addr[38413]= 574258580;
assign addr[38414]= 862265664;
assign addr[38415]= 1132798888;
assign addr[38416]= 1380375881;
assign addr[38417]= 1599979481;
assign addr[38418]= 1787159411;
assign addr[38419]= 1938122457;
assign addr[38420]= 2049809346;
assign addr[38421]= 2119956737;
assign addr[38422]= 2147143090;
assign addr[38423]= 2130817471;
assign addr[38424]= 2071310720;
assign addr[38425]= 1969828744;
assign addr[38426]= 1828428082;
assign addr[38427]= 1649974225;
assign addr[38428]= 1438083551;
assign addr[38429]= 1197050035;
assign addr[38430]= 931758235;
assign addr[38431]= 647584304;
assign addr[38432]= 350287041;
assign addr[38433]= 45891193;
assign addr[38434]= -259434643;
assign addr[38435]= -559503022;
assign addr[38436]= -848233042;
assign addr[38437]= -1119773573;
assign addr[38438]= -1368621831;
assign addr[38439]= -1589734894;
assign addr[38440]= -1778631892;
assign addr[38441]= -1931484818;
assign addr[38442]= -2045196100;
assign addr[38443]= -2117461370;
assign addr[38444]= -2146816171;
assign addr[38445]= -2132665626;
assign addr[38446]= -2075296495;
assign addr[38447]= -1975871368;
assign addr[38448]= -1836405100;
assign addr[38449]= -1659723983;
assign addr[38450]= -1449408469;
assign addr[38451]= -1209720613;
assign addr[38452]= -945517704;
assign addr[38453]= -662153826;
assign addr[38454]= -365371365;
assign addr[38455]= -61184634;
assign addr[38456]= 244242007;
assign addr[38457]= 544719071;
assign addr[38458]= 834157373;
assign addr[38459]= 1106691431;
assign addr[38460]= 1356798326;
assign addr[38461]= 1579409630;
assign addr[38462]= 1770014111;
assign addr[38463]= 1924749160;
assign addr[38464]= 2040479063;
assign addr[38465]= 2114858546;
assign addr[38466]= 2146380306;
assign addr[38467]= 2134405552;
assign addr[38468]= 2079176953;
assign addr[38469]= 1981813720;
assign addr[38470]= 1844288924;
assign addr[38471]= 1669389513;
assign addr[38472]= 1460659832;
assign addr[38473]= 1222329801;
assign addr[38474]= 959229189;
assign addr[38475]= 676689746;
assign addr[38476]= 380437148;
assign addr[38477]= 76474970;
assign addr[38478]= -229036977;
assign addr[38479]= -529907477;
assign addr[38480]= -820039373;
assign addr[38481]= -1093553126;
assign addr[38482]= -1344905966;
assign addr[38483]= -1569004214;
assign addr[38484]= -1761306505;
assign addr[38485]= -1917915825;
assign addr[38486]= -2035658475;
assign addr[38487]= -2112148396;
assign addr[38488]= -2145835515;
assign addr[38489]= -2136037160;
assign addr[38490]= -2082951896;
assign addr[38491]= -1987655498;
assign addr[38492]= -1852079154;
assign addr[38493]= -1678970324;
assign addr[38494]= -1471837070;
assign addr[38495]= -1234876957;
assign addr[38496]= -972891995;
assign addr[38497]= -691191324;
assign addr[38498]= -395483624;
assign addr[38499]= -91761426;
assign addr[38500]= 213820322;
assign addr[38501]= 515068990;
assign addr[38502]= 805879757;
assign addr[38503]= 1080359326;
assign addr[38504]= 1332945355;
assign addr[38505]= 1558519173;
assign addr[38506]= 1752509516;
assign addr[38507]= 1910985158;
assign addr[38508]= 2030734582;
assign addr[38509]= 2109331059;
assign addr[38510]= 2145181827;
assign addr[38511]= 2137560369;
assign addr[38512]= 2086621133;
assign addr[38513]= 1993396407;
assign addr[38514]= 1859775393;
assign addr[38515]= 1688465931;
assign addr[38516]= 1482939614;
assign addr[38517]= 1247361445;
assign addr[38518]= 986505429;
assign addr[38519]= 705657826;
assign addr[38520]= 410510029;
assign addr[38521]= 107043224;
assign addr[38522]= -198592817;
assign addr[38523]= -500204365;
assign addr[38524]= -791679244;
assign addr[38525]= -1067110699;
assign addr[38526]= -1320917099;
assign addr[38527]= -1547955041;
assign addr[38528]= -1743623590;
assign addr[38529]= -1903957513;
assign addr[38530]= -2025707632;
assign addr[38531]= -2106406677;
assign addr[38532]= -2144419275;
assign addr[38533]= -2138975100;
assign addr[38534]= -2090184478;
assign addr[38535]= -1999036154;
assign addr[38536]= -1867377253;
assign addr[38537]= -1697875851;
assign addr[38538]= -1493966902;
assign addr[38539]= -1259782632;
assign addr[38540]= -1000068799;
assign addr[38541]= -720088517;
assign addr[38542]= -425515602;
assign addr[38543]= -122319591;
assign addr[38544]= 183355234;
assign addr[38545]= 485314355;
assign addr[38546]= 777438554;
assign addr[38547]= 1053807919;
assign addr[38548]= 1308821808;
assign addr[38549]= 1537312353;
assign addr[38550]= 1734649179;
assign addr[38551]= 1896833245;
assign addr[38552]= 2020577882;
assign addr[38553]= 2103375398;
assign addr[38554]= 2143547897;
assign addr[38555]= 2140281282;
assign addr[38556]= 2093641749;
assign addr[38557]= 2004574453;
assign addr[38558]= 1874884346;
assign addr[38559]= 1707199606;
assign addr[38560]= 1504918373;
assign addr[38561]= 1272139887;
assign addr[38562]= 1013581418;
assign addr[38563]= 734482665;
assign addr[38564]= 440499581;
assign addr[38565]= 137589750;
assign addr[38566]= -168108346;
assign addr[38567]= -470399716;
assign addr[38568]= -763158411;
assign addr[38569]= -1040451659;
assign addr[38570]= -1296660098;
assign addr[38571]= -1526591649;
assign addr[38572]= -1725586737;
assign addr[38573]= -1889612716;
assign addr[38574]= -2015345591;
assign addr[38575]= -2100237377;
assign addr[38576]= -2142567738;
assign addr[38577]= -2141478848;
assign addr[38578]= -2096992772;
assign addr[38579]= -2010011024;
assign addr[38580]= -1882296293;
assign addr[38581]= -1716436725;
assign addr[38582]= -1515793473;
assign addr[38583]= -1284432584;
assign addr[38584]= -1027042599;
assign addr[38585]= -748839539;
assign addr[38586]= -455461206;
assign addr[38587]= -152852926;
assign addr[38588]= 152852926;
assign addr[38589]= 455461206;
assign addr[38590]= 748839539;
assign addr[38591]= 1027042599;
assign addr[38592]= 1284432584;
assign addr[38593]= 1515793473;
assign addr[38594]= 1716436725;
assign addr[38595]= 1882296293;
assign addr[38596]= 2010011024;
assign addr[38597]= 2096992772;
assign addr[38598]= 2141478848;
assign addr[38599]= 2142567738;
assign addr[38600]= 2100237377;
assign addr[38601]= 2015345591;
assign addr[38602]= 1889612716;
assign addr[38603]= 1725586737;
assign addr[38604]= 1526591649;
assign addr[38605]= 1296660098;
assign addr[38606]= 1040451659;
assign addr[38607]= 763158411;
assign addr[38608]= 470399716;
assign addr[38609]= 168108346;
assign addr[38610]= -137589750;
assign addr[38611]= -440499581;
assign addr[38612]= -734482665;
assign addr[38613]= -1013581418;
assign addr[38614]= -1272139887;
assign addr[38615]= -1504918373;
assign addr[38616]= -1707199606;
assign addr[38617]= -1874884346;
assign addr[38618]= -2004574453;
assign addr[38619]= -2093641749;
assign addr[38620]= -2140281282;
assign addr[38621]= -2143547897;
assign addr[38622]= -2103375398;
assign addr[38623]= -2020577882;
assign addr[38624]= -1896833245;
assign addr[38625]= -1734649179;
assign addr[38626]= -1537312353;
assign addr[38627]= -1308821808;
assign addr[38628]= -1053807919;
assign addr[38629]= -777438554;
assign addr[38630]= -485314355;
assign addr[38631]= -183355234;
assign addr[38632]= 122319591;
assign addr[38633]= 425515602;
assign addr[38634]= 720088517;
assign addr[38635]= 1000068799;
assign addr[38636]= 1259782632;
assign addr[38637]= 1493966902;
assign addr[38638]= 1697875851;
assign addr[38639]= 1867377253;
assign addr[38640]= 1999036154;
assign addr[38641]= 2090184478;
assign addr[38642]= 2138975100;
assign addr[38643]= 2144419275;
assign addr[38644]= 2106406677;
assign addr[38645]= 2025707632;
assign addr[38646]= 1903957513;
assign addr[38647]= 1743623590;
assign addr[38648]= 1547955041;
assign addr[38649]= 1320917099;
assign addr[38650]= 1067110699;
assign addr[38651]= 791679244;
assign addr[38652]= 500204365;
assign addr[38653]= 198592817;
assign addr[38654]= -107043224;
assign addr[38655]= -410510029;
assign addr[38656]= -705657826;
assign addr[38657]= -986505429;
assign addr[38658]= -1247361445;
assign addr[38659]= -1482939614;
assign addr[38660]= -1688465931;
assign addr[38661]= -1859775393;
assign addr[38662]= -1993396407;
assign addr[38663]= -2086621133;
assign addr[38664]= -2137560369;
assign addr[38665]= -2145181827;
assign addr[38666]= -2109331059;
assign addr[38667]= -2030734582;
assign addr[38668]= -1910985158;
assign addr[38669]= -1752509516;
assign addr[38670]= -1558519173;
assign addr[38671]= -1332945355;
assign addr[38672]= -1080359326;
assign addr[38673]= -805879757;
assign addr[38674]= -515068990;
assign addr[38675]= -213820322;
assign addr[38676]= 91761426;
assign addr[38677]= 395483624;
assign addr[38678]= 691191324;
assign addr[38679]= 972891995;
assign addr[38680]= 1234876957;
assign addr[38681]= 1471837070;
assign addr[38682]= 1678970324;
assign addr[38683]= 1852079154;
assign addr[38684]= 1987655498;
assign addr[38685]= 2082951896;
assign addr[38686]= 2136037160;
assign addr[38687]= 2145835515;
assign addr[38688]= 2112148396;
assign addr[38689]= 2035658475;
assign addr[38690]= 1917915825;
assign addr[38691]= 1761306505;
assign addr[38692]= 1569004214;
assign addr[38693]= 1344905966;
assign addr[38694]= 1093553126;
assign addr[38695]= 820039373;
assign addr[38696]= 529907477;
assign addr[38697]= 229036977;
assign addr[38698]= -76474970;
assign addr[38699]= -380437148;
assign addr[38700]= -676689746;
assign addr[38701]= -959229189;
assign addr[38702]= -1222329801;
assign addr[38703]= -1460659832;
assign addr[38704]= -1669389513;
assign addr[38705]= -1844288924;
assign addr[38706]= -1981813720;
assign addr[38707]= -2079176953;
assign addr[38708]= -2134405552;
assign addr[38709]= -2146380306;
assign addr[38710]= -2114858546;
assign addr[38711]= -2040479063;
assign addr[38712]= -1924749160;
assign addr[38713]= -1770014111;
assign addr[38714]= -1579409630;
assign addr[38715]= -1356798326;
assign addr[38716]= -1106691431;
assign addr[38717]= -834157373;
assign addr[38718]= -544719071;
assign addr[38719]= -244242007;
assign addr[38720]= 61184634;
assign addr[38721]= 365371365;
assign addr[38722]= 662153826;
assign addr[38723]= 945517704;
assign addr[38724]= 1209720613;
assign addr[38725]= 1449408469;
assign addr[38726]= 1659723983;
assign addr[38727]= 1836405100;
assign addr[38728]= 1975871368;
assign addr[38729]= 2075296495;
assign addr[38730]= 2132665626;
assign addr[38731]= 2146816171;
assign addr[38732]= 2117461370;
assign addr[38733]= 2045196100;
assign addr[38734]= 1931484818;
assign addr[38735]= 1778631892;
assign addr[38736]= 1589734894;
assign addr[38737]= 1368621831;
assign addr[38738]= 1119773573;
assign addr[38739]= 848233042;
assign addr[38740]= 559503022;
assign addr[38741]= 259434643;
assign addr[38742]= -45891193;
assign addr[38743]= -350287041;
assign addr[38744]= -647584304;
assign addr[38745]= -931758235;
assign addr[38746]= -1197050035;
assign addr[38747]= -1438083551;
assign addr[38748]= -1649974225;
assign addr[38749]= -1828428082;
assign addr[38750]= -1969828744;
assign addr[38751]= -2071310720;
assign addr[38752]= -2130817471;
assign addr[38753]= -2147143090;
assign addr[38754]= -2119956737;
assign addr[38755]= -2049809346;
assign addr[38756]= -1938122457;
assign addr[38757]= -1787159411;
assign addr[38758]= -1599979481;
assign addr[38759]= -1380375881;
assign addr[38760]= -1132798888;
assign addr[38761]= -862265664;
assign addr[38762]= -574258580;
assign addr[38763]= -274614114;
assign addr[38764]= 30595422;
assign addr[38765]= 335184940;
assign addr[38766]= 632981917;
assign addr[38767]= 917951481;
assign addr[38768]= 1184318708;
assign addr[38769]= 1426685652;
assign addr[38770]= 1640140734;
assign addr[38771]= 1820358275;
assign addr[38772]= 1963686155;
assign addr[38773]= 2067219829;
assign addr[38774]= 2128861181;
assign addr[38775]= 2147361045;
assign addr[38776]= 2122344521;
assign addr[38777]= 2054318569;
assign addr[38778]= 1944661739;
assign addr[38779]= 1795596234;
assign addr[38780]= 1610142873;
assign addr[38781]= 1392059879;
assign addr[38782]= 1145766716;
assign addr[38783]= 876254528;
assign addr[38784]= 588984994;
assign addr[38785]= 289779648;
assign addr[38786]= -15298099;
assign addr[38787]= -320065829;
assign addr[38788]= -618347408;
assign addr[38789]= -904098143;
assign addr[38790]= -1171527280;
assign addr[38791]= -1415215352;
assign addr[38792]= -1630224009;
assign addr[38793]= -1812196087;
assign addr[38794]= -1957443913;
assign addr[38795]= -2063024031;
assign addr[38796]= -2126796855;
assign addr[38797]= -2147470025;
assign addr[38798]= -2124624598;
assign addr[38799]= -2058723538;
assign addr[38800]= -1951102334;
assign addr[38801]= -1803941934;
assign addr[38802]= -1620224553;
assign addr[38803]= -1403673233;
assign addr[38804]= -1158676398;
assign addr[38805]= -890198924;
assign addr[38806]= -603681519;
assign addr[38807]= -304930476;
assign addr[38808]= 0;
assign addr[38809]= 304930476;
assign addr[38810]= 603681519;
assign addr[38811]= 890198924;
assign addr[38812]= 1158676398;
assign addr[38813]= 1403673233;
assign addr[38814]= 1620224553;
assign addr[38815]= 1803941934;
assign addr[38816]= 1951102334;
assign addr[38817]= 2058723538;
assign addr[38818]= 2124624598;
assign addr[38819]= 2147470025;
assign addr[38820]= 2126796855;
assign addr[38821]= 2063024031;
assign addr[38822]= 1957443913;
assign addr[38823]= 1812196087;
assign addr[38824]= 1630224009;
assign addr[38825]= 1415215352;
assign addr[38826]= 1171527280;
assign addr[38827]= 904098143;
assign addr[38828]= 618347408;
assign addr[38829]= 320065829;
assign addr[38830]= 15298099;
assign addr[38831]= -289779648;
assign addr[38832]= -588984994;
assign addr[38833]= -876254528;
assign addr[38834]= -1145766716;
assign addr[38835]= -1392059879;
assign addr[38836]= -1610142873;
assign addr[38837]= -1795596234;
assign addr[38838]= -1944661739;
assign addr[38839]= -2054318569;
assign addr[38840]= -2122344521;
assign addr[38841]= -2147361045;
assign addr[38842]= -2128861181;
assign addr[38843]= -2067219829;
assign addr[38844]= -1963686155;
assign addr[38845]= -1820358275;
assign addr[38846]= -1640140734;
assign addr[38847]= -1426685652;
assign addr[38848]= -1184318708;
assign addr[38849]= -917951481;
assign addr[38850]= -632981917;
assign addr[38851]= -335184940;
assign addr[38852]= -30595422;
assign addr[38853]= 274614114;
assign addr[38854]= 574258580;
assign addr[38855]= 862265664;
assign addr[38856]= 1132798888;
assign addr[38857]= 1380375881;
assign addr[38858]= 1599979481;
assign addr[38859]= 1787159411;
assign addr[38860]= 1938122457;
assign addr[38861]= 2049809346;
assign addr[38862]= 2119956737;
assign addr[38863]= 2147143090;
assign addr[38864]= 2130817471;
assign addr[38865]= 2071310720;
assign addr[38866]= 1969828744;
assign addr[38867]= 1828428082;
assign addr[38868]= 1649974225;
assign addr[38869]= 1438083551;
assign addr[38870]= 1197050035;
assign addr[38871]= 931758235;
assign addr[38872]= 647584304;
assign addr[38873]= 350287041;
assign addr[38874]= 45891193;
assign addr[38875]= -259434643;
assign addr[38876]= -559503022;
assign addr[38877]= -848233042;
assign addr[38878]= -1119773573;
assign addr[38879]= -1368621831;
assign addr[38880]= -1589734894;
assign addr[38881]= -1778631892;
assign addr[38882]= -1931484818;
assign addr[38883]= -2045196100;
assign addr[38884]= -2117461370;
assign addr[38885]= -2146816171;
assign addr[38886]= -2132665626;
assign addr[38887]= -2075296495;
assign addr[38888]= -1975871368;
assign addr[38889]= -1836405100;
assign addr[38890]= -1659723983;
assign addr[38891]= -1449408469;
assign addr[38892]= -1209720613;
assign addr[38893]= -945517704;
assign addr[38894]= -662153826;
assign addr[38895]= -365371365;
assign addr[38896]= -61184634;
assign addr[38897]= 244242007;
assign addr[38898]= 544719071;
assign addr[38899]= 834157373;
assign addr[38900]= 1106691431;
assign addr[38901]= 1356798326;
assign addr[38902]= 1579409630;
assign addr[38903]= 1770014111;
assign addr[38904]= 1924749160;
assign addr[38905]= 2040479063;
assign addr[38906]= 2114858546;
assign addr[38907]= 2146380306;
assign addr[38908]= 2134405552;
assign addr[38909]= 2079176953;
assign addr[38910]= 1981813720;
assign addr[38911]= 1844288924;
assign addr[38912]= 1669389513;
assign addr[38913]= 1460659832;
assign addr[38914]= 1222329801;
assign addr[38915]= 959229189;
assign addr[38916]= 676689746;
assign addr[38917]= 380437148;
assign addr[38918]= 76474970;
assign addr[38919]= -229036977;
assign addr[38920]= -529907477;
assign addr[38921]= -820039373;
assign addr[38922]= -1093553126;
assign addr[38923]= -1344905966;
assign addr[38924]= -1569004214;
assign addr[38925]= -1761306505;
assign addr[38926]= -1917915825;
assign addr[38927]= -2035658475;
assign addr[38928]= -2112148396;
assign addr[38929]= -2145835515;
assign addr[38930]= -2136037160;
assign addr[38931]= -2082951896;
assign addr[38932]= -1987655498;
assign addr[38933]= -1852079154;
assign addr[38934]= -1678970324;
assign addr[38935]= -1471837070;
assign addr[38936]= -1234876957;
assign addr[38937]= -972891995;
assign addr[38938]= -691191324;
assign addr[38939]= -395483624;
assign addr[38940]= -91761426;
assign addr[38941]= 213820322;
assign addr[38942]= 515068990;
assign addr[38943]= 805879757;
assign addr[38944]= 1080359326;
assign addr[38945]= 1332945355;
assign addr[38946]= 1558519173;
assign addr[38947]= 1752509516;
assign addr[38948]= 1910985158;
assign addr[38949]= 2030734582;
assign addr[38950]= 2109331059;
assign addr[38951]= 2145181827;
assign addr[38952]= 2137560369;
assign addr[38953]= 2086621133;
assign addr[38954]= 1993396407;
assign addr[38955]= 1859775393;
assign addr[38956]= 1688465931;
assign addr[38957]= 1482939614;
assign addr[38958]= 1247361445;
assign addr[38959]= 986505429;
assign addr[38960]= 705657826;
assign addr[38961]= 410510029;
assign addr[38962]= 107043224;
assign addr[38963]= -198592817;
assign addr[38964]= -500204365;
assign addr[38965]= -791679244;
assign addr[38966]= -1067110699;
assign addr[38967]= -1320917099;
assign addr[38968]= -1547955041;
assign addr[38969]= -1743623590;
assign addr[38970]= -1903957513;
assign addr[38971]= -2025707632;
assign addr[38972]= -2106406677;
assign addr[38973]= -2144419275;
assign addr[38974]= -2138975100;
assign addr[38975]= -2090184478;
assign addr[38976]= -1999036154;
assign addr[38977]= -1867377253;
assign addr[38978]= -1697875851;
assign addr[38979]= -1493966902;
assign addr[38980]= -1259782632;
assign addr[38981]= -1000068799;
assign addr[38982]= -720088517;
assign addr[38983]= -425515602;
assign addr[38984]= -122319591;
assign addr[38985]= 183355234;
assign addr[38986]= 485314355;
assign addr[38987]= 777438554;
assign addr[38988]= 1053807919;
assign addr[38989]= 1308821808;
assign addr[38990]= 1537312353;
assign addr[38991]= 1734649179;
assign addr[38992]= 1896833245;
assign addr[38993]= 2020577882;
assign addr[38994]= 2103375398;
assign addr[38995]= 2143547897;
assign addr[38996]= 2140281282;
assign addr[38997]= 2093641749;
assign addr[38998]= 2004574453;
assign addr[38999]= 1874884346;
assign addr[39000]= 1707199606;
assign addr[39001]= 1504918373;
assign addr[39002]= 1272139887;
assign addr[39003]= 1013581418;
assign addr[39004]= 734482665;
assign addr[39005]= 440499581;
assign addr[39006]= 137589750;
assign addr[39007]= -168108346;
assign addr[39008]= -470399716;
assign addr[39009]= -763158411;
assign addr[39010]= -1040451659;
assign addr[39011]= -1296660098;
assign addr[39012]= -1526591649;
assign addr[39013]= -1725586737;
assign addr[39014]= -1889612716;
assign addr[39015]= -2015345591;
assign addr[39016]= -2100237377;
assign addr[39017]= -2142567738;
assign addr[39018]= -2141478848;
assign addr[39019]= -2096992772;
assign addr[39020]= -2010011024;
assign addr[39021]= -1882296293;
assign addr[39022]= -1716436725;
assign addr[39023]= -1515793473;
assign addr[39024]= -1284432584;
assign addr[39025]= -1027042599;
assign addr[39026]= -748839539;
assign addr[39027]= -455461206;
assign addr[39028]= -152852926;
assign addr[39029]= 152852926;
assign addr[39030]= 455461206;
assign addr[39031]= 748839539;
assign addr[39032]= 1027042599;
assign addr[39033]= 1284432584;
assign addr[39034]= 1515793473;
assign addr[39035]= 1716436725;
assign addr[39036]= 1882296293;
assign addr[39037]= 2010011024;
assign addr[39038]= 2096992772;
assign addr[39039]= 2141478848;
assign addr[39040]= 2142567738;
assign addr[39041]= 2100237377;
assign addr[39042]= 2015345591;
assign addr[39043]= 1889612716;
assign addr[39044]= 1725586737;
assign addr[39045]= 1526591649;
assign addr[39046]= 1296660098;
assign addr[39047]= 1040451659;
assign addr[39048]= 763158411;
assign addr[39049]= 470399716;
assign addr[39050]= 168108346;
assign addr[39051]= -137589750;
assign addr[39052]= -440499581;
assign addr[39053]= -734482665;
assign addr[39054]= -1013581418;
assign addr[39055]= -1272139887;
assign addr[39056]= -1504918373;
assign addr[39057]= -1707199606;
assign addr[39058]= -1874884346;
assign addr[39059]= -2004574453;
assign addr[39060]= -2093641749;
assign addr[39061]= -2140281282;
assign addr[39062]= -2143547897;
assign addr[39063]= -2103375398;
assign addr[39064]= -2020577882;
assign addr[39065]= -1896833245;
assign addr[39066]= -1734649179;
assign addr[39067]= -1537312353;
assign addr[39068]= -1308821808;
assign addr[39069]= -1053807919;
assign addr[39070]= -777438554;
assign addr[39071]= -485314355;
assign addr[39072]= -183355234;
assign addr[39073]= 122319591;
assign addr[39074]= 425515602;
assign addr[39075]= 720088517;
assign addr[39076]= 1000068799;
assign addr[39077]= 1259782632;
assign addr[39078]= 1493966902;
assign addr[39079]= 1697875851;
assign addr[39080]= 1867377253;
assign addr[39081]= 1999036154;
assign addr[39082]= 2090184478;
assign addr[39083]= 2138975100;
assign addr[39084]= 2144419275;
assign addr[39085]= 2106406677;
assign addr[39086]= 2025707632;
assign addr[39087]= 1903957513;
assign addr[39088]= 1743623590;
assign addr[39089]= 1547955041;
assign addr[39090]= 1320917099;
assign addr[39091]= 1067110699;
assign addr[39092]= 791679244;
assign addr[39093]= 500204365;
assign addr[39094]= 198592817;
assign addr[39095]= -107043224;
assign addr[39096]= -410510029;
assign addr[39097]= -705657826;
assign addr[39098]= -986505429;
assign addr[39099]= -1247361445;
assign addr[39100]= -1482939614;
assign addr[39101]= -1688465931;
assign addr[39102]= -1859775393;
assign addr[39103]= -1993396407;
assign addr[39104]= -2086621133;
assign addr[39105]= -2137560369;
assign addr[39106]= -2145181827;
assign addr[39107]= -2109331059;
assign addr[39108]= -2030734582;
assign addr[39109]= -1910985158;
assign addr[39110]= -1752509516;
assign addr[39111]= -1558519173;
assign addr[39112]= -1332945355;
assign addr[39113]= -1080359326;
assign addr[39114]= -805879757;
assign addr[39115]= -515068990;
assign addr[39116]= -213820322;
assign addr[39117]= 91761426;
assign addr[39118]= 395483624;
assign addr[39119]= 691191324;
assign addr[39120]= 972891995;
assign addr[39121]= 1234876957;
assign addr[39122]= 1471837070;
assign addr[39123]= 1678970324;
assign addr[39124]= 1852079154;
assign addr[39125]= 1987655498;
assign addr[39126]= 2082951896;
assign addr[39127]= 2136037160;
assign addr[39128]= 2145835515;
assign addr[39129]= 2112148396;
assign addr[39130]= 2035658475;
assign addr[39131]= 1917915825;
assign addr[39132]= 1761306505;
assign addr[39133]= 1569004214;
assign addr[39134]= 1344905966;
assign addr[39135]= 1093553126;
assign addr[39136]= 820039373;
assign addr[39137]= 529907477;
assign addr[39138]= 229036977;
assign addr[39139]= -76474970;
assign addr[39140]= -380437148;
assign addr[39141]= -676689746;
assign addr[39142]= -959229189;
assign addr[39143]= -1222329801;
assign addr[39144]= -1460659832;
assign addr[39145]= -1669389513;
assign addr[39146]= -1844288924;
assign addr[39147]= -1981813720;
assign addr[39148]= -2079176953;
assign addr[39149]= -2134405552;
assign addr[39150]= -2146380306;
assign addr[39151]= -2114858546;
assign addr[39152]= -2040479063;
assign addr[39153]= -1924749160;
assign addr[39154]= -1770014111;
assign addr[39155]= -1579409630;
assign addr[39156]= -1356798326;
assign addr[39157]= -1106691431;
assign addr[39158]= -834157373;
assign addr[39159]= -544719071;
assign addr[39160]= -244242007;
assign addr[39161]= 61184634;
assign addr[39162]= 365371365;
assign addr[39163]= 662153826;
assign addr[39164]= 945517704;
assign addr[39165]= 1209720613;
assign addr[39166]= 1449408469;
assign addr[39167]= 1659723983;
assign addr[39168]= 1836405100;
assign addr[39169]= 1975871368;
assign addr[39170]= 2075296495;
assign addr[39171]= 2132665626;
assign addr[39172]= 2146816171;
assign addr[39173]= 2117461370;
assign addr[39174]= 2045196100;
assign addr[39175]= 1931484818;
assign addr[39176]= 1778631892;
assign addr[39177]= 1589734894;
assign addr[39178]= 1368621831;
assign addr[39179]= 1119773573;
assign addr[39180]= 848233042;
assign addr[39181]= 559503022;
assign addr[39182]= 259434643;
assign addr[39183]= -45891193;
assign addr[39184]= -350287041;
assign addr[39185]= -647584304;
assign addr[39186]= -931758235;
assign addr[39187]= -1197050035;
assign addr[39188]= -1438083551;
assign addr[39189]= -1649974225;
assign addr[39190]= -1828428082;
assign addr[39191]= -1969828744;
assign addr[39192]= -2071310720;
assign addr[39193]= -2130817471;
assign addr[39194]= -2147143090;
assign addr[39195]= -2119956737;
assign addr[39196]= -2049809346;
assign addr[39197]= -1938122457;
assign addr[39198]= -1787159411;
assign addr[39199]= -1599979481;
assign addr[39200]= -1380375881;
assign addr[39201]= -1132798888;
assign addr[39202]= -862265664;
assign addr[39203]= -574258580;
assign addr[39204]= -274614114;
assign addr[39205]= 30595422;
assign addr[39206]= 335184940;
assign addr[39207]= 632981917;
assign addr[39208]= 917951481;
assign addr[39209]= 1184318708;
assign addr[39210]= 1426685652;
assign addr[39211]= 1640140734;
assign addr[39212]= 1820358275;
assign addr[39213]= 1963686155;
assign addr[39214]= 2067219829;
assign addr[39215]= 2128861181;
assign addr[39216]= 2147361045;
assign addr[39217]= 2122344521;
assign addr[39218]= 2054318569;
assign addr[39219]= 1944661739;
assign addr[39220]= 1795596234;
assign addr[39221]= 1610142873;
assign addr[39222]= 1392059879;
assign addr[39223]= 1145766716;
assign addr[39224]= 876254528;
assign addr[39225]= 588984994;
assign addr[39226]= 289779648;
assign addr[39227]= -15298099;
assign addr[39228]= -320065829;
assign addr[39229]= -618347408;
assign addr[39230]= -904098143;
assign addr[39231]= -1171527280;
assign addr[39232]= -1415215352;
assign addr[39233]= -1630224009;
assign addr[39234]= -1812196087;
assign addr[39235]= -1957443913;
assign addr[39236]= -2063024031;
assign addr[39237]= -2126796855;
assign addr[39238]= -2147470025;
assign addr[39239]= -2124624598;
assign addr[39240]= -2058723538;
assign addr[39241]= -1951102334;
assign addr[39242]= -1803941934;
assign addr[39243]= -1620224553;
assign addr[39244]= -1403673233;
assign addr[39245]= -1158676398;
assign addr[39246]= -890198924;
assign addr[39247]= -603681519;
assign addr[39248]= -304930476;
assign addr[39249]= 0;
assign addr[39250]= 304930476;
assign addr[39251]= 603681519;
assign addr[39252]= 890198924;
assign addr[39253]= 1158676398;
assign addr[39254]= 1403673233;
assign addr[39255]= 1620224553;
assign addr[39256]= 1803941934;
assign addr[39257]= 1951102334;
assign addr[39258]= 2058723538;
assign addr[39259]= 2124624598;
assign addr[39260]= 2147470025;
assign addr[39261]= 2126796855;
assign addr[39262]= 2063024031;
assign addr[39263]= 1957443913;
assign addr[39264]= 1812196087;
assign addr[39265]= 1630224009;
assign addr[39266]= 1415215352;
assign addr[39267]= 1171527280;
assign addr[39268]= 904098143;
assign addr[39269]= 618347408;
assign addr[39270]= 320065829;
assign addr[39271]= 15298099;
assign addr[39272]= -289779648;
assign addr[39273]= -588984994;
assign addr[39274]= -876254528;
assign addr[39275]= -1145766716;
assign addr[39276]= -1392059879;
assign addr[39277]= -1610142873;
assign addr[39278]= -1795596234;
assign addr[39279]= -1944661739;
assign addr[39280]= -2054318569;
assign addr[39281]= -2122344521;
assign addr[39282]= -2147361045;
assign addr[39283]= -2128861181;
assign addr[39284]= -2067219829;
assign addr[39285]= -1963686155;
assign addr[39286]= -1820358275;
assign addr[39287]= -1640140734;
assign addr[39288]= -1426685652;
assign addr[39289]= -1184318708;
assign addr[39290]= -917951481;
assign addr[39291]= -632981917;
assign addr[39292]= -335184940;
assign addr[39293]= -30595422;
assign addr[39294]= 274614114;
assign addr[39295]= 574258580;
assign addr[39296]= 862265664;
assign addr[39297]= 1132798888;
assign addr[39298]= 1380375881;
assign addr[39299]= 1599979481;
assign addr[39300]= 1787159411;
assign addr[39301]= 1938122457;
assign addr[39302]= 2049809346;
assign addr[39303]= 2119956737;
assign addr[39304]= 2147143090;
assign addr[39305]= 2130817471;
assign addr[39306]= 2071310720;
assign addr[39307]= 1969828744;
assign addr[39308]= 1828428082;
assign addr[39309]= 1649974225;
assign addr[39310]= 1438083551;
assign addr[39311]= 1197050035;
assign addr[39312]= 931758235;
assign addr[39313]= 647584304;
assign addr[39314]= 350287041;
assign addr[39315]= 45891193;
assign addr[39316]= -259434643;
assign addr[39317]= -559503022;
assign addr[39318]= -848233042;
assign addr[39319]= -1119773573;
assign addr[39320]= -1368621831;
assign addr[39321]= -1589734894;
assign addr[39322]= -1778631892;
assign addr[39323]= -1931484818;
assign addr[39324]= -2045196100;
assign addr[39325]= -2117461370;
assign addr[39326]= -2146816171;
assign addr[39327]= -2132665626;
assign addr[39328]= -2075296495;
assign addr[39329]= -1975871368;
assign addr[39330]= -1836405100;
assign addr[39331]= -1659723983;
assign addr[39332]= -1449408469;
assign addr[39333]= -1209720613;
assign addr[39334]= -945517704;
assign addr[39335]= -662153826;
assign addr[39336]= -365371365;
assign addr[39337]= -61184634;
assign addr[39338]= 244242007;
assign addr[39339]= 544719071;
assign addr[39340]= 834157373;
assign addr[39341]= 1106691431;
assign addr[39342]= 1356798326;
assign addr[39343]= 1579409630;
assign addr[39344]= 1770014111;
assign addr[39345]= 1924749160;
assign addr[39346]= 2040479063;
assign addr[39347]= 2114858546;
assign addr[39348]= 2146380306;
assign addr[39349]= 2134405552;
assign addr[39350]= 2079176953;
assign addr[39351]= 1981813720;
assign addr[39352]= 1844288924;
assign addr[39353]= 1669389513;
assign addr[39354]= 1460659832;
assign addr[39355]= 1222329801;
assign addr[39356]= 959229189;
assign addr[39357]= 676689746;
assign addr[39358]= 380437148;
assign addr[39359]= 76474970;
assign addr[39360]= -229036977;
assign addr[39361]= -529907477;
assign addr[39362]= -820039373;
assign addr[39363]= -1093553126;
assign addr[39364]= -1344905966;
assign addr[39365]= -1569004214;
assign addr[39366]= -1761306505;
assign addr[39367]= -1917915825;
assign addr[39368]= -2035658475;
assign addr[39369]= -2112148396;
assign addr[39370]= -2145835515;
assign addr[39371]= -2136037160;
assign addr[39372]= -2082951896;
assign addr[39373]= -1987655498;
assign addr[39374]= -1852079154;
assign addr[39375]= -1678970324;
assign addr[39376]= -1471837070;
assign addr[39377]= -1234876957;
assign addr[39378]= -972891995;
assign addr[39379]= -691191324;
assign addr[39380]= -395483624;
assign addr[39381]= -91761426;
assign addr[39382]= 213820322;
assign addr[39383]= 515068990;
assign addr[39384]= 805879757;
assign addr[39385]= 1080359326;
assign addr[39386]= 1332945355;
assign addr[39387]= 1558519173;
assign addr[39388]= 1752509516;
assign addr[39389]= 1910985158;
assign addr[39390]= 2030734582;
assign addr[39391]= 2109331059;
assign addr[39392]= 2145181827;
assign addr[39393]= 2137560369;
assign addr[39394]= 2086621133;
assign addr[39395]= 1993396407;
assign addr[39396]= 1859775393;
assign addr[39397]= 1688465931;
assign addr[39398]= 1482939614;
assign addr[39399]= 1247361445;
assign addr[39400]= 986505429;
assign addr[39401]= 705657826;
assign addr[39402]= 410510029;
assign addr[39403]= 107043224;
assign addr[39404]= -198592817;
assign addr[39405]= -500204365;
assign addr[39406]= -791679244;
assign addr[39407]= -1067110699;
assign addr[39408]= -1320917099;
assign addr[39409]= -1547955041;
assign addr[39410]= -1743623590;
assign addr[39411]= -1903957513;
assign addr[39412]= -2025707632;
assign addr[39413]= -2106406677;
assign addr[39414]= -2144419275;
assign addr[39415]= -2138975100;
assign addr[39416]= -2090184478;
assign addr[39417]= -1999036154;
assign addr[39418]= -1867377253;
assign addr[39419]= -1697875851;
assign addr[39420]= -1493966902;
assign addr[39421]= -1259782632;
assign addr[39422]= -1000068799;
assign addr[39423]= -720088517;
assign addr[39424]= -425515602;
assign addr[39425]= -122319591;
assign addr[39426]= 183355234;
assign addr[39427]= 485314355;
assign addr[39428]= 777438554;
assign addr[39429]= 1053807919;
assign addr[39430]= 1308821808;
assign addr[39431]= 1537312353;
assign addr[39432]= 1734649179;
assign addr[39433]= 1896833245;
assign addr[39434]= 2020577882;
assign addr[39435]= 2103375398;
assign addr[39436]= 2143547897;
assign addr[39437]= 2140281282;
assign addr[39438]= 2093641749;
assign addr[39439]= 2004574453;
assign addr[39440]= 1874884346;
assign addr[39441]= 1707199606;
assign addr[39442]= 1504918373;
assign addr[39443]= 1272139887;
assign addr[39444]= 1013581418;
assign addr[39445]= 734482665;
assign addr[39446]= 440499581;
assign addr[39447]= 137589750;
assign addr[39448]= -168108346;
assign addr[39449]= -470399716;
assign addr[39450]= -763158411;
assign addr[39451]= -1040451659;
assign addr[39452]= -1296660098;
assign addr[39453]= -1526591649;
assign addr[39454]= -1725586737;
assign addr[39455]= -1889612716;
assign addr[39456]= -2015345591;
assign addr[39457]= -2100237377;
assign addr[39458]= -2142567738;
assign addr[39459]= -2141478848;
assign addr[39460]= -2096992772;
assign addr[39461]= -2010011024;
assign addr[39462]= -1882296293;
assign addr[39463]= -1716436725;
assign addr[39464]= -1515793473;
assign addr[39465]= -1284432584;
assign addr[39466]= -1027042599;
assign addr[39467]= -748839539;
assign addr[39468]= -455461206;
assign addr[39469]= -152852926;
assign addr[39470]= 152852926;
assign addr[39471]= 455461206;
assign addr[39472]= 748839539;
assign addr[39473]= 1027042599;
assign addr[39474]= 1284432584;
assign addr[39475]= 1515793473;
assign addr[39476]= 1716436725;
assign addr[39477]= 1882296293;
assign addr[39478]= 2010011024;
assign addr[39479]= 2096992772;
assign addr[39480]= 2141478848;
assign addr[39481]= 2142567738;
assign addr[39482]= 2100237377;
assign addr[39483]= 2015345591;
assign addr[39484]= 1889612716;
assign addr[39485]= 1725586737;
assign addr[39486]= 1526591649;
assign addr[39487]= 1296660098;
assign addr[39488]= 1040451659;
assign addr[39489]= 763158411;
assign addr[39490]= 470399716;
assign addr[39491]= 168108346;
assign addr[39492]= -137589750;
assign addr[39493]= -440499581;
assign addr[39494]= -734482665;
assign addr[39495]= -1013581418;
assign addr[39496]= -1272139887;
assign addr[39497]= -1504918373;
assign addr[39498]= -1707199606;
assign addr[39499]= -1874884346;
assign addr[39500]= -2004574453;
assign addr[39501]= -2093641749;
assign addr[39502]= -2140281282;
assign addr[39503]= -2143547897;
assign addr[39504]= -2103375398;
assign addr[39505]= -2020577882;
assign addr[39506]= -1896833245;
assign addr[39507]= -1734649179;
assign addr[39508]= -1537312353;
assign addr[39509]= -1308821808;
assign addr[39510]= -1053807919;
assign addr[39511]= -777438554;
assign addr[39512]= -485314355;
assign addr[39513]= -183355234;
assign addr[39514]= 122319591;
assign addr[39515]= 425515602;
assign addr[39516]= 720088517;
assign addr[39517]= 1000068799;
assign addr[39518]= 1259782632;
assign addr[39519]= 1493966902;
assign addr[39520]= 1697875851;
assign addr[39521]= 1867377253;
assign addr[39522]= 1999036154;
assign addr[39523]= 2090184478;
assign addr[39524]= 2138975100;
assign addr[39525]= 2144419275;
assign addr[39526]= 2106406677;
assign addr[39527]= 2025707632;
assign addr[39528]= 1903957513;
assign addr[39529]= 1743623590;
assign addr[39530]= 1547955041;
assign addr[39531]= 1320917099;
assign addr[39532]= 1067110699;
assign addr[39533]= 791679244;
assign addr[39534]= 500204365;
assign addr[39535]= 198592817;
assign addr[39536]= -107043224;
assign addr[39537]= -410510029;
assign addr[39538]= -705657826;
assign addr[39539]= -986505429;
assign addr[39540]= -1247361445;
assign addr[39541]= -1482939614;
assign addr[39542]= -1688465931;
assign addr[39543]= -1859775393;
assign addr[39544]= -1993396407;
assign addr[39545]= -2086621133;
assign addr[39546]= -2137560369;
assign addr[39547]= -2145181827;
assign addr[39548]= -2109331059;
assign addr[39549]= -2030734582;
assign addr[39550]= -1910985158;
assign addr[39551]= -1752509516;
assign addr[39552]= -1558519173;
assign addr[39553]= -1332945355;
assign addr[39554]= -1080359326;
assign addr[39555]= -805879757;
assign addr[39556]= -515068990;
assign addr[39557]= -213820322;
assign addr[39558]= 91761426;
assign addr[39559]= 395483624;
assign addr[39560]= 691191324;
assign addr[39561]= 972891995;
assign addr[39562]= 1234876957;
assign addr[39563]= 1471837070;
assign addr[39564]= 1678970324;
assign addr[39565]= 1852079154;
assign addr[39566]= 1987655498;
assign addr[39567]= 2082951896;
assign addr[39568]= 2136037160;
assign addr[39569]= 2145835515;
assign addr[39570]= 2112148396;
assign addr[39571]= 2035658475;
assign addr[39572]= 1917915825;
assign addr[39573]= 1761306505;
assign addr[39574]= 1569004214;
assign addr[39575]= 1344905966;
assign addr[39576]= 1093553126;
assign addr[39577]= 820039373;
assign addr[39578]= 529907477;
assign addr[39579]= 229036977;
assign addr[39580]= -76474970;
assign addr[39581]= -380437148;
assign addr[39582]= -676689746;
assign addr[39583]= -959229189;
assign addr[39584]= -1222329801;
assign addr[39585]= -1460659832;
assign addr[39586]= -1669389513;
assign addr[39587]= -1844288924;
assign addr[39588]= -1981813720;
assign addr[39589]= -2079176953;
assign addr[39590]= -2134405552;
assign addr[39591]= -2146380306;
assign addr[39592]= -2114858546;
assign addr[39593]= -2040479063;
assign addr[39594]= -1924749160;
assign addr[39595]= -1770014111;
assign addr[39596]= -1579409630;
assign addr[39597]= -1356798326;
assign addr[39598]= -1106691431;
assign addr[39599]= -834157373;
assign addr[39600]= -544719071;
assign addr[39601]= -244242007;
assign addr[39602]= 61184634;
assign addr[39603]= 365371365;
assign addr[39604]= 662153826;
assign addr[39605]= 945517704;
assign addr[39606]= 1209720613;
assign addr[39607]= 1449408469;
assign addr[39608]= 1659723983;
assign addr[39609]= 1836405100;
assign addr[39610]= 1975871368;
assign addr[39611]= 2075296495;
assign addr[39612]= 2132665626;
assign addr[39613]= 2146816171;
assign addr[39614]= 2117461370;
assign addr[39615]= 2045196100;
assign addr[39616]= 1931484818;
assign addr[39617]= 1778631892;
assign addr[39618]= 1589734894;
assign addr[39619]= 1368621831;
assign addr[39620]= 1119773573;
assign addr[39621]= 848233042;
assign addr[39622]= 559503022;
assign addr[39623]= 259434643;
assign addr[39624]= -45891193;
assign addr[39625]= -350287041;
assign addr[39626]= -647584304;
assign addr[39627]= -931758235;
assign addr[39628]= -1197050035;
assign addr[39629]= -1438083551;
assign addr[39630]= -1649974225;
assign addr[39631]= -1828428082;
assign addr[39632]= -1969828744;
assign addr[39633]= -2071310720;
assign addr[39634]= -2130817471;
assign addr[39635]= -2147143090;
assign addr[39636]= -2119956737;
assign addr[39637]= -2049809346;
assign addr[39638]= -1938122457;
assign addr[39639]= -1787159411;
assign addr[39640]= -1599979481;
assign addr[39641]= -1380375881;
assign addr[39642]= -1132798888;
assign addr[39643]= -862265664;
assign addr[39644]= -574258580;
assign addr[39645]= -274614114;
assign addr[39646]= 30595422;
assign addr[39647]= 335184940;
assign addr[39648]= 632981917;
assign addr[39649]= 917951481;
assign addr[39650]= 1184318708;
assign addr[39651]= 1426685652;
assign addr[39652]= 1640140734;
assign addr[39653]= 1820358275;
assign addr[39654]= 1963686155;
assign addr[39655]= 2067219829;
assign addr[39656]= 2128861181;
assign addr[39657]= 2147361045;
assign addr[39658]= 2122344521;
assign addr[39659]= 2054318569;
assign addr[39660]= 1944661739;
assign addr[39661]= 1795596234;
assign addr[39662]= 1610142873;
assign addr[39663]= 1392059879;
assign addr[39664]= 1145766716;
assign addr[39665]= 876254528;
assign addr[39666]= 588984994;
assign addr[39667]= 289779648;
assign addr[39668]= -15298099;
assign addr[39669]= -320065829;
assign addr[39670]= -618347408;
assign addr[39671]= -904098143;
assign addr[39672]= -1171527280;
assign addr[39673]= -1415215352;
assign addr[39674]= -1630224009;
assign addr[39675]= -1812196087;
assign addr[39676]= -1957443913;
assign addr[39677]= -2063024031;
assign addr[39678]= -2126796855;
assign addr[39679]= -2147470025;
assign addr[39680]= -2124624598;
assign addr[39681]= -2058723538;
assign addr[39682]= -1951102334;
assign addr[39683]= -1803941934;
assign addr[39684]= -1620224553;
assign addr[39685]= -1403673233;
assign addr[39686]= -1158676398;
assign addr[39687]= -890198924;
assign addr[39688]= -603681519;
assign addr[39689]= -304930476;
assign addr[39690]= 0;
assign addr[39691]= 304930476;
assign addr[39692]= 603681519;
assign addr[39693]= 890198924;
assign addr[39694]= 1158676398;
assign addr[39695]= 1403673233;
assign addr[39696]= 1620224553;
assign addr[39697]= 1803941934;
assign addr[39698]= 1951102334;
assign addr[39699]= 2058723538;
assign addr[39700]= 2124624598;
assign addr[39701]= 2147470025;
assign addr[39702]= 2126796855;
assign addr[39703]= 2063024031;
assign addr[39704]= 1957443913;
assign addr[39705]= 1812196087;
assign addr[39706]= 1630224009;
assign addr[39707]= 1415215352;
assign addr[39708]= 1171527280;
assign addr[39709]= 904098143;
assign addr[39710]= 618347408;
assign addr[39711]= 320065829;
assign addr[39712]= 15298099;
assign addr[39713]= -289779648;
assign addr[39714]= -588984994;
assign addr[39715]= -876254528;
assign addr[39716]= -1145766716;
assign addr[39717]= -1392059879;
assign addr[39718]= -1610142873;
assign addr[39719]= -1795596234;
assign addr[39720]= -1944661739;
assign addr[39721]= -2054318569;
assign addr[39722]= -2122344521;
assign addr[39723]= -2147361045;
assign addr[39724]= -2128861181;
assign addr[39725]= -2067219829;
assign addr[39726]= -1963686155;
assign addr[39727]= -1820358275;
assign addr[39728]= -1640140734;
assign addr[39729]= -1426685652;
assign addr[39730]= -1184318708;
assign addr[39731]= -917951481;
assign addr[39732]= -632981917;
assign addr[39733]= -335184940;
assign addr[39734]= -30595422;
assign addr[39735]= 274614114;
assign addr[39736]= 574258580;
assign addr[39737]= 862265664;
assign addr[39738]= 1132798888;
assign addr[39739]= 1380375881;
assign addr[39740]= 1599979481;
assign addr[39741]= 1787159411;
assign addr[39742]= 1938122457;
assign addr[39743]= 2049809346;
assign addr[39744]= 2119956737;
assign addr[39745]= 2147143090;
assign addr[39746]= 2130817471;
assign addr[39747]= 2071310720;
assign addr[39748]= 1969828744;
assign addr[39749]= 1828428082;
assign addr[39750]= 1649974225;
assign addr[39751]= 1438083551;
assign addr[39752]= 1197050035;
assign addr[39753]= 931758235;
assign addr[39754]= 647584304;
assign addr[39755]= 350287041;
assign addr[39756]= 45891193;
assign addr[39757]= -259434643;
assign addr[39758]= -559503022;
assign addr[39759]= -848233042;
assign addr[39760]= -1119773573;
assign addr[39761]= -1368621831;
assign addr[39762]= -1589734894;
assign addr[39763]= -1778631892;
assign addr[39764]= -1931484818;
assign addr[39765]= -2045196100;
assign addr[39766]= -2117461370;
assign addr[39767]= -2146816171;
assign addr[39768]= -2132665626;
assign addr[39769]= -2075296495;
assign addr[39770]= -1975871368;
assign addr[39771]= -1836405100;
assign addr[39772]= -1659723983;
assign addr[39773]= -1449408469;
assign addr[39774]= -1209720613;
assign addr[39775]= -945517704;
assign addr[39776]= -662153826;
assign addr[39777]= -365371365;
assign addr[39778]= -61184634;
assign addr[39779]= 244242007;
assign addr[39780]= 544719071;
assign addr[39781]= 834157373;
assign addr[39782]= 1106691431;
assign addr[39783]= 1356798326;
assign addr[39784]= 1579409630;
assign addr[39785]= 1770014111;
assign addr[39786]= 1924749160;
assign addr[39787]= 2040479063;
assign addr[39788]= 2114858546;
assign addr[39789]= 2146380306;
assign addr[39790]= 2134405552;
assign addr[39791]= 2079176953;
assign addr[39792]= 1981813720;
assign addr[39793]= 1844288924;
assign addr[39794]= 1669389513;
assign addr[39795]= 1460659832;
assign addr[39796]= 1222329801;
assign addr[39797]= 959229189;
assign addr[39798]= 676689746;
assign addr[39799]= 380437148;
assign addr[39800]= 76474970;
assign addr[39801]= -229036977;
assign addr[39802]= -529907477;
assign addr[39803]= -820039373;
assign addr[39804]= -1093553126;
assign addr[39805]= -1344905966;
assign addr[39806]= -1569004214;
assign addr[39807]= -1761306505;
assign addr[39808]= -1917915825;
assign addr[39809]= -2035658475;
assign addr[39810]= -2112148396;
assign addr[39811]= -2145835515;
assign addr[39812]= -2136037160;
assign addr[39813]= -2082951896;
assign addr[39814]= -1987655498;
assign addr[39815]= -1852079154;
assign addr[39816]= -1678970324;
assign addr[39817]= -1471837070;
assign addr[39818]= -1234876957;
assign addr[39819]= -972891995;
assign addr[39820]= -691191324;
assign addr[39821]= -395483624;
assign addr[39822]= -91761426;
assign addr[39823]= 213820322;
assign addr[39824]= 515068990;
assign addr[39825]= 805879757;
assign addr[39826]= 1080359326;
assign addr[39827]= 1332945355;
assign addr[39828]= 1558519173;
assign addr[39829]= 1752509516;
assign addr[39830]= 1910985158;
assign addr[39831]= 2030734582;
assign addr[39832]= 2109331059;
assign addr[39833]= 2145181827;
assign addr[39834]= 2137560369;
assign addr[39835]= 2086621133;
assign addr[39836]= 1993396407;
assign addr[39837]= 1859775393;
assign addr[39838]= 1688465931;
assign addr[39839]= 1482939614;
assign addr[39840]= 1247361445;
assign addr[39841]= 986505429;
assign addr[39842]= 705657826;
assign addr[39843]= 410510029;
assign addr[39844]= 107043224;
assign addr[39845]= -198592817;
assign addr[39846]= -500204365;
assign addr[39847]= -791679244;
assign addr[39848]= -1067110699;
assign addr[39849]= -1320917099;
assign addr[39850]= -1547955041;
assign addr[39851]= -1743623590;
assign addr[39852]= -1903957513;
assign addr[39853]= -2025707632;
assign addr[39854]= -2106406677;
assign addr[39855]= -2144419275;
assign addr[39856]= -2138975100;
assign addr[39857]= -2090184478;
assign addr[39858]= -1999036154;
assign addr[39859]= -1867377253;
assign addr[39860]= -1697875851;
assign addr[39861]= -1493966902;
assign addr[39862]= -1259782632;
assign addr[39863]= -1000068799;
assign addr[39864]= -720088517;
assign addr[39865]= -425515602;
assign addr[39866]= -122319591;
assign addr[39867]= 183355234;
assign addr[39868]= 485314355;
assign addr[39869]= 777438554;
assign addr[39870]= 1053807919;
assign addr[39871]= 1308821808;
assign addr[39872]= 1537312353;
assign addr[39873]= 1734649179;
assign addr[39874]= 1896833245;
assign addr[39875]= 2020577882;
assign addr[39876]= 2103375398;
assign addr[39877]= 2143547897;
assign addr[39878]= 2140281282;
assign addr[39879]= 2093641749;
assign addr[39880]= 2004574453;
assign addr[39881]= 1874884346;
assign addr[39882]= 1707199606;
assign addr[39883]= 1504918373;
assign addr[39884]= 1272139887;
assign addr[39885]= 1013581418;
assign addr[39886]= 734482665;
assign addr[39887]= 440499581;
assign addr[39888]= 137589750;
assign addr[39889]= -168108346;
assign addr[39890]= -470399716;
assign addr[39891]= -763158411;
assign addr[39892]= -1040451659;
assign addr[39893]= -1296660098;
assign addr[39894]= -1526591649;
assign addr[39895]= -1725586737;
assign addr[39896]= -1889612716;
assign addr[39897]= -2015345591;
assign addr[39898]= -2100237377;
assign addr[39899]= -2142567738;
assign addr[39900]= -2141478848;
assign addr[39901]= -2096992772;
assign addr[39902]= -2010011024;
assign addr[39903]= -1882296293;
assign addr[39904]= -1716436725;
assign addr[39905]= -1515793473;
assign addr[39906]= -1284432584;
assign addr[39907]= -1027042599;
assign addr[39908]= -748839539;
assign addr[39909]= -455461206;
assign addr[39910]= -152852926;
assign addr[39911]= 152852926;
assign addr[39912]= 455461206;
assign addr[39913]= 748839539;
assign addr[39914]= 1027042599;
assign addr[39915]= 1284432584;
assign addr[39916]= 1515793473;
assign addr[39917]= 1716436725;
assign addr[39918]= 1882296293;
assign addr[39919]= 2010011024;
assign addr[39920]= 2096992772;
assign addr[39921]= 2141478848;
assign addr[39922]= 2142567738;
assign addr[39923]= 2100237377;
assign addr[39924]= 2015345591;
assign addr[39925]= 1889612716;
assign addr[39926]= 1725586737;
assign addr[39927]= 1526591649;
assign addr[39928]= 1296660098;
assign addr[39929]= 1040451659;
assign addr[39930]= 763158411;
assign addr[39931]= 470399716;
assign addr[39932]= 168108346;
assign addr[39933]= -137589750;
assign addr[39934]= -440499581;
assign addr[39935]= -734482665;
assign addr[39936]= -1013581418;
assign addr[39937]= -1272139887;
assign addr[39938]= -1504918373;
assign addr[39939]= -1707199606;
assign addr[39940]= -1874884346;
assign addr[39941]= -2004574453;
assign addr[39942]= -2093641749;
assign addr[39943]= -2140281282;
assign addr[39944]= -2143547897;
assign addr[39945]= -2103375398;
assign addr[39946]= -2020577882;
assign addr[39947]= -1896833245;
assign addr[39948]= -1734649179;
assign addr[39949]= -1537312353;
assign addr[39950]= -1308821808;
assign addr[39951]= -1053807919;
assign addr[39952]= -777438554;
assign addr[39953]= -485314355;
assign addr[39954]= -183355234;
assign addr[39955]= 122319591;
assign addr[39956]= 425515602;
assign addr[39957]= 720088517;
assign addr[39958]= 1000068799;
assign addr[39959]= 1259782632;
assign addr[39960]= 1493966902;
assign addr[39961]= 1697875851;
assign addr[39962]= 1867377253;
assign addr[39963]= 1999036154;
assign addr[39964]= 2090184478;
assign addr[39965]= 2138975100;
assign addr[39966]= 2144419275;
assign addr[39967]= 2106406677;
assign addr[39968]= 2025707632;
assign addr[39969]= 1903957513;
assign addr[39970]= 1743623590;
assign addr[39971]= 1547955041;
assign addr[39972]= 1320917099;
assign addr[39973]= 1067110699;
assign addr[39974]= 791679244;
assign addr[39975]= 500204365;
assign addr[39976]= 198592817;
assign addr[39977]= -107043224;
assign addr[39978]= -410510029;
assign addr[39979]= -705657826;
assign addr[39980]= -986505429;
assign addr[39981]= -1247361445;
assign addr[39982]= -1482939614;
assign addr[39983]= -1688465931;
assign addr[39984]= -1859775393;
assign addr[39985]= -1993396407;
assign addr[39986]= -2086621133;
assign addr[39987]= -2137560369;
assign addr[39988]= -2145181827;
assign addr[39989]= -2109331059;
assign addr[39990]= -2030734582;
assign addr[39991]= -1910985158;
assign addr[39992]= -1752509516;
assign addr[39993]= -1558519173;
assign addr[39994]= -1332945355;
assign addr[39995]= -1080359326;
assign addr[39996]= -805879757;
assign addr[39997]= -515068990;
assign addr[39998]= -213820322;
assign addr[39999]= 91761426;
assign addr[40000]= 395483624;
assign addr[40001]= 691191324;
assign addr[40002]= 972891995;
assign addr[40003]= 1234876957;
assign addr[40004]= 1471837070;
assign addr[40005]= 1678970324;
assign addr[40006]= 1852079154;
assign addr[40007]= 1987655498;
assign addr[40008]= 2082951896;
assign addr[40009]= 2136037160;
assign addr[40010]= 2145835515;
assign addr[40011]= 2112148396;
assign addr[40012]= 2035658475;
assign addr[40013]= 1917915825;
assign addr[40014]= 1761306505;
assign addr[40015]= 1569004214;
assign addr[40016]= 1344905966;
assign addr[40017]= 1093553126;
assign addr[40018]= 820039373;
assign addr[40019]= 529907477;
assign addr[40020]= 229036977;
assign addr[40021]= -76474970;
assign addr[40022]= -380437148;
assign addr[40023]= -676689746;
assign addr[40024]= -959229189;
assign addr[40025]= -1222329801;
assign addr[40026]= -1460659832;
assign addr[40027]= -1669389513;
assign addr[40028]= -1844288924;
assign addr[40029]= -1981813720;
assign addr[40030]= -2079176953;
assign addr[40031]= -2134405552;
assign addr[40032]= -2146380306;
assign addr[40033]= -2114858546;
assign addr[40034]= -2040479063;
assign addr[40035]= -1924749160;
assign addr[40036]= -1770014111;
assign addr[40037]= -1579409630;
assign addr[40038]= -1356798326;
assign addr[40039]= -1106691431;
assign addr[40040]= -834157373;
assign addr[40041]= -544719071;
assign addr[40042]= -244242007;
assign addr[40043]= 61184634;
assign addr[40044]= 365371365;
assign addr[40045]= 662153826;
assign addr[40046]= 945517704;
assign addr[40047]= 1209720613;
assign addr[40048]= 1449408469;
assign addr[40049]= 1659723983;
assign addr[40050]= 1836405100;
assign addr[40051]= 1975871368;
assign addr[40052]= 2075296495;
assign addr[40053]= 2132665626;
assign addr[40054]= 2146816171;
assign addr[40055]= 2117461370;
assign addr[40056]= 2045196100;
assign addr[40057]= 1931484818;
assign addr[40058]= 1778631892;
assign addr[40059]= 1589734894;
assign addr[40060]= 1368621831;
assign addr[40061]= 1119773573;
assign addr[40062]= 848233042;
assign addr[40063]= 559503022;
assign addr[40064]= 259434643;
assign addr[40065]= -45891193;
assign addr[40066]= -350287041;
assign addr[40067]= -647584304;
assign addr[40068]= -931758235;
assign addr[40069]= -1197050035;
assign addr[40070]= -1438083551;
assign addr[40071]= -1649974225;
assign addr[40072]= -1828428082;
assign addr[40073]= -1969828744;
assign addr[40074]= -2071310720;
assign addr[40075]= -2130817471;
assign addr[40076]= -2147143090;
assign addr[40077]= -2119956737;
assign addr[40078]= -2049809346;
assign addr[40079]= -1938122457;
assign addr[40080]= -1787159411;
assign addr[40081]= -1599979481;
assign addr[40082]= -1380375881;
assign addr[40083]= -1132798888;
assign addr[40084]= -862265664;
assign addr[40085]= -574258580;
assign addr[40086]= -274614114;
assign addr[40087]= 30595422;
assign addr[40088]= 335184940;
assign addr[40089]= 632981917;
assign addr[40090]= 917951481;
assign addr[40091]= 1184318708;
assign addr[40092]= 1426685652;
assign addr[40093]= 1640140734;
assign addr[40094]= 1820358275;
assign addr[40095]= 1963686155;
assign addr[40096]= 2067219829;
assign addr[40097]= 2128861181;
assign addr[40098]= 2147361045;
assign addr[40099]= 2122344521;
assign addr[40100]= 2054318569;
assign addr[40101]= 1944661739;
assign addr[40102]= 1795596234;
assign addr[40103]= 1610142873;
assign addr[40104]= 1392059879;
assign addr[40105]= 1145766716;
assign addr[40106]= 876254528;
assign addr[40107]= 588984994;
assign addr[40108]= 289779648;
assign addr[40109]= -15298099;
assign addr[40110]= -320065829;
assign addr[40111]= -618347408;
assign addr[40112]= -904098143;
assign addr[40113]= -1171527280;
assign addr[40114]= -1415215352;
assign addr[40115]= -1630224009;
assign addr[40116]= -1812196087;
assign addr[40117]= -1957443913;
assign addr[40118]= -2063024031;
assign addr[40119]= -2126796855;
assign addr[40120]= -2147470025;
assign addr[40121]= -2124624598;
assign addr[40122]= -2058723538;
assign addr[40123]= -1951102334;
assign addr[40124]= -1803941934;
assign addr[40125]= -1620224553;
assign addr[40126]= -1403673233;
assign addr[40127]= -1158676398;
assign addr[40128]= -890198924;
assign addr[40129]= -603681519;
assign addr[40130]= -304930476;
assign addr[40131]= 0;
assign addr[40132]= 304930476;
assign addr[40133]= 603681519;
assign addr[40134]= 890198924;
assign addr[40135]= 1158676398;
assign addr[40136]= 1403673233;
assign addr[40137]= 1620224553;
assign addr[40138]= 1803941934;
assign addr[40139]= 1951102334;
assign addr[40140]= 2058723538;
assign addr[40141]= 2124624598;
assign addr[40142]= 2147470025;
assign addr[40143]= 2126796855;
assign addr[40144]= 2063024031;
assign addr[40145]= 1957443913;
assign addr[40146]= 1812196087;
assign addr[40147]= 1630224009;
assign addr[40148]= 1415215352;
assign addr[40149]= 1171527280;
assign addr[40150]= 904098143;
assign addr[40151]= 618347408;
assign addr[40152]= 320065829;
assign addr[40153]= 15298099;
assign addr[40154]= -289779648;
assign addr[40155]= -588984994;
assign addr[40156]= -876254528;
assign addr[40157]= -1145766716;
assign addr[40158]= -1392059879;
assign addr[40159]= -1610142873;
assign addr[40160]= -1795596234;
assign addr[40161]= -1944661739;
assign addr[40162]= -2054318569;
assign addr[40163]= -2122344521;
assign addr[40164]= -2147361045;
assign addr[40165]= -2128861181;
assign addr[40166]= -2067219829;
assign addr[40167]= -1963686155;
assign addr[40168]= -1820358275;
assign addr[40169]= -1640140734;
assign addr[40170]= -1426685652;
assign addr[40171]= -1184318708;
assign addr[40172]= -917951481;
assign addr[40173]= -632981917;
assign addr[40174]= -335184940;
assign addr[40175]= -30595422;
assign addr[40176]= 274614114;
assign addr[40177]= 574258580;
assign addr[40178]= 862265664;
assign addr[40179]= 1132798888;
assign addr[40180]= 1380375881;
assign addr[40181]= 1599979481;
assign addr[40182]= 1787159411;
assign addr[40183]= 1938122457;
assign addr[40184]= 2049809346;
assign addr[40185]= 2119956737;
assign addr[40186]= 2147143090;
assign addr[40187]= 2130817471;
assign addr[40188]= 2071310720;
assign addr[40189]= 1969828744;
assign addr[40190]= 1828428082;
assign addr[40191]= 1649974225;
assign addr[40192]= 1438083551;
assign addr[40193]= 1197050035;
assign addr[40194]= 931758235;
assign addr[40195]= 647584304;
assign addr[40196]= 350287041;
assign addr[40197]= 45891193;
assign addr[40198]= -259434643;
assign addr[40199]= -559503022;
assign addr[40200]= -848233042;
assign addr[40201]= -1119773573;
assign addr[40202]= -1368621831;
assign addr[40203]= -1589734894;
assign addr[40204]= -1778631892;
assign addr[40205]= -1931484818;
assign addr[40206]= -2045196100;
assign addr[40207]= -2117461370;
assign addr[40208]= -2146816171;
assign addr[40209]= -2132665626;
assign addr[40210]= -2075296495;
assign addr[40211]= -1975871368;
assign addr[40212]= -1836405100;
assign addr[40213]= -1659723983;
assign addr[40214]= -1449408469;
assign addr[40215]= -1209720613;
assign addr[40216]= -945517704;
assign addr[40217]= -662153826;
assign addr[40218]= -365371365;
assign addr[40219]= -61184634;
assign addr[40220]= 244242007;
assign addr[40221]= 544719071;
assign addr[40222]= 834157373;
assign addr[40223]= 1106691431;
assign addr[40224]= 1356798326;
assign addr[40225]= 1579409630;
assign addr[40226]= 1770014111;
assign addr[40227]= 1924749160;
assign addr[40228]= 2040479063;
assign addr[40229]= 2114858546;
assign addr[40230]= 2146380306;
assign addr[40231]= 2134405552;
assign addr[40232]= 2079176953;
assign addr[40233]= 1981813720;
assign addr[40234]= 1844288924;
assign addr[40235]= 1669389513;
assign addr[40236]= 1460659832;
assign addr[40237]= 1222329801;
assign addr[40238]= 959229189;
assign addr[40239]= 676689746;
assign addr[40240]= 380437148;
assign addr[40241]= 76474970;
assign addr[40242]= -229036977;
assign addr[40243]= -529907477;
assign addr[40244]= -820039373;
assign addr[40245]= -1093553126;
assign addr[40246]= -1344905966;
assign addr[40247]= -1569004214;
assign addr[40248]= -1761306505;
assign addr[40249]= -1917915825;
assign addr[40250]= -2035658475;
assign addr[40251]= -2112148396;
assign addr[40252]= -2145835515;
assign addr[40253]= -2136037160;
assign addr[40254]= -2082951896;
assign addr[40255]= -1987655498;
assign addr[40256]= -1852079154;
assign addr[40257]= -1678970324;
assign addr[40258]= -1471837070;
assign addr[40259]= -1234876957;
assign addr[40260]= -972891995;
assign addr[40261]= -691191324;
assign addr[40262]= -395483624;
assign addr[40263]= -91761426;
assign addr[40264]= 213820322;
assign addr[40265]= 515068990;
assign addr[40266]= 805879757;
assign addr[40267]= 1080359326;
assign addr[40268]= 1332945355;
assign addr[40269]= 1558519173;
assign addr[40270]= 1752509516;
assign addr[40271]= 1910985158;
assign addr[40272]= 2030734582;
assign addr[40273]= 2109331059;
assign addr[40274]= 2145181827;
assign addr[40275]= 2137560369;
assign addr[40276]= 2086621133;
assign addr[40277]= 1993396407;
assign addr[40278]= 1859775393;
assign addr[40279]= 1688465931;
assign addr[40280]= 1482939614;
assign addr[40281]= 1247361445;
assign addr[40282]= 986505429;
assign addr[40283]= 705657826;
assign addr[40284]= 410510029;
assign addr[40285]= 107043224;
assign addr[40286]= -198592817;
assign addr[40287]= -500204365;
assign addr[40288]= -791679244;
assign addr[40289]= -1067110699;
assign addr[40290]= -1320917099;
assign addr[40291]= -1547955041;
assign addr[40292]= -1743623590;
assign addr[40293]= -1903957513;
assign addr[40294]= -2025707632;
assign addr[40295]= -2106406677;
assign addr[40296]= -2144419275;
assign addr[40297]= -2138975100;
assign addr[40298]= -2090184478;
assign addr[40299]= -1999036154;
assign addr[40300]= -1867377253;
assign addr[40301]= -1697875851;
assign addr[40302]= -1493966902;
assign addr[40303]= -1259782632;
assign addr[40304]= -1000068799;
assign addr[40305]= -720088517;
assign addr[40306]= -425515602;
assign addr[40307]= -122319591;
assign addr[40308]= 183355234;
assign addr[40309]= 485314355;
assign addr[40310]= 777438554;
assign addr[40311]= 1053807919;
assign addr[40312]= 1308821808;
assign addr[40313]= 1537312353;
assign addr[40314]= 1734649179;
assign addr[40315]= 1896833245;
assign addr[40316]= 2020577882;
assign addr[40317]= 2103375398;
assign addr[40318]= 2143547897;
assign addr[40319]= 2140281282;
assign addr[40320]= 2093641749;
assign addr[40321]= 2004574453;
assign addr[40322]= 1874884346;
assign addr[40323]= 1707199606;
assign addr[40324]= 1504918373;
assign addr[40325]= 1272139887;
assign addr[40326]= 1013581418;
assign addr[40327]= 734482665;
assign addr[40328]= 440499581;
assign addr[40329]= 137589750;
assign addr[40330]= -168108346;
assign addr[40331]= -470399716;
assign addr[40332]= -763158411;
assign addr[40333]= -1040451659;
assign addr[40334]= -1296660098;
assign addr[40335]= -1526591649;
assign addr[40336]= -1725586737;
assign addr[40337]= -1889612716;
assign addr[40338]= -2015345591;
assign addr[40339]= -2100237377;
assign addr[40340]= -2142567738;
assign addr[40341]= -2141478848;
assign addr[40342]= -2096992772;
assign addr[40343]= -2010011024;
assign addr[40344]= -1882296293;
assign addr[40345]= -1716436725;
assign addr[40346]= -1515793473;
assign addr[40347]= -1284432584;
assign addr[40348]= -1027042599;
assign addr[40349]= -748839539;
assign addr[40350]= -455461206;
assign addr[40351]= -152852926;
assign addr[40352]= 152852926;
assign addr[40353]= 455461206;
assign addr[40354]= 748839539;
assign addr[40355]= 1027042599;
assign addr[40356]= 1284432584;
assign addr[40357]= 1515793473;
assign addr[40358]= 1716436725;
assign addr[40359]= 1882296293;
assign addr[40360]= 2010011024;
assign addr[40361]= 2096992772;
assign addr[40362]= 2141478848;
assign addr[40363]= 2142567738;
assign addr[40364]= 2100237377;
assign addr[40365]= 2015345591;
assign addr[40366]= 1889612716;
assign addr[40367]= 1725586737;
assign addr[40368]= 1526591649;
assign addr[40369]= 1296660098;
assign addr[40370]= 1040451659;
assign addr[40371]= 763158411;
assign addr[40372]= 470399716;
assign addr[40373]= 168108346;
assign addr[40374]= -137589750;
assign addr[40375]= -440499581;
assign addr[40376]= -734482665;
assign addr[40377]= -1013581418;
assign addr[40378]= -1272139887;
assign addr[40379]= -1504918373;
assign addr[40380]= -1707199606;
assign addr[40381]= -1874884346;
assign addr[40382]= -2004574453;
assign addr[40383]= -2093641749;
assign addr[40384]= -2140281282;
assign addr[40385]= -2143547897;
assign addr[40386]= -2103375398;
assign addr[40387]= -2020577882;
assign addr[40388]= -1896833245;
assign addr[40389]= -1734649179;
assign addr[40390]= -1537312353;
assign addr[40391]= -1308821808;
assign addr[40392]= -1053807919;
assign addr[40393]= -777438554;
assign addr[40394]= -485314355;
assign addr[40395]= -183355234;
assign addr[40396]= 122319591;
assign addr[40397]= 425515602;
assign addr[40398]= 720088517;
assign addr[40399]= 1000068799;
assign addr[40400]= 1259782632;
assign addr[40401]= 1493966902;
assign addr[40402]= 1697875851;
assign addr[40403]= 1867377253;
assign addr[40404]= 1999036154;
assign addr[40405]= 2090184478;
assign addr[40406]= 2138975100;
assign addr[40407]= 2144419275;
assign addr[40408]= 2106406677;
assign addr[40409]= 2025707632;
assign addr[40410]= 1903957513;
assign addr[40411]= 1743623590;
assign addr[40412]= 1547955041;
assign addr[40413]= 1320917099;
assign addr[40414]= 1067110699;
assign addr[40415]= 791679244;
assign addr[40416]= 500204365;
assign addr[40417]= 198592817;
assign addr[40418]= -107043224;
assign addr[40419]= -410510029;
assign addr[40420]= -705657826;
assign addr[40421]= -986505429;
assign addr[40422]= -1247361445;
assign addr[40423]= -1482939614;
assign addr[40424]= -1688465931;
assign addr[40425]= -1859775393;
assign addr[40426]= -1993396407;
assign addr[40427]= -2086621133;
assign addr[40428]= -2137560369;
assign addr[40429]= -2145181827;
assign addr[40430]= -2109331059;
assign addr[40431]= -2030734582;
assign addr[40432]= -1910985158;
assign addr[40433]= -1752509516;
assign addr[40434]= -1558519173;
assign addr[40435]= -1332945355;
assign addr[40436]= -1080359326;
assign addr[40437]= -805879757;
assign addr[40438]= -515068990;
assign addr[40439]= -213820322;
assign addr[40440]= 91761426;
assign addr[40441]= 395483624;
assign addr[40442]= 691191324;
assign addr[40443]= 972891995;
assign addr[40444]= 1234876957;
assign addr[40445]= 1471837070;
assign addr[40446]= 1678970324;
assign addr[40447]= 1852079154;
assign addr[40448]= 1987655498;
assign addr[40449]= 2082951896;
assign addr[40450]= 2136037160;
assign addr[40451]= 2145835515;
assign addr[40452]= 2112148396;
assign addr[40453]= 2035658475;
assign addr[40454]= 1917915825;
assign addr[40455]= 1761306505;
assign addr[40456]= 1569004214;
assign addr[40457]= 1344905966;
assign addr[40458]= 1093553126;
assign addr[40459]= 820039373;
assign addr[40460]= 529907477;
assign addr[40461]= 229036977;
assign addr[40462]= -76474970;
assign addr[40463]= -380437148;
assign addr[40464]= -676689746;
assign addr[40465]= -959229189;
assign addr[40466]= -1222329801;
assign addr[40467]= -1460659832;
assign addr[40468]= -1669389513;
assign addr[40469]= -1844288924;
assign addr[40470]= -1981813720;
assign addr[40471]= -2079176953;
assign addr[40472]= -2134405552;
assign addr[40473]= -2146380306;
assign addr[40474]= -2114858546;
assign addr[40475]= -2040479063;
assign addr[40476]= -1924749160;
assign addr[40477]= -1770014111;
assign addr[40478]= -1579409630;
assign addr[40479]= -1356798326;
assign addr[40480]= -1106691431;
assign addr[40481]= -834157373;
assign addr[40482]= -544719071;
assign addr[40483]= -244242007;
assign addr[40484]= 61184634;
assign addr[40485]= 365371365;
assign addr[40486]= 662153826;
assign addr[40487]= 945517704;
assign addr[40488]= 1209720613;
assign addr[40489]= 1449408469;
assign addr[40490]= 1659723983;
assign addr[40491]= 1836405100;
assign addr[40492]= 1975871368;
assign addr[40493]= 2075296495;
assign addr[40494]= 2132665626;
assign addr[40495]= 2146816171;
assign addr[40496]= 2117461370;
assign addr[40497]= 2045196100;
assign addr[40498]= 1931484818;
assign addr[40499]= 1778631892;
assign addr[40500]= 1589734894;
assign addr[40501]= 1368621831;
assign addr[40502]= 1119773573;
assign addr[40503]= 848233042;
assign addr[40504]= 559503022;
assign addr[40505]= 259434643;
assign addr[40506]= -45891193;
assign addr[40507]= -350287041;
assign addr[40508]= -647584304;
assign addr[40509]= -931758235;
assign addr[40510]= -1197050035;
assign addr[40511]= -1438083551;
assign addr[40512]= -1649974225;
assign addr[40513]= -1828428082;
assign addr[40514]= -1969828744;
assign addr[40515]= -2071310720;
assign addr[40516]= -2130817471;
assign addr[40517]= -2147143090;
assign addr[40518]= -2119956737;
assign addr[40519]= -2049809346;
assign addr[40520]= -1938122457;
assign addr[40521]= -1787159411;
assign addr[40522]= -1599979481;
assign addr[40523]= -1380375881;
assign addr[40524]= -1132798888;
assign addr[40525]= -862265664;
assign addr[40526]= -574258580;
assign addr[40527]= -274614114;
assign addr[40528]= 30595422;
assign addr[40529]= 335184940;
assign addr[40530]= 632981917;
assign addr[40531]= 917951481;
assign addr[40532]= 1184318708;
assign addr[40533]= 1426685652;
assign addr[40534]= 1640140734;
assign addr[40535]= 1820358275;
assign addr[40536]= 1963686155;
assign addr[40537]= 2067219829;
assign addr[40538]= 2128861181;
assign addr[40539]= 2147361045;
assign addr[40540]= 2122344521;
assign addr[40541]= 2054318569;
assign addr[40542]= 1944661739;
assign addr[40543]= 1795596234;
assign addr[40544]= 1610142873;
assign addr[40545]= 1392059879;
assign addr[40546]= 1145766716;
assign addr[40547]= 876254528;
assign addr[40548]= 588984994;
assign addr[40549]= 289779648;
assign addr[40550]= -15298099;
assign addr[40551]= -320065829;
assign addr[40552]= -618347408;
assign addr[40553]= -904098143;
assign addr[40554]= -1171527280;
assign addr[40555]= -1415215352;
assign addr[40556]= -1630224009;
assign addr[40557]= -1812196087;
assign addr[40558]= -1957443913;
assign addr[40559]= -2063024031;
assign addr[40560]= -2126796855;
assign addr[40561]= -2147470025;
assign addr[40562]= -2124624598;
assign addr[40563]= -2058723538;
assign addr[40564]= -1951102334;
assign addr[40565]= -1803941934;
assign addr[40566]= -1620224553;
assign addr[40567]= -1403673233;
assign addr[40568]= -1158676398;
assign addr[40569]= -890198924;
assign addr[40570]= -603681519;
assign addr[40571]= -304930476;
assign addr[40572]= 0;
assign addr[40573]= 304930476;
assign addr[40574]= 603681519;
assign addr[40575]= 890198924;
assign addr[40576]= 1158676398;
assign addr[40577]= 1403673233;
assign addr[40578]= 1620224553;
assign addr[40579]= 1803941934;
assign addr[40580]= 1951102334;
assign addr[40581]= 2058723538;
assign addr[40582]= 2124624598;
assign addr[40583]= 2147470025;
assign addr[40584]= 2126796855;
assign addr[40585]= 2063024031;
assign addr[40586]= 1957443913;
assign addr[40587]= 1812196087;
assign addr[40588]= 1630224009;
assign addr[40589]= 1415215352;
assign addr[40590]= 1171527280;
assign addr[40591]= 904098143;
assign addr[40592]= 618347408;
assign addr[40593]= 320065829;
assign addr[40594]= 15298099;
assign addr[40595]= -289779648;
assign addr[40596]= -588984994;
assign addr[40597]= -876254528;
assign addr[40598]= -1145766716;
assign addr[40599]= -1392059879;
assign addr[40600]= -1610142873;
assign addr[40601]= -1795596234;
assign addr[40602]= -1944661739;
assign addr[40603]= -2054318569;
assign addr[40604]= -2122344521;
assign addr[40605]= -2147361045;
assign addr[40606]= -2128861181;
assign addr[40607]= -2067219829;
assign addr[40608]= -1963686155;
assign addr[40609]= -1820358275;
assign addr[40610]= -1640140734;
assign addr[40611]= -1426685652;
assign addr[40612]= -1184318708;
assign addr[40613]= -917951481;
assign addr[40614]= -632981917;
assign addr[40615]= -335184940;
assign addr[40616]= -30595422;
assign addr[40617]= 274614114;
assign addr[40618]= 574258580;
assign addr[40619]= 862265664;
assign addr[40620]= 1132798888;
assign addr[40621]= 1380375881;
assign addr[40622]= 1599979481;
assign addr[40623]= 1787159411;
assign addr[40624]= 1938122457;
assign addr[40625]= 2049809346;
assign addr[40626]= 2119956737;
assign addr[40627]= 2147143090;
assign addr[40628]= 2130817471;
assign addr[40629]= 2071310720;
assign addr[40630]= 1969828744;
assign addr[40631]= 1828428082;
assign addr[40632]= 1649974225;
assign addr[40633]= 1438083551;
assign addr[40634]= 1197050035;
assign addr[40635]= 931758235;
assign addr[40636]= 647584304;
assign addr[40637]= 350287041;
assign addr[40638]= 45891193;
assign addr[40639]= -259434643;
assign addr[40640]= -559503022;
assign addr[40641]= -848233042;
assign addr[40642]= -1119773573;
assign addr[40643]= -1368621831;
assign addr[40644]= -1589734894;
assign addr[40645]= -1778631892;
assign addr[40646]= -1931484818;
assign addr[40647]= -2045196100;
assign addr[40648]= -2117461370;
assign addr[40649]= -2146816171;
assign addr[40650]= -2132665626;
assign addr[40651]= -2075296495;
assign addr[40652]= -1975871368;
assign addr[40653]= -1836405100;
assign addr[40654]= -1659723983;
assign addr[40655]= -1449408469;
assign addr[40656]= -1209720613;
assign addr[40657]= -945517704;
assign addr[40658]= -662153826;
assign addr[40659]= -365371365;
assign addr[40660]= -61184634;
assign addr[40661]= 244242007;
assign addr[40662]= 544719071;
assign addr[40663]= 834157373;
assign addr[40664]= 1106691431;
assign addr[40665]= 1356798326;
assign addr[40666]= 1579409630;
assign addr[40667]= 1770014111;
assign addr[40668]= 1924749160;
assign addr[40669]= 2040479063;
assign addr[40670]= 2114858546;
assign addr[40671]= 2146380306;
assign addr[40672]= 2134405552;
assign addr[40673]= 2079176953;
assign addr[40674]= 1981813720;
assign addr[40675]= 1844288924;
assign addr[40676]= 1669389513;
assign addr[40677]= 1460659832;
assign addr[40678]= 1222329801;
assign addr[40679]= 959229189;
assign addr[40680]= 676689746;
assign addr[40681]= 380437148;
assign addr[40682]= 76474970;
assign addr[40683]= -229036977;
assign addr[40684]= -529907477;
assign addr[40685]= -820039373;
assign addr[40686]= -1093553126;
assign addr[40687]= -1344905966;
assign addr[40688]= -1569004214;
assign addr[40689]= -1761306505;
assign addr[40690]= -1917915825;
assign addr[40691]= -2035658475;
assign addr[40692]= -2112148396;
assign addr[40693]= -2145835515;
assign addr[40694]= -2136037160;
assign addr[40695]= -2082951896;
assign addr[40696]= -1987655498;
assign addr[40697]= -1852079154;
assign addr[40698]= -1678970324;
assign addr[40699]= -1471837070;
assign addr[40700]= -1234876957;
assign addr[40701]= -972891995;
assign addr[40702]= -691191324;
assign addr[40703]= -395483624;
assign addr[40704]= -91761426;
assign addr[40705]= 213820322;
assign addr[40706]= 515068990;
assign addr[40707]= 805879757;
assign addr[40708]= 1080359326;
assign addr[40709]= 1332945355;
assign addr[40710]= 1558519173;
assign addr[40711]= 1752509516;
assign addr[40712]= 1910985158;
assign addr[40713]= 2030734582;
assign addr[40714]= 2109331059;
assign addr[40715]= 2145181827;
assign addr[40716]= 2137560369;
assign addr[40717]= 2086621133;
assign addr[40718]= 1993396407;
assign addr[40719]= 1859775393;
assign addr[40720]= 1688465931;
assign addr[40721]= 1482939614;
assign addr[40722]= 1247361445;
assign addr[40723]= 986505429;
assign addr[40724]= 705657826;
assign addr[40725]= 410510029;
assign addr[40726]= 107043224;
assign addr[40727]= -198592817;
assign addr[40728]= -500204365;
assign addr[40729]= -791679244;
assign addr[40730]= -1067110699;
assign addr[40731]= -1320917099;
assign addr[40732]= -1547955041;
assign addr[40733]= -1743623590;
assign addr[40734]= -1903957513;
assign addr[40735]= -2025707632;
assign addr[40736]= -2106406677;
assign addr[40737]= -2144419275;
assign addr[40738]= -2138975100;
assign addr[40739]= -2090184478;
assign addr[40740]= -1999036154;
assign addr[40741]= -1867377253;
assign addr[40742]= -1697875851;
assign addr[40743]= -1493966902;
assign addr[40744]= -1259782632;
assign addr[40745]= -1000068799;
assign addr[40746]= -720088517;
assign addr[40747]= -425515602;
assign addr[40748]= -122319591;
assign addr[40749]= 183355234;
assign addr[40750]= 485314355;
assign addr[40751]= 777438554;
assign addr[40752]= 1053807919;
assign addr[40753]= 1308821808;
assign addr[40754]= 1537312353;
assign addr[40755]= 1734649179;
assign addr[40756]= 1896833245;
assign addr[40757]= 2020577882;
assign addr[40758]= 2103375398;
assign addr[40759]= 2143547897;
assign addr[40760]= 2140281282;
assign addr[40761]= 2093641749;
assign addr[40762]= 2004574453;
assign addr[40763]= 1874884346;
assign addr[40764]= 1707199606;
assign addr[40765]= 1504918373;
assign addr[40766]= 1272139887;
assign addr[40767]= 1013581418;
assign addr[40768]= 734482665;
assign addr[40769]= 440499581;
assign addr[40770]= 137589750;
assign addr[40771]= -168108346;
assign addr[40772]= -470399716;
assign addr[40773]= -763158411;
assign addr[40774]= -1040451659;
assign addr[40775]= -1296660098;
assign addr[40776]= -1526591649;
assign addr[40777]= -1725586737;
assign addr[40778]= -1889612716;
assign addr[40779]= -2015345591;
assign addr[40780]= -2100237377;
assign addr[40781]= -2142567738;
assign addr[40782]= -2141478848;
assign addr[40783]= -2096992772;
assign addr[40784]= -2010011024;
assign addr[40785]= -1882296293;
assign addr[40786]= -1716436725;
assign addr[40787]= -1515793473;
assign addr[40788]= -1284432584;
assign addr[40789]= -1027042599;
assign addr[40790]= -748839539;
assign addr[40791]= -455461206;
assign addr[40792]= -152852926;
assign addr[40793]= 152852926;
assign addr[40794]= 455461206;
assign addr[40795]= 748839539;
assign addr[40796]= 1027042599;
assign addr[40797]= 1284432584;
assign addr[40798]= 1515793473;
assign addr[40799]= 1716436725;
assign addr[40800]= 1882296293;
assign addr[40801]= 2010011024;
assign addr[40802]= 2096992772;
assign addr[40803]= 2141478848;
assign addr[40804]= 2142567738;
assign addr[40805]= 2100237377;
assign addr[40806]= 2015345591;
assign addr[40807]= 1889612716;
assign addr[40808]= 1725586737;
assign addr[40809]= 1526591649;
assign addr[40810]= 1296660098;
assign addr[40811]= 1040451659;
assign addr[40812]= 763158411;
assign addr[40813]= 470399716;
assign addr[40814]= 168108346;
assign addr[40815]= -137589750;
assign addr[40816]= -440499581;
assign addr[40817]= -734482665;
assign addr[40818]= -1013581418;
assign addr[40819]= -1272139887;
assign addr[40820]= -1504918373;
assign addr[40821]= -1707199606;
assign addr[40822]= -1874884346;
assign addr[40823]= -2004574453;
assign addr[40824]= -2093641749;
assign addr[40825]= -2140281282;
assign addr[40826]= -2143547897;
assign addr[40827]= -2103375398;
assign addr[40828]= -2020577882;
assign addr[40829]= -1896833245;
assign addr[40830]= -1734649179;
assign addr[40831]= -1537312353;
assign addr[40832]= -1308821808;
assign addr[40833]= -1053807919;
assign addr[40834]= -777438554;
assign addr[40835]= -485314355;
assign addr[40836]= -183355234;
assign addr[40837]= 122319591;
assign addr[40838]= 425515602;
assign addr[40839]= 720088517;
assign addr[40840]= 1000068799;
assign addr[40841]= 1259782632;
assign addr[40842]= 1493966902;
assign addr[40843]= 1697875851;
assign addr[40844]= 1867377253;
assign addr[40845]= 1999036154;
assign addr[40846]= 2090184478;
assign addr[40847]= 2138975100;
assign addr[40848]= 2144419275;
assign addr[40849]= 2106406677;
assign addr[40850]= 2025707632;
assign addr[40851]= 1903957513;
assign addr[40852]= 1743623590;
assign addr[40853]= 1547955041;
assign addr[40854]= 1320917099;
assign addr[40855]= 1067110699;
assign addr[40856]= 791679244;
assign addr[40857]= 500204365;
assign addr[40858]= 198592817;
assign addr[40859]= -107043224;
assign addr[40860]= -410510029;
assign addr[40861]= -705657826;
assign addr[40862]= -986505429;
assign addr[40863]= -1247361445;
assign addr[40864]= -1482939614;
assign addr[40865]= -1688465931;
assign addr[40866]= -1859775393;
assign addr[40867]= -1993396407;
assign addr[40868]= -2086621133;
assign addr[40869]= -2137560369;
assign addr[40870]= -2145181827;
assign addr[40871]= -2109331059;
assign addr[40872]= -2030734582;
assign addr[40873]= -1910985158;
assign addr[40874]= -1752509516;
assign addr[40875]= -1558519173;
assign addr[40876]= -1332945355;
assign addr[40877]= -1080359326;
assign addr[40878]= -805879757;
assign addr[40879]= -515068990;
assign addr[40880]= -213820322;
assign addr[40881]= 91761426;
assign addr[40882]= 395483624;
assign addr[40883]= 691191324;
assign addr[40884]= 972891995;
assign addr[40885]= 1234876957;
assign addr[40886]= 1471837070;
assign addr[40887]= 1678970324;
assign addr[40888]= 1852079154;
assign addr[40889]= 1987655498;
assign addr[40890]= 2082951896;
assign addr[40891]= 2136037160;
assign addr[40892]= 2145835515;
assign addr[40893]= 2112148396;
assign addr[40894]= 2035658475;
assign addr[40895]= 1917915825;
assign addr[40896]= 1761306505;
assign addr[40897]= 1569004214;
assign addr[40898]= 1344905966;
assign addr[40899]= 1093553126;
assign addr[40900]= 820039373;
assign addr[40901]= 529907477;
assign addr[40902]= 229036977;
assign addr[40903]= -76474970;
assign addr[40904]= -380437148;
assign addr[40905]= -676689746;
assign addr[40906]= -959229189;
assign addr[40907]= -1222329801;
assign addr[40908]= -1460659832;
assign addr[40909]= -1669389513;
assign addr[40910]= -1844288924;
assign addr[40911]= -1981813720;
assign addr[40912]= -2079176953;
assign addr[40913]= -2134405552;
assign addr[40914]= -2146380306;
assign addr[40915]= -2114858546;
assign addr[40916]= -2040479063;
assign addr[40917]= -1924749160;
assign addr[40918]= -1770014111;
assign addr[40919]= -1579409630;
assign addr[40920]= -1356798326;
assign addr[40921]= -1106691431;
assign addr[40922]= -834157373;
assign addr[40923]= -544719071;
assign addr[40924]= -244242007;
assign addr[40925]= 61184634;
assign addr[40926]= 365371365;
assign addr[40927]= 662153826;
assign addr[40928]= 945517704;
assign addr[40929]= 1209720613;
assign addr[40930]= 1449408469;
assign addr[40931]= 1659723983;
assign addr[40932]= 1836405100;
assign addr[40933]= 1975871368;
assign addr[40934]= 2075296495;
assign addr[40935]= 2132665626;
assign addr[40936]= 2146816171;
assign addr[40937]= 2117461370;
assign addr[40938]= 2045196100;
assign addr[40939]= 1931484818;
assign addr[40940]= 1778631892;
assign addr[40941]= 1589734894;
assign addr[40942]= 1368621831;
assign addr[40943]= 1119773573;
assign addr[40944]= 848233042;
assign addr[40945]= 559503022;
assign addr[40946]= 259434643;
assign addr[40947]= -45891193;
assign addr[40948]= -350287041;
assign addr[40949]= -647584304;
assign addr[40950]= -931758235;
assign addr[40951]= -1197050035;
assign addr[40952]= -1438083551;
assign addr[40953]= -1649974225;
assign addr[40954]= -1828428082;
assign addr[40955]= -1969828744;
assign addr[40956]= -2071310720;
assign addr[40957]= -2130817471;
assign addr[40958]= -2147143090;
assign addr[40959]= -2119956737;
assign addr[40960]= -2049809346;
assign addr[40961]= -1938122457;
assign addr[40962]= -1787159411;
assign addr[40963]= -1599979481;
assign addr[40964]= -1380375881;
assign addr[40965]= -1132798888;
assign addr[40966]= -862265664;
assign addr[40967]= -574258580;
assign addr[40968]= -274614114;
assign addr[40969]= 30595422;
assign addr[40970]= 335184940;
assign addr[40971]= 632981917;
assign addr[40972]= 917951481;
assign addr[40973]= 1184318708;
assign addr[40974]= 1426685652;
assign addr[40975]= 1640140734;
assign addr[40976]= 1820358275;
assign addr[40977]= 1963686155;
assign addr[40978]= 2067219829;
assign addr[40979]= 2128861181;
assign addr[40980]= 2147361045;
assign addr[40981]= 2122344521;
assign addr[40982]= 2054318569;
assign addr[40983]= 1944661739;
assign addr[40984]= 1795596234;
assign addr[40985]= 1610142873;
assign addr[40986]= 1392059879;
assign addr[40987]= 1145766716;
assign addr[40988]= 876254528;
assign addr[40989]= 588984994;
assign addr[40990]= 289779648;
assign addr[40991]= -15298099;
assign addr[40992]= -320065829;
assign addr[40993]= -618347408;
assign addr[40994]= -904098143;
assign addr[40995]= -1171527280;
assign addr[40996]= -1415215352;
assign addr[40997]= -1630224009;
assign addr[40998]= -1812196087;
assign addr[40999]= -1957443913;
assign addr[41000]= -2063024031;
assign addr[41001]= -2126796855;
assign addr[41002]= -2147470025;
assign addr[41003]= -2124624598;
assign addr[41004]= -2058723538;
assign addr[41005]= -1951102334;
assign addr[41006]= -1803941934;
assign addr[41007]= -1620224553;
assign addr[41008]= -1403673233;
assign addr[41009]= -1158676398;
assign addr[41010]= -890198924;
assign addr[41011]= -603681519;
assign addr[41012]= -304930476;
assign addr[41013]= 0;
assign addr[41014]= 304930476;
assign addr[41015]= 603681519;
assign addr[41016]= 890198924;
assign addr[41017]= 1158676398;
assign addr[41018]= 1403673233;
assign addr[41019]= 1620224553;
assign addr[41020]= 1803941934;
assign addr[41021]= 1951102334;
assign addr[41022]= 2058723538;
assign addr[41023]= 2124624598;
assign addr[41024]= 2147470025;
assign addr[41025]= 2126796855;
assign addr[41026]= 2063024031;
assign addr[41027]= 1957443913;
assign addr[41028]= 1812196087;
assign addr[41029]= 1630224009;
assign addr[41030]= 1415215352;
assign addr[41031]= 1171527280;
assign addr[41032]= 904098143;
assign addr[41033]= 618347408;
assign addr[41034]= 320065829;
assign addr[41035]= 15298099;
assign addr[41036]= -289779648;
assign addr[41037]= -588984994;
assign addr[41038]= -876254528;
assign addr[41039]= -1145766716;
assign addr[41040]= -1392059879;
assign addr[41041]= -1610142873;
assign addr[41042]= -1795596234;
assign addr[41043]= -1944661739;
assign addr[41044]= -2054318569;
assign addr[41045]= -2122344521;
assign addr[41046]= -2147361045;
assign addr[41047]= -2128861181;
assign addr[41048]= -2067219829;
assign addr[41049]= -1963686155;
assign addr[41050]= -1820358275;
assign addr[41051]= -1640140734;
assign addr[41052]= -1426685652;
assign addr[41053]= -1184318708;
assign addr[41054]= -917951481;
assign addr[41055]= -632981917;
assign addr[41056]= -335184940;
assign addr[41057]= -30595422;
assign addr[41058]= 274614114;
assign addr[41059]= 574258580;
assign addr[41060]= 862265664;
assign addr[41061]= 1132798888;
assign addr[41062]= 1380375881;
assign addr[41063]= 1599979481;
assign addr[41064]= 1787159411;
assign addr[41065]= 1938122457;
assign addr[41066]= 2049809346;
assign addr[41067]= 2119956737;
assign addr[41068]= 2147143090;
assign addr[41069]= 2130817471;
assign addr[41070]= 2071310720;
assign addr[41071]= 1969828744;
assign addr[41072]= 1828428082;
assign addr[41073]= 1649974225;
assign addr[41074]= 1438083551;
assign addr[41075]= 1197050035;
assign addr[41076]= 931758235;
assign addr[41077]= 647584304;
assign addr[41078]= 350287041;
assign addr[41079]= 45891193;
assign addr[41080]= -259434643;
assign addr[41081]= -559503022;
assign addr[41082]= -848233042;
assign addr[41083]= -1119773573;
assign addr[41084]= -1368621831;
assign addr[41085]= -1589734894;
assign addr[41086]= -1778631892;
assign addr[41087]= -1931484818;
assign addr[41088]= -2045196100;
assign addr[41089]= -2117461370;
assign addr[41090]= -2146816171;
assign addr[41091]= -2132665626;
assign addr[41092]= -2075296495;
assign addr[41093]= -1975871368;
assign addr[41094]= -1836405100;
assign addr[41095]= -1659723983;
assign addr[41096]= -1449408469;
assign addr[41097]= -1209720613;
assign addr[41098]= -945517704;
assign addr[41099]= -662153826;
assign addr[41100]= -365371365;
assign addr[41101]= -61184634;
assign addr[41102]= 244242007;
assign addr[41103]= 544719071;
assign addr[41104]= 834157373;
assign addr[41105]= 1106691431;
assign addr[41106]= 1356798326;
assign addr[41107]= 1579409630;
assign addr[41108]= 1770014111;
assign addr[41109]= 1924749160;
assign addr[41110]= 2040479063;
assign addr[41111]= 2114858546;
assign addr[41112]= 2146380306;
assign addr[41113]= 2134405552;
assign addr[41114]= 2079176953;
assign addr[41115]= 1981813720;
assign addr[41116]= 1844288924;
assign addr[41117]= 1669389513;
assign addr[41118]= 1460659832;
assign addr[41119]= 1222329801;
assign addr[41120]= 959229189;
assign addr[41121]= 676689746;
assign addr[41122]= 380437148;
assign addr[41123]= 76474970;
assign addr[41124]= -229036977;
assign addr[41125]= -529907477;
assign addr[41126]= -820039373;
assign addr[41127]= -1093553126;
assign addr[41128]= -1344905966;
assign addr[41129]= -1569004214;
assign addr[41130]= -1761306505;
assign addr[41131]= -1917915825;
assign addr[41132]= -2035658475;
assign addr[41133]= -2112148396;
assign addr[41134]= -2145835515;
assign addr[41135]= -2136037160;
assign addr[41136]= -2082951896;
assign addr[41137]= -1987655498;
assign addr[41138]= -1852079154;
assign addr[41139]= -1678970324;
assign addr[41140]= -1471837070;
assign addr[41141]= -1234876957;
assign addr[41142]= -972891995;
assign addr[41143]= -691191324;
assign addr[41144]= -395483624;
assign addr[41145]= -91761426;
assign addr[41146]= 213820322;
assign addr[41147]= 515068990;
assign addr[41148]= 805879757;
assign addr[41149]= 1080359326;
assign addr[41150]= 1332945355;
assign addr[41151]= 1558519173;
assign addr[41152]= 1752509516;
assign addr[41153]= 1910985158;
assign addr[41154]= 2030734582;
assign addr[41155]= 2109331059;
assign addr[41156]= 2145181827;
assign addr[41157]= 2137560369;
assign addr[41158]= 2086621133;
assign addr[41159]= 1993396407;
assign addr[41160]= 1859775393;
assign addr[41161]= 1688465931;
assign addr[41162]= 1482939614;
assign addr[41163]= 1247361445;
assign addr[41164]= 986505429;
assign addr[41165]= 705657826;
assign addr[41166]= 410510029;
assign addr[41167]= 107043224;
assign addr[41168]= -198592817;
assign addr[41169]= -500204365;
assign addr[41170]= -791679244;
assign addr[41171]= -1067110699;
assign addr[41172]= -1320917099;
assign addr[41173]= -1547955041;
assign addr[41174]= -1743623590;
assign addr[41175]= -1903957513;
assign addr[41176]= -2025707632;
assign addr[41177]= -2106406677;
assign addr[41178]= -2144419275;
assign addr[41179]= -2138975100;
assign addr[41180]= -2090184478;
assign addr[41181]= -1999036154;
assign addr[41182]= -1867377253;
assign addr[41183]= -1697875851;
assign addr[41184]= -1493966902;
assign addr[41185]= -1259782632;
assign addr[41186]= -1000068799;
assign addr[41187]= -720088517;
assign addr[41188]= -425515602;
assign addr[41189]= -122319591;
assign addr[41190]= 183355234;
assign addr[41191]= 485314355;
assign addr[41192]= 777438554;
assign addr[41193]= 1053807919;
assign addr[41194]= 1308821808;
assign addr[41195]= 1537312353;
assign addr[41196]= 1734649179;
assign addr[41197]= 1896833245;
assign addr[41198]= 2020577882;
assign addr[41199]= 2103375398;
assign addr[41200]= 2143547897;
assign addr[41201]= 2140281282;
assign addr[41202]= 2093641749;
assign addr[41203]= 2004574453;
assign addr[41204]= 1874884346;
assign addr[41205]= 1707199606;
assign addr[41206]= 1504918373;
assign addr[41207]= 1272139887;
assign addr[41208]= 1013581418;
assign addr[41209]= 734482665;
assign addr[41210]= 440499581;
assign addr[41211]= 137589750;
assign addr[41212]= -168108346;
assign addr[41213]= -470399716;
assign addr[41214]= -763158411;
assign addr[41215]= -1040451659;
assign addr[41216]= -1296660098;
assign addr[41217]= -1526591649;
assign addr[41218]= -1725586737;
assign addr[41219]= -1889612716;
assign addr[41220]= -2015345591;
assign addr[41221]= -2100237377;
assign addr[41222]= -2142567738;
assign addr[41223]= -2141478848;
assign addr[41224]= -2096992772;
assign addr[41225]= -2010011024;
assign addr[41226]= -1882296293;
assign addr[41227]= -1716436725;
assign addr[41228]= -1515793473;
assign addr[41229]= -1284432584;
assign addr[41230]= -1027042599;
assign addr[41231]= -748839539;
assign addr[41232]= -455461206;
assign addr[41233]= -152852926;
assign addr[41234]= 152852926;
assign addr[41235]= 455461206;
assign addr[41236]= 748839539;
assign addr[41237]= 1027042599;
assign addr[41238]= 1284432584;
assign addr[41239]= 1515793473;
assign addr[41240]= 1716436725;
assign addr[41241]= 1882296293;
assign addr[41242]= 2010011024;
assign addr[41243]= 2096992772;
assign addr[41244]= 2141478848;
assign addr[41245]= 2142567738;
assign addr[41246]= 2100237377;
assign addr[41247]= 2015345591;
assign addr[41248]= 1889612716;
assign addr[41249]= 1725586737;
assign addr[41250]= 1526591649;
assign addr[41251]= 1296660098;
assign addr[41252]= 1040451659;
assign addr[41253]= 763158411;
assign addr[41254]= 470399716;
assign addr[41255]= 168108346;
assign addr[41256]= -137589750;
assign addr[41257]= -440499581;
assign addr[41258]= -734482665;
assign addr[41259]= -1013581418;
assign addr[41260]= -1272139887;
assign addr[41261]= -1504918373;
assign addr[41262]= -1707199606;
assign addr[41263]= -1874884346;
assign addr[41264]= -2004574453;
assign addr[41265]= -2093641749;
assign addr[41266]= -2140281282;
assign addr[41267]= -2143547897;
assign addr[41268]= -2103375398;
assign addr[41269]= -2020577882;
assign addr[41270]= -1896833245;
assign addr[41271]= -1734649179;
assign addr[41272]= -1537312353;
assign addr[41273]= -1308821808;
assign addr[41274]= -1053807919;
assign addr[41275]= -777438554;
assign addr[41276]= -485314355;
assign addr[41277]= -183355234;
assign addr[41278]= 122319591;
assign addr[41279]= 425515602;
assign addr[41280]= 720088517;
assign addr[41281]= 1000068799;
assign addr[41282]= 1259782632;
assign addr[41283]= 1493966902;
assign addr[41284]= 1697875851;
assign addr[41285]= 1867377253;
assign addr[41286]= 1999036154;
assign addr[41287]= 2090184478;
assign addr[41288]= 2138975100;
assign addr[41289]= 2144419275;
assign addr[41290]= 2106406677;
assign addr[41291]= 2025707632;
assign addr[41292]= 1903957513;
assign addr[41293]= 1743623590;
assign addr[41294]= 1547955041;
assign addr[41295]= 1320917099;
assign addr[41296]= 1067110699;
assign addr[41297]= 791679244;
assign addr[41298]= 500204365;
assign addr[41299]= 198592817;
assign addr[41300]= -107043224;
assign addr[41301]= -410510029;
assign addr[41302]= -705657826;
assign addr[41303]= -986505429;
assign addr[41304]= -1247361445;
assign addr[41305]= -1482939614;
assign addr[41306]= -1688465931;
assign addr[41307]= -1859775393;
assign addr[41308]= -1993396407;
assign addr[41309]= -2086621133;
assign addr[41310]= -2137560369;
assign addr[41311]= -2145181827;
assign addr[41312]= -2109331059;
assign addr[41313]= -2030734582;
assign addr[41314]= -1910985158;
assign addr[41315]= -1752509516;
assign addr[41316]= -1558519173;
assign addr[41317]= -1332945355;
assign addr[41318]= -1080359326;
assign addr[41319]= -805879757;
assign addr[41320]= -515068990;
assign addr[41321]= -213820322;
assign addr[41322]= 91761426;
assign addr[41323]= 395483624;
assign addr[41324]= 691191324;
assign addr[41325]= 972891995;
assign addr[41326]= 1234876957;
assign addr[41327]= 1471837070;
assign addr[41328]= 1678970324;
assign addr[41329]= 1852079154;
assign addr[41330]= 1987655498;
assign addr[41331]= 2082951896;
assign addr[41332]= 2136037160;
assign addr[41333]= 2145835515;
assign addr[41334]= 2112148396;
assign addr[41335]= 2035658475;
assign addr[41336]= 1917915825;
assign addr[41337]= 1761306505;
assign addr[41338]= 1569004214;
assign addr[41339]= 1344905966;
assign addr[41340]= 1093553126;
assign addr[41341]= 820039373;
assign addr[41342]= 529907477;
assign addr[41343]= 229036977;
assign addr[41344]= -76474970;
assign addr[41345]= -380437148;
assign addr[41346]= -676689746;
assign addr[41347]= -959229189;
assign addr[41348]= -1222329801;
assign addr[41349]= -1460659832;
assign addr[41350]= -1669389513;
assign addr[41351]= -1844288924;
assign addr[41352]= -1981813720;
assign addr[41353]= -2079176953;
assign addr[41354]= -2134405552;
assign addr[41355]= -2146380306;
assign addr[41356]= -2114858546;
assign addr[41357]= -2040479063;
assign addr[41358]= -1924749160;
assign addr[41359]= -1770014111;
assign addr[41360]= -1579409630;
assign addr[41361]= -1356798326;
assign addr[41362]= -1106691431;
assign addr[41363]= -834157373;
assign addr[41364]= -544719071;
assign addr[41365]= -244242007;
assign addr[41366]= 61184634;
assign addr[41367]= 365371365;
assign addr[41368]= 662153826;
assign addr[41369]= 945517704;
assign addr[41370]= 1209720613;
assign addr[41371]= 1449408469;
assign addr[41372]= 1659723983;
assign addr[41373]= 1836405100;
assign addr[41374]= 1975871368;
assign addr[41375]= 2075296495;
assign addr[41376]= 2132665626;
assign addr[41377]= 2146816171;
assign addr[41378]= 2117461370;
assign addr[41379]= 2045196100;
assign addr[41380]= 1931484818;
assign addr[41381]= 1778631892;
assign addr[41382]= 1589734894;
assign addr[41383]= 1368621831;
assign addr[41384]= 1119773573;
assign addr[41385]= 848233042;
assign addr[41386]= 559503022;
assign addr[41387]= 259434643;
assign addr[41388]= -45891193;
assign addr[41389]= -350287041;
assign addr[41390]= -647584304;
assign addr[41391]= -931758235;
assign addr[41392]= -1197050035;
assign addr[41393]= -1438083551;
assign addr[41394]= -1649974225;
assign addr[41395]= -1828428082;
assign addr[41396]= -1969828744;
assign addr[41397]= -2071310720;
assign addr[41398]= -2130817471;
assign addr[41399]= -2147143090;
assign addr[41400]= -2119956737;
assign addr[41401]= -2049809346;
assign addr[41402]= -1938122457;
assign addr[41403]= -1787159411;
assign addr[41404]= -1599979481;
assign addr[41405]= -1380375881;
assign addr[41406]= -1132798888;
assign addr[41407]= -862265664;
assign addr[41408]= -574258580;
assign addr[41409]= -274614114;
assign addr[41410]= 30595422;
assign addr[41411]= 335184940;
assign addr[41412]= 632981917;
assign addr[41413]= 917951481;
assign addr[41414]= 1184318708;
assign addr[41415]= 1426685652;
assign addr[41416]= 1640140734;
assign addr[41417]= 1820358275;
assign addr[41418]= 1963686155;
assign addr[41419]= 2067219829;
assign addr[41420]= 2128861181;
assign addr[41421]= 2147361045;
assign addr[41422]= 2122344521;
assign addr[41423]= 2054318569;
assign addr[41424]= 1944661739;
assign addr[41425]= 1795596234;
assign addr[41426]= 1610142873;
assign addr[41427]= 1392059879;
assign addr[41428]= 1145766716;
assign addr[41429]= 876254528;
assign addr[41430]= 588984994;
assign addr[41431]= 289779648;
assign addr[41432]= -15298099;
assign addr[41433]= -320065829;
assign addr[41434]= -618347408;
assign addr[41435]= -904098143;
assign addr[41436]= -1171527280;
assign addr[41437]= -1415215352;
assign addr[41438]= -1630224009;
assign addr[41439]= -1812196087;
assign addr[41440]= -1957443913;
assign addr[41441]= -2063024031;
assign addr[41442]= -2126796855;
assign addr[41443]= -2147470025;
assign addr[41444]= -2124624598;
assign addr[41445]= -2058723538;
assign addr[41446]= -1951102334;
assign addr[41447]= -1803941934;
assign addr[41448]= -1620224553;
assign addr[41449]= -1403673233;
assign addr[41450]= -1158676398;
assign addr[41451]= -890198924;
assign addr[41452]= -603681519;
assign addr[41453]= -304930476;
assign addr[41454]= 0;
assign addr[41455]= 304930476;
assign addr[41456]= 603681519;
assign addr[41457]= 890198924;
assign addr[41458]= 1158676398;
assign addr[41459]= 1403673233;
assign addr[41460]= 1620224553;
assign addr[41461]= 1803941934;
assign addr[41462]= 1951102334;
assign addr[41463]= 2058723538;
assign addr[41464]= 2124624598;
assign addr[41465]= 2147470025;
assign addr[41466]= 2126796855;
assign addr[41467]= 2063024031;
assign addr[41468]= 1957443913;
assign addr[41469]= 1812196087;
assign addr[41470]= 1630224009;
assign addr[41471]= 1415215352;
assign addr[41472]= 1171527280;
assign addr[41473]= 904098143;
assign addr[41474]= 618347408;
assign addr[41475]= 320065829;
assign addr[41476]= 15298099;
assign addr[41477]= -289779648;
assign addr[41478]= -588984994;
assign addr[41479]= -876254528;
assign addr[41480]= -1145766716;
assign addr[41481]= -1392059879;
assign addr[41482]= -1610142873;
assign addr[41483]= -1795596234;
assign addr[41484]= -1944661739;
assign addr[41485]= -2054318569;
assign addr[41486]= -2122344521;
assign addr[41487]= -2147361045;
assign addr[41488]= -2128861181;
assign addr[41489]= -2067219829;
assign addr[41490]= -1963686155;
assign addr[41491]= -1820358275;
assign addr[41492]= -1640140734;
assign addr[41493]= -1426685652;
assign addr[41494]= -1184318708;
assign addr[41495]= -917951481;
assign addr[41496]= -632981917;
assign addr[41497]= -335184940;
assign addr[41498]= -30595422;
assign addr[41499]= 274614114;
assign addr[41500]= 574258580;
assign addr[41501]= 862265664;
assign addr[41502]= 1132798888;
assign addr[41503]= 1380375881;
assign addr[41504]= 1599979481;
assign addr[41505]= 1787159411;
assign addr[41506]= 1938122457;
assign addr[41507]= 2049809346;
assign addr[41508]= 2119956737;
assign addr[41509]= 2147143090;
assign addr[41510]= 2130817471;
assign addr[41511]= 2071310720;
assign addr[41512]= 1969828744;
assign addr[41513]= 1828428082;
assign addr[41514]= 1649974225;
assign addr[41515]= 1438083551;
assign addr[41516]= 1197050035;
assign addr[41517]= 931758235;
assign addr[41518]= 647584304;
assign addr[41519]= 350287041;
assign addr[41520]= 45891193;
assign addr[41521]= -259434643;
assign addr[41522]= -559503022;
assign addr[41523]= -848233042;
assign addr[41524]= -1119773573;
assign addr[41525]= -1368621831;
assign addr[41526]= -1589734894;
assign addr[41527]= -1778631892;
assign addr[41528]= -1931484818;
assign addr[41529]= -2045196100;
assign addr[41530]= -2117461370;
assign addr[41531]= -2146816171;
assign addr[41532]= -2132665626;
assign addr[41533]= -2075296495;
assign addr[41534]= -1975871368;
assign addr[41535]= -1836405100;
assign addr[41536]= -1659723983;
assign addr[41537]= -1449408469;
assign addr[41538]= -1209720613;
assign addr[41539]= -945517704;
assign addr[41540]= -662153826;
assign addr[41541]= -365371365;
assign addr[41542]= -61184634;
assign addr[41543]= 244242007;
assign addr[41544]= 544719071;
assign addr[41545]= 834157373;
assign addr[41546]= 1106691431;
assign addr[41547]= 1356798326;
assign addr[41548]= 1579409630;
assign addr[41549]= 1770014111;
assign addr[41550]= 1924749160;
assign addr[41551]= 2040479063;
assign addr[41552]= 2114858546;
assign addr[41553]= 2146380306;
assign addr[41554]= 2134405552;
assign addr[41555]= 2079176953;
assign addr[41556]= 1981813720;
assign addr[41557]= 1844288924;
assign addr[41558]= 1669389513;
assign addr[41559]= 1460659832;
assign addr[41560]= 1222329801;
assign addr[41561]= 959229189;
assign addr[41562]= 676689746;
assign addr[41563]= 380437148;
assign addr[41564]= 76474970;
assign addr[41565]= -229036977;
assign addr[41566]= -529907477;
assign addr[41567]= -820039373;
assign addr[41568]= -1093553126;
assign addr[41569]= -1344905966;
assign addr[41570]= -1569004214;
assign addr[41571]= -1761306505;
assign addr[41572]= -1917915825;
assign addr[41573]= -2035658475;
assign addr[41574]= -2112148396;
assign addr[41575]= -2145835515;
assign addr[41576]= -2136037160;
assign addr[41577]= -2082951896;
assign addr[41578]= -1987655498;
assign addr[41579]= -1852079154;
assign addr[41580]= -1678970324;
assign addr[41581]= -1471837070;
assign addr[41582]= -1234876957;
assign addr[41583]= -972891995;
assign addr[41584]= -691191324;
assign addr[41585]= -395483624;
assign addr[41586]= -91761426;
assign addr[41587]= 213820322;
assign addr[41588]= 515068990;
assign addr[41589]= 805879757;
assign addr[41590]= 1080359326;
assign addr[41591]= 1332945355;
assign addr[41592]= 1558519173;
assign addr[41593]= 1752509516;
assign addr[41594]= 1910985158;
assign addr[41595]= 2030734582;
assign addr[41596]= 2109331059;
assign addr[41597]= 2145181827;
assign addr[41598]= 2137560369;
assign addr[41599]= 2086621133;
assign addr[41600]= 1993396407;
assign addr[41601]= 1859775393;
assign addr[41602]= 1688465931;
assign addr[41603]= 1482939614;
assign addr[41604]= 1247361445;
assign addr[41605]= 986505429;
assign addr[41606]= 705657826;
assign addr[41607]= 410510029;
assign addr[41608]= 107043224;
assign addr[41609]= -198592817;
assign addr[41610]= -500204365;
assign addr[41611]= -791679244;
assign addr[41612]= -1067110699;
assign addr[41613]= -1320917099;
assign addr[41614]= -1547955041;
assign addr[41615]= -1743623590;
assign addr[41616]= -1903957513;
assign addr[41617]= -2025707632;
assign addr[41618]= -2106406677;
assign addr[41619]= -2144419275;
assign addr[41620]= -2138975100;
assign addr[41621]= -2090184478;
assign addr[41622]= -1999036154;
assign addr[41623]= -1867377253;
assign addr[41624]= -1697875851;
assign addr[41625]= -1493966902;
assign addr[41626]= -1259782632;
assign addr[41627]= -1000068799;
assign addr[41628]= -720088517;
assign addr[41629]= -425515602;
assign addr[41630]= -122319591;
assign addr[41631]= 183355234;
assign addr[41632]= 485314355;
assign addr[41633]= 777438554;
assign addr[41634]= 1053807919;
assign addr[41635]= 1308821808;
assign addr[41636]= 1537312353;
assign addr[41637]= 1734649179;
assign addr[41638]= 1896833245;
assign addr[41639]= 2020577882;
assign addr[41640]= 2103375398;
assign addr[41641]= 2143547897;
assign addr[41642]= 2140281282;
assign addr[41643]= 2093641749;
assign addr[41644]= 2004574453;
assign addr[41645]= 1874884346;
assign addr[41646]= 1707199606;
assign addr[41647]= 1504918373;
assign addr[41648]= 1272139887;
assign addr[41649]= 1013581418;
assign addr[41650]= 734482665;
assign addr[41651]= 440499581;
assign addr[41652]= 137589750;
assign addr[41653]= -168108346;
assign addr[41654]= -470399716;
assign addr[41655]= -763158411;
assign addr[41656]= -1040451659;
assign addr[41657]= -1296660098;
assign addr[41658]= -1526591649;
assign addr[41659]= -1725586737;
assign addr[41660]= -1889612716;
assign addr[41661]= -2015345591;
assign addr[41662]= -2100237377;
assign addr[41663]= -2142567738;
assign addr[41664]= -2141478848;
assign addr[41665]= -2096992772;
assign addr[41666]= -2010011024;
assign addr[41667]= -1882296293;
assign addr[41668]= -1716436725;
assign addr[41669]= -1515793473;
assign addr[41670]= -1284432584;
assign addr[41671]= -1027042599;
assign addr[41672]= -748839539;
assign addr[41673]= -455461206;
assign addr[41674]= -152852926;
assign addr[41675]= 152852926;
assign addr[41676]= 455461206;
assign addr[41677]= 748839539;
assign addr[41678]= 1027042599;
assign addr[41679]= 1284432584;
assign addr[41680]= 1515793473;
assign addr[41681]= 1716436725;
assign addr[41682]= 1882296293;
assign addr[41683]= 2010011024;
assign addr[41684]= 2096992772;
assign addr[41685]= 2141478848;
assign addr[41686]= 2142567738;
assign addr[41687]= 2100237377;
assign addr[41688]= 2015345591;
assign addr[41689]= 1889612716;
assign addr[41690]= 1725586737;
assign addr[41691]= 1526591649;
assign addr[41692]= 1296660098;
assign addr[41693]= 1040451659;
assign addr[41694]= 763158411;
assign addr[41695]= 470399716;
assign addr[41696]= 168108346;
assign addr[41697]= -137589750;
assign addr[41698]= -440499581;
assign addr[41699]= -734482665;
assign addr[41700]= -1013581418;
assign addr[41701]= -1272139887;
assign addr[41702]= -1504918373;
assign addr[41703]= -1707199606;
assign addr[41704]= -1874884346;
assign addr[41705]= -2004574453;
assign addr[41706]= -2093641749;
assign addr[41707]= -2140281282;
assign addr[41708]= -2143547897;
assign addr[41709]= -2103375398;
assign addr[41710]= -2020577882;
assign addr[41711]= -1896833245;
assign addr[41712]= -1734649179;
assign addr[41713]= -1537312353;
assign addr[41714]= -1308821808;
assign addr[41715]= -1053807919;
assign addr[41716]= -777438554;
assign addr[41717]= -485314355;
assign addr[41718]= -183355234;
assign addr[41719]= 122319591;
assign addr[41720]= 425515602;
assign addr[41721]= 720088517;
assign addr[41722]= 1000068799;
assign addr[41723]= 1259782632;
assign addr[41724]= 1493966902;
assign addr[41725]= 1697875851;
assign addr[41726]= 1867377253;
assign addr[41727]= 1999036154;
assign addr[41728]= 2090184478;
assign addr[41729]= 2138975100;
assign addr[41730]= 2144419275;
assign addr[41731]= 2106406677;
assign addr[41732]= 2025707632;
assign addr[41733]= 1903957513;
assign addr[41734]= 1743623590;
assign addr[41735]= 1547955041;
assign addr[41736]= 1320917099;
assign addr[41737]= 1067110699;
assign addr[41738]= 791679244;
assign addr[41739]= 500204365;
assign addr[41740]= 198592817;
assign addr[41741]= -107043224;
assign addr[41742]= -410510029;
assign addr[41743]= -705657826;
assign addr[41744]= -986505429;
assign addr[41745]= -1247361445;
assign addr[41746]= -1482939614;
assign addr[41747]= -1688465931;
assign addr[41748]= -1859775393;
assign addr[41749]= -1993396407;
assign addr[41750]= -2086621133;
assign addr[41751]= -2137560369;
assign addr[41752]= -2145181827;
assign addr[41753]= -2109331059;
assign addr[41754]= -2030734582;
assign addr[41755]= -1910985158;
assign addr[41756]= -1752509516;
assign addr[41757]= -1558519173;
assign addr[41758]= -1332945355;
assign addr[41759]= -1080359326;
assign addr[41760]= -805879757;
assign addr[41761]= -515068990;
assign addr[41762]= -213820322;
assign addr[41763]= 91761426;
assign addr[41764]= 395483624;
assign addr[41765]= 691191324;
assign addr[41766]= 972891995;
assign addr[41767]= 1234876957;
assign addr[41768]= 1471837070;
assign addr[41769]= 1678970324;
assign addr[41770]= 1852079154;
assign addr[41771]= 1987655498;
assign addr[41772]= 2082951896;
assign addr[41773]= 2136037160;
assign addr[41774]= 2145835515;
assign addr[41775]= 2112148396;
assign addr[41776]= 2035658475;
assign addr[41777]= 1917915825;
assign addr[41778]= 1761306505;
assign addr[41779]= 1569004214;
assign addr[41780]= 1344905966;
assign addr[41781]= 1093553126;
assign addr[41782]= 820039373;
assign addr[41783]= 529907477;
assign addr[41784]= 229036977;
assign addr[41785]= -76474970;
assign addr[41786]= -380437148;
assign addr[41787]= -676689746;
assign addr[41788]= -959229189;
assign addr[41789]= -1222329801;
assign addr[41790]= -1460659832;
assign addr[41791]= -1669389513;
assign addr[41792]= -1844288924;
assign addr[41793]= -1981813720;
assign addr[41794]= -2079176953;
assign addr[41795]= -2134405552;
assign addr[41796]= -2146380306;
assign addr[41797]= -2114858546;
assign addr[41798]= -2040479063;
assign addr[41799]= -1924749160;
assign addr[41800]= -1770014111;
assign addr[41801]= -1579409630;
assign addr[41802]= -1356798326;
assign addr[41803]= -1106691431;
assign addr[41804]= -834157373;
assign addr[41805]= -544719071;
assign addr[41806]= -244242007;
assign addr[41807]= 61184634;
assign addr[41808]= 365371365;
assign addr[41809]= 662153826;
assign addr[41810]= 945517704;
assign addr[41811]= 1209720613;
assign addr[41812]= 1449408469;
assign addr[41813]= 1659723983;
assign addr[41814]= 1836405100;
assign addr[41815]= 1975871368;
assign addr[41816]= 2075296495;
assign addr[41817]= 2132665626;
assign addr[41818]= 2146816171;
assign addr[41819]= 2117461370;
assign addr[41820]= 2045196100;
assign addr[41821]= 1931484818;
assign addr[41822]= 1778631892;
assign addr[41823]= 1589734894;
assign addr[41824]= 1368621831;
assign addr[41825]= 1119773573;
assign addr[41826]= 848233042;
assign addr[41827]= 559503022;
assign addr[41828]= 259434643;
assign addr[41829]= -45891193;
assign addr[41830]= -350287041;
assign addr[41831]= -647584304;
assign addr[41832]= -931758235;
assign addr[41833]= -1197050035;
assign addr[41834]= -1438083551;
assign addr[41835]= -1649974225;
assign addr[41836]= -1828428082;
assign addr[41837]= -1969828744;
assign addr[41838]= -2071310720;
assign addr[41839]= -2130817471;
assign addr[41840]= -2147143090;
assign addr[41841]= -2119956737;
assign addr[41842]= -2049809346;
assign addr[41843]= -1938122457;
assign addr[41844]= -1787159411;
assign addr[41845]= -1599979481;
assign addr[41846]= -1380375881;
assign addr[41847]= -1132798888;
assign addr[41848]= -862265664;
assign addr[41849]= -574258580;
assign addr[41850]= -274614114;
assign addr[41851]= 30595422;
assign addr[41852]= 335184940;
assign addr[41853]= 632981917;
assign addr[41854]= 917951481;
assign addr[41855]= 1184318708;
assign addr[41856]= 1426685652;
assign addr[41857]= 1640140734;
assign addr[41858]= 1820358275;
assign addr[41859]= 1963686155;
assign addr[41860]= 2067219829;
assign addr[41861]= 2128861181;
assign addr[41862]= 2147361045;
assign addr[41863]= 2122344521;
assign addr[41864]= 2054318569;
assign addr[41865]= 1944661739;
assign addr[41866]= 1795596234;
assign addr[41867]= 1610142873;
assign addr[41868]= 1392059879;
assign addr[41869]= 1145766716;
assign addr[41870]= 876254528;
assign addr[41871]= 588984994;
assign addr[41872]= 289779648;
assign addr[41873]= -15298099;
assign addr[41874]= -320065829;
assign addr[41875]= -618347408;
assign addr[41876]= -904098143;
assign addr[41877]= -1171527280;
assign addr[41878]= -1415215352;
assign addr[41879]= -1630224009;
assign addr[41880]= -1812196087;
assign addr[41881]= -1957443913;
assign addr[41882]= -2063024031;
assign addr[41883]= -2126796855;
assign addr[41884]= -2147470025;
assign addr[41885]= -2124624598;
assign addr[41886]= -2058723538;
assign addr[41887]= -1951102334;
assign addr[41888]= -1803941934;
assign addr[41889]= -1620224553;
assign addr[41890]= -1403673233;
assign addr[41891]= -1158676398;
assign addr[41892]= -890198924;
assign addr[41893]= -603681519;
assign addr[41894]= -304930476;
assign addr[41895]= 0;
assign addr[41896]= 304930476;
assign addr[41897]= 603681519;
assign addr[41898]= 890198924;
assign addr[41899]= 1158676398;
assign addr[41900]= 1403673233;
assign addr[41901]= 1620224553;
assign addr[41902]= 1803941934;
assign addr[41903]= 1951102334;
assign addr[41904]= 2058723538;
assign addr[41905]= 2124624598;
assign addr[41906]= 2147470025;
assign addr[41907]= 2126796855;
assign addr[41908]= 2063024031;
assign addr[41909]= 1957443913;
assign addr[41910]= 1812196087;
assign addr[41911]= 1630224009;
assign addr[41912]= 1415215352;
assign addr[41913]= 1171527280;
assign addr[41914]= 904098143;
assign addr[41915]= 618347408;
assign addr[41916]= 320065829;
assign addr[41917]= 15298099;
assign addr[41918]= -289779648;
assign addr[41919]= -588984994;
assign addr[41920]= -876254528;
assign addr[41921]= -1145766716;
assign addr[41922]= -1392059879;
assign addr[41923]= -1610142873;
assign addr[41924]= -1795596234;
assign addr[41925]= -1944661739;
assign addr[41926]= -2054318569;
assign addr[41927]= -2122344521;
assign addr[41928]= -2147361045;
assign addr[41929]= -2128861181;
assign addr[41930]= -2067219829;
assign addr[41931]= -1963686155;
assign addr[41932]= -1820358275;
assign addr[41933]= -1640140734;
assign addr[41934]= -1426685652;
assign addr[41935]= -1184318708;
assign addr[41936]= -917951481;
assign addr[41937]= -632981917;
assign addr[41938]= -335184940;
assign addr[41939]= -30595422;
assign addr[41940]= 274614114;
assign addr[41941]= 574258580;
assign addr[41942]= 862265664;
assign addr[41943]= 1132798888;
assign addr[41944]= 1380375881;
assign addr[41945]= 1599979481;
assign addr[41946]= 1787159411;
assign addr[41947]= 1938122457;
assign addr[41948]= 2049809346;
assign addr[41949]= 2119956737;
assign addr[41950]= 2147143090;
assign addr[41951]= 2130817471;
assign addr[41952]= 2071310720;
assign addr[41953]= 1969828744;
assign addr[41954]= 1828428082;
assign addr[41955]= 1649974225;
assign addr[41956]= 1438083551;
assign addr[41957]= 1197050035;
assign addr[41958]= 931758235;
assign addr[41959]= 647584304;
assign addr[41960]= 350287041;
assign addr[41961]= 45891193;
assign addr[41962]= -259434643;
assign addr[41963]= -559503022;
assign addr[41964]= -848233042;
assign addr[41965]= -1119773573;
assign addr[41966]= -1368621831;
assign addr[41967]= -1589734894;
assign addr[41968]= -1778631892;
assign addr[41969]= -1931484818;
assign addr[41970]= -2045196100;
assign addr[41971]= -2117461370;
assign addr[41972]= -2146816171;
assign addr[41973]= -2132665626;
assign addr[41974]= -2075296495;
assign addr[41975]= -1975871368;
assign addr[41976]= -1836405100;
assign addr[41977]= -1659723983;
assign addr[41978]= -1449408469;
assign addr[41979]= -1209720613;
assign addr[41980]= -945517704;
assign addr[41981]= -662153826;
assign addr[41982]= -365371365;
assign addr[41983]= -61184634;
assign addr[41984]= 244242007;
assign addr[41985]= 544719071;
assign addr[41986]= 834157373;
assign addr[41987]= 1106691431;
assign addr[41988]= 1356798326;
assign addr[41989]= 1579409630;
assign addr[41990]= 1770014111;
assign addr[41991]= 1924749160;
assign addr[41992]= 2040479063;
assign addr[41993]= 2114858546;
assign addr[41994]= 2146380306;
assign addr[41995]= 2134405552;
assign addr[41996]= 2079176953;
assign addr[41997]= 1981813720;
assign addr[41998]= 1844288924;
assign addr[41999]= 1669389513;
assign addr[42000]= 1460659832;
assign addr[42001]= 1222329801;
assign addr[42002]= 959229189;
assign addr[42003]= 676689746;
assign addr[42004]= 380437148;
assign addr[42005]= 76474970;
assign addr[42006]= -229036977;
assign addr[42007]= -529907477;
assign addr[42008]= -820039373;
assign addr[42009]= -1093553126;
assign addr[42010]= -1344905966;
assign addr[42011]= -1569004214;
assign addr[42012]= -1761306505;
assign addr[42013]= -1917915825;
assign addr[42014]= -2035658475;
assign addr[42015]= -2112148396;
assign addr[42016]= -2145835515;
assign addr[42017]= -2136037160;
assign addr[42018]= -2082951896;
assign addr[42019]= -1987655498;
assign addr[42020]= -1852079154;
assign addr[42021]= -1678970324;
assign addr[42022]= -1471837070;
assign addr[42023]= -1234876957;
assign addr[42024]= -972891995;
assign addr[42025]= -691191324;
assign addr[42026]= -395483624;
assign addr[42027]= -91761426;
assign addr[42028]= 213820322;
assign addr[42029]= 515068990;
assign addr[42030]= 805879757;
assign addr[42031]= 1080359326;
assign addr[42032]= 1332945355;
assign addr[42033]= 1558519173;
assign addr[42034]= 1752509516;
assign addr[42035]= 1910985158;
assign addr[42036]= 2030734582;
assign addr[42037]= 2109331059;
assign addr[42038]= 2145181827;
assign addr[42039]= 2137560369;
assign addr[42040]= 2086621133;
assign addr[42041]= 1993396407;
assign addr[42042]= 1859775393;
assign addr[42043]= 1688465931;
assign addr[42044]= 1482939614;
assign addr[42045]= 1247361445;
assign addr[42046]= 986505429;
assign addr[42047]= 705657826;
assign addr[42048]= 410510029;
assign addr[42049]= 107043224;
assign addr[42050]= -198592817;
assign addr[42051]= -500204365;
assign addr[42052]= -791679244;
assign addr[42053]= -1067110699;
assign addr[42054]= -1320917099;
assign addr[42055]= -1547955041;
assign addr[42056]= -1743623590;
assign addr[42057]= -1903957513;
assign addr[42058]= -2025707632;
assign addr[42059]= -2106406677;
assign addr[42060]= -2144419275;
assign addr[42061]= -2138975100;
assign addr[42062]= -2090184478;
assign addr[42063]= -1999036154;
assign addr[42064]= -1867377253;
assign addr[42065]= -1697875851;
assign addr[42066]= -1493966902;
assign addr[42067]= -1259782632;
assign addr[42068]= -1000068799;
assign addr[42069]= -720088517;
assign addr[42070]= -425515602;
assign addr[42071]= -122319591;
assign addr[42072]= 183355234;
assign addr[42073]= 485314355;
assign addr[42074]= 777438554;
assign addr[42075]= 1053807919;
assign addr[42076]= 1308821808;
assign addr[42077]= 1537312353;
assign addr[42078]= 1734649179;
assign addr[42079]= 1896833245;
assign addr[42080]= 2020577882;
assign addr[42081]= 2103375398;
assign addr[42082]= 2143547897;
assign addr[42083]= 2140281282;
assign addr[42084]= 2093641749;
assign addr[42085]= 2004574453;
assign addr[42086]= 1874884346;
assign addr[42087]= 1707199606;
assign addr[42088]= 1504918373;
assign addr[42089]= 1272139887;
assign addr[42090]= 1013581418;
assign addr[42091]= 734482665;
assign addr[42092]= 440499581;
assign addr[42093]= 137589750;
assign addr[42094]= -168108346;
assign addr[42095]= -470399716;
assign addr[42096]= -763158411;
assign addr[42097]= -1040451659;
assign addr[42098]= -1296660098;
assign addr[42099]= -1526591649;
assign addr[42100]= -1725586737;
assign addr[42101]= -1889612716;
assign addr[42102]= -2015345591;
assign addr[42103]= -2100237377;
assign addr[42104]= -2142567738;
assign addr[42105]= -2141478848;
assign addr[42106]= -2096992772;
assign addr[42107]= -2010011024;
assign addr[42108]= -1882296293;
assign addr[42109]= -1716436725;
assign addr[42110]= -1515793473;
assign addr[42111]= -1284432584;
assign addr[42112]= -1027042599;
assign addr[42113]= -748839539;
assign addr[42114]= -455461206;
assign addr[42115]= -152852926;
assign addr[42116]= 152852926;
assign addr[42117]= 455461206;
assign addr[42118]= 748839539;
assign addr[42119]= 1027042599;
assign addr[42120]= 1284432584;
assign addr[42121]= 1515793473;
assign addr[42122]= 1716436725;
assign addr[42123]= 1882296293;
assign addr[42124]= 2010011024;
assign addr[42125]= 2096992772;
assign addr[42126]= 2141478848;
assign addr[42127]= 2142567738;
assign addr[42128]= 2100237377;
assign addr[42129]= 2015345591;
assign addr[42130]= 1889612716;
assign addr[42131]= 1725586737;
assign addr[42132]= 1526591649;
assign addr[42133]= 1296660098;
assign addr[42134]= 1040451659;
assign addr[42135]= 763158411;
assign addr[42136]= 470399716;
assign addr[42137]= 168108346;
assign addr[42138]= -137589750;
assign addr[42139]= -440499581;
assign addr[42140]= -734482665;
assign addr[42141]= -1013581418;
assign addr[42142]= -1272139887;
assign addr[42143]= -1504918373;
assign addr[42144]= -1707199606;
assign addr[42145]= -1874884346;
assign addr[42146]= -2004574453;
assign addr[42147]= -2093641749;
assign addr[42148]= -2140281282;
assign addr[42149]= -2143547897;
assign addr[42150]= -2103375398;
assign addr[42151]= -2020577882;
assign addr[42152]= -1896833245;
assign addr[42153]= -1734649179;
assign addr[42154]= -1537312353;
assign addr[42155]= -1308821808;
assign addr[42156]= -1053807919;
assign addr[42157]= -777438554;
assign addr[42158]= -485314355;
assign addr[42159]= -183355234;
assign addr[42160]= 122319591;
assign addr[42161]= 425515602;
assign addr[42162]= 720088517;
assign addr[42163]= 1000068799;
assign addr[42164]= 1259782632;
assign addr[42165]= 1493966902;
assign addr[42166]= 1697875851;
assign addr[42167]= 1867377253;
assign addr[42168]= 1999036154;
assign addr[42169]= 2090184478;
assign addr[42170]= 2138975100;
assign addr[42171]= 2144419275;
assign addr[42172]= 2106406677;
assign addr[42173]= 2025707632;
assign addr[42174]= 1903957513;
assign addr[42175]= 1743623590;
assign addr[42176]= 1547955041;
assign addr[42177]= 1320917099;
assign addr[42178]= 1067110699;
assign addr[42179]= 791679244;
assign addr[42180]= 500204365;
assign addr[42181]= 198592817;
assign addr[42182]= -107043224;
assign addr[42183]= -410510029;
assign addr[42184]= -705657826;
assign addr[42185]= -986505429;
assign addr[42186]= -1247361445;
assign addr[42187]= -1482939614;
assign addr[42188]= -1688465931;
assign addr[42189]= -1859775393;
assign addr[42190]= -1993396407;
assign addr[42191]= -2086621133;
assign addr[42192]= -2137560369;
assign addr[42193]= -2145181827;
assign addr[42194]= -2109331059;
assign addr[42195]= -2030734582;
assign addr[42196]= -1910985158;
assign addr[42197]= -1752509516;
assign addr[42198]= -1558519173;
assign addr[42199]= -1332945355;
assign addr[42200]= -1080359326;
assign addr[42201]= -805879757;
assign addr[42202]= -515068990;
assign addr[42203]= -213820322;
assign addr[42204]= 91761426;
assign addr[42205]= 395483624;
assign addr[42206]= 691191324;
assign addr[42207]= 972891995;
assign addr[42208]= 1234876957;
assign addr[42209]= 1471837070;
assign addr[42210]= 1678970324;
assign addr[42211]= 1852079154;
assign addr[42212]= 1987655498;
assign addr[42213]= 2082951896;
assign addr[42214]= 2136037160;
assign addr[42215]= 2145835515;
assign addr[42216]= 2112148396;
assign addr[42217]= 2035658475;
assign addr[42218]= 1917915825;
assign addr[42219]= 1761306505;
assign addr[42220]= 1569004214;
assign addr[42221]= 1344905966;
assign addr[42222]= 1093553126;
assign addr[42223]= 820039373;
assign addr[42224]= 529907477;
assign addr[42225]= 229036977;
assign addr[42226]= -76474970;
assign addr[42227]= -380437148;
assign addr[42228]= -676689746;
assign addr[42229]= -959229189;
assign addr[42230]= -1222329801;
assign addr[42231]= -1460659832;
assign addr[42232]= -1669389513;
assign addr[42233]= -1844288924;
assign addr[42234]= -1981813720;
assign addr[42235]= -2079176953;
assign addr[42236]= -2134405552;
assign addr[42237]= -2146380306;
assign addr[42238]= -2114858546;
assign addr[42239]= -2040479063;
assign addr[42240]= -1924749160;
assign addr[42241]= -1770014111;
assign addr[42242]= -1579409630;
assign addr[42243]= -1356798326;
assign addr[42244]= -1106691431;
assign addr[42245]= -834157373;
assign addr[42246]= -544719071;
assign addr[42247]= -244242007;
assign addr[42248]= 61184634;
assign addr[42249]= 365371365;
assign addr[42250]= 662153826;
assign addr[42251]= 945517704;
assign addr[42252]= 1209720613;
assign addr[42253]= 1449408469;
assign addr[42254]= 1659723983;
assign addr[42255]= 1836405100;
assign addr[42256]= 1975871368;
assign addr[42257]= 2075296495;
assign addr[42258]= 2132665626;
assign addr[42259]= 2146816171;
assign addr[42260]= 2117461370;
assign addr[42261]= 2045196100;
assign addr[42262]= 1931484818;
assign addr[42263]= 1778631892;
assign addr[42264]= 1589734894;
assign addr[42265]= 1368621831;
assign addr[42266]= 1119773573;
assign addr[42267]= 848233042;
assign addr[42268]= 559503022;
assign addr[42269]= 259434643;
assign addr[42270]= -45891193;
assign addr[42271]= -350287041;
assign addr[42272]= -647584304;
assign addr[42273]= -931758235;
assign addr[42274]= -1197050035;
assign addr[42275]= -1438083551;
assign addr[42276]= -1649974225;
assign addr[42277]= -1828428082;
assign addr[42278]= -1969828744;
assign addr[42279]= -2071310720;
assign addr[42280]= -2130817471;
assign addr[42281]= -2147143090;
assign addr[42282]= -2119956737;
assign addr[42283]= -2049809346;
assign addr[42284]= -1938122457;
assign addr[42285]= -1787159411;
assign addr[42286]= -1599979481;
assign addr[42287]= -1380375881;
assign addr[42288]= -1132798888;
assign addr[42289]= -862265664;
assign addr[42290]= -574258580;
assign addr[42291]= -274614114;
assign addr[42292]= 30595422;
assign addr[42293]= 335184940;
assign addr[42294]= 632981917;
assign addr[42295]= 917951481;
assign addr[42296]= 1184318708;
assign addr[42297]= 1426685652;
assign addr[42298]= 1640140734;
assign addr[42299]= 1820358275;
assign addr[42300]= 1963686155;
assign addr[42301]= 2067219829;
assign addr[42302]= 2128861181;
assign addr[42303]= 2147361045;
assign addr[42304]= 2122344521;
assign addr[42305]= 2054318569;
assign addr[42306]= 1944661739;
assign addr[42307]= 1795596234;
assign addr[42308]= 1610142873;
assign addr[42309]= 1392059879;
assign addr[42310]= 1145766716;
assign addr[42311]= 876254528;
assign addr[42312]= 588984994;
assign addr[42313]= 289779648;
assign addr[42314]= -15298099;
assign addr[42315]= -320065829;
assign addr[42316]= -618347408;
assign addr[42317]= -904098143;
assign addr[42318]= -1171527280;
assign addr[42319]= -1415215352;
assign addr[42320]= -1630224009;
assign addr[42321]= -1812196087;
assign addr[42322]= -1957443913;
assign addr[42323]= -2063024031;
assign addr[42324]= -2126796855;
assign addr[42325]= -2147470025;
assign addr[42326]= -2124624598;
assign addr[42327]= -2058723538;
assign addr[42328]= -1951102334;
assign addr[42329]= -1803941934;
assign addr[42330]= -1620224553;
assign addr[42331]= -1403673233;
assign addr[42332]= -1158676398;
assign addr[42333]= -890198924;
assign addr[42334]= -603681519;
assign addr[42335]= -304930476;
assign addr[42336]= 0;
assign addr[42337]= 304930476;
assign addr[42338]= 603681519;
assign addr[42339]= 890198924;
assign addr[42340]= 1158676398;
assign addr[42341]= 1403673233;
assign addr[42342]= 1620224553;
assign addr[42343]= 1803941934;
assign addr[42344]= 1951102334;
assign addr[42345]= 2058723538;
assign addr[42346]= 2124624598;
assign addr[42347]= 2147470025;
assign addr[42348]= 2126796855;
assign addr[42349]= 2063024031;
assign addr[42350]= 1957443913;
assign addr[42351]= 1812196087;
assign addr[42352]= 1630224009;
assign addr[42353]= 1415215352;
assign addr[42354]= 1171527280;
assign addr[42355]= 904098143;
assign addr[42356]= 618347408;
assign addr[42357]= 320065829;
assign addr[42358]= 15298099;
assign addr[42359]= -289779648;
assign addr[42360]= -588984994;
assign addr[42361]= -876254528;
assign addr[42362]= -1145766716;
assign addr[42363]= -1392059879;
assign addr[42364]= -1610142873;
assign addr[42365]= -1795596234;
assign addr[42366]= -1944661739;
assign addr[42367]= -2054318569;
assign addr[42368]= -2122344521;
assign addr[42369]= -2147361045;
assign addr[42370]= -2128861181;
assign addr[42371]= -2067219829;
assign addr[42372]= -1963686155;
assign addr[42373]= -1820358275;
assign addr[42374]= -1640140734;
assign addr[42375]= -1426685652;
assign addr[42376]= -1184318708;
assign addr[42377]= -917951481;
assign addr[42378]= -632981917;
assign addr[42379]= -335184940;
assign addr[42380]= -30595422;
assign addr[42381]= 274614114;
assign addr[42382]= 574258580;
assign addr[42383]= 862265664;
assign addr[42384]= 1132798888;
assign addr[42385]= 1380375881;
assign addr[42386]= 1599979481;
assign addr[42387]= 1787159411;
assign addr[42388]= 1938122457;
assign addr[42389]= 2049809346;
assign addr[42390]= 2119956737;
assign addr[42391]= 2147143090;
assign addr[42392]= 2130817471;
assign addr[42393]= 2071310720;
assign addr[42394]= 1969828744;
assign addr[42395]= 1828428082;
assign addr[42396]= 1649974225;
assign addr[42397]= 1438083551;
assign addr[42398]= 1197050035;
assign addr[42399]= 931758235;
assign addr[42400]= 647584304;
assign addr[42401]= 350287041;
assign addr[42402]= 45891193;
assign addr[42403]= -259434643;
assign addr[42404]= -559503022;
assign addr[42405]= -848233042;
assign addr[42406]= -1119773573;
assign addr[42407]= -1368621831;
assign addr[42408]= -1589734894;
assign addr[42409]= -1778631892;
assign addr[42410]= -1931484818;
assign addr[42411]= -2045196100;
assign addr[42412]= -2117461370;
assign addr[42413]= -2146816171;
assign addr[42414]= -2132665626;
assign addr[42415]= -2075296495;
assign addr[42416]= -1975871368;
assign addr[42417]= -1836405100;
assign addr[42418]= -1659723983;
assign addr[42419]= -1449408469;
assign addr[42420]= -1209720613;
assign addr[42421]= -945517704;
assign addr[42422]= -662153826;
assign addr[42423]= -365371365;
assign addr[42424]= -61184634;
assign addr[42425]= 244242007;
assign addr[42426]= 544719071;
assign addr[42427]= 834157373;
assign addr[42428]= 1106691431;
assign addr[42429]= 1356798326;
assign addr[42430]= 1579409630;
assign addr[42431]= 1770014111;
assign addr[42432]= 1924749160;
assign addr[42433]= 2040479063;
assign addr[42434]= 2114858546;
assign addr[42435]= 2146380306;
assign addr[42436]= 2134405552;
assign addr[42437]= 2079176953;
assign addr[42438]= 1981813720;
assign addr[42439]= 1844288924;
assign addr[42440]= 1669389513;
assign addr[42441]= 1460659832;
assign addr[42442]= 1222329801;
assign addr[42443]= 959229189;
assign addr[42444]= 676689746;
assign addr[42445]= 380437148;
assign addr[42446]= 76474970;
assign addr[42447]= -229036977;
assign addr[42448]= -529907477;
assign addr[42449]= -820039373;
assign addr[42450]= -1093553126;
assign addr[42451]= -1344905966;
assign addr[42452]= -1569004214;
assign addr[42453]= -1761306505;
assign addr[42454]= -1917915825;
assign addr[42455]= -2035658475;
assign addr[42456]= -2112148396;
assign addr[42457]= -2145835515;
assign addr[42458]= -2136037160;
assign addr[42459]= -2082951896;
assign addr[42460]= -1987655498;
assign addr[42461]= -1852079154;
assign addr[42462]= -1678970324;
assign addr[42463]= -1471837070;
assign addr[42464]= -1234876957;
assign addr[42465]= -972891995;
assign addr[42466]= -691191324;
assign addr[42467]= -395483624;
assign addr[42468]= -91761426;
assign addr[42469]= 213820322;
assign addr[42470]= 515068990;
assign addr[42471]= 805879757;
assign addr[42472]= 1080359326;
assign addr[42473]= 1332945355;
assign addr[42474]= 1558519173;
assign addr[42475]= 1752509516;
assign addr[42476]= 1910985158;
assign addr[42477]= 2030734582;
assign addr[42478]= 2109331059;
assign addr[42479]= 2145181827;
assign addr[42480]= 2137560369;
assign addr[42481]= 2086621133;
assign addr[42482]= 1993396407;
assign addr[42483]= 1859775393;
assign addr[42484]= 1688465931;
assign addr[42485]= 1482939614;
assign addr[42486]= 1247361445;
assign addr[42487]= 986505429;
assign addr[42488]= 705657826;
assign addr[42489]= 410510029;
assign addr[42490]= 107043224;
assign addr[42491]= -198592817;
assign addr[42492]= -500204365;
assign addr[42493]= -791679244;
assign addr[42494]= -1067110699;
assign addr[42495]= -1320917099;
assign addr[42496]= -1547955041;
assign addr[42497]= -1743623590;
assign addr[42498]= -1903957513;
assign addr[42499]= -2025707632;
assign addr[42500]= -2106406677;
assign addr[42501]= -2144419275;
assign addr[42502]= -2138975100;
assign addr[42503]= -2090184478;
assign addr[42504]= -1999036154;
assign addr[42505]= -1867377253;
assign addr[42506]= -1697875851;
assign addr[42507]= -1493966902;
assign addr[42508]= -1259782632;
assign addr[42509]= -1000068799;
assign addr[42510]= -720088517;
assign addr[42511]= -425515602;
assign addr[42512]= -122319591;
assign addr[42513]= 183355234;
assign addr[42514]= 485314355;
assign addr[42515]= 777438554;
assign addr[42516]= 1053807919;
assign addr[42517]= 1308821808;
assign addr[42518]= 1537312353;
assign addr[42519]= 1734649179;
assign addr[42520]= 1896833245;
assign addr[42521]= 2020577882;
assign addr[42522]= 2103375398;
assign addr[42523]= 2143547897;
assign addr[42524]= 2140281282;
assign addr[42525]= 2093641749;
assign addr[42526]= 2004574453;
assign addr[42527]= 1874884346;
assign addr[42528]= 1707199606;
assign addr[42529]= 1504918373;
assign addr[42530]= 1272139887;
assign addr[42531]= 1013581418;
assign addr[42532]= 734482665;
assign addr[42533]= 440499581;
assign addr[42534]= 137589750;
assign addr[42535]= -168108346;
assign addr[42536]= -470399716;
assign addr[42537]= -763158411;
assign addr[42538]= -1040451659;
assign addr[42539]= -1296660098;
assign addr[42540]= -1526591649;
assign addr[42541]= -1725586737;
assign addr[42542]= -1889612716;
assign addr[42543]= -2015345591;
assign addr[42544]= -2100237377;
assign addr[42545]= -2142567738;
assign addr[42546]= -2141478848;
assign addr[42547]= -2096992772;
assign addr[42548]= -2010011024;
assign addr[42549]= -1882296293;
assign addr[42550]= -1716436725;
assign addr[42551]= -1515793473;
assign addr[42552]= -1284432584;
assign addr[42553]= -1027042599;
assign addr[42554]= -748839539;
assign addr[42555]= -455461206;
assign addr[42556]= -152852926;
assign addr[42557]= 152852926;
assign addr[42558]= 455461206;
assign addr[42559]= 748839539;
assign addr[42560]= 1027042599;
assign addr[42561]= 1284432584;
assign addr[42562]= 1515793473;
assign addr[42563]= 1716436725;
assign addr[42564]= 1882296293;
assign addr[42565]= 2010011024;
assign addr[42566]= 2096992772;
assign addr[42567]= 2141478848;
assign addr[42568]= 2142567738;
assign addr[42569]= 2100237377;
assign addr[42570]= 2015345591;
assign addr[42571]= 1889612716;
assign addr[42572]= 1725586737;
assign addr[42573]= 1526591649;
assign addr[42574]= 1296660098;
assign addr[42575]= 1040451659;
assign addr[42576]= 763158411;
assign addr[42577]= 470399716;
assign addr[42578]= 168108346;
assign addr[42579]= -137589750;
assign addr[42580]= -440499581;
assign addr[42581]= -734482665;
assign addr[42582]= -1013581418;
assign addr[42583]= -1272139887;
assign addr[42584]= -1504918373;
assign addr[42585]= -1707199606;
assign addr[42586]= -1874884346;
assign addr[42587]= -2004574453;
assign addr[42588]= -2093641749;
assign addr[42589]= -2140281282;
assign addr[42590]= -2143547897;
assign addr[42591]= -2103375398;
assign addr[42592]= -2020577882;
assign addr[42593]= -1896833245;
assign addr[42594]= -1734649179;
assign addr[42595]= -1537312353;
assign addr[42596]= -1308821808;
assign addr[42597]= -1053807919;
assign addr[42598]= -777438554;
assign addr[42599]= -485314355;
assign addr[42600]= -183355234;
assign addr[42601]= 122319591;
assign addr[42602]= 425515602;
assign addr[42603]= 720088517;
assign addr[42604]= 1000068799;
assign addr[42605]= 1259782632;
assign addr[42606]= 1493966902;
assign addr[42607]= 1697875851;
assign addr[42608]= 1867377253;
assign addr[42609]= 1999036154;
assign addr[42610]= 2090184478;
assign addr[42611]= 2138975100;
assign addr[42612]= 2144419275;
assign addr[42613]= 2106406677;
assign addr[42614]= 2025707632;
assign addr[42615]= 1903957513;
assign addr[42616]= 1743623590;
assign addr[42617]= 1547955041;
assign addr[42618]= 1320917099;
assign addr[42619]= 1067110699;
assign addr[42620]= 791679244;
assign addr[42621]= 500204365;
assign addr[42622]= 198592817;
assign addr[42623]= -107043224;
assign addr[42624]= -410510029;
assign addr[42625]= -705657826;
assign addr[42626]= -986505429;
assign addr[42627]= -1247361445;
assign addr[42628]= -1482939614;
assign addr[42629]= -1688465931;
assign addr[42630]= -1859775393;
assign addr[42631]= -1993396407;
assign addr[42632]= -2086621133;
assign addr[42633]= -2137560369;
assign addr[42634]= -2145181827;
assign addr[42635]= -2109331059;
assign addr[42636]= -2030734582;
assign addr[42637]= -1910985158;
assign addr[42638]= -1752509516;
assign addr[42639]= -1558519173;
assign addr[42640]= -1332945355;
assign addr[42641]= -1080359326;
assign addr[42642]= -805879757;
assign addr[42643]= -515068990;
assign addr[42644]= -213820322;
assign addr[42645]= 91761426;
assign addr[42646]= 395483624;
assign addr[42647]= 691191324;
assign addr[42648]= 972891995;
assign addr[42649]= 1234876957;
assign addr[42650]= 1471837070;
assign addr[42651]= 1678970324;
assign addr[42652]= 1852079154;
assign addr[42653]= 1987655498;
assign addr[42654]= 2082951896;
assign addr[42655]= 2136037160;
assign addr[42656]= 2145835515;
assign addr[42657]= 2112148396;
assign addr[42658]= 2035658475;
assign addr[42659]= 1917915825;
assign addr[42660]= 1761306505;
assign addr[42661]= 1569004214;
assign addr[42662]= 1344905966;
assign addr[42663]= 1093553126;
assign addr[42664]= 820039373;
assign addr[42665]= 529907477;
assign addr[42666]= 229036977;
assign addr[42667]= -76474970;
assign addr[42668]= -380437148;
assign addr[42669]= -676689746;
assign addr[42670]= -959229189;
assign addr[42671]= -1222329801;
assign addr[42672]= -1460659832;
assign addr[42673]= -1669389513;
assign addr[42674]= -1844288924;
assign addr[42675]= -1981813720;
assign addr[42676]= -2079176953;
assign addr[42677]= -2134405552;
assign addr[42678]= -2146380306;
assign addr[42679]= -2114858546;
assign addr[42680]= -2040479063;
assign addr[42681]= -1924749160;
assign addr[42682]= -1770014111;
assign addr[42683]= -1579409630;
assign addr[42684]= -1356798326;
assign addr[42685]= -1106691431;
assign addr[42686]= -834157373;
assign addr[42687]= -544719071;
assign addr[42688]= -244242007;
assign addr[42689]= 61184634;
assign addr[42690]= 365371365;
assign addr[42691]= 662153826;
assign addr[42692]= 945517704;
assign addr[42693]= 1209720613;
assign addr[42694]= 1449408469;
assign addr[42695]= 1659723983;
assign addr[42696]= 1836405100;
assign addr[42697]= 1975871368;
assign addr[42698]= 2075296495;
assign addr[42699]= 2132665626;
assign addr[42700]= 2146816171;
assign addr[42701]= 2117461370;
assign addr[42702]= 2045196100;
assign addr[42703]= 1931484818;
assign addr[42704]= 1778631892;
assign addr[42705]= 1589734894;
assign addr[42706]= 1368621831;
assign addr[42707]= 1119773573;
assign addr[42708]= 848233042;
assign addr[42709]= 559503022;
assign addr[42710]= 259434643;
assign addr[42711]= -45891193;
assign addr[42712]= -350287041;
assign addr[42713]= -647584304;
assign addr[42714]= -931758235;
assign addr[42715]= -1197050035;
assign addr[42716]= -1438083551;
assign addr[42717]= -1649974225;
assign addr[42718]= -1828428082;
assign addr[42719]= -1969828744;
assign addr[42720]= -2071310720;
assign addr[42721]= -2130817471;
assign addr[42722]= -2147143090;
assign addr[42723]= -2119956737;
assign addr[42724]= -2049809346;
assign addr[42725]= -1938122457;
assign addr[42726]= -1787159411;
assign addr[42727]= -1599979481;
assign addr[42728]= -1380375881;
assign addr[42729]= -1132798888;
assign addr[42730]= -862265664;
assign addr[42731]= -574258580;
assign addr[42732]= -274614114;
assign addr[42733]= 30595422;
assign addr[42734]= 335184940;
assign addr[42735]= 632981917;
assign addr[42736]= 917951481;
assign addr[42737]= 1184318708;
assign addr[42738]= 1426685652;
assign addr[42739]= 1640140734;
assign addr[42740]= 1820358275;
assign addr[42741]= 1963686155;
assign addr[42742]= 2067219829;
assign addr[42743]= 2128861181;
assign addr[42744]= 2147361045;
assign addr[42745]= 2122344521;
assign addr[42746]= 2054318569;
assign addr[42747]= 1944661739;
assign addr[42748]= 1795596234;
assign addr[42749]= 1610142873;
assign addr[42750]= 1392059879;
assign addr[42751]= 1145766716;
assign addr[42752]= 876254528;
assign addr[42753]= 588984994;
assign addr[42754]= 289779648;
assign addr[42755]= -15298099;
assign addr[42756]= -320065829;
assign addr[42757]= -618347408;
assign addr[42758]= -904098143;
assign addr[42759]= -1171527280;
assign addr[42760]= -1415215352;
assign addr[42761]= -1630224009;
assign addr[42762]= -1812196087;
assign addr[42763]= -1957443913;
assign addr[42764]= -2063024031;
assign addr[42765]= -2126796855;
assign addr[42766]= -2147470025;
assign addr[42767]= -2124624598;
assign addr[42768]= -2058723538;
assign addr[42769]= -1951102334;
assign addr[42770]= -1803941934;
assign addr[42771]= -1620224553;
assign addr[42772]= -1403673233;
assign addr[42773]= -1158676398;
assign addr[42774]= -890198924;
assign addr[42775]= -603681519;
assign addr[42776]= -304930476;
assign addr[42777]= 0;
assign addr[42778]= 304930476;
assign addr[42779]= 603681519;
assign addr[42780]= 890198924;
assign addr[42781]= 1158676398;
assign addr[42782]= 1403673233;
assign addr[42783]= 1620224553;
assign addr[42784]= 1803941934;
assign addr[42785]= 1951102334;
assign addr[42786]= 2058723538;
assign addr[42787]= 2124624598;
assign addr[42788]= 2147470025;
assign addr[42789]= 2126796855;
assign addr[42790]= 2063024031;
assign addr[42791]= 1957443913;
assign addr[42792]= 1812196087;
assign addr[42793]= 1630224009;
assign addr[42794]= 1415215352;
assign addr[42795]= 1171527280;
assign addr[42796]= 904098143;
assign addr[42797]= 618347408;
assign addr[42798]= 320065829;
assign addr[42799]= 15298099;
assign addr[42800]= -289779648;
assign addr[42801]= -588984994;
assign addr[42802]= -876254528;
assign addr[42803]= -1145766716;
assign addr[42804]= -1392059879;
assign addr[42805]= -1610142873;
assign addr[42806]= -1795596234;
assign addr[42807]= -1944661739;
assign addr[42808]= -2054318569;
assign addr[42809]= -2122344521;
assign addr[42810]= -2147361045;
assign addr[42811]= -2128861181;
assign addr[42812]= -2067219829;
assign addr[42813]= -1963686155;
assign addr[42814]= -1820358275;
assign addr[42815]= -1640140734;
assign addr[42816]= -1426685652;
assign addr[42817]= -1184318708;
assign addr[42818]= -917951481;
assign addr[42819]= -632981917;
assign addr[42820]= -335184940;
assign addr[42821]= -30595422;
assign addr[42822]= 274614114;
assign addr[42823]= 574258580;
assign addr[42824]= 862265664;
assign addr[42825]= 1132798888;
assign addr[42826]= 1380375881;
assign addr[42827]= 1599979481;
assign addr[42828]= 1787159411;
assign addr[42829]= 1938122457;
assign addr[42830]= 2049809346;
assign addr[42831]= 2119956737;
assign addr[42832]= 2147143090;
assign addr[42833]= 2130817471;
assign addr[42834]= 2071310720;
assign addr[42835]= 1969828744;
assign addr[42836]= 1828428082;
assign addr[42837]= 1649974225;
assign addr[42838]= 1438083551;
assign addr[42839]= 1197050035;
assign addr[42840]= 931758235;
assign addr[42841]= 647584304;
assign addr[42842]= 350287041;
assign addr[42843]= 45891193;
assign addr[42844]= -259434643;
assign addr[42845]= -559503022;
assign addr[42846]= -848233042;
assign addr[42847]= -1119773573;
assign addr[42848]= -1368621831;
assign addr[42849]= -1589734894;
assign addr[42850]= -1778631892;
assign addr[42851]= -1931484818;
assign addr[42852]= -2045196100;
assign addr[42853]= -2117461370;
assign addr[42854]= -2146816171;
assign addr[42855]= -2132665626;
assign addr[42856]= -2075296495;
assign addr[42857]= -1975871368;
assign addr[42858]= -1836405100;
assign addr[42859]= -1659723983;
assign addr[42860]= -1449408469;
assign addr[42861]= -1209720613;
assign addr[42862]= -945517704;
assign addr[42863]= -662153826;
assign addr[42864]= -365371365;
assign addr[42865]= -61184634;
assign addr[42866]= 244242007;
assign addr[42867]= 544719071;
assign addr[42868]= 834157373;
assign addr[42869]= 1106691431;
assign addr[42870]= 1356798326;
assign addr[42871]= 1579409630;
assign addr[42872]= 1770014111;
assign addr[42873]= 1924749160;
assign addr[42874]= 2040479063;
assign addr[42875]= 2114858546;
assign addr[42876]= 2146380306;
assign addr[42877]= 2134405552;
assign addr[42878]= 2079176953;
assign addr[42879]= 1981813720;
assign addr[42880]= 1844288924;
assign addr[42881]= 1669389513;
assign addr[42882]= 1460659832;
assign addr[42883]= 1222329801;
assign addr[42884]= 959229189;
assign addr[42885]= 676689746;
assign addr[42886]= 380437148;
assign addr[42887]= 76474970;
assign addr[42888]= -229036977;
assign addr[42889]= -529907477;
assign addr[42890]= -820039373;
assign addr[42891]= -1093553126;
assign addr[42892]= -1344905966;
assign addr[42893]= -1569004214;
assign addr[42894]= -1761306505;
assign addr[42895]= -1917915825;
assign addr[42896]= -2035658475;
assign addr[42897]= -2112148396;
assign addr[42898]= -2145835515;
assign addr[42899]= -2136037160;
assign addr[42900]= -2082951896;
assign addr[42901]= -1987655498;
assign addr[42902]= -1852079154;
assign addr[42903]= -1678970324;
assign addr[42904]= -1471837070;
assign addr[42905]= -1234876957;
assign addr[42906]= -972891995;
assign addr[42907]= -691191324;
assign addr[42908]= -395483624;
assign addr[42909]= -91761426;
assign addr[42910]= 213820322;
assign addr[42911]= 515068990;
assign addr[42912]= 805879757;
assign addr[42913]= 1080359326;
assign addr[42914]= 1332945355;
assign addr[42915]= 1558519173;
assign addr[42916]= 1752509516;
assign addr[42917]= 1910985158;
assign addr[42918]= 2030734582;
assign addr[42919]= 2109331059;
assign addr[42920]= 2145181827;
assign addr[42921]= 2137560369;
assign addr[42922]= 2086621133;
assign addr[42923]= 1993396407;
assign addr[42924]= 1859775393;
assign addr[42925]= 1688465931;
assign addr[42926]= 1482939614;
assign addr[42927]= 1247361445;
assign addr[42928]= 986505429;
assign addr[42929]= 705657826;
assign addr[42930]= 410510029;
assign addr[42931]= 107043224;
assign addr[42932]= -198592817;
assign addr[42933]= -500204365;
assign addr[42934]= -791679244;
assign addr[42935]= -1067110699;
assign addr[42936]= -1320917099;
assign addr[42937]= -1547955041;
assign addr[42938]= -1743623590;
assign addr[42939]= -1903957513;
assign addr[42940]= -2025707632;
assign addr[42941]= -2106406677;
assign addr[42942]= -2144419275;
assign addr[42943]= -2138975100;
assign addr[42944]= -2090184478;
assign addr[42945]= -1999036154;
assign addr[42946]= -1867377253;
assign addr[42947]= -1697875851;
assign addr[42948]= -1493966902;
assign addr[42949]= -1259782632;
assign addr[42950]= -1000068799;
assign addr[42951]= -720088517;
assign addr[42952]= -425515602;
assign addr[42953]= -122319591;
assign addr[42954]= 183355234;
assign addr[42955]= 485314355;
assign addr[42956]= 777438554;
assign addr[42957]= 1053807919;
assign addr[42958]= 1308821808;
assign addr[42959]= 1537312353;
assign addr[42960]= 1734649179;
assign addr[42961]= 1896833245;
assign addr[42962]= 2020577882;
assign addr[42963]= 2103375398;
assign addr[42964]= 2143547897;
assign addr[42965]= 2140281282;
assign addr[42966]= 2093641749;
assign addr[42967]= 2004574453;
assign addr[42968]= 1874884346;
assign addr[42969]= 1707199606;
assign addr[42970]= 1504918373;
assign addr[42971]= 1272139887;
assign addr[42972]= 1013581418;
assign addr[42973]= 734482665;
assign addr[42974]= 440499581;
assign addr[42975]= 137589750;
assign addr[42976]= -168108346;
assign addr[42977]= -470399716;
assign addr[42978]= -763158411;
assign addr[42979]= -1040451659;
assign addr[42980]= -1296660098;
assign addr[42981]= -1526591649;
assign addr[42982]= -1725586737;
assign addr[42983]= -1889612716;
assign addr[42984]= -2015345591;
assign addr[42985]= -2100237377;
assign addr[42986]= -2142567738;
assign addr[42987]= -2141478848;
assign addr[42988]= -2096992772;
assign addr[42989]= -2010011024;
assign addr[42990]= -1882296293;
assign addr[42991]= -1716436725;
assign addr[42992]= -1515793473;
assign addr[42993]= -1284432584;
assign addr[42994]= -1027042599;
assign addr[42995]= -748839539;
assign addr[42996]= -455461206;
assign addr[42997]= -152852926;
assign addr[42998]= 152852926;
assign addr[42999]= 455461206;
assign addr[43000]= 748839539;
assign addr[43001]= 1027042599;
assign addr[43002]= 1284432584;
assign addr[43003]= 1515793473;
assign addr[43004]= 1716436725;
assign addr[43005]= 1882296293;
assign addr[43006]= 2010011024;
assign addr[43007]= 2096992772;
assign addr[43008]= 2141478848;
assign addr[43009]= 2142567738;
assign addr[43010]= 2100237377;
assign addr[43011]= 2015345591;
assign addr[43012]= 1889612716;
assign addr[43013]= 1725586737;
assign addr[43014]= 1526591649;
assign addr[43015]= 1296660098;
assign addr[43016]= 1040451659;
assign addr[43017]= 763158411;
assign addr[43018]= 470399716;
assign addr[43019]= 168108346;
assign addr[43020]= -137589750;
assign addr[43021]= -440499581;
assign addr[43022]= -734482665;
assign addr[43023]= -1013581418;
assign addr[43024]= -1272139887;
assign addr[43025]= -1504918373;
assign addr[43026]= -1707199606;
assign addr[43027]= -1874884346;
assign addr[43028]= -2004574453;
assign addr[43029]= -2093641749;
assign addr[43030]= -2140281282;
assign addr[43031]= -2143547897;
assign addr[43032]= -2103375398;
assign addr[43033]= -2020577882;
assign addr[43034]= -1896833245;
assign addr[43035]= -1734649179;
assign addr[43036]= -1537312353;
assign addr[43037]= -1308821808;
assign addr[43038]= -1053807919;
assign addr[43039]= -777438554;
assign addr[43040]= -485314355;
assign addr[43041]= -183355234;
assign addr[43042]= 122319591;
assign addr[43043]= 425515602;
assign addr[43044]= 720088517;
assign addr[43045]= 1000068799;
assign addr[43046]= 1259782632;
assign addr[43047]= 1493966902;
assign addr[43048]= 1697875851;
assign addr[43049]= 1867377253;
assign addr[43050]= 1999036154;
assign addr[43051]= 2090184478;
assign addr[43052]= 2138975100;
assign addr[43053]= 2144419275;
assign addr[43054]= 2106406677;
assign addr[43055]= 2025707632;
assign addr[43056]= 1903957513;
assign addr[43057]= 1743623590;
assign addr[43058]= 1547955041;
assign addr[43059]= 1320917099;
assign addr[43060]= 1067110699;
assign addr[43061]= 791679244;
assign addr[43062]= 500204365;
assign addr[43063]= 198592817;
assign addr[43064]= -107043224;
assign addr[43065]= -410510029;
assign addr[43066]= -705657826;
assign addr[43067]= -986505429;
assign addr[43068]= -1247361445;
assign addr[43069]= -1482939614;
assign addr[43070]= -1688465931;
assign addr[43071]= -1859775393;
assign addr[43072]= -1993396407;
assign addr[43073]= -2086621133;
assign addr[43074]= -2137560369;
assign addr[43075]= -2145181827;
assign addr[43076]= -2109331059;
assign addr[43077]= -2030734582;
assign addr[43078]= -1910985158;
assign addr[43079]= -1752509516;
assign addr[43080]= -1558519173;
assign addr[43081]= -1332945355;
assign addr[43082]= -1080359326;
assign addr[43083]= -805879757;
assign addr[43084]= -515068990;
assign addr[43085]= -213820322;
assign addr[43086]= 91761426;
assign addr[43087]= 395483624;
assign addr[43088]= 691191324;
assign addr[43089]= 972891995;
assign addr[43090]= 1234876957;
assign addr[43091]= 1471837070;
assign addr[43092]= 1678970324;
assign addr[43093]= 1852079154;
assign addr[43094]= 1987655498;
assign addr[43095]= 2082951896;
assign addr[43096]= 2136037160;
assign addr[43097]= 2145835515;
assign addr[43098]= 2112148396;
assign addr[43099]= 2035658475;
assign addr[43100]= 1917915825;
assign addr[43101]= 1761306505;
assign addr[43102]= 1569004214;
assign addr[43103]= 1344905966;
assign addr[43104]= 1093553126;
assign addr[43105]= 820039373;
assign addr[43106]= 529907477;
assign addr[43107]= 229036977;
assign addr[43108]= -76474970;
assign addr[43109]= -380437148;
assign addr[43110]= -676689746;
assign addr[43111]= -959229189;
assign addr[43112]= -1222329801;
assign addr[43113]= -1460659832;
assign addr[43114]= -1669389513;
assign addr[43115]= -1844288924;
assign addr[43116]= -1981813720;
assign addr[43117]= -2079176953;
assign addr[43118]= -2134405552;
assign addr[43119]= -2146380306;
assign addr[43120]= -2114858546;
assign addr[43121]= -2040479063;
assign addr[43122]= -1924749160;
assign addr[43123]= -1770014111;
assign addr[43124]= -1579409630;
assign addr[43125]= -1356798326;
assign addr[43126]= -1106691431;
assign addr[43127]= -834157373;
assign addr[43128]= -544719071;
assign addr[43129]= -244242007;
assign addr[43130]= 61184634;
assign addr[43131]= 365371365;
assign addr[43132]= 662153826;
assign addr[43133]= 945517704;
assign addr[43134]= 1209720613;
assign addr[43135]= 1449408469;
assign addr[43136]= 1659723983;
assign addr[43137]= 1836405100;
assign addr[43138]= 1975871368;
assign addr[43139]= 2075296495;
assign addr[43140]= 2132665626;
assign addr[43141]= 2146816171;
assign addr[43142]= 2117461370;
assign addr[43143]= 2045196100;
assign addr[43144]= 1931484818;
assign addr[43145]= 1778631892;
assign addr[43146]= 1589734894;
assign addr[43147]= 1368621831;
assign addr[43148]= 1119773573;
assign addr[43149]= 848233042;
assign addr[43150]= 559503022;
assign addr[43151]= 259434643;
assign addr[43152]= -45891193;
assign addr[43153]= -350287041;
assign addr[43154]= -647584304;
assign addr[43155]= -931758235;
assign addr[43156]= -1197050035;
assign addr[43157]= -1438083551;
assign addr[43158]= -1649974225;
assign addr[43159]= -1828428082;
assign addr[43160]= -1969828744;
assign addr[43161]= -2071310720;
assign addr[43162]= -2130817471;
assign addr[43163]= -2147143090;
assign addr[43164]= -2119956737;
assign addr[43165]= -2049809346;
assign addr[43166]= -1938122457;
assign addr[43167]= -1787159411;
assign addr[43168]= -1599979481;
assign addr[43169]= -1380375881;
assign addr[43170]= -1132798888;
assign addr[43171]= -862265664;
assign addr[43172]= -574258580;
assign addr[43173]= -274614114;
assign addr[43174]= 30595422;
assign addr[43175]= 335184940;
assign addr[43176]= 632981917;
assign addr[43177]= 917951481;
assign addr[43178]= 1184318708;
assign addr[43179]= 1426685652;
assign addr[43180]= 1640140734;
assign addr[43181]= 1820358275;
assign addr[43182]= 1963686155;
assign addr[43183]= 2067219829;
assign addr[43184]= 2128861181;
assign addr[43185]= 2147361045;
assign addr[43186]= 2122344521;
assign addr[43187]= 2054318569;
assign addr[43188]= 1944661739;
assign addr[43189]= 1795596234;
assign addr[43190]= 1610142873;
assign addr[43191]= 1392059879;
assign addr[43192]= 1145766716;
assign addr[43193]= 876254528;
assign addr[43194]= 588984994;
assign addr[43195]= 289779648;
assign addr[43196]= -15298099;
assign addr[43197]= -320065829;
assign addr[43198]= -618347408;
assign addr[43199]= -904098143;
assign addr[43200]= -1171527280;
assign addr[43201]= -1415215352;
assign addr[43202]= -1630224009;
assign addr[43203]= -1812196087;
assign addr[43204]= -1957443913;
assign addr[43205]= -2063024031;
assign addr[43206]= -2126796855;
assign addr[43207]= -2147470025;
assign addr[43208]= -2124624598;
assign addr[43209]= -2058723538;
assign addr[43210]= -1951102334;
assign addr[43211]= -1803941934;
assign addr[43212]= -1620224553;
assign addr[43213]= -1403673233;
assign addr[43214]= -1158676398;
assign addr[43215]= -890198924;
assign addr[43216]= -603681519;
assign addr[43217]= -304930476;
assign addr[43218]= 0;
assign addr[43219]= 304930476;
assign addr[43220]= 603681519;
assign addr[43221]= 890198924;
assign addr[43222]= 1158676398;
assign addr[43223]= 1403673233;
assign addr[43224]= 1620224553;
assign addr[43225]= 1803941934;
assign addr[43226]= 1951102334;
assign addr[43227]= 2058723538;
assign addr[43228]= 2124624598;
assign addr[43229]= 2147470025;
assign addr[43230]= 2126796855;
assign addr[43231]= 2063024031;
assign addr[43232]= 1957443913;
assign addr[43233]= 1812196087;
assign addr[43234]= 1630224009;
assign addr[43235]= 1415215352;
assign addr[43236]= 1171527280;
assign addr[43237]= 904098143;
assign addr[43238]= 618347408;
assign addr[43239]= 320065829;
assign addr[43240]= 15298099;
assign addr[43241]= -289779648;
assign addr[43242]= -588984994;
assign addr[43243]= -876254528;
assign addr[43244]= -1145766716;
assign addr[43245]= -1392059879;
assign addr[43246]= -1610142873;
assign addr[43247]= -1795596234;
assign addr[43248]= -1944661739;
assign addr[43249]= -2054318569;
assign addr[43250]= -2122344521;
assign addr[43251]= -2147361045;
assign addr[43252]= -2128861181;
assign addr[43253]= -2067219829;
assign addr[43254]= -1963686155;
assign addr[43255]= -1820358275;
assign addr[43256]= -1640140734;
assign addr[43257]= -1426685652;
assign addr[43258]= -1184318708;
assign addr[43259]= -917951481;
assign addr[43260]= -632981917;
assign addr[43261]= -335184940;
assign addr[43262]= -30595422;
assign addr[43263]= 274614114;
assign addr[43264]= 574258580;
assign addr[43265]= 862265664;
assign addr[43266]= 1132798888;
assign addr[43267]= 1380375881;
assign addr[43268]= 1599979481;
assign addr[43269]= 1787159411;
assign addr[43270]= 1938122457;
assign addr[43271]= 2049809346;
assign addr[43272]= 2119956737;
assign addr[43273]= 2147143090;
assign addr[43274]= 2130817471;
assign addr[43275]= 2071310720;
assign addr[43276]= 1969828744;
assign addr[43277]= 1828428082;
assign addr[43278]= 1649974225;
assign addr[43279]= 1438083551;
assign addr[43280]= 1197050035;
assign addr[43281]= 931758235;
assign addr[43282]= 647584304;
assign addr[43283]= 350287041;
assign addr[43284]= 45891193;
assign addr[43285]= -259434643;
assign addr[43286]= -559503022;
assign addr[43287]= -848233042;
assign addr[43288]= -1119773573;
assign addr[43289]= -1368621831;
assign addr[43290]= -1589734894;
assign addr[43291]= -1778631892;
assign addr[43292]= -1931484818;
assign addr[43293]= -2045196100;
assign addr[43294]= -2117461370;
assign addr[43295]= -2146816171;
assign addr[43296]= -2132665626;
assign addr[43297]= -2075296495;
assign addr[43298]= -1975871368;
assign addr[43299]= -1836405100;
assign addr[43300]= -1659723983;
assign addr[43301]= -1449408469;
assign addr[43302]= -1209720613;
assign addr[43303]= -945517704;
assign addr[43304]= -662153826;
assign addr[43305]= -365371365;
assign addr[43306]= -61184634;
assign addr[43307]= 244242007;
assign addr[43308]= 544719071;
assign addr[43309]= 834157373;
assign addr[43310]= 1106691431;
assign addr[43311]= 1356798326;
assign addr[43312]= 1579409630;
assign addr[43313]= 1770014111;
assign addr[43314]= 1924749160;
assign addr[43315]= 2040479063;
assign addr[43316]= 2114858546;
assign addr[43317]= 2146380306;
assign addr[43318]= 2134405552;
assign addr[43319]= 2079176953;
assign addr[43320]= 1981813720;
assign addr[43321]= 1844288924;
assign addr[43322]= 1669389513;
assign addr[43323]= 1460659832;
assign addr[43324]= 1222329801;
assign addr[43325]= 959229189;
assign addr[43326]= 676689746;
assign addr[43327]= 380437148;
assign addr[43328]= 76474970;
assign addr[43329]= -229036977;
assign addr[43330]= -529907477;
assign addr[43331]= -820039373;
assign addr[43332]= -1093553126;
assign addr[43333]= -1344905966;
assign addr[43334]= -1569004214;
assign addr[43335]= -1761306505;
assign addr[43336]= -1917915825;
assign addr[43337]= -2035658475;
assign addr[43338]= -2112148396;
assign addr[43339]= -2145835515;
assign addr[43340]= -2136037160;
assign addr[43341]= -2082951896;
assign addr[43342]= -1987655498;
assign addr[43343]= -1852079154;
assign addr[43344]= -1678970324;
assign addr[43345]= -1471837070;
assign addr[43346]= -1234876957;
assign addr[43347]= -972891995;
assign addr[43348]= -691191324;
assign addr[43349]= -395483624;
assign addr[43350]= -91761426;
assign addr[43351]= 213820322;
assign addr[43352]= 515068990;
assign addr[43353]= 805879757;
assign addr[43354]= 1080359326;
assign addr[43355]= 1332945355;
assign addr[43356]= 1558519173;
assign addr[43357]= 1752509516;
assign addr[43358]= 1910985158;
assign addr[43359]= 2030734582;
assign addr[43360]= 2109331059;
assign addr[43361]= 2145181827;
assign addr[43362]= 2137560369;
assign addr[43363]= 2086621133;
assign addr[43364]= 1993396407;
assign addr[43365]= 1859775393;
assign addr[43366]= 1688465931;
assign addr[43367]= 1482939614;
assign addr[43368]= 1247361445;
assign addr[43369]= 986505429;
assign addr[43370]= 705657826;
assign addr[43371]= 410510029;
assign addr[43372]= 107043224;
assign addr[43373]= -198592817;
assign addr[43374]= -500204365;
assign addr[43375]= -791679244;
assign addr[43376]= -1067110699;
assign addr[43377]= -1320917099;
assign addr[43378]= -1547955041;
assign addr[43379]= -1743623590;
assign addr[43380]= -1903957513;
assign addr[43381]= -2025707632;
assign addr[43382]= -2106406677;
assign addr[43383]= -2144419275;
assign addr[43384]= -2138975100;
assign addr[43385]= -2090184478;
assign addr[43386]= -1999036154;
assign addr[43387]= -1867377253;
assign addr[43388]= -1697875851;
assign addr[43389]= -1493966902;
assign addr[43390]= -1259782632;
assign addr[43391]= -1000068799;
assign addr[43392]= -720088517;
assign addr[43393]= -425515602;
assign addr[43394]= -122319591;
assign addr[43395]= 183355234;
assign addr[43396]= 485314355;
assign addr[43397]= 777438554;
assign addr[43398]= 1053807919;
assign addr[43399]= 1308821808;
assign addr[43400]= 1537312353;
assign addr[43401]= 1734649179;
assign addr[43402]= 1896833245;
assign addr[43403]= 2020577882;
assign addr[43404]= 2103375398;
assign addr[43405]= 2143547897;
assign addr[43406]= 2140281282;
assign addr[43407]= 2093641749;
assign addr[43408]= 2004574453;
assign addr[43409]= 1874884346;
assign addr[43410]= 1707199606;
assign addr[43411]= 1504918373;
assign addr[43412]= 1272139887;
assign addr[43413]= 1013581418;
assign addr[43414]= 734482665;
assign addr[43415]= 440499581;
assign addr[43416]= 137589750;
assign addr[43417]= -168108346;
assign addr[43418]= -470399716;
assign addr[43419]= -763158411;
assign addr[43420]= -1040451659;
assign addr[43421]= -1296660098;
assign addr[43422]= -1526591649;
assign addr[43423]= -1725586737;
assign addr[43424]= -1889612716;
assign addr[43425]= -2015345591;
assign addr[43426]= -2100237377;
assign addr[43427]= -2142567738;
assign addr[43428]= -2141478848;
assign addr[43429]= -2096992772;
assign addr[43430]= -2010011024;
assign addr[43431]= -1882296293;
assign addr[43432]= -1716436725;
assign addr[43433]= -1515793473;
assign addr[43434]= -1284432584;
assign addr[43435]= -1027042599;
assign addr[43436]= -748839539;
assign addr[43437]= -455461206;
assign addr[43438]= -152852926;
assign addr[43439]= 152852926;
assign addr[43440]= 455461206;
assign addr[43441]= 748839539;
assign addr[43442]= 1027042599;
assign addr[43443]= 1284432584;
assign addr[43444]= 1515793473;
assign addr[43445]= 1716436725;
assign addr[43446]= 1882296293;
assign addr[43447]= 2010011024;
assign addr[43448]= 2096992772;
assign addr[43449]= 2141478848;
assign addr[43450]= 2142567738;
assign addr[43451]= 2100237377;
assign addr[43452]= 2015345591;
assign addr[43453]= 1889612716;
assign addr[43454]= 1725586737;
assign addr[43455]= 1526591649;
assign addr[43456]= 1296660098;
assign addr[43457]= 1040451659;
assign addr[43458]= 763158411;
assign addr[43459]= 470399716;
assign addr[43460]= 168108346;
assign addr[43461]= -137589750;
assign addr[43462]= -440499581;
assign addr[43463]= -734482665;
assign addr[43464]= -1013581418;
assign addr[43465]= -1272139887;
assign addr[43466]= -1504918373;
assign addr[43467]= -1707199606;
assign addr[43468]= -1874884346;
assign addr[43469]= -2004574453;
assign addr[43470]= -2093641749;
assign addr[43471]= -2140281282;
assign addr[43472]= -2143547897;
assign addr[43473]= -2103375398;
assign addr[43474]= -2020577882;
assign addr[43475]= -1896833245;
assign addr[43476]= -1734649179;
assign addr[43477]= -1537312353;
assign addr[43478]= -1308821808;
assign addr[43479]= -1053807919;
assign addr[43480]= -777438554;
assign addr[43481]= -485314355;
assign addr[43482]= -183355234;
assign addr[43483]= 122319591;
assign addr[43484]= 425515602;
assign addr[43485]= 720088517;
assign addr[43486]= 1000068799;
assign addr[43487]= 1259782632;
assign addr[43488]= 1493966902;
assign addr[43489]= 1697875851;
assign addr[43490]= 1867377253;
assign addr[43491]= 1999036154;
assign addr[43492]= 2090184478;
assign addr[43493]= 2138975100;
assign addr[43494]= 2144419275;
assign addr[43495]= 2106406677;
assign addr[43496]= 2025707632;
assign addr[43497]= 1903957513;
assign addr[43498]= 1743623590;
assign addr[43499]= 1547955041;
assign addr[43500]= 1320917099;
assign addr[43501]= 1067110699;
assign addr[43502]= 791679244;
assign addr[43503]= 500204365;
assign addr[43504]= 198592817;
assign addr[43505]= -107043224;
assign addr[43506]= -410510029;
assign addr[43507]= -705657826;
assign addr[43508]= -986505429;
assign addr[43509]= -1247361445;
assign addr[43510]= -1482939614;
assign addr[43511]= -1688465931;
assign addr[43512]= -1859775393;
assign addr[43513]= -1993396407;
assign addr[43514]= -2086621133;
assign addr[43515]= -2137560369;
assign addr[43516]= -2145181827;
assign addr[43517]= -2109331059;
assign addr[43518]= -2030734582;
assign addr[43519]= -1910985158;
assign addr[43520]= -1752509516;
assign addr[43521]= -1558519173;
assign addr[43522]= -1332945355;
assign addr[43523]= -1080359326;
assign addr[43524]= -805879757;
assign addr[43525]= -515068990;
assign addr[43526]= -213820322;
assign addr[43527]= 91761426;
assign addr[43528]= 395483624;
assign addr[43529]= 691191324;
assign addr[43530]= 972891995;
assign addr[43531]= 1234876957;
assign addr[43532]= 1471837070;
assign addr[43533]= 1678970324;
assign addr[43534]= 1852079154;
assign addr[43535]= 1987655498;
assign addr[43536]= 2082951896;
assign addr[43537]= 2136037160;
assign addr[43538]= 2145835515;
assign addr[43539]= 2112148396;
assign addr[43540]= 2035658475;
assign addr[43541]= 1917915825;
assign addr[43542]= 1761306505;
assign addr[43543]= 1569004214;
assign addr[43544]= 1344905966;
assign addr[43545]= 1093553126;
assign addr[43546]= 820039373;
assign addr[43547]= 529907477;
assign addr[43548]= 229036977;
assign addr[43549]= -76474970;
assign addr[43550]= -380437148;
assign addr[43551]= -676689746;
assign addr[43552]= -959229189;
assign addr[43553]= -1222329801;
assign addr[43554]= -1460659832;
assign addr[43555]= -1669389513;
assign addr[43556]= -1844288924;
assign addr[43557]= -1981813720;
assign addr[43558]= -2079176953;
assign addr[43559]= -2134405552;
assign addr[43560]= -2146380306;
assign addr[43561]= -2114858546;
assign addr[43562]= -2040479063;
assign addr[43563]= -1924749160;
assign addr[43564]= -1770014111;
assign addr[43565]= -1579409630;
assign addr[43566]= -1356798326;
assign addr[43567]= -1106691431;
assign addr[43568]= -834157373;
assign addr[43569]= -544719071;
assign addr[43570]= -244242007;
assign addr[43571]= 61184634;
assign addr[43572]= 365371365;
assign addr[43573]= 662153826;
assign addr[43574]= 945517704;
assign addr[43575]= 1209720613;
assign addr[43576]= 1449408469;
assign addr[43577]= 1659723983;
assign addr[43578]= 1836405100;
assign addr[43579]= 1975871368;
assign addr[43580]= 2075296495;
assign addr[43581]= 2132665626;
assign addr[43582]= 2146816171;
assign addr[43583]= 2117461370;
assign addr[43584]= 2045196100;
assign addr[43585]= 1931484818;
assign addr[43586]= 1778631892;
assign addr[43587]= 1589734894;
assign addr[43588]= 1368621831;
assign addr[43589]= 1119773573;
assign addr[43590]= 848233042;
assign addr[43591]= 559503022;
assign addr[43592]= 259434643;
assign addr[43593]= -45891193;
assign addr[43594]= -350287041;
assign addr[43595]= -647584304;
assign addr[43596]= -931758235;
assign addr[43597]= -1197050035;
assign addr[43598]= -1438083551;
assign addr[43599]= -1649974225;
assign addr[43600]= -1828428082;
assign addr[43601]= -1969828744;
assign addr[43602]= -2071310720;
assign addr[43603]= -2130817471;
assign addr[43604]= -2147143090;
assign addr[43605]= -2119956737;
assign addr[43606]= -2049809346;
assign addr[43607]= -1938122457;
assign addr[43608]= -1787159411;
assign addr[43609]= -1599979481;
assign addr[43610]= -1380375881;
assign addr[43611]= -1132798888;
assign addr[43612]= -862265664;
assign addr[43613]= -574258580;
assign addr[43614]= -274614114;
assign addr[43615]= 30595422;
assign addr[43616]= 335184940;
assign addr[43617]= 632981917;
assign addr[43618]= 917951481;
assign addr[43619]= 1184318708;
assign addr[43620]= 1426685652;
assign addr[43621]= 1640140734;
assign addr[43622]= 1820358275;
assign addr[43623]= 1963686155;
assign addr[43624]= 2067219829;
assign addr[43625]= 2128861181;
assign addr[43626]= 2147361045;
assign addr[43627]= 2122344521;
assign addr[43628]= 2054318569;
assign addr[43629]= 1944661739;
assign addr[43630]= 1795596234;
assign addr[43631]= 1610142873;
assign addr[43632]= 1392059879;
assign addr[43633]= 1145766716;
assign addr[43634]= 876254528;
assign addr[43635]= 588984994;
assign addr[43636]= 289779648;
assign addr[43637]= -15298099;
assign addr[43638]= -320065829;
assign addr[43639]= -618347408;
assign addr[43640]= -904098143;
assign addr[43641]= -1171527280;
assign addr[43642]= -1415215352;
assign addr[43643]= -1630224009;
assign addr[43644]= -1812196087;
assign addr[43645]= -1957443913;
assign addr[43646]= -2063024031;
assign addr[43647]= -2126796855;
assign addr[43648]= -2147470025;
assign addr[43649]= -2124624598;
assign addr[43650]= -2058723538;
assign addr[43651]= -1951102334;
assign addr[43652]= -1803941934;
assign addr[43653]= -1620224553;
assign addr[43654]= -1403673233;
assign addr[43655]= -1158676398;
assign addr[43656]= -890198924;
assign addr[43657]= -603681519;
assign addr[43658]= -304930476;
assign addr[43659]= 0;
assign addr[43660]= 304930476;
assign addr[43661]= 603681519;
assign addr[43662]= 890198924;
assign addr[43663]= 1158676398;
assign addr[43664]= 1403673233;
assign addr[43665]= 1620224553;
assign addr[43666]= 1803941934;
assign addr[43667]= 1951102334;
assign addr[43668]= 2058723538;
assign addr[43669]= 2124624598;
assign addr[43670]= 2147470025;
assign addr[43671]= 2126796855;
assign addr[43672]= 2063024031;
assign addr[43673]= 1957443913;
assign addr[43674]= 1812196087;
assign addr[43675]= 1630224009;
assign addr[43676]= 1415215352;
assign addr[43677]= 1171527280;
assign addr[43678]= 904098143;
assign addr[43679]= 618347408;
assign addr[43680]= 320065829;
assign addr[43681]= 15298099;
assign addr[43682]= -289779648;
assign addr[43683]= -588984994;
assign addr[43684]= -876254528;
assign addr[43685]= -1145766716;
assign addr[43686]= -1392059879;
assign addr[43687]= -1610142873;
assign addr[43688]= -1795596234;
assign addr[43689]= -1944661739;
assign addr[43690]= -2054318569;
assign addr[43691]= -2122344521;
assign addr[43692]= -2147361045;
assign addr[43693]= -2128861181;
assign addr[43694]= -2067219829;
assign addr[43695]= -1963686155;
assign addr[43696]= -1820358275;
assign addr[43697]= -1640140734;
assign addr[43698]= -1426685652;
assign addr[43699]= -1184318708;
assign addr[43700]= -917951481;
assign addr[43701]= -632981917;
assign addr[43702]= -335184940;
assign addr[43703]= -30595422;
assign addr[43704]= 274614114;
assign addr[43705]= 574258580;
assign addr[43706]= 862265664;
assign addr[43707]= 1132798888;
assign addr[43708]= 1380375881;
assign addr[43709]= 1599979481;
assign addr[43710]= 1787159411;
assign addr[43711]= 1938122457;
assign addr[43712]= 2049809346;
assign addr[43713]= 2119956737;
assign addr[43714]= 2147143090;
assign addr[43715]= 2130817471;
assign addr[43716]= 2071310720;
assign addr[43717]= 1969828744;
assign addr[43718]= 1828428082;
assign addr[43719]= 1649974225;
assign addr[43720]= 1438083551;
assign addr[43721]= 1197050035;
assign addr[43722]= 931758235;
assign addr[43723]= 647584304;
assign addr[43724]= 350287041;
assign addr[43725]= 45891193;
assign addr[43726]= -259434643;
assign addr[43727]= -559503022;
assign addr[43728]= -848233042;
assign addr[43729]= -1119773573;
assign addr[43730]= -1368621831;
assign addr[43731]= -1589734894;
assign addr[43732]= -1778631892;
assign addr[43733]= -1931484818;
assign addr[43734]= -2045196100;
assign addr[43735]= -2117461370;
assign addr[43736]= -2146816171;
assign addr[43737]= -2132665626;
assign addr[43738]= -2075296495;
assign addr[43739]= -1975871368;
assign addr[43740]= -1836405100;
assign addr[43741]= -1659723983;
assign addr[43742]= -1449408469;
assign addr[43743]= -1209720613;
assign addr[43744]= -945517704;
assign addr[43745]= -662153826;
assign addr[43746]= -365371365;
assign addr[43747]= -61184634;
assign addr[43748]= 244242007;
assign addr[43749]= 544719071;
assign addr[43750]= 834157373;
assign addr[43751]= 1106691431;
assign addr[43752]= 1356798326;
assign addr[43753]= 1579409630;
assign addr[43754]= 1770014111;
assign addr[43755]= 1924749160;
assign addr[43756]= 2040479063;
assign addr[43757]= 2114858546;
assign addr[43758]= 2146380306;
assign addr[43759]= 2134405552;
assign addr[43760]= 2079176953;
assign addr[43761]= 1981813720;
assign addr[43762]= 1844288924;
assign addr[43763]= 1669389513;
assign addr[43764]= 1460659832;
assign addr[43765]= 1222329801;
assign addr[43766]= 959229189;
assign addr[43767]= 676689746;
assign addr[43768]= 380437148;
assign addr[43769]= 76474970;
assign addr[43770]= -229036977;
assign addr[43771]= -529907477;
assign addr[43772]= -820039373;
assign addr[43773]= -1093553126;
assign addr[43774]= -1344905966;
assign addr[43775]= -1569004214;
assign addr[43776]= -1761306505;
assign addr[43777]= -1917915825;
assign addr[43778]= -2035658475;
assign addr[43779]= -2112148396;
assign addr[43780]= -2145835515;
assign addr[43781]= -2136037160;
assign addr[43782]= -2082951896;
assign addr[43783]= -1987655498;
assign addr[43784]= -1852079154;
assign addr[43785]= -1678970324;
assign addr[43786]= -1471837070;
assign addr[43787]= -1234876957;
assign addr[43788]= -972891995;
assign addr[43789]= -691191324;
assign addr[43790]= -395483624;
assign addr[43791]= -91761426;
assign addr[43792]= 213820322;
assign addr[43793]= 515068990;
assign addr[43794]= 805879757;
assign addr[43795]= 1080359326;
assign addr[43796]= 1332945355;
assign addr[43797]= 1558519173;
assign addr[43798]= 1752509516;
assign addr[43799]= 1910985158;
assign addr[43800]= 2030734582;
assign addr[43801]= 2109331059;
assign addr[43802]= 2145181827;
assign addr[43803]= 2137560369;
assign addr[43804]= 2086621133;
assign addr[43805]= 1993396407;
assign addr[43806]= 1859775393;
assign addr[43807]= 1688465931;
assign addr[43808]= 1482939614;
assign addr[43809]= 1247361445;
assign addr[43810]= 986505429;
assign addr[43811]= 705657826;
assign addr[43812]= 410510029;
assign addr[43813]= 107043224;
assign addr[43814]= -198592817;
assign addr[43815]= -500204365;
assign addr[43816]= -791679244;
assign addr[43817]= -1067110699;
assign addr[43818]= -1320917099;
assign addr[43819]= -1547955041;
assign addr[43820]= -1743623590;
assign addr[43821]= -1903957513;
assign addr[43822]= -2025707632;
assign addr[43823]= -2106406677;
assign addr[43824]= -2144419275;
assign addr[43825]= -2138975100;
assign addr[43826]= -2090184478;
assign addr[43827]= -1999036154;
assign addr[43828]= -1867377253;
assign addr[43829]= -1697875851;
assign addr[43830]= -1493966902;
assign addr[43831]= -1259782632;
assign addr[43832]= -1000068799;
assign addr[43833]= -720088517;
assign addr[43834]= -425515602;
assign addr[43835]= -122319591;
assign addr[43836]= 183355234;
assign addr[43837]= 485314355;
assign addr[43838]= 777438554;
assign addr[43839]= 1053807919;
assign addr[43840]= 1308821808;
assign addr[43841]= 1537312353;
assign addr[43842]= 1734649179;
assign addr[43843]= 1896833245;
assign addr[43844]= 2020577882;
assign addr[43845]= 2103375398;
assign addr[43846]= 2143547897;
assign addr[43847]= 2140281282;
assign addr[43848]= 2093641749;
assign addr[43849]= 2004574453;
assign addr[43850]= 1874884346;
assign addr[43851]= 1707199606;
assign addr[43852]= 1504918373;
assign addr[43853]= 1272139887;
assign addr[43854]= 1013581418;
assign addr[43855]= 734482665;
assign addr[43856]= 440499581;
assign addr[43857]= 137589750;
assign addr[43858]= -168108346;
assign addr[43859]= -470399716;
assign addr[43860]= -763158411;
assign addr[43861]= -1040451659;
assign addr[43862]= -1296660098;
assign addr[43863]= -1526591649;
assign addr[43864]= -1725586737;
assign addr[43865]= -1889612716;
assign addr[43866]= -2015345591;
assign addr[43867]= -2100237377;
assign addr[43868]= -2142567738;
assign addr[43869]= -2141478848;
assign addr[43870]= -2096992772;
assign addr[43871]= -2010011024;
assign addr[43872]= -1882296293;
assign addr[43873]= -1716436725;
assign addr[43874]= -1515793473;
assign addr[43875]= -1284432584;
assign addr[43876]= -1027042599;
assign addr[43877]= -748839539;
assign addr[43878]= -455461206;
assign addr[43879]= -152852926;
assign addr[43880]= 152852926;
assign addr[43881]= 455461206;
assign addr[43882]= 748839539;
assign addr[43883]= 1027042599;
assign addr[43884]= 1284432584;
assign addr[43885]= 1515793473;
assign addr[43886]= 1716436725;
assign addr[43887]= 1882296293;
assign addr[43888]= 2010011024;
assign addr[43889]= 2096992772;
assign addr[43890]= 2141478848;
assign addr[43891]= 2142567738;
assign addr[43892]= 2100237377;
assign addr[43893]= 2015345591;
assign addr[43894]= 1889612716;
assign addr[43895]= 1725586737;
assign addr[43896]= 1526591649;
assign addr[43897]= 1296660098;
assign addr[43898]= 1040451659;
assign addr[43899]= 763158411;
assign addr[43900]= 470399716;
assign addr[43901]= 168108346;
assign addr[43902]= -137589750;
assign addr[43903]= -440499581;
assign addr[43904]= -734482665;
assign addr[43905]= -1013581418;
assign addr[43906]= -1272139887;
assign addr[43907]= -1504918373;
assign addr[43908]= -1707199606;
assign addr[43909]= -1874884346;
assign addr[43910]= -2004574453;
assign addr[43911]= -2093641749;
assign addr[43912]= -2140281282;
assign addr[43913]= -2143547897;
assign addr[43914]= -2103375398;
assign addr[43915]= -2020577882;
assign addr[43916]= -1896833245;
assign addr[43917]= -1734649179;
assign addr[43918]= -1537312353;
assign addr[43919]= -1308821808;
assign addr[43920]= -1053807919;
assign addr[43921]= -777438554;
assign addr[43922]= -485314355;
assign addr[43923]= -183355234;
assign addr[43924]= 122319591;
assign addr[43925]= 425515602;
assign addr[43926]= 720088517;
assign addr[43927]= 1000068799;
assign addr[43928]= 1259782632;
assign addr[43929]= 1493966902;
assign addr[43930]= 1697875851;
assign addr[43931]= 1867377253;
assign addr[43932]= 1999036154;
assign addr[43933]= 2090184478;
assign addr[43934]= 2138975100;
assign addr[43935]= 2144419275;
assign addr[43936]= 2106406677;
assign addr[43937]= 2025707632;
assign addr[43938]= 1903957513;
assign addr[43939]= 1743623590;
assign addr[43940]= 1547955041;
assign addr[43941]= 1320917099;
assign addr[43942]= 1067110699;
assign addr[43943]= 791679244;
assign addr[43944]= 500204365;
assign addr[43945]= 198592817;
assign addr[43946]= -107043224;
assign addr[43947]= -410510029;
assign addr[43948]= -705657826;
assign addr[43949]= -986505429;
assign addr[43950]= -1247361445;
assign addr[43951]= -1482939614;
assign addr[43952]= -1688465931;
assign addr[43953]= -1859775393;
assign addr[43954]= -1993396407;
assign addr[43955]= -2086621133;
assign addr[43956]= -2137560369;
assign addr[43957]= -2145181827;
assign addr[43958]= -2109331059;
assign addr[43959]= -2030734582;
assign addr[43960]= -1910985158;
assign addr[43961]= -1752509516;
assign addr[43962]= -1558519173;
assign addr[43963]= -1332945355;
assign addr[43964]= -1080359326;
assign addr[43965]= -805879757;
assign addr[43966]= -515068990;
assign addr[43967]= -213820322;
assign addr[43968]= 91761426;
assign addr[43969]= 395483624;
assign addr[43970]= 691191324;
assign addr[43971]= 972891995;
assign addr[43972]= 1234876957;
assign addr[43973]= 1471837070;
assign addr[43974]= 1678970324;
assign addr[43975]= 1852079154;
assign addr[43976]= 1987655498;
assign addr[43977]= 2082951896;
assign addr[43978]= 2136037160;
assign addr[43979]= 2145835515;
assign addr[43980]= 2112148396;
assign addr[43981]= 2035658475;
assign addr[43982]= 1917915825;
assign addr[43983]= 1761306505;
assign addr[43984]= 1569004214;
assign addr[43985]= 1344905966;
assign addr[43986]= 1093553126;
assign addr[43987]= 820039373;
assign addr[43988]= 529907477;
assign addr[43989]= 229036977;
assign addr[43990]= -76474970;
assign addr[43991]= -380437148;
assign addr[43992]= -676689746;
assign addr[43993]= -959229189;
assign addr[43994]= -1222329801;
assign addr[43995]= -1460659832;
assign addr[43996]= -1669389513;
assign addr[43997]= -1844288924;
assign addr[43998]= -1981813720;
assign addr[43999]= -2079176953;
assign addr[44000]= -2134405552;
assign addr[44001]= -2146380306;
assign addr[44002]= -2114858546;
assign addr[44003]= -2040479063;
assign addr[44004]= -1924749160;
assign addr[44005]= -1770014111;
assign addr[44006]= -1579409630;
assign addr[44007]= -1356798326;
assign addr[44008]= -1106691431;
assign addr[44009]= -834157373;
assign addr[44010]= -544719071;
assign addr[44011]= -244242007;
assign addr[44012]= 61184634;
assign addr[44013]= 365371365;
assign addr[44014]= 662153826;
assign addr[44015]= 945517704;
assign addr[44016]= 1209720613;
assign addr[44017]= 1449408469;
assign addr[44018]= 1659723983;
assign addr[44019]= 1836405100;
assign addr[44020]= 1975871368;
assign addr[44021]= 2075296495;
assign addr[44022]= 2132665626;
assign addr[44023]= 2146816171;
assign addr[44024]= 2117461370;
assign addr[44025]= 2045196100;
assign addr[44026]= 1931484818;
assign addr[44027]= 1778631892;
assign addr[44028]= 1589734894;
assign addr[44029]= 1368621831;
assign addr[44030]= 1119773573;
assign addr[44031]= 848233042;
assign addr[44032]= 559503022;
assign addr[44033]= 259434643;
assign addr[44034]= -45891193;
assign addr[44035]= -350287041;
assign addr[44036]= -647584304;
assign addr[44037]= -931758235;
assign addr[44038]= -1197050035;
assign addr[44039]= -1438083551;
assign addr[44040]= -1649974225;
assign addr[44041]= -1828428082;
assign addr[44042]= -1969828744;
assign addr[44043]= -2071310720;
assign addr[44044]= -2130817471;
assign addr[44045]= -2147143090;
assign addr[44046]= -2119956737;
assign addr[44047]= -2049809346;
assign addr[44048]= -1938122457;
assign addr[44049]= -1787159411;
assign addr[44050]= -1599979481;
assign addr[44051]= -1380375881;
assign addr[44052]= -1132798888;
assign addr[44053]= -862265664;
assign addr[44054]= -574258580;
assign addr[44055]= -274614114;
assign addr[44056]= 30595422;
assign addr[44057]= 335184940;
assign addr[44058]= 632981917;
assign addr[44059]= 917951481;
assign addr[44060]= 1184318708;
assign addr[44061]= 1426685652;
assign addr[44062]= 1640140734;
assign addr[44063]= 1820358275;
assign addr[44064]= 1963686155;
assign addr[44065]= 2067219829;
assign addr[44066]= 2128861181;
assign addr[44067]= 2147361045;
assign addr[44068]= 2122344521;
assign addr[44069]= 2054318569;
assign addr[44070]= 1944661739;
assign addr[44071]= 1795596234;
assign addr[44072]= 1610142873;
assign addr[44073]= 1392059879;
assign addr[44074]= 1145766716;
assign addr[44075]= 876254528;
assign addr[44076]= 588984994;
assign addr[44077]= 289779648;
assign addr[44078]= -15298099;
assign addr[44079]= -320065829;
assign addr[44080]= -618347408;
assign addr[44081]= -904098143;
assign addr[44082]= -1171527280;
assign addr[44083]= -1415215352;
assign addr[44084]= -1630224009;
assign addr[44085]= -1812196087;
assign addr[44086]= -1957443913;
assign addr[44087]= -2063024031;
assign addr[44088]= -2126796855;
assign addr[44089]= -2147470025;
assign addr[44090]= -2124624598;
assign addr[44091]= -2058723538;
assign addr[44092]= -1951102334;
assign addr[44093]= -1803941934;
assign addr[44094]= -1620224553;
assign addr[44095]= -1403673233;
assign addr[44096]= -1158676398;
assign addr[44097]= -890198924;
assign addr[44098]= -603681519;
assign addr[44099]= -304930476;
assign addr[44100]= 0;
assign addr[44101]= 304930476;
assign addr[44102]= 603681519;
assign addr[44103]= 890198924;
assign addr[44104]= 1158676398;
assign addr[44105]= 1403673233;
assign addr[44106]= 1620224553;
assign addr[44107]= 1803941934;
assign addr[44108]= 1951102334;
assign addr[44109]= 2058723538;
assign addr[44110]= 2124624598;
assign addr[44111]= 2147470025;
assign addr[44112]= 2126796855;
assign addr[44113]= 2063024031;
assign addr[44114]= 1957443913;
assign addr[44115]= 1812196087;
assign addr[44116]= 1630224009;
assign addr[44117]= 1415215352;
assign addr[44118]= 1171527280;
assign addr[44119]= 904098143;
assign addr[44120]= 618347408;
assign addr[44121]= 320065829;
assign addr[44122]= 15298099;
assign addr[44123]= -289779648;
assign addr[44124]= -588984994;
assign addr[44125]= -876254528;
assign addr[44126]= -1145766716;
assign addr[44127]= -1392059879;
assign addr[44128]= -1610142873;
assign addr[44129]= -1795596234;
assign addr[44130]= -1944661739;
assign addr[44131]= -2054318569;
assign addr[44132]= -2122344521;
assign addr[44133]= -2147361045;
assign addr[44134]= -2128861181;
assign addr[44135]= -2067219829;
assign addr[44136]= -1963686155;
assign addr[44137]= -1820358275;
assign addr[44138]= -1640140734;
assign addr[44139]= -1426685652;
assign addr[44140]= -1184318708;
assign addr[44141]= -917951481;
assign addr[44142]= -632981917;
assign addr[44143]= -335184940;
assign addr[44144]= -30595422;
assign addr[44145]= 274614114;
assign addr[44146]= 574258580;
assign addr[44147]= 862265664;
assign addr[44148]= 1132798888;
assign addr[44149]= 1380375881;
assign addr[44150]= 1599979481;
assign addr[44151]= 1787159411;
assign addr[44152]= 1938122457;
assign addr[44153]= 2049809346;
assign addr[44154]= 2119956737;
assign addr[44155]= 2147143090;
assign addr[44156]= 2130817471;
assign addr[44157]= 2071310720;
assign addr[44158]= 1969828744;
assign addr[44159]= 1828428082;
assign addr[44160]= 1649974225;
assign addr[44161]= 1438083551;
assign addr[44162]= 1197050035;
assign addr[44163]= 931758235;
assign addr[44164]= 647584304;
assign addr[44165]= 350287041;
assign addr[44166]= 45891193;
assign addr[44167]= -259434643;
assign addr[44168]= -559503022;
assign addr[44169]= -848233042;
assign addr[44170]= -1119773573;
assign addr[44171]= -1368621831;
assign addr[44172]= -1589734894;
assign addr[44173]= -1778631892;
assign addr[44174]= -1931484818;
assign addr[44175]= -2045196100;
assign addr[44176]= -2117461370;
assign addr[44177]= -2146816171;
assign addr[44178]= -2132665626;
assign addr[44179]= -2075296495;
assign addr[44180]= -1975871368;
assign addr[44181]= -1836405100;
assign addr[44182]= -1659723983;
assign addr[44183]= -1449408469;
assign addr[44184]= -1209720613;
assign addr[44185]= -945517704;
assign addr[44186]= -662153826;
assign addr[44187]= -365371365;
assign addr[44188]= -61184634;
assign addr[44189]= 244242007;
assign addr[44190]= 544719071;
assign addr[44191]= 834157373;
assign addr[44192]= 1106691431;
assign addr[44193]= 1356798326;
assign addr[44194]= 1579409630;
assign addr[44195]= 1770014111;
assign addr[44196]= 1924749160;
assign addr[44197]= 2040479063;
assign addr[44198]= 2114858546;
assign addr[44199]= 2146380306;
assign addr[44200]= 2134405552;
assign addr[44201]= 2079176953;
assign addr[44202]= 1981813720;
assign addr[44203]= 1844288924;
assign addr[44204]= 1669389513;
assign addr[44205]= 1460659832;
assign addr[44206]= 1222329801;
assign addr[44207]= 959229189;
assign addr[44208]= 676689746;
assign addr[44209]= 380437148;
assign addr[44210]= 76474970;
assign addr[44211]= -229036977;
assign addr[44212]= -529907477;
assign addr[44213]= -820039373;
assign addr[44214]= -1093553126;
assign addr[44215]= -1344905966;
assign addr[44216]= -1569004214;
assign addr[44217]= -1761306505;
assign addr[44218]= -1917915825;
assign addr[44219]= -2035658475;
assign addr[44220]= -2112148396;
assign addr[44221]= -2145835515;
assign addr[44222]= -2136037160;
assign addr[44223]= -2082951896;
assign addr[44224]= -1987655498;
assign addr[44225]= -1852079154;
assign addr[44226]= -1678970324;
assign addr[44227]= -1471837070;
assign addr[44228]= -1234876957;
assign addr[44229]= -972891995;
assign addr[44230]= -691191324;
assign addr[44231]= -395483624;
assign addr[44232]= -91761426;
assign addr[44233]= 213820322;
assign addr[44234]= 515068990;
assign addr[44235]= 805879757;
assign addr[44236]= 1080359326;
assign addr[44237]= 1332945355;
assign addr[44238]= 1558519173;
assign addr[44239]= 1752509516;
assign addr[44240]= 1910985158;
assign addr[44241]= 2030734582;
assign addr[44242]= 2109331059;
assign addr[44243]= 2145181827;
assign addr[44244]= 2137560369;
assign addr[44245]= 2086621133;
assign addr[44246]= 1993396407;
assign addr[44247]= 1859775393;
assign addr[44248]= 1688465931;
assign addr[44249]= 1482939614;
assign addr[44250]= 1247361445;
assign addr[44251]= 986505429;
assign addr[44252]= 705657826;
assign addr[44253]= 410510029;
assign addr[44254]= 107043224;
assign addr[44255]= -198592817;
assign addr[44256]= -500204365;
assign addr[44257]= -791679244;
assign addr[44258]= -1067110699;
assign addr[44259]= -1320917099;
assign addr[44260]= -1547955041;
assign addr[44261]= -1743623590;
assign addr[44262]= -1903957513;
assign addr[44263]= -2025707632;
assign addr[44264]= -2106406677;
assign addr[44265]= -2144419275;
assign addr[44266]= -2138975100;
assign addr[44267]= -2090184478;
assign addr[44268]= -1999036154;
assign addr[44269]= -1867377253;
assign addr[44270]= -1697875851;
assign addr[44271]= -1493966902;
assign addr[44272]= -1259782632;
assign addr[44273]= -1000068799;
assign addr[44274]= -720088517;
assign addr[44275]= -425515602;
assign addr[44276]= -122319591;
assign addr[44277]= 183355234;
assign addr[44278]= 485314355;
assign addr[44279]= 777438554;
assign addr[44280]= 1053807919;
assign addr[44281]= 1308821808;
assign addr[44282]= 1537312353;
assign addr[44283]= 1734649179;
assign addr[44284]= 1896833245;
assign addr[44285]= 2020577882;
assign addr[44286]= 2103375398;
assign addr[44287]= 2143547897;
assign addr[44288]= 2140281282;
assign addr[44289]= 2093641749;
assign addr[44290]= 2004574453;
assign addr[44291]= 1874884346;
assign addr[44292]= 1707199606;
assign addr[44293]= 1504918373;
assign addr[44294]= 1272139887;
assign addr[44295]= 1013581418;
assign addr[44296]= 734482665;
assign addr[44297]= 440499581;
assign addr[44298]= 137589750;
assign addr[44299]= -168108346;
assign addr[44300]= -470399716;
assign addr[44301]= -763158411;
assign addr[44302]= -1040451659;
assign addr[44303]= -1296660098;
assign addr[44304]= -1526591649;
assign addr[44305]= -1725586737;
assign addr[44306]= -1889612716;
assign addr[44307]= -2015345591;
assign addr[44308]= -2100237377;
assign addr[44309]= -2142567738;
assign addr[44310]= -2141478848;
assign addr[44311]= -2096992772;
assign addr[44312]= -2010011024;
assign addr[44313]= -1882296293;
assign addr[44314]= -1716436725;
assign addr[44315]= -1515793473;
assign addr[44316]= -1284432584;
assign addr[44317]= -1027042599;
assign addr[44318]= -748839539;
assign addr[44319]= -455461206;
assign addr[44320]= -152852926;
assign addr[44321]= 152852926;
assign addr[44322]= 455461206;
assign addr[44323]= 748839539;
assign addr[44324]= 1027042599;
assign addr[44325]= 1284432584;
assign addr[44326]= 1515793473;
assign addr[44327]= 1716436725;
assign addr[44328]= 1882296293;
assign addr[44329]= 2010011024;
assign addr[44330]= 2096992772;
assign addr[44331]= 2141478848;
assign addr[44332]= 2142567738;
assign addr[44333]= 2100237377;
assign addr[44334]= 2015345591;
assign addr[44335]= 1889612716;
assign addr[44336]= 1725586737;
assign addr[44337]= 1526591649;
assign addr[44338]= 1296660098;
assign addr[44339]= 1040451659;
assign addr[44340]= 763158411;
assign addr[44341]= 470399716;
assign addr[44342]= 168108346;
assign addr[44343]= -137589750;
assign addr[44344]= -440499581;
assign addr[44345]= -734482665;
assign addr[44346]= -1013581418;
assign addr[44347]= -1272139887;
assign addr[44348]= -1504918373;
assign addr[44349]= -1707199606;
assign addr[44350]= -1874884346;
assign addr[44351]= -2004574453;
assign addr[44352]= -2093641749;
assign addr[44353]= -2140281282;
assign addr[44354]= -2143547897;
assign addr[44355]= -2103375398;
assign addr[44356]= -2020577882;
assign addr[44357]= -1896833245;
assign addr[44358]= -1734649179;
assign addr[44359]= -1537312353;
assign addr[44360]= -1308821808;
assign addr[44361]= -1053807919;
assign addr[44362]= -777438554;
assign addr[44363]= -485314355;
assign addr[44364]= -183355234;
assign addr[44365]= 122319591;
assign addr[44366]= 425515602;
assign addr[44367]= 720088517;
assign addr[44368]= 1000068799;
assign addr[44369]= 1259782632;
assign addr[44370]= 1493966902;
assign addr[44371]= 1697875851;
assign addr[44372]= 1867377253;
assign addr[44373]= 1999036154;
assign addr[44374]= 2090184478;
assign addr[44375]= 2138975100;
assign addr[44376]= 2144419275;
assign addr[44377]= 2106406677;
assign addr[44378]= 2025707632;
assign addr[44379]= 1903957513;
assign addr[44380]= 1743623590;
assign addr[44381]= 1547955041;
assign addr[44382]= 1320917099;
assign addr[44383]= 1067110699;
assign addr[44384]= 791679244;
assign addr[44385]= 500204365;
assign addr[44386]= 198592817;
assign addr[44387]= -107043224;
assign addr[44388]= -410510029;
assign addr[44389]= -705657826;
assign addr[44390]= -986505429;
assign addr[44391]= -1247361445;
assign addr[44392]= -1482939614;
assign addr[44393]= -1688465931;
assign addr[44394]= -1859775393;
assign addr[44395]= -1993396407;
assign addr[44396]= -2086621133;
assign addr[44397]= -2137560369;
assign addr[44398]= -2145181827;
assign addr[44399]= -2109331059;
assign addr[44400]= -2030734582;
assign addr[44401]= -1910985158;
assign addr[44402]= -1752509516;
assign addr[44403]= -1558519173;
assign addr[44404]= -1332945355;
assign addr[44405]= -1080359326;
assign addr[44406]= -805879757;
assign addr[44407]= -515068990;
assign addr[44408]= -213820322;
assign addr[44409]= 91761426;
assign addr[44410]= 395483624;
assign addr[44411]= 691191324;
assign addr[44412]= 972891995;
assign addr[44413]= 1234876957;
assign addr[44414]= 1471837070;
assign addr[44415]= 1678970324;
assign addr[44416]= 1852079154;
assign addr[44417]= 1987655498;
assign addr[44418]= 2082951896;
assign addr[44419]= 2136037160;
assign addr[44420]= 2145835515;
assign addr[44421]= 2112148396;
assign addr[44422]= 2035658475;
assign addr[44423]= 1917915825;
assign addr[44424]= 1761306505;
assign addr[44425]= 1569004214;
assign addr[44426]= 1344905966;
assign addr[44427]= 1093553126;
assign addr[44428]= 820039373;
assign addr[44429]= 529907477;
assign addr[44430]= 229036977;
assign addr[44431]= -76474970;
assign addr[44432]= -380437148;
assign addr[44433]= -676689746;
assign addr[44434]= -959229189;
assign addr[44435]= -1222329801;
assign addr[44436]= -1460659832;
assign addr[44437]= -1669389513;
assign addr[44438]= -1844288924;
assign addr[44439]= -1981813720;
assign addr[44440]= -2079176953;
assign addr[44441]= -2134405552;
assign addr[44442]= -2146380306;
assign addr[44443]= -2114858546;
assign addr[44444]= -2040479063;
assign addr[44445]= -1924749160;
assign addr[44446]= -1770014111;
assign addr[44447]= -1579409630;
assign addr[44448]= -1356798326;
assign addr[44449]= -1106691431;
assign addr[44450]= -834157373;
assign addr[44451]= -544719071;
assign addr[44452]= -244242007;
assign addr[44453]= 61184634;
assign addr[44454]= 365371365;
assign addr[44455]= 662153826;
assign addr[44456]= 945517704;
assign addr[44457]= 1209720613;
assign addr[44458]= 1449408469;
assign addr[44459]= 1659723983;
assign addr[44460]= 1836405100;
assign addr[44461]= 1975871368;
assign addr[44462]= 2075296495;
assign addr[44463]= 2132665626;
assign addr[44464]= 2146816171;
assign addr[44465]= 2117461370;
assign addr[44466]= 2045196100;
assign addr[44467]= 1931484818;
assign addr[44468]= 1778631892;
assign addr[44469]= 1589734894;
assign addr[44470]= 1368621831;
assign addr[44471]= 1119773573;
assign addr[44472]= 848233042;
assign addr[44473]= 559503022;
assign addr[44474]= 259434643;
assign addr[44475]= -45891193;
assign addr[44476]= -350287041;
assign addr[44477]= -647584304;
assign addr[44478]= -931758235;
assign addr[44479]= -1197050035;
assign addr[44480]= -1438083551;
assign addr[44481]= -1649974225;
assign addr[44482]= -1828428082;
assign addr[44483]= -1969828744;
assign addr[44484]= -2071310720;
assign addr[44485]= -2130817471;
assign addr[44486]= -2147143090;
assign addr[44487]= -2119956737;
assign addr[44488]= -2049809346;
assign addr[44489]= -1938122457;
assign addr[44490]= -1787159411;
assign addr[44491]= -1599979481;
assign addr[44492]= -1380375881;
assign addr[44493]= -1132798888;
assign addr[44494]= -862265664;
assign addr[44495]= -574258580;
assign addr[44496]= -274614114;
assign addr[44497]= 30595422;
assign addr[44498]= 335184940;
assign addr[44499]= 632981917;
assign addr[44500]= 917951481;
assign addr[44501]= 1184318708;
assign addr[44502]= 1426685652;
assign addr[44503]= 1640140734;
assign addr[44504]= 1820358275;
assign addr[44505]= 1963686155;
assign addr[44506]= 2067219829;
assign addr[44507]= 2128861181;
assign addr[44508]= 2147361045;
assign addr[44509]= 2122344521;
assign addr[44510]= 2054318569;
assign addr[44511]= 1944661739;
assign addr[44512]= 1795596234;
assign addr[44513]= 1610142873;
assign addr[44514]= 1392059879;
assign addr[44515]= 1145766716;
assign addr[44516]= 876254528;
assign addr[44517]= 588984994;
assign addr[44518]= 289779648;
assign addr[44519]= -15298099;
assign addr[44520]= -320065829;
assign addr[44521]= -618347408;
assign addr[44522]= -904098143;
assign addr[44523]= -1171527280;
assign addr[44524]= -1415215352;
assign addr[44525]= -1630224009;
assign addr[44526]= -1812196087;
assign addr[44527]= -1957443913;
assign addr[44528]= -2063024031;
assign addr[44529]= -2126796855;
assign addr[44530]= -2147470025;
assign addr[44531]= -2124624598;
assign addr[44532]= -2058723538;
assign addr[44533]= -1951102334;
assign addr[44534]= -1803941934;
assign addr[44535]= -1620224553;
assign addr[44536]= -1403673233;
assign addr[44537]= -1158676398;
assign addr[44538]= -890198924;
assign addr[44539]= -603681519;
assign addr[44540]= -304930476;
assign addr[44541]= 0;
assign addr[44542]= 304930476;
assign addr[44543]= 603681519;
assign addr[44544]= 890198924;
assign addr[44545]= 1158676398;
assign addr[44546]= 1403673233;
assign addr[44547]= 1620224553;
assign addr[44548]= 1803941934;
assign addr[44549]= 1951102334;
assign addr[44550]= 2058723538;
assign addr[44551]= 2124624598;
assign addr[44552]= 2147470025;
assign addr[44553]= 2126796855;
assign addr[44554]= 2063024031;
assign addr[44555]= 1957443913;
assign addr[44556]= 1812196087;
assign addr[44557]= 1630224009;
assign addr[44558]= 1415215352;
assign addr[44559]= 1171527280;
assign addr[44560]= 904098143;
assign addr[44561]= 618347408;
assign addr[44562]= 320065829;
assign addr[44563]= 15298099;
assign addr[44564]= -289779648;
assign addr[44565]= -588984994;
assign addr[44566]= -876254528;
assign addr[44567]= -1145766716;
assign addr[44568]= -1392059879;
assign addr[44569]= -1610142873;
assign addr[44570]= -1795596234;
assign addr[44571]= -1944661739;
assign addr[44572]= -2054318569;
assign addr[44573]= -2122344521;
assign addr[44574]= -2147361045;
assign addr[44575]= -2128861181;
assign addr[44576]= -2067219829;
assign addr[44577]= -1963686155;
assign addr[44578]= -1820358275;
assign addr[44579]= -1640140734;
assign addr[44580]= -1426685652;
assign addr[44581]= -1184318708;
assign addr[44582]= -917951481;
assign addr[44583]= -632981917;
assign addr[44584]= -335184940;
assign addr[44585]= -30595422;
assign addr[44586]= 274614114;
assign addr[44587]= 574258580;
assign addr[44588]= 862265664;
assign addr[44589]= 1132798888;
assign addr[44590]= 1380375881;
assign addr[44591]= 1599979481;
assign addr[44592]= 1787159411;
assign addr[44593]= 1938122457;
assign addr[44594]= 2049809346;
assign addr[44595]= 2119956737;
assign addr[44596]= 2147143090;
assign addr[44597]= 2130817471;
assign addr[44598]= 2071310720;
assign addr[44599]= 1969828744;
assign addr[44600]= 1828428082;
assign addr[44601]= 1649974225;
assign addr[44602]= 1438083551;
assign addr[44603]= 1197050035;
assign addr[44604]= 931758235;
assign addr[44605]= 647584304;
assign addr[44606]= 350287041;
assign addr[44607]= 45891193;
assign addr[44608]= -259434643;
assign addr[44609]= -559503022;
assign addr[44610]= -848233042;
assign addr[44611]= -1119773573;
assign addr[44612]= -1368621831;
assign addr[44613]= -1589734894;
assign addr[44614]= -1778631892;
assign addr[44615]= -1931484818;
assign addr[44616]= -2045196100;
assign addr[44617]= -2117461370;
assign addr[44618]= -2146816171;
assign addr[44619]= -2132665626;
assign addr[44620]= -2075296495;
assign addr[44621]= -1975871368;
assign addr[44622]= -1836405100;
assign addr[44623]= -1659723983;
assign addr[44624]= -1449408469;
assign addr[44625]= -1209720613;
assign addr[44626]= -945517704;
assign addr[44627]= -662153826;
assign addr[44628]= -365371365;
assign addr[44629]= -61184634;
assign addr[44630]= 244242007;
assign addr[44631]= 544719071;
assign addr[44632]= 834157373;
assign addr[44633]= 1106691431;
assign addr[44634]= 1356798326;
assign addr[44635]= 1579409630;
assign addr[44636]= 1770014111;
assign addr[44637]= 1924749160;
assign addr[44638]= 2040479063;
assign addr[44639]= 2114858546;
assign addr[44640]= 2146380306;
assign addr[44641]= 2134405552;
assign addr[44642]= 2079176953;
assign addr[44643]= 1981813720;
assign addr[44644]= 1844288924;
assign addr[44645]= 1669389513;
assign addr[44646]= 1460659832;
assign addr[44647]= 1222329801;
assign addr[44648]= 959229189;
assign addr[44649]= 676689746;
assign addr[44650]= 380437148;
assign addr[44651]= 76474970;
assign addr[44652]= -229036977;
assign addr[44653]= -529907477;
assign addr[44654]= -820039373;
assign addr[44655]= -1093553126;
assign addr[44656]= -1344905966;
assign addr[44657]= -1569004214;
assign addr[44658]= -1761306505;
assign addr[44659]= -1917915825;
assign addr[44660]= -2035658475;
assign addr[44661]= -2112148396;
assign addr[44662]= -2145835515;
assign addr[44663]= -2136037160;
assign addr[44664]= -2082951896;
assign addr[44665]= -1987655498;
assign addr[44666]= -1852079154;
assign addr[44667]= -1678970324;
assign addr[44668]= -1471837070;
assign addr[44669]= -1234876957;
assign addr[44670]= -972891995;
assign addr[44671]= -691191324;
assign addr[44672]= -395483624;
assign addr[44673]= -91761426;
assign addr[44674]= 213820322;
assign addr[44675]= 515068990;
assign addr[44676]= 805879757;
assign addr[44677]= 1080359326;
assign addr[44678]= 1332945355;
assign addr[44679]= 1558519173;
assign addr[44680]= 1752509516;
assign addr[44681]= 1910985158;
assign addr[44682]= 2030734582;
assign addr[44683]= 2109331059;
assign addr[44684]= 2145181827;
assign addr[44685]= 2137560369;
assign addr[44686]= 2086621133;
assign addr[44687]= 1993396407;
assign addr[44688]= 1859775393;
assign addr[44689]= 1688465931;
assign addr[44690]= 1482939614;
assign addr[44691]= 1247361445;
assign addr[44692]= 986505429;
assign addr[44693]= 705657826;
assign addr[44694]= 410510029;
assign addr[44695]= 107043224;
assign addr[44696]= -198592817;
assign addr[44697]= -500204365;
assign addr[44698]= -791679244;
assign addr[44699]= -1067110699;
assign addr[44700]= -1320917099;
assign addr[44701]= -1547955041;
assign addr[44702]= -1743623590;
assign addr[44703]= -1903957513;
assign addr[44704]= -2025707632;
assign addr[44705]= -2106406677;
assign addr[44706]= -2144419275;
assign addr[44707]= -2138975100;
assign addr[44708]= -2090184478;
assign addr[44709]= -1999036154;
assign addr[44710]= -1867377253;
assign addr[44711]= -1697875851;
assign addr[44712]= -1493966902;
assign addr[44713]= -1259782632;
assign addr[44714]= -1000068799;
assign addr[44715]= -720088517;
assign addr[44716]= -425515602;
assign addr[44717]= -122319591;
assign addr[44718]= 183355234;
assign addr[44719]= 485314355;
assign addr[44720]= 777438554;
assign addr[44721]= 1053807919;
assign addr[44722]= 1308821808;
assign addr[44723]= 1537312353;
assign addr[44724]= 1734649179;
assign addr[44725]= 1896833245;
assign addr[44726]= 2020577882;
assign addr[44727]= 2103375398;
assign addr[44728]= 2143547897;
assign addr[44729]= 2140281282;
assign addr[44730]= 2093641749;
assign addr[44731]= 2004574453;
assign addr[44732]= 1874884346;
assign addr[44733]= 1707199606;
assign addr[44734]= 1504918373;
assign addr[44735]= 1272139887;
assign addr[44736]= 1013581418;
assign addr[44737]= 734482665;
assign addr[44738]= 440499581;
assign addr[44739]= 137589750;
assign addr[44740]= -168108346;
assign addr[44741]= -470399716;
assign addr[44742]= -763158411;
assign addr[44743]= -1040451659;
assign addr[44744]= -1296660098;
assign addr[44745]= -1526591649;
assign addr[44746]= -1725586737;
assign addr[44747]= -1889612716;
assign addr[44748]= -2015345591;
assign addr[44749]= -2100237377;
assign addr[44750]= -2142567738;
assign addr[44751]= -2141478848;
assign addr[44752]= -2096992772;
assign addr[44753]= -2010011024;
assign addr[44754]= -1882296293;
assign addr[44755]= -1716436725;
assign addr[44756]= -1515793473;
assign addr[44757]= -1284432584;
assign addr[44758]= -1027042599;
assign addr[44759]= -748839539;
assign addr[44760]= -455461206;
assign addr[44761]= -152852926;
assign addr[44762]= 152852926;
assign addr[44763]= 455461206;
assign addr[44764]= 748839539;
assign addr[44765]= 1027042599;
assign addr[44766]= 1284432584;
assign addr[44767]= 1515793473;
assign addr[44768]= 1716436725;
assign addr[44769]= 1882296293;
assign addr[44770]= 2010011024;
assign addr[44771]= 2096992772;
assign addr[44772]= 2141478848;
assign addr[44773]= 2142567738;
assign addr[44774]= 2100237377;
assign addr[44775]= 2015345591;
assign addr[44776]= 1889612716;
assign addr[44777]= 1725586737;
assign addr[44778]= 1526591649;
assign addr[44779]= 1296660098;
assign addr[44780]= 1040451659;
assign addr[44781]= 763158411;
assign addr[44782]= 470399716;
assign addr[44783]= 168108346;
assign addr[44784]= -137589750;
assign addr[44785]= -440499581;
assign addr[44786]= -734482665;
assign addr[44787]= -1013581418;
assign addr[44788]= -1272139887;
assign addr[44789]= -1504918373;
assign addr[44790]= -1707199606;
assign addr[44791]= -1874884346;
assign addr[44792]= -2004574453;
assign addr[44793]= -2093641749;
assign addr[44794]= -2140281282;
assign addr[44795]= -2143547897;
assign addr[44796]= -2103375398;
assign addr[44797]= -2020577882;
assign addr[44798]= -1896833245;
assign addr[44799]= -1734649179;
assign addr[44800]= -1537312353;
assign addr[44801]= -1308821808;
assign addr[44802]= -1053807919;
assign addr[44803]= -777438554;
assign addr[44804]= -485314355;
assign addr[44805]= -183355234;
assign addr[44806]= 122319591;
assign addr[44807]= 425515602;
assign addr[44808]= 720088517;
assign addr[44809]= 1000068799;
assign addr[44810]= 1259782632;
assign addr[44811]= 1493966902;
assign addr[44812]= 1697875851;
assign addr[44813]= 1867377253;
assign addr[44814]= 1999036154;
assign addr[44815]= 2090184478;
assign addr[44816]= 2138975100;
assign addr[44817]= 2144419275;
assign addr[44818]= 2106406677;
assign addr[44819]= 2025707632;
assign addr[44820]= 1903957513;
assign addr[44821]= 1743623590;
assign addr[44822]= 1547955041;
assign addr[44823]= 1320917099;
assign addr[44824]= 1067110699;
assign addr[44825]= 791679244;
assign addr[44826]= 500204365;
assign addr[44827]= 198592817;
assign addr[44828]= -107043224;
assign addr[44829]= -410510029;
assign addr[44830]= -705657826;
assign addr[44831]= -986505429;
assign addr[44832]= -1247361445;
assign addr[44833]= -1482939614;
assign addr[44834]= -1688465931;
assign addr[44835]= -1859775393;
assign addr[44836]= -1993396407;
assign addr[44837]= -2086621133;
assign addr[44838]= -2137560369;
assign addr[44839]= -2145181827;
assign addr[44840]= -2109331059;
assign addr[44841]= -2030734582;
assign addr[44842]= -1910985158;
assign addr[44843]= -1752509516;
assign addr[44844]= -1558519173;
assign addr[44845]= -1332945355;
assign addr[44846]= -1080359326;
assign addr[44847]= -805879757;
assign addr[44848]= -515068990;
assign addr[44849]= -213820322;
assign addr[44850]= 91761426;
assign addr[44851]= 395483624;
assign addr[44852]= 691191324;
assign addr[44853]= 972891995;
assign addr[44854]= 1234876957;
assign addr[44855]= 1471837070;
assign addr[44856]= 1678970324;
assign addr[44857]= 1852079154;
assign addr[44858]= 1987655498;
assign addr[44859]= 2082951896;
assign addr[44860]= 2136037160;
assign addr[44861]= 2145835515;
assign addr[44862]= 2112148396;
assign addr[44863]= 2035658475;
assign addr[44864]= 1917915825;
assign addr[44865]= 1761306505;
assign addr[44866]= 1569004214;
assign addr[44867]= 1344905966;
assign addr[44868]= 1093553126;
assign addr[44869]= 820039373;
assign addr[44870]= 529907477;
assign addr[44871]= 229036977;
assign addr[44872]= -76474970;
assign addr[44873]= -380437148;
assign addr[44874]= -676689746;
assign addr[44875]= -959229189;
assign addr[44876]= -1222329801;
assign addr[44877]= -1460659832;
assign addr[44878]= -1669389513;
assign addr[44879]= -1844288924;
assign addr[44880]= -1981813720;
assign addr[44881]= -2079176953;
assign addr[44882]= -2134405552;
assign addr[44883]= -2146380306;
assign addr[44884]= -2114858546;
assign addr[44885]= -2040479063;
assign addr[44886]= -1924749160;
assign addr[44887]= -1770014111;
assign addr[44888]= -1579409630;
assign addr[44889]= -1356798326;
assign addr[44890]= -1106691431;
assign addr[44891]= -834157373;
assign addr[44892]= -544719071;
assign addr[44893]= -244242007;
assign addr[44894]= 61184634;
assign addr[44895]= 365371365;
assign addr[44896]= 662153826;
assign addr[44897]= 945517704;
assign addr[44898]= 1209720613;
assign addr[44899]= 1449408469;
assign addr[44900]= 1659723983;
assign addr[44901]= 1836405100;
assign addr[44902]= 1975871368;
assign addr[44903]= 2075296495;
assign addr[44904]= 2132665626;
assign addr[44905]= 2146816171;
assign addr[44906]= 2117461370;
assign addr[44907]= 2045196100;
assign addr[44908]= 1931484818;
assign addr[44909]= 1778631892;
assign addr[44910]= 1589734894;
assign addr[44911]= 1368621831;
assign addr[44912]= 1119773573;
assign addr[44913]= 848233042;
assign addr[44914]= 559503022;
assign addr[44915]= 259434643;
assign addr[44916]= -45891193;
assign addr[44917]= -350287041;
assign addr[44918]= -647584304;
assign addr[44919]= -931758235;
assign addr[44920]= -1197050035;
assign addr[44921]= -1438083551;
assign addr[44922]= -1649974225;
assign addr[44923]= -1828428082;
assign addr[44924]= -1969828744;
assign addr[44925]= -2071310720;
assign addr[44926]= -2130817471;
assign addr[44927]= -2147143090;
assign addr[44928]= -2119956737;
assign addr[44929]= -2049809346;
assign addr[44930]= -1938122457;
assign addr[44931]= -1787159411;
assign addr[44932]= -1599979481;
assign addr[44933]= -1380375881;
assign addr[44934]= -1132798888;
assign addr[44935]= -862265664;
assign addr[44936]= -574258580;
assign addr[44937]= -274614114;
assign addr[44938]= 30595422;
assign addr[44939]= 335184940;
assign addr[44940]= 632981917;
assign addr[44941]= 917951481;
assign addr[44942]= 1184318708;
assign addr[44943]= 1426685652;
assign addr[44944]= 1640140734;
assign addr[44945]= 1820358275;
assign addr[44946]= 1963686155;
assign addr[44947]= 2067219829;
assign addr[44948]= 2128861181;
assign addr[44949]= 2147361045;
assign addr[44950]= 2122344521;
assign addr[44951]= 2054318569;
assign addr[44952]= 1944661739;
assign addr[44953]= 1795596234;
assign addr[44954]= 1610142873;
assign addr[44955]= 1392059879;
assign addr[44956]= 1145766716;
assign addr[44957]= 876254528;
assign addr[44958]= 588984994;
assign addr[44959]= 289779648;
assign addr[44960]= -15298099;
assign addr[44961]= -320065829;
assign addr[44962]= -618347408;
assign addr[44963]= -904098143;
assign addr[44964]= -1171527280;
assign addr[44965]= -1415215352;
assign addr[44966]= -1630224009;
assign addr[44967]= -1812196087;
assign addr[44968]= -1957443913;
assign addr[44969]= -2063024031;
assign addr[44970]= -2126796855;
assign addr[44971]= -2147470025;
assign addr[44972]= -2124624598;
assign addr[44973]= -2058723538;
assign addr[44974]= -1951102334;
assign addr[44975]= -1803941934;
assign addr[44976]= -1620224553;
assign addr[44977]= -1403673233;
assign addr[44978]= -1158676398;
assign addr[44979]= -890198924;
assign addr[44980]= -603681519;
assign addr[44981]= -304930476;
assign addr[44982]= 0;
assign addr[44983]= 304930476;
assign addr[44984]= 603681519;
assign addr[44985]= 890198924;
assign addr[44986]= 1158676398;
assign addr[44987]= 1403673233;
assign addr[44988]= 1620224553;
assign addr[44989]= 1803941934;
assign addr[44990]= 1951102334;
assign addr[44991]= 2058723538;
assign addr[44992]= 2124624598;
assign addr[44993]= 2147470025;
assign addr[44994]= 2126796855;
assign addr[44995]= 2063024031;
assign addr[44996]= 1957443913;
assign addr[44997]= 1812196087;
assign addr[44998]= 1630224009;
assign addr[44999]= 1415215352;
assign addr[45000]= 1171527280;
assign addr[45001]= 904098143;
assign addr[45002]= 618347408;
assign addr[45003]= 320065829;
assign addr[45004]= 15298099;
assign addr[45005]= -289779648;
assign addr[45006]= -588984994;
assign addr[45007]= -876254528;
assign addr[45008]= -1145766716;
assign addr[45009]= -1392059879;
assign addr[45010]= -1610142873;
assign addr[45011]= -1795596234;
assign addr[45012]= -1944661739;
assign addr[45013]= -2054318569;
assign addr[45014]= -2122344521;
assign addr[45015]= -2147361045;
assign addr[45016]= -2128861181;
assign addr[45017]= -2067219829;
assign addr[45018]= -1963686155;
assign addr[45019]= -1820358275;
assign addr[45020]= -1640140734;
assign addr[45021]= -1426685652;
assign addr[45022]= -1184318708;
assign addr[45023]= -917951481;
assign addr[45024]= -632981917;
assign addr[45025]= -335184940;
assign addr[45026]= -30595422;
assign addr[45027]= 274614114;
assign addr[45028]= 574258580;
assign addr[45029]= 862265664;
assign addr[45030]= 1132798888;
assign addr[45031]= 1380375881;
assign addr[45032]= 1599979481;
assign addr[45033]= 1787159411;
assign addr[45034]= 1938122457;
assign addr[45035]= 2049809346;
assign addr[45036]= 2119956737;
assign addr[45037]= 2147143090;
assign addr[45038]= 2130817471;
assign addr[45039]= 2071310720;
assign addr[45040]= 1969828744;
assign addr[45041]= 1828428082;
assign addr[45042]= 1649974225;
assign addr[45043]= 1438083551;
assign addr[45044]= 1197050035;
assign addr[45045]= 931758235;
assign addr[45046]= 647584304;
assign addr[45047]= 350287041;
assign addr[45048]= 45891193;
assign addr[45049]= -259434643;
assign addr[45050]= -559503022;
assign addr[45051]= -848233042;
assign addr[45052]= -1119773573;
assign addr[45053]= -1368621831;
assign addr[45054]= -1589734894;
assign addr[45055]= -1778631892;
assign addr[45056]= -1931484818;
assign addr[45057]= -2045196100;
assign addr[45058]= -2117461370;
assign addr[45059]= -2146816171;
assign addr[45060]= -2132665626;
assign addr[45061]= -2075296495;
assign addr[45062]= -1975871368;
assign addr[45063]= -1836405100;
assign addr[45064]= -1659723983;
assign addr[45065]= -1449408469;
assign addr[45066]= -1209720613;
assign addr[45067]= -945517704;
assign addr[45068]= -662153826;
assign addr[45069]= -365371365;
assign addr[45070]= -61184634;
assign addr[45071]= 244242007;
assign addr[45072]= 544719071;
assign addr[45073]= 834157373;
assign addr[45074]= 1106691431;
assign addr[45075]= 1356798326;
assign addr[45076]= 1579409630;
assign addr[45077]= 1770014111;
assign addr[45078]= 1924749160;
assign addr[45079]= 2040479063;
assign addr[45080]= 2114858546;
assign addr[45081]= 2146380306;
assign addr[45082]= 2134405552;
assign addr[45083]= 2079176953;
assign addr[45084]= 1981813720;
assign addr[45085]= 1844288924;
assign addr[45086]= 1669389513;
assign addr[45087]= 1460659832;
assign addr[45088]= 1222329801;
assign addr[45089]= 959229189;
assign addr[45090]= 676689746;
assign addr[45091]= 380437148;
assign addr[45092]= 76474970;
assign addr[45093]= -229036977;
assign addr[45094]= -529907477;
assign addr[45095]= -820039373;
assign addr[45096]= -1093553126;
assign addr[45097]= -1344905966;
assign addr[45098]= -1569004214;
assign addr[45099]= -1761306505;
assign addr[45100]= -1917915825;
assign addr[45101]= -2035658475;
assign addr[45102]= -2112148396;
assign addr[45103]= -2145835515;
assign addr[45104]= -2136037160;
assign addr[45105]= -2082951896;
assign addr[45106]= -1987655498;
assign addr[45107]= -1852079154;
assign addr[45108]= -1678970324;
assign addr[45109]= -1471837070;
assign addr[45110]= -1234876957;
assign addr[45111]= -972891995;
assign addr[45112]= -691191324;
assign addr[45113]= -395483624;
assign addr[45114]= -91761426;
assign addr[45115]= 213820322;
assign addr[45116]= 515068990;
assign addr[45117]= 805879757;
assign addr[45118]= 1080359326;
assign addr[45119]= 1332945355;
assign addr[45120]= 1558519173;
assign addr[45121]= 1752509516;
assign addr[45122]= 1910985158;
assign addr[45123]= 2030734582;
assign addr[45124]= 2109331059;
assign addr[45125]= 2145181827;
assign addr[45126]= 2137560369;
assign addr[45127]= 2086621133;
assign addr[45128]= 1993396407;
assign addr[45129]= 1859775393;
assign addr[45130]= 1688465931;
assign addr[45131]= 1482939614;
assign addr[45132]= 1247361445;
assign addr[45133]= 986505429;
assign addr[45134]= 705657826;
assign addr[45135]= 410510029;
assign addr[45136]= 107043224;
assign addr[45137]= -198592817;
assign addr[45138]= -500204365;
assign addr[45139]= -791679244;
assign addr[45140]= -1067110699;
assign addr[45141]= -1320917099;
assign addr[45142]= -1547955041;
assign addr[45143]= -1743623590;
assign addr[45144]= -1903957513;
assign addr[45145]= -2025707632;
assign addr[45146]= -2106406677;
assign addr[45147]= -2144419275;
assign addr[45148]= -2138975100;
assign addr[45149]= -2090184478;
assign addr[45150]= -1999036154;
assign addr[45151]= -1867377253;
assign addr[45152]= -1697875851;
assign addr[45153]= -1493966902;
assign addr[45154]= -1259782632;
assign addr[45155]= -1000068799;
assign addr[45156]= -720088517;
assign addr[45157]= -425515602;
assign addr[45158]= -122319591;
assign addr[45159]= 183355234;
assign addr[45160]= 485314355;
assign addr[45161]= 777438554;
assign addr[45162]= 1053807919;
assign addr[45163]= 1308821808;
assign addr[45164]= 1537312353;
assign addr[45165]= 1734649179;
assign addr[45166]= 1896833245;
assign addr[45167]= 2020577882;
assign addr[45168]= 2103375398;
assign addr[45169]= 2143547897;
assign addr[45170]= 2140281282;
assign addr[45171]= 2093641749;
assign addr[45172]= 2004574453;
assign addr[45173]= 1874884346;
assign addr[45174]= 1707199606;
assign addr[45175]= 1504918373;
assign addr[45176]= 1272139887;
assign addr[45177]= 1013581418;
assign addr[45178]= 734482665;
assign addr[45179]= 440499581;
assign addr[45180]= 137589750;
assign addr[45181]= -168108346;
assign addr[45182]= -470399716;
assign addr[45183]= -763158411;
assign addr[45184]= -1040451659;
assign addr[45185]= -1296660098;
assign addr[45186]= -1526591649;
assign addr[45187]= -1725586737;
assign addr[45188]= -1889612716;
assign addr[45189]= -2015345591;
assign addr[45190]= -2100237377;
assign addr[45191]= -2142567738;
assign addr[45192]= -2141478848;
assign addr[45193]= -2096992772;
assign addr[45194]= -2010011024;
assign addr[45195]= -1882296293;
assign addr[45196]= -1716436725;
assign addr[45197]= -1515793473;
assign addr[45198]= -1284432584;
assign addr[45199]= -1027042599;
assign addr[45200]= -748839539;
assign addr[45201]= -455461206;
assign addr[45202]= -152852926;
assign addr[45203]= 152852926;
assign addr[45204]= 455461206;
assign addr[45205]= 748839539;
assign addr[45206]= 1027042599;
assign addr[45207]= 1284432584;
assign addr[45208]= 1515793473;
assign addr[45209]= 1716436725;
assign addr[45210]= 1882296293;
assign addr[45211]= 2010011024;
assign addr[45212]= 2096992772;
assign addr[45213]= 2141478848;
assign addr[45214]= 2142567738;
assign addr[45215]= 2100237377;
assign addr[45216]= 2015345591;
assign addr[45217]= 1889612716;
assign addr[45218]= 1725586737;
assign addr[45219]= 1526591649;
assign addr[45220]= 1296660098;
assign addr[45221]= 1040451659;
assign addr[45222]= 763158411;
assign addr[45223]= 470399716;
assign addr[45224]= 168108346;
assign addr[45225]= -137589750;
assign addr[45226]= -440499581;
assign addr[45227]= -734482665;
assign addr[45228]= -1013581418;
assign addr[45229]= -1272139887;
assign addr[45230]= -1504918373;
assign addr[45231]= -1707199606;
assign addr[45232]= -1874884346;
assign addr[45233]= -2004574453;
assign addr[45234]= -2093641749;
assign addr[45235]= -2140281282;
assign addr[45236]= -2143547897;
assign addr[45237]= -2103375398;
assign addr[45238]= -2020577882;
assign addr[45239]= -1896833245;
assign addr[45240]= -1734649179;
assign addr[45241]= -1537312353;
assign addr[45242]= -1308821808;
assign addr[45243]= -1053807919;
assign addr[45244]= -777438554;
assign addr[45245]= -485314355;
assign addr[45246]= -183355234;
assign addr[45247]= 122319591;
assign addr[45248]= 425515602;
assign addr[45249]= 720088517;
assign addr[45250]= 1000068799;
assign addr[45251]= 1259782632;
assign addr[45252]= 1493966902;
assign addr[45253]= 1697875851;
assign addr[45254]= 1867377253;
assign addr[45255]= 1999036154;
assign addr[45256]= 2090184478;
assign addr[45257]= 2138975100;
assign addr[45258]= 2144419275;
assign addr[45259]= 2106406677;
assign addr[45260]= 2025707632;
assign addr[45261]= 1903957513;
assign addr[45262]= 1743623590;
assign addr[45263]= 1547955041;
assign addr[45264]= 1320917099;
assign addr[45265]= 1067110699;
assign addr[45266]= 791679244;
assign addr[45267]= 500204365;
assign addr[45268]= 198592817;
assign addr[45269]= -107043224;
assign addr[45270]= -410510029;
assign addr[45271]= -705657826;
assign addr[45272]= -986505429;
assign addr[45273]= -1247361445;
assign addr[45274]= -1482939614;
assign addr[45275]= -1688465931;
assign addr[45276]= -1859775393;
assign addr[45277]= -1993396407;
assign addr[45278]= -2086621133;
assign addr[45279]= -2137560369;
assign addr[45280]= -2145181827;
assign addr[45281]= -2109331059;
assign addr[45282]= -2030734582;
assign addr[45283]= -1910985158;
assign addr[45284]= -1752509516;
assign addr[45285]= -1558519173;
assign addr[45286]= -1332945355;
assign addr[45287]= -1080359326;
assign addr[45288]= -805879757;
assign addr[45289]= -515068990;
assign addr[45290]= -213820322;
assign addr[45291]= 91761426;
assign addr[45292]= 395483624;
assign addr[45293]= 691191324;
assign addr[45294]= 972891995;
assign addr[45295]= 1234876957;
assign addr[45296]= 1471837070;
assign addr[45297]= 1678970324;
assign addr[45298]= 1852079154;
assign addr[45299]= 1987655498;
assign addr[45300]= 2082951896;
assign addr[45301]= 2136037160;
assign addr[45302]= 2145835515;
assign addr[45303]= 2112148396;
assign addr[45304]= 2035658475;
assign addr[45305]= 1917915825;
assign addr[45306]= 1761306505;
assign addr[45307]= 1569004214;
assign addr[45308]= 1344905966;
assign addr[45309]= 1093553126;
assign addr[45310]= 820039373;
assign addr[45311]= 529907477;
assign addr[45312]= 229036977;
assign addr[45313]= -76474970;
assign addr[45314]= -380437148;
assign addr[45315]= -676689746;
assign addr[45316]= -959229189;
assign addr[45317]= -1222329801;
assign addr[45318]= -1460659832;
assign addr[45319]= -1669389513;
assign addr[45320]= -1844288924;
assign addr[45321]= -1981813720;
assign addr[45322]= -2079176953;
assign addr[45323]= -2134405552;
assign addr[45324]= -2146380306;
assign addr[45325]= -2114858546;
assign addr[45326]= -2040479063;
assign addr[45327]= -1924749160;
assign addr[45328]= -1770014111;
assign addr[45329]= -1579409630;
assign addr[45330]= -1356798326;
assign addr[45331]= -1106691431;
assign addr[45332]= -834157373;
assign addr[45333]= -544719071;
assign addr[45334]= -244242007;
assign addr[45335]= 61184634;
assign addr[45336]= 365371365;
assign addr[45337]= 662153826;
assign addr[45338]= 945517704;
assign addr[45339]= 1209720613;
assign addr[45340]= 1449408469;
assign addr[45341]= 1659723983;
assign addr[45342]= 1836405100;
assign addr[45343]= 1975871368;
assign addr[45344]= 2075296495;
assign addr[45345]= 2132665626;
assign addr[45346]= 2146816171;
assign addr[45347]= 2117461370;
assign addr[45348]= 2045196100;
assign addr[45349]= 1931484818;
assign addr[45350]= 1778631892;
assign addr[45351]= 1589734894;
assign addr[45352]= 1368621831;
assign addr[45353]= 1119773573;
assign addr[45354]= 848233042;
assign addr[45355]= 559503022;
assign addr[45356]= 259434643;
assign addr[45357]= -45891193;
assign addr[45358]= -350287041;
assign addr[45359]= -647584304;
assign addr[45360]= -931758235;
assign addr[45361]= -1197050035;
assign addr[45362]= -1438083551;
assign addr[45363]= -1649974225;
assign addr[45364]= -1828428082;
assign addr[45365]= -1969828744;
assign addr[45366]= -2071310720;
assign addr[45367]= -2130817471;
assign addr[45368]= -2147143090;
assign addr[45369]= -2119956737;
assign addr[45370]= -2049809346;
assign addr[45371]= -1938122457;
assign addr[45372]= -1787159411;
assign addr[45373]= -1599979481;
assign addr[45374]= -1380375881;
assign addr[45375]= -1132798888;
assign addr[45376]= -862265664;
assign addr[45377]= -574258580;
assign addr[45378]= -274614114;
assign addr[45379]= 30595422;
assign addr[45380]= 335184940;
assign addr[45381]= 632981917;
assign addr[45382]= 917951481;
assign addr[45383]= 1184318708;
assign addr[45384]= 1426685652;
assign addr[45385]= 1640140734;
assign addr[45386]= 1820358275;
assign addr[45387]= 1963686155;
assign addr[45388]= 2067219829;
assign addr[45389]= 2128861181;
assign addr[45390]= 2147361045;
assign addr[45391]= 2122344521;
assign addr[45392]= 2054318569;
assign addr[45393]= 1944661739;
assign addr[45394]= 1795596234;
assign addr[45395]= 1610142873;
assign addr[45396]= 1392059879;
assign addr[45397]= 1145766716;
assign addr[45398]= 876254528;
assign addr[45399]= 588984994;
assign addr[45400]= 289779648;
assign addr[45401]= -15298099;
assign addr[45402]= -320065829;
assign addr[45403]= -618347408;
assign addr[45404]= -904098143;
assign addr[45405]= -1171527280;
assign addr[45406]= -1415215352;
assign addr[45407]= -1630224009;
assign addr[45408]= -1812196087;
assign addr[45409]= -1957443913;
assign addr[45410]= -2063024031;
assign addr[45411]= -2126796855;
assign addr[45412]= -2147470025;
assign addr[45413]= -2124624598;
assign addr[45414]= -2058723538;
assign addr[45415]= -1951102334;
assign addr[45416]= -1803941934;
assign addr[45417]= -1620224553;
assign addr[45418]= -1403673233;
assign addr[45419]= -1158676398;
assign addr[45420]= -890198924;
assign addr[45421]= -603681519;
assign addr[45422]= -304930476;
assign addr[45423]= 0;
assign addr[45424]= 304930476;
assign addr[45425]= 603681519;
assign addr[45426]= 890198924;
assign addr[45427]= 1158676398;
assign addr[45428]= 1403673233;
assign addr[45429]= 1620224553;
assign addr[45430]= 1803941934;
assign addr[45431]= 1951102334;
assign addr[45432]= 2058723538;
assign addr[45433]= 2124624598;
assign addr[45434]= 2147470025;
assign addr[45435]= 2126796855;
assign addr[45436]= 2063024031;
assign addr[45437]= 1957443913;
assign addr[45438]= 1812196087;
assign addr[45439]= 1630224009;
assign addr[45440]= 1415215352;
assign addr[45441]= 1171527280;
assign addr[45442]= 904098143;
assign addr[45443]= 618347408;
assign addr[45444]= 320065829;
assign addr[45445]= 15298099;
assign addr[45446]= -289779648;
assign addr[45447]= -588984994;
assign addr[45448]= -876254528;
assign addr[45449]= -1145766716;
assign addr[45450]= -1392059879;
assign addr[45451]= -1610142873;
assign addr[45452]= -1795596234;
assign addr[45453]= -1944661739;
assign addr[45454]= -2054318569;
assign addr[45455]= -2122344521;
assign addr[45456]= -2147361045;
assign addr[45457]= -2128861181;
assign addr[45458]= -2067219829;
assign addr[45459]= -1963686155;
assign addr[45460]= -1820358275;
assign addr[45461]= -1640140734;
assign addr[45462]= -1426685652;
assign addr[45463]= -1184318708;
assign addr[45464]= -917951481;
assign addr[45465]= -632981917;
assign addr[45466]= -335184940;
assign addr[45467]= -30595422;
assign addr[45468]= 274614114;
assign addr[45469]= 574258580;
assign addr[45470]= 862265664;
assign addr[45471]= 1132798888;
assign addr[45472]= 1380375881;
assign addr[45473]= 1599979481;
assign addr[45474]= 1787159411;
assign addr[45475]= 1938122457;
assign addr[45476]= 2049809346;
assign addr[45477]= 2119956737;
assign addr[45478]= 2147143090;
assign addr[45479]= 2130817471;
assign addr[45480]= 2071310720;
assign addr[45481]= 1969828744;
assign addr[45482]= 1828428082;
assign addr[45483]= 1649974225;
assign addr[45484]= 1438083551;
assign addr[45485]= 1197050035;
assign addr[45486]= 931758235;
assign addr[45487]= 647584304;
assign addr[45488]= 350287041;
assign addr[45489]= 45891193;
assign addr[45490]= -259434643;
assign addr[45491]= -559503022;
assign addr[45492]= -848233042;
assign addr[45493]= -1119773573;
assign addr[45494]= -1368621831;
assign addr[45495]= -1589734894;
assign addr[45496]= -1778631892;
assign addr[45497]= -1931484818;
assign addr[45498]= -2045196100;
assign addr[45499]= -2117461370;
assign addr[45500]= -2146816171;
assign addr[45501]= -2132665626;
assign addr[45502]= -2075296495;
assign addr[45503]= -1975871368;
assign addr[45504]= -1836405100;
assign addr[45505]= -1659723983;
assign addr[45506]= -1449408469;
assign addr[45507]= -1209720613;
assign addr[45508]= -945517704;
assign addr[45509]= -662153826;
assign addr[45510]= -365371365;
assign addr[45511]= -61184634;
assign addr[45512]= 244242007;
assign addr[45513]= 544719071;
assign addr[45514]= 834157373;
assign addr[45515]= 1106691431;
assign addr[45516]= 1356798326;
assign addr[45517]= 1579409630;
assign addr[45518]= 1770014111;
assign addr[45519]= 1924749160;
assign addr[45520]= 2040479063;
assign addr[45521]= 2114858546;
assign addr[45522]= 2146380306;
assign addr[45523]= 2134405552;
assign addr[45524]= 2079176953;
assign addr[45525]= 1981813720;
assign addr[45526]= 1844288924;
assign addr[45527]= 1669389513;
assign addr[45528]= 1460659832;
assign addr[45529]= 1222329801;
assign addr[45530]= 959229189;
assign addr[45531]= 676689746;
assign addr[45532]= 380437148;
assign addr[45533]= 76474970;
assign addr[45534]= -229036977;
assign addr[45535]= -529907477;
assign addr[45536]= -820039373;
assign addr[45537]= -1093553126;
assign addr[45538]= -1344905966;
assign addr[45539]= -1569004214;
assign addr[45540]= -1761306505;
assign addr[45541]= -1917915825;
assign addr[45542]= -2035658475;
assign addr[45543]= -2112148396;
assign addr[45544]= -2145835515;
assign addr[45545]= -2136037160;
assign addr[45546]= -2082951896;
assign addr[45547]= -1987655498;
assign addr[45548]= -1852079154;
assign addr[45549]= -1678970324;
assign addr[45550]= -1471837070;
assign addr[45551]= -1234876957;
assign addr[45552]= -972891995;
assign addr[45553]= -691191324;
assign addr[45554]= -395483624;
assign addr[45555]= -91761426;
assign addr[45556]= 213820322;
assign addr[45557]= 515068990;
assign addr[45558]= 805879757;
assign addr[45559]= 1080359326;
assign addr[45560]= 1332945355;
assign addr[45561]= 1558519173;
assign addr[45562]= 1752509516;
assign addr[45563]= 1910985158;
assign addr[45564]= 2030734582;
assign addr[45565]= 2109331059;
assign addr[45566]= 2145181827;
assign addr[45567]= 2137560369;
assign addr[45568]= 2086621133;
assign addr[45569]= 1993396407;
assign addr[45570]= 1859775393;
assign addr[45571]= 1688465931;
assign addr[45572]= 1482939614;
assign addr[45573]= 1247361445;
assign addr[45574]= 986505429;
assign addr[45575]= 705657826;
assign addr[45576]= 410510029;
assign addr[45577]= 107043224;
assign addr[45578]= -198592817;
assign addr[45579]= -500204365;
assign addr[45580]= -791679244;
assign addr[45581]= -1067110699;
assign addr[45582]= -1320917099;
assign addr[45583]= -1547955041;
assign addr[45584]= -1743623590;
assign addr[45585]= -1903957513;
assign addr[45586]= -2025707632;
assign addr[45587]= -2106406677;
assign addr[45588]= -2144419275;
assign addr[45589]= -2138975100;
assign addr[45590]= -2090184478;
assign addr[45591]= -1999036154;
assign addr[45592]= -1867377253;
assign addr[45593]= -1697875851;
assign addr[45594]= -1493966902;
assign addr[45595]= -1259782632;
assign addr[45596]= -1000068799;
assign addr[45597]= -720088517;
assign addr[45598]= -425515602;
assign addr[45599]= -122319591;
assign addr[45600]= 183355234;
assign addr[45601]= 485314355;
assign addr[45602]= 777438554;
assign addr[45603]= 1053807919;
assign addr[45604]= 1308821808;
assign addr[45605]= 1537312353;
assign addr[45606]= 1734649179;
assign addr[45607]= 1896833245;
assign addr[45608]= 2020577882;
assign addr[45609]= 2103375398;
assign addr[45610]= 2143547897;
assign addr[45611]= 2140281282;
assign addr[45612]= 2093641749;
assign addr[45613]= 2004574453;
assign addr[45614]= 1874884346;
assign addr[45615]= 1707199606;
assign addr[45616]= 1504918373;
assign addr[45617]= 1272139887;
assign addr[45618]= 1013581418;
assign addr[45619]= 734482665;
assign addr[45620]= 440499581;
assign addr[45621]= 137589750;
assign addr[45622]= -168108346;
assign addr[45623]= -470399716;
assign addr[45624]= -763158411;
assign addr[45625]= -1040451659;
assign addr[45626]= -1296660098;
assign addr[45627]= -1526591649;
assign addr[45628]= -1725586737;
assign addr[45629]= -1889612716;
assign addr[45630]= -2015345591;
assign addr[45631]= -2100237377;
assign addr[45632]= -2142567738;
assign addr[45633]= -2141478848;
assign addr[45634]= -2096992772;
assign addr[45635]= -2010011024;
assign addr[45636]= -1882296293;
assign addr[45637]= -1716436725;
assign addr[45638]= -1515793473;
assign addr[45639]= -1284432584;
assign addr[45640]= -1027042599;
assign addr[45641]= -748839539;
assign addr[45642]= -455461206;
assign addr[45643]= -152852926;
assign addr[45644]= 152852926;
assign addr[45645]= 455461206;
assign addr[45646]= 748839539;
assign addr[45647]= 1027042599;
assign addr[45648]= 1284432584;
assign addr[45649]= 1515793473;
assign addr[45650]= 1716436725;
assign addr[45651]= 1882296293;
assign addr[45652]= 2010011024;
assign addr[45653]= 2096992772;
assign addr[45654]= 2141478848;
assign addr[45655]= 2142567738;
assign addr[45656]= 2100237377;
assign addr[45657]= 2015345591;
assign addr[45658]= 1889612716;
assign addr[45659]= 1725586737;
assign addr[45660]= 1526591649;
assign addr[45661]= 1296660098;
assign addr[45662]= 1040451659;
assign addr[45663]= 763158411;
assign addr[45664]= 470399716;
assign addr[45665]= 168108346;
assign addr[45666]= -137589750;
assign addr[45667]= -440499581;
assign addr[45668]= -734482665;
assign addr[45669]= -1013581418;
assign addr[45670]= -1272139887;
assign addr[45671]= -1504918373;
assign addr[45672]= -1707199606;
assign addr[45673]= -1874884346;
assign addr[45674]= -2004574453;
assign addr[45675]= -2093641749;
assign addr[45676]= -2140281282;
assign addr[45677]= -2143547897;
assign addr[45678]= -2103375398;
assign addr[45679]= -2020577882;
assign addr[45680]= -1896833245;
assign addr[45681]= -1734649179;
assign addr[45682]= -1537312353;
assign addr[45683]= -1308821808;
assign addr[45684]= -1053807919;
assign addr[45685]= -777438554;
assign addr[45686]= -485314355;
assign addr[45687]= -183355234;
assign addr[45688]= 122319591;
assign addr[45689]= 425515602;
assign addr[45690]= 720088517;
assign addr[45691]= 1000068799;
assign addr[45692]= 1259782632;
assign addr[45693]= 1493966902;
assign addr[45694]= 1697875851;
assign addr[45695]= 1867377253;
assign addr[45696]= 1999036154;
assign addr[45697]= 2090184478;
assign addr[45698]= 2138975100;
assign addr[45699]= 2144419275;
assign addr[45700]= 2106406677;
assign addr[45701]= 2025707632;
assign addr[45702]= 1903957513;
assign addr[45703]= 1743623590;
assign addr[45704]= 1547955041;
assign addr[45705]= 1320917099;
assign addr[45706]= 1067110699;
assign addr[45707]= 791679244;
assign addr[45708]= 500204365;
assign addr[45709]= 198592817;
assign addr[45710]= -107043224;
assign addr[45711]= -410510029;
assign addr[45712]= -705657826;
assign addr[45713]= -986505429;
assign addr[45714]= -1247361445;
assign addr[45715]= -1482939614;
assign addr[45716]= -1688465931;
assign addr[45717]= -1859775393;
assign addr[45718]= -1993396407;
assign addr[45719]= -2086621133;
assign addr[45720]= -2137560369;
assign addr[45721]= -2145181827;
assign addr[45722]= -2109331059;
assign addr[45723]= -2030734582;
assign addr[45724]= -1910985158;
assign addr[45725]= -1752509516;
assign addr[45726]= -1558519173;
assign addr[45727]= -1332945355;
assign addr[45728]= -1080359326;
assign addr[45729]= -805879757;
assign addr[45730]= -515068990;
assign addr[45731]= -213820322;
assign addr[45732]= 91761426;
assign addr[45733]= 395483624;
assign addr[45734]= 691191324;
assign addr[45735]= 972891995;
assign addr[45736]= 1234876957;
assign addr[45737]= 1471837070;
assign addr[45738]= 1678970324;
assign addr[45739]= 1852079154;
assign addr[45740]= 1987655498;
assign addr[45741]= 2082951896;
assign addr[45742]= 2136037160;
assign addr[45743]= 2145835515;
assign addr[45744]= 2112148396;
assign addr[45745]= 2035658475;
assign addr[45746]= 1917915825;
assign addr[45747]= 1761306505;
assign addr[45748]= 1569004214;
assign addr[45749]= 1344905966;
assign addr[45750]= 1093553126;
assign addr[45751]= 820039373;
assign addr[45752]= 529907477;
assign addr[45753]= 229036977;
assign addr[45754]= -76474970;
assign addr[45755]= -380437148;
assign addr[45756]= -676689746;
assign addr[45757]= -959229189;
assign addr[45758]= -1222329801;
assign addr[45759]= -1460659832;
assign addr[45760]= -1669389513;
assign addr[45761]= -1844288924;
assign addr[45762]= -1981813720;
assign addr[45763]= -2079176953;
assign addr[45764]= -2134405552;
assign addr[45765]= -2146380306;
assign addr[45766]= -2114858546;
assign addr[45767]= -2040479063;
assign addr[45768]= -1924749160;
assign addr[45769]= -1770014111;
assign addr[45770]= -1579409630;
assign addr[45771]= -1356798326;
assign addr[45772]= -1106691431;
assign addr[45773]= -834157373;
assign addr[45774]= -544719071;
assign addr[45775]= -244242007;
assign addr[45776]= 61184634;
assign addr[45777]= 365371365;
assign addr[45778]= 662153826;
assign addr[45779]= 945517704;
assign addr[45780]= 1209720613;
assign addr[45781]= 1449408469;
assign addr[45782]= 1659723983;
assign addr[45783]= 1836405100;
assign addr[45784]= 1975871368;
assign addr[45785]= 2075296495;
assign addr[45786]= 2132665626;
assign addr[45787]= 2146816171;
assign addr[45788]= 2117461370;
assign addr[45789]= 2045196100;
assign addr[45790]= 1931484818;
assign addr[45791]= 1778631892;
assign addr[45792]= 1589734894;
assign addr[45793]= 1368621831;
assign addr[45794]= 1119773573;
assign addr[45795]= 848233042;
assign addr[45796]= 559503022;
assign addr[45797]= 259434643;
assign addr[45798]= -45891193;
assign addr[45799]= -350287041;
assign addr[45800]= -647584304;
assign addr[45801]= -931758235;
assign addr[45802]= -1197050035;
assign addr[45803]= -1438083551;
assign addr[45804]= -1649974225;
assign addr[45805]= -1828428082;
assign addr[45806]= -1969828744;
assign addr[45807]= -2071310720;
assign addr[45808]= -2130817471;
assign addr[45809]= -2147143090;
assign addr[45810]= -2119956737;
assign addr[45811]= -2049809346;
assign addr[45812]= -1938122457;
assign addr[45813]= -1787159411;
assign addr[45814]= -1599979481;
assign addr[45815]= -1380375881;
assign addr[45816]= -1132798888;
assign addr[45817]= -862265664;
assign addr[45818]= -574258580;
assign addr[45819]= -274614114;
assign addr[45820]= 30595422;
assign addr[45821]= 335184940;
assign addr[45822]= 632981917;
assign addr[45823]= 917951481;
assign addr[45824]= 1184318708;
assign addr[45825]= 1426685652;
assign addr[45826]= 1640140734;
assign addr[45827]= 1820358275;
assign addr[45828]= 1963686155;
assign addr[45829]= 2067219829;
assign addr[45830]= 2128861181;
assign addr[45831]= 2147361045;
assign addr[45832]= 2122344521;
assign addr[45833]= 2054318569;
assign addr[45834]= 1944661739;
assign addr[45835]= 1795596234;
assign addr[45836]= 1610142873;
assign addr[45837]= 1392059879;
assign addr[45838]= 1145766716;
assign addr[45839]= 876254528;
assign addr[45840]= 588984994;
assign addr[45841]= 289779648;
assign addr[45842]= -15298099;
assign addr[45843]= -320065829;
assign addr[45844]= -618347408;
assign addr[45845]= -904098143;
assign addr[45846]= -1171527280;
assign addr[45847]= -1415215352;
assign addr[45848]= -1630224009;
assign addr[45849]= -1812196087;
assign addr[45850]= -1957443913;
assign addr[45851]= -2063024031;
assign addr[45852]= -2126796855;
assign addr[45853]= -2147470025;
assign addr[45854]= -2124624598;
assign addr[45855]= -2058723538;
assign addr[45856]= -1951102334;
assign addr[45857]= -1803941934;
assign addr[45858]= -1620224553;
assign addr[45859]= -1403673233;
assign addr[45860]= -1158676398;
assign addr[45861]= -890198924;
assign addr[45862]= -603681519;
assign addr[45863]= -304930476;
assign addr[45864]= 0;
assign addr[45865]= 304930476;
assign addr[45866]= 603681519;
assign addr[45867]= 890198924;
assign addr[45868]= 1158676398;
assign addr[45869]= 1403673233;
assign addr[45870]= 1620224553;
assign addr[45871]= 1803941934;
assign addr[45872]= 1951102334;
assign addr[45873]= 2058723538;
assign addr[45874]= 2124624598;
assign addr[45875]= 2147470025;
assign addr[45876]= 2126796855;
assign addr[45877]= 2063024031;
assign addr[45878]= 1957443913;
assign addr[45879]= 1812196087;
assign addr[45880]= 1630224009;
assign addr[45881]= 1415215352;
assign addr[45882]= 1171527280;
assign addr[45883]= 904098143;
assign addr[45884]= 618347408;
assign addr[45885]= 320065829;
assign addr[45886]= 15298099;
assign addr[45887]= -289779648;
assign addr[45888]= -588984994;
assign addr[45889]= -876254528;
assign addr[45890]= -1145766716;
assign addr[45891]= -1392059879;
assign addr[45892]= -1610142873;
assign addr[45893]= -1795596234;
assign addr[45894]= -1944661739;
assign addr[45895]= -2054318569;
assign addr[45896]= -2122344521;
assign addr[45897]= -2147361045;
assign addr[45898]= -2128861181;
assign addr[45899]= -2067219829;
assign addr[45900]= -1963686155;
assign addr[45901]= -1820358275;
assign addr[45902]= -1640140734;
assign addr[45903]= -1426685652;
assign addr[45904]= -1184318708;
assign addr[45905]= -917951481;
assign addr[45906]= -632981917;
assign addr[45907]= -335184940;
assign addr[45908]= -30595422;
assign addr[45909]= 274614114;
assign addr[45910]= 574258580;
assign addr[45911]= 862265664;
assign addr[45912]= 1132798888;
assign addr[45913]= 1380375881;
assign addr[45914]= 1599979481;
assign addr[45915]= 1787159411;
assign addr[45916]= 1938122457;
assign addr[45917]= 2049809346;
assign addr[45918]= 2119956737;
assign addr[45919]= 2147143090;
assign addr[45920]= 2130817471;
assign addr[45921]= 2071310720;
assign addr[45922]= 1969828744;
assign addr[45923]= 1828428082;
assign addr[45924]= 1649974225;
assign addr[45925]= 1438083551;
assign addr[45926]= 1197050035;
assign addr[45927]= 931758235;
assign addr[45928]= 647584304;
assign addr[45929]= 350287041;
assign addr[45930]= 45891193;
assign addr[45931]= -259434643;
assign addr[45932]= -559503022;
assign addr[45933]= -848233042;
assign addr[45934]= -1119773573;
assign addr[45935]= -1368621831;
assign addr[45936]= -1589734894;
assign addr[45937]= -1778631892;
assign addr[45938]= -1931484818;
assign addr[45939]= -2045196100;
assign addr[45940]= -2117461370;
assign addr[45941]= -2146816171;
assign addr[45942]= -2132665626;
assign addr[45943]= -2075296495;
assign addr[45944]= -1975871368;
assign addr[45945]= -1836405100;
assign addr[45946]= -1659723983;
assign addr[45947]= -1449408469;
assign addr[45948]= -1209720613;
assign addr[45949]= -945517704;
assign addr[45950]= -662153826;
assign addr[45951]= -365371365;
assign addr[45952]= -61184634;
assign addr[45953]= 244242007;
assign addr[45954]= 544719071;
assign addr[45955]= 834157373;
assign addr[45956]= 1106691431;
assign addr[45957]= 1356798326;
assign addr[45958]= 1579409630;
assign addr[45959]= 1770014111;
assign addr[45960]= 1924749160;
assign addr[45961]= 2040479063;
assign addr[45962]= 2114858546;
assign addr[45963]= 2146380306;
assign addr[45964]= 2134405552;
assign addr[45965]= 2079176953;
assign addr[45966]= 1981813720;
assign addr[45967]= 1844288924;
assign addr[45968]= 1669389513;
assign addr[45969]= 1460659832;
assign addr[45970]= 1222329801;
assign addr[45971]= 959229189;
assign addr[45972]= 676689746;
assign addr[45973]= 380437148;
assign addr[45974]= 76474970;
assign addr[45975]= -229036977;
assign addr[45976]= -529907477;
assign addr[45977]= -820039373;
assign addr[45978]= -1093553126;
assign addr[45979]= -1344905966;
assign addr[45980]= -1569004214;
assign addr[45981]= -1761306505;
assign addr[45982]= -1917915825;
assign addr[45983]= -2035658475;
assign addr[45984]= -2112148396;
assign addr[45985]= -2145835515;
assign addr[45986]= -2136037160;
assign addr[45987]= -2082951896;
assign addr[45988]= -1987655498;
assign addr[45989]= -1852079154;
assign addr[45990]= -1678970324;
assign addr[45991]= -1471837070;
assign addr[45992]= -1234876957;
assign addr[45993]= -972891995;
assign addr[45994]= -691191324;
assign addr[45995]= -395483624;
assign addr[45996]= -91761426;
assign addr[45997]= 213820322;
assign addr[45998]= 515068990;
assign addr[45999]= 805879757;
assign addr[46000]= 1080359326;
assign addr[46001]= 1332945355;
assign addr[46002]= 1558519173;
assign addr[46003]= 1752509516;
assign addr[46004]= 1910985158;
assign addr[46005]= 2030734582;
assign addr[46006]= 2109331059;
assign addr[46007]= 2145181827;
assign addr[46008]= 2137560369;
assign addr[46009]= 2086621133;
assign addr[46010]= 1993396407;
assign addr[46011]= 1859775393;
assign addr[46012]= 1688465931;
assign addr[46013]= 1482939614;
assign addr[46014]= 1247361445;
assign addr[46015]= 986505429;
assign addr[46016]= 705657826;
assign addr[46017]= 410510029;
assign addr[46018]= 107043224;
assign addr[46019]= -198592817;
assign addr[46020]= -500204365;
assign addr[46021]= -791679244;
assign addr[46022]= -1067110699;
assign addr[46023]= -1320917099;
assign addr[46024]= -1547955041;
assign addr[46025]= -1743623590;
assign addr[46026]= -1903957513;
assign addr[46027]= -2025707632;
assign addr[46028]= -2106406677;
assign addr[46029]= -2144419275;
assign addr[46030]= -2138975100;
assign addr[46031]= -2090184478;
assign addr[46032]= -1999036154;
assign addr[46033]= -1867377253;
assign addr[46034]= -1697875851;
assign addr[46035]= -1493966902;
assign addr[46036]= -1259782632;
assign addr[46037]= -1000068799;
assign addr[46038]= -720088517;
assign addr[46039]= -425515602;
assign addr[46040]= -122319591;
assign addr[46041]= 183355234;
assign addr[46042]= 485314355;
assign addr[46043]= 777438554;
assign addr[46044]= 1053807919;
assign addr[46045]= 1308821808;
assign addr[46046]= 1537312353;
assign addr[46047]= 1734649179;
assign addr[46048]= 1896833245;
assign addr[46049]= 2020577882;
assign addr[46050]= 2103375398;
assign addr[46051]= 2143547897;
assign addr[46052]= 2140281282;
assign addr[46053]= 2093641749;
assign addr[46054]= 2004574453;
assign addr[46055]= 1874884346;
assign addr[46056]= 1707199606;
assign addr[46057]= 1504918373;
assign addr[46058]= 1272139887;
assign addr[46059]= 1013581418;
assign addr[46060]= 734482665;
assign addr[46061]= 440499581;
assign addr[46062]= 137589750;
assign addr[46063]= -168108346;
assign addr[46064]= -470399716;
assign addr[46065]= -763158411;
assign addr[46066]= -1040451659;
assign addr[46067]= -1296660098;
assign addr[46068]= -1526591649;
assign addr[46069]= -1725586737;
assign addr[46070]= -1889612716;
assign addr[46071]= -2015345591;
assign addr[46072]= -2100237377;
assign addr[46073]= -2142567738;
assign addr[46074]= -2141478848;
assign addr[46075]= -2096992772;
assign addr[46076]= -2010011024;
assign addr[46077]= -1882296293;
assign addr[46078]= -1716436725;
assign addr[46079]= -1515793473;
assign addr[46080]= -1284432584;
assign addr[46081]= -1027042599;
assign addr[46082]= -748839539;
assign addr[46083]= -455461206;
assign addr[46084]= -152852926;
assign addr[46085]= 152852926;
assign addr[46086]= 455461206;
assign addr[46087]= 748839539;
assign addr[46088]= 1027042599;
assign addr[46089]= 1284432584;
assign addr[46090]= 1515793473;
assign addr[46091]= 1716436725;
assign addr[46092]= 1882296293;
assign addr[46093]= 2010011024;
assign addr[46094]= 2096992772;
assign addr[46095]= 2141478848;
assign addr[46096]= 2142567738;
assign addr[46097]= 2100237377;
assign addr[46098]= 2015345591;
assign addr[46099]= 1889612716;
assign addr[46100]= 1725586737;
assign addr[46101]= 1526591649;
assign addr[46102]= 1296660098;
assign addr[46103]= 1040451659;
assign addr[46104]= 763158411;
assign addr[46105]= 470399716;
assign addr[46106]= 168108346;
assign addr[46107]= -137589750;
assign addr[46108]= -440499581;
assign addr[46109]= -734482665;
assign addr[46110]= -1013581418;
assign addr[46111]= -1272139887;
assign addr[46112]= -1504918373;
assign addr[46113]= -1707199606;
assign addr[46114]= -1874884346;
assign addr[46115]= -2004574453;
assign addr[46116]= -2093641749;
assign addr[46117]= -2140281282;
assign addr[46118]= -2143547897;
assign addr[46119]= -2103375398;
assign addr[46120]= -2020577882;
assign addr[46121]= -1896833245;
assign addr[46122]= -1734649179;
assign addr[46123]= -1537312353;
assign addr[46124]= -1308821808;
assign addr[46125]= -1053807919;
assign addr[46126]= -777438554;
assign addr[46127]= -485314355;
assign addr[46128]= -183355234;
assign addr[46129]= 122319591;
assign addr[46130]= 425515602;
assign addr[46131]= 720088517;
assign addr[46132]= 1000068799;
assign addr[46133]= 1259782632;
assign addr[46134]= 1493966902;
assign addr[46135]= 1697875851;
assign addr[46136]= 1867377253;
assign addr[46137]= 1999036154;
assign addr[46138]= 2090184478;
assign addr[46139]= 2138975100;
assign addr[46140]= 2144419275;
assign addr[46141]= 2106406677;
assign addr[46142]= 2025707632;
assign addr[46143]= 1903957513;
assign addr[46144]= 1743623590;
assign addr[46145]= 1547955041;
assign addr[46146]= 1320917099;
assign addr[46147]= 1067110699;
assign addr[46148]= 791679244;
assign addr[46149]= 500204365;
assign addr[46150]= 198592817;
assign addr[46151]= -107043224;
assign addr[46152]= -410510029;
assign addr[46153]= -705657826;
assign addr[46154]= -986505429;
assign addr[46155]= -1247361445;
assign addr[46156]= -1482939614;
assign addr[46157]= -1688465931;
assign addr[46158]= -1859775393;
assign addr[46159]= -1993396407;
assign addr[46160]= -2086621133;
assign addr[46161]= -2137560369;
assign addr[46162]= -2145181827;
assign addr[46163]= -2109331059;
assign addr[46164]= -2030734582;
assign addr[46165]= -1910985158;
assign addr[46166]= -1752509516;
assign addr[46167]= -1558519173;
assign addr[46168]= -1332945355;
assign addr[46169]= -1080359326;
assign addr[46170]= -805879757;
assign addr[46171]= -515068990;
assign addr[46172]= -213820322;
assign addr[46173]= 91761426;
assign addr[46174]= 395483624;
assign addr[46175]= 691191324;
assign addr[46176]= 972891995;
assign addr[46177]= 1234876957;
assign addr[46178]= 1471837070;
assign addr[46179]= 1678970324;
assign addr[46180]= 1852079154;
assign addr[46181]= 1987655498;
assign addr[46182]= 2082951896;
assign addr[46183]= 2136037160;
assign addr[46184]= 2145835515;
assign addr[46185]= 2112148396;
assign addr[46186]= 2035658475;
assign addr[46187]= 1917915825;
assign addr[46188]= 1761306505;
assign addr[46189]= 1569004214;
assign addr[46190]= 1344905966;
assign addr[46191]= 1093553126;
assign addr[46192]= 820039373;
assign addr[46193]= 529907477;
assign addr[46194]= 229036977;
assign addr[46195]= -76474970;
assign addr[46196]= -380437148;
assign addr[46197]= -676689746;
assign addr[46198]= -959229189;
assign addr[46199]= -1222329801;
assign addr[46200]= -1460659832;
assign addr[46201]= -1669389513;
assign addr[46202]= -1844288924;
assign addr[46203]= -1981813720;
assign addr[46204]= -2079176953;
assign addr[46205]= -2134405552;
assign addr[46206]= -2146380306;
assign addr[46207]= -2114858546;
assign addr[46208]= -2040479063;
assign addr[46209]= -1924749160;
assign addr[46210]= -1770014111;
assign addr[46211]= -1579409630;
assign addr[46212]= -1356798326;
assign addr[46213]= -1106691431;
assign addr[46214]= -834157373;
assign addr[46215]= -544719071;
assign addr[46216]= -244242007;
assign addr[46217]= 61184634;
assign addr[46218]= 365371365;
assign addr[46219]= 662153826;
assign addr[46220]= 945517704;
assign addr[46221]= 1209720613;
assign addr[46222]= 1449408469;
assign addr[46223]= 1659723983;
assign addr[46224]= 1836405100;
assign addr[46225]= 1975871368;
assign addr[46226]= 2075296495;
assign addr[46227]= 2132665626;
assign addr[46228]= 2146816171;
assign addr[46229]= 2117461370;
assign addr[46230]= 2045196100;
assign addr[46231]= 1931484818;
assign addr[46232]= 1778631892;
assign addr[46233]= 1589734894;
assign addr[46234]= 1368621831;
assign addr[46235]= 1119773573;
assign addr[46236]= 848233042;
assign addr[46237]= 559503022;
assign addr[46238]= 259434643;
assign addr[46239]= -45891193;
assign addr[46240]= -350287041;
assign addr[46241]= -647584304;
assign addr[46242]= -931758235;
assign addr[46243]= -1197050035;
assign addr[46244]= -1438083551;
assign addr[46245]= -1649974225;
assign addr[46246]= -1828428082;
assign addr[46247]= -1969828744;
assign addr[46248]= -2071310720;
assign addr[46249]= -2130817471;
assign addr[46250]= -2147143090;
assign addr[46251]= -2119956737;
assign addr[46252]= -2049809346;
assign addr[46253]= -1938122457;
assign addr[46254]= -1787159411;
assign addr[46255]= -1599979481;
assign addr[46256]= -1380375881;
assign addr[46257]= -1132798888;
assign addr[46258]= -862265664;
assign addr[46259]= -574258580;
assign addr[46260]= -274614114;
assign addr[46261]= 30595422;
assign addr[46262]= 335184940;
assign addr[46263]= 632981917;
assign addr[46264]= 917951481;
assign addr[46265]= 1184318708;
assign addr[46266]= 1426685652;
assign addr[46267]= 1640140734;
assign addr[46268]= 1820358275;
assign addr[46269]= 1963686155;
assign addr[46270]= 2067219829;
assign addr[46271]= 2128861181;
assign addr[46272]= 2147361045;
assign addr[46273]= 2122344521;
assign addr[46274]= 2054318569;
assign addr[46275]= 1944661739;
assign addr[46276]= 1795596234;
assign addr[46277]= 1610142873;
assign addr[46278]= 1392059879;
assign addr[46279]= 1145766716;
assign addr[46280]= 876254528;
assign addr[46281]= 588984994;
assign addr[46282]= 289779648;
assign addr[46283]= -15298099;
assign addr[46284]= -320065829;
assign addr[46285]= -618347408;
assign addr[46286]= -904098143;
assign addr[46287]= -1171527280;
assign addr[46288]= -1415215352;
assign addr[46289]= -1630224009;
assign addr[46290]= -1812196087;
assign addr[46291]= -1957443913;
assign addr[46292]= -2063024031;
assign addr[46293]= -2126796855;
assign addr[46294]= -2147470025;
assign addr[46295]= -2124624598;
assign addr[46296]= -2058723538;
assign addr[46297]= -1951102334;
assign addr[46298]= -1803941934;
assign addr[46299]= -1620224553;
assign addr[46300]= -1403673233;
assign addr[46301]= -1158676398;
assign addr[46302]= -890198924;
assign addr[46303]= -603681519;
assign addr[46304]= -304930476;
assign addr[46305]= 0;
assign addr[46306]= 304930476;
assign addr[46307]= 603681519;
assign addr[46308]= 890198924;
assign addr[46309]= 1158676398;
assign addr[46310]= 1403673233;
assign addr[46311]= 1620224553;
assign addr[46312]= 1803941934;
assign addr[46313]= 1951102334;
assign addr[46314]= 2058723538;
assign addr[46315]= 2124624598;
assign addr[46316]= 2147470025;
assign addr[46317]= 2126796855;
assign addr[46318]= 2063024031;
assign addr[46319]= 1957443913;
assign addr[46320]= 1812196087;
assign addr[46321]= 1630224009;
assign addr[46322]= 1415215352;
assign addr[46323]= 1171527280;
assign addr[46324]= 904098143;
assign addr[46325]= 618347408;
assign addr[46326]= 320065829;
assign addr[46327]= 15298099;
assign addr[46328]= -289779648;
assign addr[46329]= -588984994;
assign addr[46330]= -876254528;
assign addr[46331]= -1145766716;
assign addr[46332]= -1392059879;
assign addr[46333]= -1610142873;
assign addr[46334]= -1795596234;
assign addr[46335]= -1944661739;
assign addr[46336]= -2054318569;
assign addr[46337]= -2122344521;
assign addr[46338]= -2147361045;
assign addr[46339]= -2128861181;
assign addr[46340]= -2067219829;
assign addr[46341]= -1963686155;
assign addr[46342]= -1820358275;
assign addr[46343]= -1640140734;
assign addr[46344]= -1426685652;
assign addr[46345]= -1184318708;
assign addr[46346]= -917951481;
assign addr[46347]= -632981917;
assign addr[46348]= -335184940;
assign addr[46349]= -30595422;
assign addr[46350]= 274614114;
assign addr[46351]= 574258580;
assign addr[46352]= 862265664;
assign addr[46353]= 1132798888;
assign addr[46354]= 1380375881;
assign addr[46355]= 1599979481;
assign addr[46356]= 1787159411;
assign addr[46357]= 1938122457;
assign addr[46358]= 2049809346;
assign addr[46359]= 2119956737;
assign addr[46360]= 2147143090;
assign addr[46361]= 2130817471;
assign addr[46362]= 2071310720;
assign addr[46363]= 1969828744;
assign addr[46364]= 1828428082;
assign addr[46365]= 1649974225;
assign addr[46366]= 1438083551;
assign addr[46367]= 1197050035;
assign addr[46368]= 931758235;
assign addr[46369]= 647584304;
assign addr[46370]= 350287041;
assign addr[46371]= 45891193;
assign addr[46372]= -259434643;
assign addr[46373]= -559503022;
assign addr[46374]= -848233042;
assign addr[46375]= -1119773573;
assign addr[46376]= -1368621831;
assign addr[46377]= -1589734894;
assign addr[46378]= -1778631892;
assign addr[46379]= -1931484818;
assign addr[46380]= -2045196100;
assign addr[46381]= -2117461370;
assign addr[46382]= -2146816171;
assign addr[46383]= -2132665626;
assign addr[46384]= -2075296495;
assign addr[46385]= -1975871368;
assign addr[46386]= -1836405100;
assign addr[46387]= -1659723983;
assign addr[46388]= -1449408469;
assign addr[46389]= -1209720613;
assign addr[46390]= -945517704;
assign addr[46391]= -662153826;
assign addr[46392]= -365371365;
assign addr[46393]= -61184634;
assign addr[46394]= 244242007;
assign addr[46395]= 544719071;
assign addr[46396]= 834157373;
assign addr[46397]= 1106691431;
assign addr[46398]= 1356798326;
assign addr[46399]= 1579409630;
assign addr[46400]= 1770014111;
assign addr[46401]= 1924749160;
assign addr[46402]= 2040479063;
assign addr[46403]= 2114858546;
assign addr[46404]= 2146380306;
assign addr[46405]= 2134405552;
assign addr[46406]= 2079176953;
assign addr[46407]= 1981813720;
assign addr[46408]= 1844288924;
assign addr[46409]= 1669389513;
assign addr[46410]= 1460659832;
assign addr[46411]= 1222329801;
assign addr[46412]= 959229189;
assign addr[46413]= 676689746;
assign addr[46414]= 380437148;
assign addr[46415]= 76474970;
assign addr[46416]= -229036977;
assign addr[46417]= -529907477;
assign addr[46418]= -820039373;
assign addr[46419]= -1093553126;
assign addr[46420]= -1344905966;
assign addr[46421]= -1569004214;
assign addr[46422]= -1761306505;
assign addr[46423]= -1917915825;
assign addr[46424]= -2035658475;
assign addr[46425]= -2112148396;
assign addr[46426]= -2145835515;
assign addr[46427]= -2136037160;
assign addr[46428]= -2082951896;
assign addr[46429]= -1987655498;
assign addr[46430]= -1852079154;
assign addr[46431]= -1678970324;
assign addr[46432]= -1471837070;
assign addr[46433]= -1234876957;
assign addr[46434]= -972891995;
assign addr[46435]= -691191324;
assign addr[46436]= -395483624;
assign addr[46437]= -91761426;
assign addr[46438]= 213820322;
assign addr[46439]= 515068990;
assign addr[46440]= 805879757;
assign addr[46441]= 1080359326;
assign addr[46442]= 1332945355;
assign addr[46443]= 1558519173;
assign addr[46444]= 1752509516;
assign addr[46445]= 1910985158;
assign addr[46446]= 2030734582;
assign addr[46447]= 2109331059;
assign addr[46448]= 2145181827;
assign addr[46449]= 2137560369;
assign addr[46450]= 2086621133;
assign addr[46451]= 1993396407;
assign addr[46452]= 1859775393;
assign addr[46453]= 1688465931;
assign addr[46454]= 1482939614;
assign addr[46455]= 1247361445;
assign addr[46456]= 986505429;
assign addr[46457]= 705657826;
assign addr[46458]= 410510029;
assign addr[46459]= 107043224;
assign addr[46460]= -198592817;
assign addr[46461]= -500204365;
assign addr[46462]= -791679244;
assign addr[46463]= -1067110699;
assign addr[46464]= -1320917099;
assign addr[46465]= -1547955041;
assign addr[46466]= -1743623590;
assign addr[46467]= -1903957513;
assign addr[46468]= -2025707632;
assign addr[46469]= -2106406677;
assign addr[46470]= -2144419275;
assign addr[46471]= -2138975100;
assign addr[46472]= -2090184478;
assign addr[46473]= -1999036154;
assign addr[46474]= -1867377253;
assign addr[46475]= -1697875851;
assign addr[46476]= -1493966902;
assign addr[46477]= -1259782632;
assign addr[46478]= -1000068799;
assign addr[46479]= -720088517;
assign addr[46480]= -425515602;
assign addr[46481]= -122319591;
assign addr[46482]= 183355234;
assign addr[46483]= 485314355;
assign addr[46484]= 777438554;
assign addr[46485]= 1053807919;
assign addr[46486]= 1308821808;
assign addr[46487]= 1537312353;
assign addr[46488]= 1734649179;
assign addr[46489]= 1896833245;
assign addr[46490]= 2020577882;
assign addr[46491]= 2103375398;
assign addr[46492]= 2143547897;
assign addr[46493]= 2140281282;
assign addr[46494]= 2093641749;
assign addr[46495]= 2004574453;
assign addr[46496]= 1874884346;
assign addr[46497]= 1707199606;
assign addr[46498]= 1504918373;
assign addr[46499]= 1272139887;
assign addr[46500]= 1013581418;
assign addr[46501]= 734482665;
assign addr[46502]= 440499581;
assign addr[46503]= 137589750;
assign addr[46504]= -168108346;
assign addr[46505]= -470399716;
assign addr[46506]= -763158411;
assign addr[46507]= -1040451659;
assign addr[46508]= -1296660098;
assign addr[46509]= -1526591649;
assign addr[46510]= -1725586737;
assign addr[46511]= -1889612716;
assign addr[46512]= -2015345591;
assign addr[46513]= -2100237377;
assign addr[46514]= -2142567738;
assign addr[46515]= -2141478848;
assign addr[46516]= -2096992772;
assign addr[46517]= -2010011024;
assign addr[46518]= -1882296293;
assign addr[46519]= -1716436725;
assign addr[46520]= -1515793473;
assign addr[46521]= -1284432584;
assign addr[46522]= -1027042599;
assign addr[46523]= -748839539;
assign addr[46524]= -455461206;
assign addr[46525]= -152852926;
assign addr[46526]= 152852926;
assign addr[46527]= 455461206;
assign addr[46528]= 748839539;
assign addr[46529]= 1027042599;
assign addr[46530]= 1284432584;
assign addr[46531]= 1515793473;
assign addr[46532]= 1716436725;
assign addr[46533]= 1882296293;
assign addr[46534]= 2010011024;
assign addr[46535]= 2096992772;
assign addr[46536]= 2141478848;
assign addr[46537]= 2142567738;
assign addr[46538]= 2100237377;
assign addr[46539]= 2015345591;
assign addr[46540]= 1889612716;
assign addr[46541]= 1725586737;
assign addr[46542]= 1526591649;
assign addr[46543]= 1296660098;
assign addr[46544]= 1040451659;
assign addr[46545]= 763158411;
assign addr[46546]= 470399716;
assign addr[46547]= 168108346;
assign addr[46548]= -137589750;
assign addr[46549]= -440499581;
assign addr[46550]= -734482665;
assign addr[46551]= -1013581418;
assign addr[46552]= -1272139887;
assign addr[46553]= -1504918373;
assign addr[46554]= -1707199606;
assign addr[46555]= -1874884346;
assign addr[46556]= -2004574453;
assign addr[46557]= -2093641749;
assign addr[46558]= -2140281282;
assign addr[46559]= -2143547897;
assign addr[46560]= -2103375398;
assign addr[46561]= -2020577882;
assign addr[46562]= -1896833245;
assign addr[46563]= -1734649179;
assign addr[46564]= -1537312353;
assign addr[46565]= -1308821808;
assign addr[46566]= -1053807919;
assign addr[46567]= -777438554;
assign addr[46568]= -485314355;
assign addr[46569]= -183355234;
assign addr[46570]= 122319591;
assign addr[46571]= 425515602;
assign addr[46572]= 720088517;
assign addr[46573]= 1000068799;
assign addr[46574]= 1259782632;
assign addr[46575]= 1493966902;
assign addr[46576]= 1697875851;
assign addr[46577]= 1867377253;
assign addr[46578]= 1999036154;
assign addr[46579]= 2090184478;
assign addr[46580]= 2138975100;
assign addr[46581]= 2144419275;
assign addr[46582]= 2106406677;
assign addr[46583]= 2025707632;
assign addr[46584]= 1903957513;
assign addr[46585]= 1743623590;
assign addr[46586]= 1547955041;
assign addr[46587]= 1320917099;
assign addr[46588]= 1067110699;
assign addr[46589]= 791679244;
assign addr[46590]= 500204365;
assign addr[46591]= 198592817;
assign addr[46592]= -107043224;
assign addr[46593]= -410510029;
assign addr[46594]= -705657826;
assign addr[46595]= -986505429;
assign addr[46596]= -1247361445;
assign addr[46597]= -1482939614;
assign addr[46598]= -1688465931;
assign addr[46599]= -1859775393;
assign addr[46600]= -1993396407;
assign addr[46601]= -2086621133;
assign addr[46602]= -2137560369;
assign addr[46603]= -2145181827;
assign addr[46604]= -2109331059;
assign addr[46605]= -2030734582;
assign addr[46606]= -1910985158;
assign addr[46607]= -1752509516;
assign addr[46608]= -1558519173;
assign addr[46609]= -1332945355;
assign addr[46610]= -1080359326;
assign addr[46611]= -805879757;
assign addr[46612]= -515068990;
assign addr[46613]= -213820322;
assign addr[46614]= 91761426;
assign addr[46615]= 395483624;
assign addr[46616]= 691191324;
assign addr[46617]= 972891995;
assign addr[46618]= 1234876957;
assign addr[46619]= 1471837070;
assign addr[46620]= 1678970324;
assign addr[46621]= 1852079154;
assign addr[46622]= 1987655498;
assign addr[46623]= 2082951896;
assign addr[46624]= 2136037160;
assign addr[46625]= 2145835515;
assign addr[46626]= 2112148396;
assign addr[46627]= 2035658475;
assign addr[46628]= 1917915825;
assign addr[46629]= 1761306505;
assign addr[46630]= 1569004214;
assign addr[46631]= 1344905966;
assign addr[46632]= 1093553126;
assign addr[46633]= 820039373;
assign addr[46634]= 529907477;
assign addr[46635]= 229036977;
assign addr[46636]= -76474970;
assign addr[46637]= -380437148;
assign addr[46638]= -676689746;
assign addr[46639]= -959229189;
assign addr[46640]= -1222329801;
assign addr[46641]= -1460659832;
assign addr[46642]= -1669389513;
assign addr[46643]= -1844288924;
assign addr[46644]= -1981813720;
assign addr[46645]= -2079176953;
assign addr[46646]= -2134405552;
assign addr[46647]= -2146380306;
assign addr[46648]= -2114858546;
assign addr[46649]= -2040479063;
assign addr[46650]= -1924749160;
assign addr[46651]= -1770014111;
assign addr[46652]= -1579409630;
assign addr[46653]= -1356798326;
assign addr[46654]= -1106691431;
assign addr[46655]= -834157373;
assign addr[46656]= -544719071;
assign addr[46657]= -244242007;
assign addr[46658]= 61184634;
assign addr[46659]= 365371365;
assign addr[46660]= 662153826;
assign addr[46661]= 945517704;
assign addr[46662]= 1209720613;
assign addr[46663]= 1449408469;
assign addr[46664]= 1659723983;
assign addr[46665]= 1836405100;
assign addr[46666]= 1975871368;
assign addr[46667]= 2075296495;
assign addr[46668]= 2132665626;
assign addr[46669]= 2146816171;
assign addr[46670]= 2117461370;
assign addr[46671]= 2045196100;
assign addr[46672]= 1931484818;
assign addr[46673]= 1778631892;
assign addr[46674]= 1589734894;
assign addr[46675]= 1368621831;
assign addr[46676]= 1119773573;
assign addr[46677]= 848233042;
assign addr[46678]= 559503022;
assign addr[46679]= 259434643;
assign addr[46680]= -45891193;
assign addr[46681]= -350287041;
assign addr[46682]= -647584304;
assign addr[46683]= -931758235;
assign addr[46684]= -1197050035;
assign addr[46685]= -1438083551;
assign addr[46686]= -1649974225;
assign addr[46687]= -1828428082;
assign addr[46688]= -1969828744;
assign addr[46689]= -2071310720;
assign addr[46690]= -2130817471;
assign addr[46691]= -2147143090;
assign addr[46692]= -2119956737;
assign addr[46693]= -2049809346;
assign addr[46694]= -1938122457;
assign addr[46695]= -1787159411;
assign addr[46696]= -1599979481;
assign addr[46697]= -1380375881;
assign addr[46698]= -1132798888;
assign addr[46699]= -862265664;
assign addr[46700]= -574258580;
assign addr[46701]= -274614114;
assign addr[46702]= 30595422;
assign addr[46703]= 335184940;
assign addr[46704]= 632981917;
assign addr[46705]= 917951481;
assign addr[46706]= 1184318708;
assign addr[46707]= 1426685652;
assign addr[46708]= 1640140734;
assign addr[46709]= 1820358275;
assign addr[46710]= 1963686155;
assign addr[46711]= 2067219829;
assign addr[46712]= 2128861181;
assign addr[46713]= 2147361045;
assign addr[46714]= 2122344521;
assign addr[46715]= 2054318569;
assign addr[46716]= 1944661739;
assign addr[46717]= 1795596234;
assign addr[46718]= 1610142873;
assign addr[46719]= 1392059879;
assign addr[46720]= 1145766716;
assign addr[46721]= 876254528;
assign addr[46722]= 588984994;
assign addr[46723]= 289779648;
assign addr[46724]= -15298099;
assign addr[46725]= -320065829;
assign addr[46726]= -618347408;
assign addr[46727]= -904098143;
assign addr[46728]= -1171527280;
assign addr[46729]= -1415215352;
assign addr[46730]= -1630224009;
assign addr[46731]= -1812196087;
assign addr[46732]= -1957443913;
assign addr[46733]= -2063024031;
assign addr[46734]= -2126796855;
assign addr[46735]= -2147470025;
assign addr[46736]= -2124624598;
assign addr[46737]= -2058723538;
assign addr[46738]= -1951102334;
assign addr[46739]= -1803941934;
assign addr[46740]= -1620224553;
assign addr[46741]= -1403673233;
assign addr[46742]= -1158676398;
assign addr[46743]= -890198924;
assign addr[46744]= -603681519;
assign addr[46745]= -304930476;
assign addr[46746]= 0;
assign addr[46747]= 304930476;
assign addr[46748]= 603681519;
assign addr[46749]= 890198924;
assign addr[46750]= 1158676398;
assign addr[46751]= 1403673233;
assign addr[46752]= 1620224553;
assign addr[46753]= 1803941934;
assign addr[46754]= 1951102334;
assign addr[46755]= 2058723538;
assign addr[46756]= 2124624598;
assign addr[46757]= 2147470025;
assign addr[46758]= 2126796855;
assign addr[46759]= 2063024031;
assign addr[46760]= 1957443913;
assign addr[46761]= 1812196087;
assign addr[46762]= 1630224009;
assign addr[46763]= 1415215352;
assign addr[46764]= 1171527280;
assign addr[46765]= 904098143;
assign addr[46766]= 618347408;
assign addr[46767]= 320065829;
assign addr[46768]= 15298099;
assign addr[46769]= -289779648;
assign addr[46770]= -588984994;
assign addr[46771]= -876254528;
assign addr[46772]= -1145766716;
assign addr[46773]= -1392059879;
assign addr[46774]= -1610142873;
assign addr[46775]= -1795596234;
assign addr[46776]= -1944661739;
assign addr[46777]= -2054318569;
assign addr[46778]= -2122344521;
assign addr[46779]= -2147361045;
assign addr[46780]= -2128861181;
assign addr[46781]= -2067219829;
assign addr[46782]= -1963686155;
assign addr[46783]= -1820358275;
assign addr[46784]= -1640140734;
assign addr[46785]= -1426685652;
assign addr[46786]= -1184318708;
assign addr[46787]= -917951481;
assign addr[46788]= -632981917;
assign addr[46789]= -335184940;
assign addr[46790]= -30595422;
assign addr[46791]= 274614114;
assign addr[46792]= 574258580;
assign addr[46793]= 862265664;
assign addr[46794]= 1132798888;
assign addr[46795]= 1380375881;
assign addr[46796]= 1599979481;
assign addr[46797]= 1787159411;
assign addr[46798]= 1938122457;
assign addr[46799]= 2049809346;
assign addr[46800]= 2119956737;
assign addr[46801]= 2147143090;
assign addr[46802]= 2130817471;
assign addr[46803]= 2071310720;
assign addr[46804]= 1969828744;
assign addr[46805]= 1828428082;
assign addr[46806]= 1649974225;
assign addr[46807]= 1438083551;
assign addr[46808]= 1197050035;
assign addr[46809]= 931758235;
assign addr[46810]= 647584304;
assign addr[46811]= 350287041;
assign addr[46812]= 45891193;
assign addr[46813]= -259434643;
assign addr[46814]= -559503022;
assign addr[46815]= -848233042;
assign addr[46816]= -1119773573;
assign addr[46817]= -1368621831;
assign addr[46818]= -1589734894;
assign addr[46819]= -1778631892;
assign addr[46820]= -1931484818;
assign addr[46821]= -2045196100;
assign addr[46822]= -2117461370;
assign addr[46823]= -2146816171;
assign addr[46824]= -2132665626;
assign addr[46825]= -2075296495;
assign addr[46826]= -1975871368;
assign addr[46827]= -1836405100;
assign addr[46828]= -1659723983;
assign addr[46829]= -1449408469;
assign addr[46830]= -1209720613;
assign addr[46831]= -945517704;
assign addr[46832]= -662153826;
assign addr[46833]= -365371365;
assign addr[46834]= -61184634;
assign addr[46835]= 244242007;
assign addr[46836]= 544719071;
assign addr[46837]= 834157373;
assign addr[46838]= 1106691431;
assign addr[46839]= 1356798326;
assign addr[46840]= 1579409630;
assign addr[46841]= 1770014111;
assign addr[46842]= 1924749160;
assign addr[46843]= 2040479063;
assign addr[46844]= 2114858546;
assign addr[46845]= 2146380306;
assign addr[46846]= 2134405552;
assign addr[46847]= 2079176953;
assign addr[46848]= 1981813720;
assign addr[46849]= 1844288924;
assign addr[46850]= 1669389513;
assign addr[46851]= 1460659832;
assign addr[46852]= 1222329801;
assign addr[46853]= 959229189;
assign addr[46854]= 676689746;
assign addr[46855]= 380437148;
assign addr[46856]= 76474970;
assign addr[46857]= -229036977;
assign addr[46858]= -529907477;
assign addr[46859]= -820039373;
assign addr[46860]= -1093553126;
assign addr[46861]= -1344905966;
assign addr[46862]= -1569004214;
assign addr[46863]= -1761306505;
assign addr[46864]= -1917915825;
assign addr[46865]= -2035658475;
assign addr[46866]= -2112148396;
assign addr[46867]= -2145835515;
assign addr[46868]= -2136037160;
assign addr[46869]= -2082951896;
assign addr[46870]= -1987655498;
assign addr[46871]= -1852079154;
assign addr[46872]= -1678970324;
assign addr[46873]= -1471837070;
assign addr[46874]= -1234876957;
assign addr[46875]= -972891995;
assign addr[46876]= -691191324;
assign addr[46877]= -395483624;
assign addr[46878]= -91761426;
assign addr[46879]= 213820322;
assign addr[46880]= 515068990;
assign addr[46881]= 805879757;
assign addr[46882]= 1080359326;
assign addr[46883]= 1332945355;
assign addr[46884]= 1558519173;
assign addr[46885]= 1752509516;
assign addr[46886]= 1910985158;
assign addr[46887]= 2030734582;
assign addr[46888]= 2109331059;
assign addr[46889]= 2145181827;
assign addr[46890]= 2137560369;
assign addr[46891]= 2086621133;
assign addr[46892]= 1993396407;
assign addr[46893]= 1859775393;
assign addr[46894]= 1688465931;
assign addr[46895]= 1482939614;
assign addr[46896]= 1247361445;
assign addr[46897]= 986505429;
assign addr[46898]= 705657826;
assign addr[46899]= 410510029;
assign addr[46900]= 107043224;
assign addr[46901]= -198592817;
assign addr[46902]= -500204365;
assign addr[46903]= -791679244;
assign addr[46904]= -1067110699;
assign addr[46905]= -1320917099;
assign addr[46906]= -1547955041;
assign addr[46907]= -1743623590;
assign addr[46908]= -1903957513;
assign addr[46909]= -2025707632;
assign addr[46910]= -2106406677;
assign addr[46911]= -2144419275;
assign addr[46912]= -2138975100;
assign addr[46913]= -2090184478;
assign addr[46914]= -1999036154;
assign addr[46915]= -1867377253;
assign addr[46916]= -1697875851;
assign addr[46917]= -1493966902;
assign addr[46918]= -1259782632;
assign addr[46919]= -1000068799;
assign addr[46920]= -720088517;
assign addr[46921]= -425515602;
assign addr[46922]= -122319591;
assign addr[46923]= 183355234;
assign addr[46924]= 485314355;
assign addr[46925]= 777438554;
assign addr[46926]= 1053807919;
assign addr[46927]= 1308821808;
assign addr[46928]= 1537312353;
assign addr[46929]= 1734649179;
assign addr[46930]= 1896833245;
assign addr[46931]= 2020577882;
assign addr[46932]= 2103375398;
assign addr[46933]= 2143547897;
assign addr[46934]= 2140281282;
assign addr[46935]= 2093641749;
assign addr[46936]= 2004574453;
assign addr[46937]= 1874884346;
assign addr[46938]= 1707199606;
assign addr[46939]= 1504918373;
assign addr[46940]= 1272139887;
assign addr[46941]= 1013581418;
assign addr[46942]= 734482665;
assign addr[46943]= 440499581;
assign addr[46944]= 137589750;
assign addr[46945]= -168108346;
assign addr[46946]= -470399716;
assign addr[46947]= -763158411;
assign addr[46948]= -1040451659;
assign addr[46949]= -1296660098;
assign addr[46950]= -1526591649;
assign addr[46951]= -1725586737;
assign addr[46952]= -1889612716;
assign addr[46953]= -2015345591;
assign addr[46954]= -2100237377;
assign addr[46955]= -2142567738;
assign addr[46956]= -2141478848;
assign addr[46957]= -2096992772;
assign addr[46958]= -2010011024;
assign addr[46959]= -1882296293;
assign addr[46960]= -1716436725;
assign addr[46961]= -1515793473;
assign addr[46962]= -1284432584;
assign addr[46963]= -1027042599;
assign addr[46964]= -748839539;
assign addr[46965]= -455461206;
assign addr[46966]= -152852926;
assign addr[46967]= 152852926;
assign addr[46968]= 455461206;
assign addr[46969]= 748839539;
assign addr[46970]= 1027042599;
assign addr[46971]= 1284432584;
assign addr[46972]= 1515793473;
assign addr[46973]= 1716436725;
assign addr[46974]= 1882296293;
assign addr[46975]= 2010011024;
assign addr[46976]= 2096992772;
assign addr[46977]= 2141478848;
assign addr[46978]= 2142567738;
assign addr[46979]= 2100237377;
assign addr[46980]= 2015345591;
assign addr[46981]= 1889612716;
assign addr[46982]= 1725586737;
assign addr[46983]= 1526591649;
assign addr[46984]= 1296660098;
assign addr[46985]= 1040451659;
assign addr[46986]= 763158411;
assign addr[46987]= 470399716;
assign addr[46988]= 168108346;
assign addr[46989]= -137589750;
assign addr[46990]= -440499581;
assign addr[46991]= -734482665;
assign addr[46992]= -1013581418;
assign addr[46993]= -1272139887;
assign addr[46994]= -1504918373;
assign addr[46995]= -1707199606;
assign addr[46996]= -1874884346;
assign addr[46997]= -2004574453;
assign addr[46998]= -2093641749;
assign addr[46999]= -2140281282;
assign addr[47000]= -2143547897;
assign addr[47001]= -2103375398;
assign addr[47002]= -2020577882;
assign addr[47003]= -1896833245;
assign addr[47004]= -1734649179;
assign addr[47005]= -1537312353;
assign addr[47006]= -1308821808;
assign addr[47007]= -1053807919;
assign addr[47008]= -777438554;
assign addr[47009]= -485314355;
assign addr[47010]= -183355234;
assign addr[47011]= 122319591;
assign addr[47012]= 425515602;
assign addr[47013]= 720088517;
assign addr[47014]= 1000068799;
assign addr[47015]= 1259782632;
assign addr[47016]= 1493966902;
assign addr[47017]= 1697875851;
assign addr[47018]= 1867377253;
assign addr[47019]= 1999036154;
assign addr[47020]= 2090184478;
assign addr[47021]= 2138975100;
assign addr[47022]= 2144419275;
assign addr[47023]= 2106406677;
assign addr[47024]= 2025707632;
assign addr[47025]= 1903957513;
assign addr[47026]= 1743623590;
assign addr[47027]= 1547955041;
assign addr[47028]= 1320917099;
assign addr[47029]= 1067110699;
assign addr[47030]= 791679244;
assign addr[47031]= 500204365;
assign addr[47032]= 198592817;
assign addr[47033]= -107043224;
assign addr[47034]= -410510029;
assign addr[47035]= -705657826;
assign addr[47036]= -986505429;
assign addr[47037]= -1247361445;
assign addr[47038]= -1482939614;
assign addr[47039]= -1688465931;
assign addr[47040]= -1859775393;
assign addr[47041]= -1993396407;
assign addr[47042]= -2086621133;
assign addr[47043]= -2137560369;
assign addr[47044]= -2145181827;
assign addr[47045]= -2109331059;
assign addr[47046]= -2030734582;
assign addr[47047]= -1910985158;
assign addr[47048]= -1752509516;
assign addr[47049]= -1558519173;
assign addr[47050]= -1332945355;
assign addr[47051]= -1080359326;
assign addr[47052]= -805879757;
assign addr[47053]= -515068990;
assign addr[47054]= -213820322;
assign addr[47055]= 91761426;
assign addr[47056]= 395483624;
assign addr[47057]= 691191324;
assign addr[47058]= 972891995;
assign addr[47059]= 1234876957;
assign addr[47060]= 1471837070;
assign addr[47061]= 1678970324;
assign addr[47062]= 1852079154;
assign addr[47063]= 1987655498;
assign addr[47064]= 2082951896;
assign addr[47065]= 2136037160;
assign addr[47066]= 2145835515;
assign addr[47067]= 2112148396;
assign addr[47068]= 2035658475;
assign addr[47069]= 1917915825;
assign addr[47070]= 1761306505;
assign addr[47071]= 1569004214;
assign addr[47072]= 1344905966;
assign addr[47073]= 1093553126;
assign addr[47074]= 820039373;
assign addr[47075]= 529907477;
assign addr[47076]= 229036977;
assign addr[47077]= -76474970;
assign addr[47078]= -380437148;
assign addr[47079]= -676689746;
assign addr[47080]= -959229189;
assign addr[47081]= -1222329801;
assign addr[47082]= -1460659832;
assign addr[47083]= -1669389513;
assign addr[47084]= -1844288924;
assign addr[47085]= -1981813720;
assign addr[47086]= -2079176953;
assign addr[47087]= -2134405552;
assign addr[47088]= -2146380306;
assign addr[47089]= -2114858546;
assign addr[47090]= -2040479063;
assign addr[47091]= -1924749160;
assign addr[47092]= -1770014111;
assign addr[47093]= -1579409630;
assign addr[47094]= -1356798326;
assign addr[47095]= -1106691431;
assign addr[47096]= -834157373;
assign addr[47097]= -544719071;
assign addr[47098]= -244242007;
assign addr[47099]= 61184634;
assign addr[47100]= 365371365;
assign addr[47101]= 662153826;
assign addr[47102]= 945517704;
assign addr[47103]= 1209720613;
assign addr[47104]= 1449408469;
assign addr[47105]= 1659723983;
assign addr[47106]= 1836405100;
assign addr[47107]= 1975871368;
assign addr[47108]= 2075296495;
assign addr[47109]= 2132665626;
assign addr[47110]= 2146816171;
assign addr[47111]= 2117461370;
assign addr[47112]= 2045196100;
assign addr[47113]= 1931484818;
assign addr[47114]= 1778631892;
assign addr[47115]= 1589734894;
assign addr[47116]= 1368621831;
assign addr[47117]= 1119773573;
assign addr[47118]= 848233042;
assign addr[47119]= 559503022;
assign addr[47120]= 259434643;
assign addr[47121]= -45891193;
assign addr[47122]= -350287041;
assign addr[47123]= -647584304;
assign addr[47124]= -931758235;
assign addr[47125]= -1197050035;
assign addr[47126]= -1438083551;
assign addr[47127]= -1649974225;
assign addr[47128]= -1828428082;
assign addr[47129]= -1969828744;
assign addr[47130]= -2071310720;
assign addr[47131]= -2130817471;
assign addr[47132]= -2147143090;
assign addr[47133]= -2119956737;
assign addr[47134]= -2049809346;
assign addr[47135]= -1938122457;
assign addr[47136]= -1787159411;
assign addr[47137]= -1599979481;
assign addr[47138]= -1380375881;
assign addr[47139]= -1132798888;
assign addr[47140]= -862265664;
assign addr[47141]= -574258580;
assign addr[47142]= -274614114;
assign addr[47143]= 30595422;
assign addr[47144]= 335184940;
assign addr[47145]= 632981917;
assign addr[47146]= 917951481;
assign addr[47147]= 1184318708;
assign addr[47148]= 1426685652;
assign addr[47149]= 1640140734;
assign addr[47150]= 1820358275;
assign addr[47151]= 1963686155;
assign addr[47152]= 2067219829;
assign addr[47153]= 2128861181;
assign addr[47154]= 2147361045;
assign addr[47155]= 2122344521;
assign addr[47156]= 2054318569;
assign addr[47157]= 1944661739;
assign addr[47158]= 1795596234;
assign addr[47159]= 1610142873;
assign addr[47160]= 1392059879;
assign addr[47161]= 1145766716;
assign addr[47162]= 876254528;
assign addr[47163]= 588984994;
assign addr[47164]= 289779648;
assign addr[47165]= -15298099;
assign addr[47166]= -320065829;
assign addr[47167]= -618347408;
assign addr[47168]= -904098143;
assign addr[47169]= -1171527280;
assign addr[47170]= -1415215352;
assign addr[47171]= -1630224009;
assign addr[47172]= -1812196087;
assign addr[47173]= -1957443913;
assign addr[47174]= -2063024031;
assign addr[47175]= -2126796855;
assign addr[47176]= -2147470025;
assign addr[47177]= -2124624598;
assign addr[47178]= -2058723538;
assign addr[47179]= -1951102334;
assign addr[47180]= -1803941934;
assign addr[47181]= -1620224553;
assign addr[47182]= -1403673233;
assign addr[47183]= -1158676398;
assign addr[47184]= -890198924;
assign addr[47185]= -603681519;
assign addr[47186]= -304930476;
assign addr[47187]= 0;
assign addr[47188]= 304930476;
assign addr[47189]= 603681519;
assign addr[47190]= 890198924;
assign addr[47191]= 1158676398;
assign addr[47192]= 1403673233;
assign addr[47193]= 1620224553;
assign addr[47194]= 1803941934;
assign addr[47195]= 1951102334;
assign addr[47196]= 2058723538;
assign addr[47197]= 2124624598;
assign addr[47198]= 2147470025;
assign addr[47199]= 2126796855;
assign addr[47200]= 2063024031;
assign addr[47201]= 1957443913;
assign addr[47202]= 1812196087;
assign addr[47203]= 1630224009;
assign addr[47204]= 1415215352;
assign addr[47205]= 1171527280;
assign addr[47206]= 904098143;
assign addr[47207]= 618347408;
assign addr[47208]= 320065829;
assign addr[47209]= 15298099;
assign addr[47210]= -289779648;
assign addr[47211]= -588984994;
assign addr[47212]= -876254528;
assign addr[47213]= -1145766716;
assign addr[47214]= -1392059879;
assign addr[47215]= -1610142873;
assign addr[47216]= -1795596234;
assign addr[47217]= -1944661739;
assign addr[47218]= -2054318569;
assign addr[47219]= -2122344521;
assign addr[47220]= -2147361045;
assign addr[47221]= -2128861181;
assign addr[47222]= -2067219829;
assign addr[47223]= -1963686155;
assign addr[47224]= -1820358275;
assign addr[47225]= -1640140734;
assign addr[47226]= -1426685652;
assign addr[47227]= -1184318708;
assign addr[47228]= -917951481;
assign addr[47229]= -632981917;
assign addr[47230]= -335184940;
assign addr[47231]= -30595422;
assign addr[47232]= 274614114;
assign addr[47233]= 574258580;
assign addr[47234]= 862265664;
assign addr[47235]= 1132798888;
assign addr[47236]= 1380375881;
assign addr[47237]= 1599979481;
assign addr[47238]= 1787159411;
assign addr[47239]= 1938122457;
assign addr[47240]= 2049809346;
assign addr[47241]= 2119956737;
assign addr[47242]= 2147143090;
assign addr[47243]= 2130817471;
assign addr[47244]= 2071310720;
assign addr[47245]= 1969828744;
assign addr[47246]= 1828428082;
assign addr[47247]= 1649974225;
assign addr[47248]= 1438083551;
assign addr[47249]= 1197050035;
assign addr[47250]= 931758235;
assign addr[47251]= 647584304;
assign addr[47252]= 350287041;
assign addr[47253]= 45891193;
assign addr[47254]= -259434643;
assign addr[47255]= -559503022;
assign addr[47256]= -848233042;
assign addr[47257]= -1119773573;
assign addr[47258]= -1368621831;
assign addr[47259]= -1589734894;
assign addr[47260]= -1778631892;
assign addr[47261]= -1931484818;
assign addr[47262]= -2045196100;
assign addr[47263]= -2117461370;
assign addr[47264]= -2146816171;
assign addr[47265]= -2132665626;
assign addr[47266]= -2075296495;
assign addr[47267]= -1975871368;
assign addr[47268]= -1836405100;
assign addr[47269]= -1659723983;
assign addr[47270]= -1449408469;
assign addr[47271]= -1209720613;
assign addr[47272]= -945517704;
assign addr[47273]= -662153826;
assign addr[47274]= -365371365;
assign addr[47275]= -61184634;
assign addr[47276]= 244242007;
assign addr[47277]= 544719071;
assign addr[47278]= 834157373;
assign addr[47279]= 1106691431;
assign addr[47280]= 1356798326;
assign addr[47281]= 1579409630;
assign addr[47282]= 1770014111;
assign addr[47283]= 1924749160;
assign addr[47284]= 2040479063;
assign addr[47285]= 2114858546;
assign addr[47286]= 2146380306;
assign addr[47287]= 2134405552;
assign addr[47288]= 2079176953;
assign addr[47289]= 1981813720;
assign addr[47290]= 1844288924;
assign addr[47291]= 1669389513;
assign addr[47292]= 1460659832;
assign addr[47293]= 1222329801;
assign addr[47294]= 959229189;
assign addr[47295]= 676689746;
assign addr[47296]= 380437148;
assign addr[47297]= 76474970;
assign addr[47298]= -229036977;
assign addr[47299]= -529907477;
assign addr[47300]= -820039373;
assign addr[47301]= -1093553126;
assign addr[47302]= -1344905966;
assign addr[47303]= -1569004214;
assign addr[47304]= -1761306505;
assign addr[47305]= -1917915825;
assign addr[47306]= -2035658475;
assign addr[47307]= -2112148396;
assign addr[47308]= -2145835515;
assign addr[47309]= -2136037160;
assign addr[47310]= -2082951896;
assign addr[47311]= -1987655498;
assign addr[47312]= -1852079154;
assign addr[47313]= -1678970324;
assign addr[47314]= -1471837070;
assign addr[47315]= -1234876957;
assign addr[47316]= -972891995;
assign addr[47317]= -691191324;
assign addr[47318]= -395483624;
assign addr[47319]= -91761426;
assign addr[47320]= 213820322;
assign addr[47321]= 515068990;
assign addr[47322]= 805879757;
assign addr[47323]= 1080359326;
assign addr[47324]= 1332945355;
assign addr[47325]= 1558519173;
assign addr[47326]= 1752509516;
assign addr[47327]= 1910985158;
assign addr[47328]= 2030734582;
assign addr[47329]= 2109331059;
assign addr[47330]= 2145181827;
assign addr[47331]= 2137560369;
assign addr[47332]= 2086621133;
assign addr[47333]= 1993396407;
assign addr[47334]= 1859775393;
assign addr[47335]= 1688465931;
assign addr[47336]= 1482939614;
assign addr[47337]= 1247361445;
assign addr[47338]= 986505429;
assign addr[47339]= 705657826;
assign addr[47340]= 410510029;
assign addr[47341]= 107043224;
assign addr[47342]= -198592817;
assign addr[47343]= -500204365;
assign addr[47344]= -791679244;
assign addr[47345]= -1067110699;
assign addr[47346]= -1320917099;
assign addr[47347]= -1547955041;
assign addr[47348]= -1743623590;
assign addr[47349]= -1903957513;
assign addr[47350]= -2025707632;
assign addr[47351]= -2106406677;
assign addr[47352]= -2144419275;
assign addr[47353]= -2138975100;
assign addr[47354]= -2090184478;
assign addr[47355]= -1999036154;
assign addr[47356]= -1867377253;
assign addr[47357]= -1697875851;
assign addr[47358]= -1493966902;
assign addr[47359]= -1259782632;
assign addr[47360]= -1000068799;
assign addr[47361]= -720088517;
assign addr[47362]= -425515602;
assign addr[47363]= -122319591;
assign addr[47364]= 183355234;
assign addr[47365]= 485314355;
assign addr[47366]= 777438554;
assign addr[47367]= 1053807919;
assign addr[47368]= 1308821808;
assign addr[47369]= 1537312353;
assign addr[47370]= 1734649179;
assign addr[47371]= 1896833245;
assign addr[47372]= 2020577882;
assign addr[47373]= 2103375398;
assign addr[47374]= 2143547897;
assign addr[47375]= 2140281282;
assign addr[47376]= 2093641749;
assign addr[47377]= 2004574453;
assign addr[47378]= 1874884346;
assign addr[47379]= 1707199606;
assign addr[47380]= 1504918373;
assign addr[47381]= 1272139887;
assign addr[47382]= 1013581418;
assign addr[47383]= 734482665;
assign addr[47384]= 440499581;
assign addr[47385]= 137589750;
assign addr[47386]= -168108346;
assign addr[47387]= -470399716;
assign addr[47388]= -763158411;
assign addr[47389]= -1040451659;
assign addr[47390]= -1296660098;
assign addr[47391]= -1526591649;
assign addr[47392]= -1725586737;
assign addr[47393]= -1889612716;
assign addr[47394]= -2015345591;
assign addr[47395]= -2100237377;
assign addr[47396]= -2142567738;
assign addr[47397]= -2141478848;
assign addr[47398]= -2096992772;
assign addr[47399]= -2010011024;
assign addr[47400]= -1882296293;
assign addr[47401]= -1716436725;
assign addr[47402]= -1515793473;
assign addr[47403]= -1284432584;
assign addr[47404]= -1027042599;
assign addr[47405]= -748839539;
assign addr[47406]= -455461206;
assign addr[47407]= -152852926;
assign addr[47408]= 152852926;
assign addr[47409]= 455461206;
assign addr[47410]= 748839539;
assign addr[47411]= 1027042599;
assign addr[47412]= 1284432584;
assign addr[47413]= 1515793473;
assign addr[47414]= 1716436725;
assign addr[47415]= 1882296293;
assign addr[47416]= 2010011024;
assign addr[47417]= 2096992772;
assign addr[47418]= 2141478848;
assign addr[47419]= 2142567738;
assign addr[47420]= 2100237377;
assign addr[47421]= 2015345591;
assign addr[47422]= 1889612716;
assign addr[47423]= 1725586737;
assign addr[47424]= 1526591649;
assign addr[47425]= 1296660098;
assign addr[47426]= 1040451659;
assign addr[47427]= 763158411;
assign addr[47428]= 470399716;
assign addr[47429]= 168108346;
assign addr[47430]= -137589750;
assign addr[47431]= -440499581;
assign addr[47432]= -734482665;
assign addr[47433]= -1013581418;
assign addr[47434]= -1272139887;
assign addr[47435]= -1504918373;
assign addr[47436]= -1707199606;
assign addr[47437]= -1874884346;
assign addr[47438]= -2004574453;
assign addr[47439]= -2093641749;
assign addr[47440]= -2140281282;
assign addr[47441]= -2143547897;
assign addr[47442]= -2103375398;
assign addr[47443]= -2020577882;
assign addr[47444]= -1896833245;
assign addr[47445]= -1734649179;
assign addr[47446]= -1537312353;
assign addr[47447]= -1308821808;
assign addr[47448]= -1053807919;
assign addr[47449]= -777438554;
assign addr[47450]= -485314355;
assign addr[47451]= -183355234;
assign addr[47452]= 122319591;
assign addr[47453]= 425515602;
assign addr[47454]= 720088517;
assign addr[47455]= 1000068799;
assign addr[47456]= 1259782632;
assign addr[47457]= 1493966902;
assign addr[47458]= 1697875851;
assign addr[47459]= 1867377253;
assign addr[47460]= 1999036154;
assign addr[47461]= 2090184478;
assign addr[47462]= 2138975100;
assign addr[47463]= 2144419275;
assign addr[47464]= 2106406677;
assign addr[47465]= 2025707632;
assign addr[47466]= 1903957513;
assign addr[47467]= 1743623590;
assign addr[47468]= 1547955041;
assign addr[47469]= 1320917099;
assign addr[47470]= 1067110699;
assign addr[47471]= 791679244;
assign addr[47472]= 500204365;
assign addr[47473]= 198592817;
assign addr[47474]= -107043224;
assign addr[47475]= -410510029;
assign addr[47476]= -705657826;
assign addr[47477]= -986505429;
assign addr[47478]= -1247361445;
assign addr[47479]= -1482939614;
assign addr[47480]= -1688465931;
assign addr[47481]= -1859775393;
assign addr[47482]= -1993396407;
assign addr[47483]= -2086621133;
assign addr[47484]= -2137560369;
assign addr[47485]= -2145181827;
assign addr[47486]= -2109331059;
assign addr[47487]= -2030734582;
assign addr[47488]= -1910985158;
assign addr[47489]= -1752509516;
assign addr[47490]= -1558519173;
assign addr[47491]= -1332945355;
assign addr[47492]= -1080359326;
assign addr[47493]= -805879757;
assign addr[47494]= -515068990;
assign addr[47495]= -213820322;
assign addr[47496]= 91761426;
assign addr[47497]= 395483624;
assign addr[47498]= 691191324;
assign addr[47499]= 972891995;
assign addr[47500]= 1234876957;
assign addr[47501]= 1471837070;
assign addr[47502]= 1678970324;
assign addr[47503]= 1852079154;
assign addr[47504]= 1987655498;
assign addr[47505]= 2082951896;
assign addr[47506]= 2136037160;
assign addr[47507]= 2145835515;
assign addr[47508]= 2112148396;
assign addr[47509]= 2035658475;
assign addr[47510]= 1917915825;
assign addr[47511]= 1761306505;
assign addr[47512]= 1569004214;
assign addr[47513]= 1344905966;
assign addr[47514]= 1093553126;
assign addr[47515]= 820039373;
assign addr[47516]= 529907477;
assign addr[47517]= 229036977;
assign addr[47518]= -76474970;
assign addr[47519]= -380437148;
assign addr[47520]= -676689746;
assign addr[47521]= -959229189;
assign addr[47522]= -1222329801;
assign addr[47523]= -1460659832;
assign addr[47524]= -1669389513;
assign addr[47525]= -1844288924;
assign addr[47526]= -1981813720;
assign addr[47527]= -2079176953;
assign addr[47528]= -2134405552;
assign addr[47529]= -2146380306;
assign addr[47530]= -2114858546;
assign addr[47531]= -2040479063;
assign addr[47532]= -1924749160;
assign addr[47533]= -1770014111;
assign addr[47534]= -1579409630;
assign addr[47535]= -1356798326;
assign addr[47536]= -1106691431;
assign addr[47537]= -834157373;
assign addr[47538]= -544719071;
assign addr[47539]= -244242007;
assign addr[47540]= 61184634;
assign addr[47541]= 365371365;
assign addr[47542]= 662153826;
assign addr[47543]= 945517704;
assign addr[47544]= 1209720613;
assign addr[47545]= 1449408469;
assign addr[47546]= 1659723983;
assign addr[47547]= 1836405100;
assign addr[47548]= 1975871368;
assign addr[47549]= 2075296495;
assign addr[47550]= 2132665626;
assign addr[47551]= 2146816171;
assign addr[47552]= 2117461370;
assign addr[47553]= 2045196100;
assign addr[47554]= 1931484818;
assign addr[47555]= 1778631892;
assign addr[47556]= 1589734894;
assign addr[47557]= 1368621831;
assign addr[47558]= 1119773573;
assign addr[47559]= 848233042;
assign addr[47560]= 559503022;
assign addr[47561]= 259434643;
assign addr[47562]= -45891193;
assign addr[47563]= -350287041;
assign addr[47564]= -647584304;
assign addr[47565]= -931758235;
assign addr[47566]= -1197050035;
assign addr[47567]= -1438083551;
assign addr[47568]= -1649974225;
assign addr[47569]= -1828428082;
assign addr[47570]= -1969828744;
assign addr[47571]= -2071310720;
assign addr[47572]= -2130817471;
assign addr[47573]= -2147143090;
assign addr[47574]= -2119956737;
assign addr[47575]= -2049809346;
assign addr[47576]= -1938122457;
assign addr[47577]= -1787159411;
assign addr[47578]= -1599979481;
assign addr[47579]= -1380375881;
assign addr[47580]= -1132798888;
assign addr[47581]= -862265664;
assign addr[47582]= -574258580;
assign addr[47583]= -274614114;
assign addr[47584]= 30595422;
assign addr[47585]= 335184940;
assign addr[47586]= 632981917;
assign addr[47587]= 917951481;
assign addr[47588]= 1184318708;
assign addr[47589]= 1426685652;
assign addr[47590]= 1640140734;
assign addr[47591]= 1820358275;
assign addr[47592]= 1963686155;
assign addr[47593]= 2067219829;
assign addr[47594]= 2128861181;
assign addr[47595]= 2147361045;
assign addr[47596]= 2122344521;
assign addr[47597]= 2054318569;
assign addr[47598]= 1944661739;
assign addr[47599]= 1795596234;
assign addr[47600]= 1610142873;
assign addr[47601]= 1392059879;
assign addr[47602]= 1145766716;
assign addr[47603]= 876254528;
assign addr[47604]= 588984994;
assign addr[47605]= 289779648;
assign addr[47606]= -15298099;
assign addr[47607]= -320065829;
assign addr[47608]= -618347408;
assign addr[47609]= -904098143;
assign addr[47610]= -1171527280;
assign addr[47611]= -1415215352;
assign addr[47612]= -1630224009;
assign addr[47613]= -1812196087;
assign addr[47614]= -1957443913;
assign addr[47615]= -2063024031;
assign addr[47616]= -2126796855;
assign addr[47617]= -2147470025;
assign addr[47618]= -2124624598;
assign addr[47619]= -2058723538;
assign addr[47620]= -1951102334;
assign addr[47621]= -1803941934;
assign addr[47622]= -1620224553;
assign addr[47623]= -1403673233;
assign addr[47624]= -1158676398;
assign addr[47625]= -890198924;
assign addr[47626]= -603681519;
assign addr[47627]= -304930476;
assign addr[47628]= 0;
assign addr[47629]= 304930476;
assign addr[47630]= 603681519;
assign addr[47631]= 890198924;
assign addr[47632]= 1158676398;
assign addr[47633]= 1403673233;
assign addr[47634]= 1620224553;
assign addr[47635]= 1803941934;
assign addr[47636]= 1951102334;
assign addr[47637]= 2058723538;
assign addr[47638]= 2124624598;
assign addr[47639]= 2147470025;
assign addr[47640]= 2126796855;
assign addr[47641]= 2063024031;
assign addr[47642]= 1957443913;
assign addr[47643]= 1812196087;
assign addr[47644]= 1630224009;
assign addr[47645]= 1415215352;
assign addr[47646]= 1171527280;
assign addr[47647]= 904098143;
assign addr[47648]= 618347408;
assign addr[47649]= 320065829;
assign addr[47650]= 15298099;
assign addr[47651]= -289779648;
assign addr[47652]= -588984994;
assign addr[47653]= -876254528;
assign addr[47654]= -1145766716;
assign addr[47655]= -1392059879;
assign addr[47656]= -1610142873;
assign addr[47657]= -1795596234;
assign addr[47658]= -1944661739;
assign addr[47659]= -2054318569;
assign addr[47660]= -2122344521;
assign addr[47661]= -2147361045;
assign addr[47662]= -2128861181;
assign addr[47663]= -2067219829;
assign addr[47664]= -1963686155;
assign addr[47665]= -1820358275;
assign addr[47666]= -1640140734;
assign addr[47667]= -1426685652;
assign addr[47668]= -1184318708;
assign addr[47669]= -917951481;
assign addr[47670]= -632981917;
assign addr[47671]= -335184940;
assign addr[47672]= -30595422;
assign addr[47673]= 274614114;
assign addr[47674]= 574258580;
assign addr[47675]= 862265664;
assign addr[47676]= 1132798888;
assign addr[47677]= 1380375881;
assign addr[47678]= 1599979481;
assign addr[47679]= 1787159411;
assign addr[47680]= 1938122457;
assign addr[47681]= 2049809346;
assign addr[47682]= 2119956737;
assign addr[47683]= 2147143090;
assign addr[47684]= 2130817471;
assign addr[47685]= 2071310720;
assign addr[47686]= 1969828744;
assign addr[47687]= 1828428082;
assign addr[47688]= 1649974225;
assign addr[47689]= 1438083551;
assign addr[47690]= 1197050035;
assign addr[47691]= 931758235;
assign addr[47692]= 647584304;
assign addr[47693]= 350287041;
assign addr[47694]= 45891193;
assign addr[47695]= -259434643;
assign addr[47696]= -559503022;
assign addr[47697]= -848233042;
assign addr[47698]= -1119773573;
assign addr[47699]= -1368621831;
assign addr[47700]= -1589734894;
assign addr[47701]= -1778631892;
assign addr[47702]= -1931484818;
assign addr[47703]= -2045196100;
assign addr[47704]= -2117461370;
assign addr[47705]= -2146816171;
assign addr[47706]= -2132665626;
assign addr[47707]= -2075296495;
assign addr[47708]= -1975871368;
assign addr[47709]= -1836405100;
assign addr[47710]= -1659723983;
assign addr[47711]= -1449408469;
assign addr[47712]= -1209720613;
assign addr[47713]= -945517704;
assign addr[47714]= -662153826;
assign addr[47715]= -365371365;
assign addr[47716]= -61184634;
assign addr[47717]= 244242007;
assign addr[47718]= 544719071;
assign addr[47719]= 834157373;
assign addr[47720]= 1106691431;
assign addr[47721]= 1356798326;
assign addr[47722]= 1579409630;
assign addr[47723]= 1770014111;
assign addr[47724]= 1924749160;
assign addr[47725]= 2040479063;
assign addr[47726]= 2114858546;
assign addr[47727]= 2146380306;
assign addr[47728]= 2134405552;
assign addr[47729]= 2079176953;
assign addr[47730]= 1981813720;
assign addr[47731]= 1844288924;
assign addr[47732]= 1669389513;
assign addr[47733]= 1460659832;
assign addr[47734]= 1222329801;
assign addr[47735]= 959229189;
assign addr[47736]= 676689746;
assign addr[47737]= 380437148;
assign addr[47738]= 76474970;
assign addr[47739]= -229036977;
assign addr[47740]= -529907477;
assign addr[47741]= -820039373;
assign addr[47742]= -1093553126;
assign addr[47743]= -1344905966;
assign addr[47744]= -1569004214;
assign addr[47745]= -1761306505;
assign addr[47746]= -1917915825;
assign addr[47747]= -2035658475;
assign addr[47748]= -2112148396;
assign addr[47749]= -2145835515;
assign addr[47750]= -2136037160;
assign addr[47751]= -2082951896;
assign addr[47752]= -1987655498;
assign addr[47753]= -1852079154;
assign addr[47754]= -1678970324;
assign addr[47755]= -1471837070;
assign addr[47756]= -1234876957;
assign addr[47757]= -972891995;
assign addr[47758]= -691191324;
assign addr[47759]= -395483624;
assign addr[47760]= -91761426;
assign addr[47761]= 213820322;
assign addr[47762]= 515068990;
assign addr[47763]= 805879757;
assign addr[47764]= 1080359326;
assign addr[47765]= 1332945355;
assign addr[47766]= 1558519173;
assign addr[47767]= 1752509516;
assign addr[47768]= 1910985158;
assign addr[47769]= 2030734582;
assign addr[47770]= 2109331059;
assign addr[47771]= 2145181827;
assign addr[47772]= 2137560369;
assign addr[47773]= 2086621133;
assign addr[47774]= 1993396407;
assign addr[47775]= 1859775393;
assign addr[47776]= 1688465931;
assign addr[47777]= 1482939614;
assign addr[47778]= 1247361445;
assign addr[47779]= 986505429;
assign addr[47780]= 705657826;
assign addr[47781]= 410510029;
assign addr[47782]= 107043224;
assign addr[47783]= -198592817;
assign addr[47784]= -500204365;
assign addr[47785]= -791679244;
assign addr[47786]= -1067110699;
assign addr[47787]= -1320917099;
assign addr[47788]= -1547955041;
assign addr[47789]= -1743623590;
assign addr[47790]= -1903957513;
assign addr[47791]= -2025707632;
assign addr[47792]= -2106406677;
assign addr[47793]= -2144419275;
assign addr[47794]= -2138975100;
assign addr[47795]= -2090184478;
assign addr[47796]= -1999036154;
assign addr[47797]= -1867377253;
assign addr[47798]= -1697875851;
assign addr[47799]= -1493966902;
assign addr[47800]= -1259782632;
assign addr[47801]= -1000068799;
assign addr[47802]= -720088517;
assign addr[47803]= -425515602;
assign addr[47804]= -122319591;
assign addr[47805]= 183355234;
assign addr[47806]= 485314355;
assign addr[47807]= 777438554;
assign addr[47808]= 1053807919;
assign addr[47809]= 1308821808;
assign addr[47810]= 1537312353;
assign addr[47811]= 1734649179;
assign addr[47812]= 1896833245;
assign addr[47813]= 2020577882;
assign addr[47814]= 2103375398;
assign addr[47815]= 2143547897;
assign addr[47816]= 2140281282;
assign addr[47817]= 2093641749;
assign addr[47818]= 2004574453;
assign addr[47819]= 1874884346;
assign addr[47820]= 1707199606;
assign addr[47821]= 1504918373;
assign addr[47822]= 1272139887;
assign addr[47823]= 1013581418;
assign addr[47824]= 734482665;
assign addr[47825]= 440499581;
assign addr[47826]= 137589750;
assign addr[47827]= -168108346;
assign addr[47828]= -470399716;
assign addr[47829]= -763158411;
assign addr[47830]= -1040451659;
assign addr[47831]= -1296660098;
assign addr[47832]= -1526591649;
assign addr[47833]= -1725586737;
assign addr[47834]= -1889612716;
assign addr[47835]= -2015345591;
assign addr[47836]= -2100237377;
assign addr[47837]= -2142567738;
assign addr[47838]= -2141478848;
assign addr[47839]= -2096992772;
assign addr[47840]= -2010011024;
assign addr[47841]= -1882296293;
assign addr[47842]= -1716436725;
assign addr[47843]= -1515793473;
assign addr[47844]= -1284432584;
assign addr[47845]= -1027042599;
assign addr[47846]= -748839539;
assign addr[47847]= -455461206;
assign addr[47848]= -152852926;
assign addr[47849]= 152852926;
assign addr[47850]= 455461206;
assign addr[47851]= 748839539;
assign addr[47852]= 1027042599;
assign addr[47853]= 1284432584;
assign addr[47854]= 1515793473;
assign addr[47855]= 1716436725;
assign addr[47856]= 1882296293;
assign addr[47857]= 2010011024;
assign addr[47858]= 2096992772;
assign addr[47859]= 2141478848;
assign addr[47860]= 2142567738;
assign addr[47861]= 2100237377;
assign addr[47862]= 2015345591;
assign addr[47863]= 1889612716;
assign addr[47864]= 1725586737;
assign addr[47865]= 1526591649;
assign addr[47866]= 1296660098;
assign addr[47867]= 1040451659;
assign addr[47868]= 763158411;
assign addr[47869]= 470399716;
assign addr[47870]= 168108346;
assign addr[47871]= -137589750;
assign addr[47872]= -440499581;
assign addr[47873]= -734482665;
assign addr[47874]= -1013581418;
assign addr[47875]= -1272139887;
assign addr[47876]= -1504918373;
assign addr[47877]= -1707199606;
assign addr[47878]= -1874884346;
assign addr[47879]= -2004574453;
assign addr[47880]= -2093641749;
assign addr[47881]= -2140281282;
assign addr[47882]= -2143547897;
assign addr[47883]= -2103375398;
assign addr[47884]= -2020577882;
assign addr[47885]= -1896833245;
assign addr[47886]= -1734649179;
assign addr[47887]= -1537312353;
assign addr[47888]= -1308821808;
assign addr[47889]= -1053807919;
assign addr[47890]= -777438554;
assign addr[47891]= -485314355;
assign addr[47892]= -183355234;
assign addr[47893]= 122319591;
assign addr[47894]= 425515602;
assign addr[47895]= 720088517;
assign addr[47896]= 1000068799;
assign addr[47897]= 1259782632;
assign addr[47898]= 1493966902;
assign addr[47899]= 1697875851;
assign addr[47900]= 1867377253;
assign addr[47901]= 1999036154;
assign addr[47902]= 2090184478;
assign addr[47903]= 2138975100;
assign addr[47904]= 2144419275;
assign addr[47905]= 2106406677;
assign addr[47906]= 2025707632;
assign addr[47907]= 1903957513;
assign addr[47908]= 1743623590;
assign addr[47909]= 1547955041;
assign addr[47910]= 1320917099;
assign addr[47911]= 1067110699;
assign addr[47912]= 791679244;
assign addr[47913]= 500204365;
assign addr[47914]= 198592817;
assign addr[47915]= -107043224;
assign addr[47916]= -410510029;
assign addr[47917]= -705657826;
assign addr[47918]= -986505429;
assign addr[47919]= -1247361445;
assign addr[47920]= -1482939614;
assign addr[47921]= -1688465931;
assign addr[47922]= -1859775393;
assign addr[47923]= -1993396407;
assign addr[47924]= -2086621133;
assign addr[47925]= -2137560369;
assign addr[47926]= -2145181827;
assign addr[47927]= -2109331059;
assign addr[47928]= -2030734582;
assign addr[47929]= -1910985158;
assign addr[47930]= -1752509516;
assign addr[47931]= -1558519173;
assign addr[47932]= -1332945355;
assign addr[47933]= -1080359326;
assign addr[47934]= -805879757;
assign addr[47935]= -515068990;
assign addr[47936]= -213820322;
assign addr[47937]= 91761426;
assign addr[47938]= 395483624;
assign addr[47939]= 691191324;
assign addr[47940]= 972891995;
assign addr[47941]= 1234876957;
assign addr[47942]= 1471837070;
assign addr[47943]= 1678970324;
assign addr[47944]= 1852079154;
assign addr[47945]= 1987655498;
assign addr[47946]= 2082951896;
assign addr[47947]= 2136037160;
assign addr[47948]= 2145835515;
assign addr[47949]= 2112148396;
assign addr[47950]= 2035658475;
assign addr[47951]= 1917915825;
assign addr[47952]= 1761306505;
assign addr[47953]= 1569004214;
assign addr[47954]= 1344905966;
assign addr[47955]= 1093553126;
assign addr[47956]= 820039373;
assign addr[47957]= 529907477;
assign addr[47958]= 229036977;
assign addr[47959]= -76474970;
assign addr[47960]= -380437148;
assign addr[47961]= -676689746;
assign addr[47962]= -959229189;
assign addr[47963]= -1222329801;
assign addr[47964]= -1460659832;
assign addr[47965]= -1669389513;
assign addr[47966]= -1844288924;
assign addr[47967]= -1981813720;
assign addr[47968]= -2079176953;
assign addr[47969]= -2134405552;
assign addr[47970]= -2146380306;
assign addr[47971]= -2114858546;
assign addr[47972]= -2040479063;
assign addr[47973]= -1924749160;
assign addr[47974]= -1770014111;
assign addr[47975]= -1579409630;
assign addr[47976]= -1356798326;
assign addr[47977]= -1106691431;
assign addr[47978]= -834157373;
assign addr[47979]= -544719071;
assign addr[47980]= -244242007;
assign addr[47981]= 61184634;
assign addr[47982]= 365371365;
assign addr[47983]= 662153826;
assign addr[47984]= 945517704;
assign addr[47985]= 1209720613;
assign addr[47986]= 1449408469;
assign addr[47987]= 1659723983;
assign addr[47988]= 1836405100;
assign addr[47989]= 1975871368;
assign addr[47990]= 2075296495;
assign addr[47991]= 2132665626;
assign addr[47992]= 2146816171;
assign addr[47993]= 2117461370;
assign addr[47994]= 2045196100;
assign addr[47995]= 1931484818;
assign addr[47996]= 1778631892;
assign addr[47997]= 1589734894;
assign addr[47998]= 1368621831;
assign addr[47999]= 1119773573;
assign addr[48000]= 848233042;
assign addr[48001]= 559503022;
assign addr[48002]= 259434643;
assign addr[48003]= -45891193;
assign addr[48004]= -350287041;
assign addr[48005]= -647584304;
assign addr[48006]= -931758235;
assign addr[48007]= -1197050035;
assign addr[48008]= -1438083551;
assign addr[48009]= -1649974225;
assign addr[48010]= -1828428082;
assign addr[48011]= -1969828744;
assign addr[48012]= -2071310720;
assign addr[48013]= -2130817471;
assign addr[48014]= -2147143090;
assign addr[48015]= -2119956737;
assign addr[48016]= -2049809346;
assign addr[48017]= -1938122457;
assign addr[48018]= -1787159411;
assign addr[48019]= -1599979481;
assign addr[48020]= -1380375881;
assign addr[48021]= -1132798888;
assign addr[48022]= -862265664;
assign addr[48023]= -574258580;
assign addr[48024]= -274614114;
assign addr[48025]= 30595422;
assign addr[48026]= 335184940;
assign addr[48027]= 632981917;
assign addr[48028]= 917951481;
assign addr[48029]= 1184318708;
assign addr[48030]= 1426685652;
assign addr[48031]= 1640140734;
assign addr[48032]= 1820358275;
assign addr[48033]= 1963686155;
assign addr[48034]= 2067219829;
assign addr[48035]= 2128861181;
assign addr[48036]= 2147361045;
assign addr[48037]= 2122344521;
assign addr[48038]= 2054318569;
assign addr[48039]= 1944661739;
assign addr[48040]= 1795596234;
assign addr[48041]= 1610142873;
assign addr[48042]= 1392059879;
assign addr[48043]= 1145766716;
assign addr[48044]= 876254528;
assign addr[48045]= 588984994;
assign addr[48046]= 289779648;
assign addr[48047]= -15298099;
assign addr[48048]= -320065829;
assign addr[48049]= -618347408;
assign addr[48050]= -904098143;
assign addr[48051]= -1171527280;
assign addr[48052]= -1415215352;
assign addr[48053]= -1630224009;
assign addr[48054]= -1812196087;
assign addr[48055]= -1957443913;
assign addr[48056]= -2063024031;
assign addr[48057]= -2126796855;
assign addr[48058]= -2147470025;
assign addr[48059]= -2124624598;
assign addr[48060]= -2058723538;
assign addr[48061]= -1951102334;
assign addr[48062]= -1803941934;
assign addr[48063]= -1620224553;
assign addr[48064]= -1403673233;
assign addr[48065]= -1158676398;
assign addr[48066]= -890198924;
assign addr[48067]= -603681519;
assign addr[48068]= -304930476;
assign addr[48069]= 0;
assign addr[48070]= 304930476;
assign addr[48071]= 603681519;
assign addr[48072]= 890198924;
assign addr[48073]= 1158676398;
assign addr[48074]= 1403673233;
assign addr[48075]= 1620224553;
assign addr[48076]= 1803941934;
assign addr[48077]= 1951102334;
assign addr[48078]= 2058723538;
assign addr[48079]= 2124624598;
assign addr[48080]= 2147470025;
assign addr[48081]= 2126796855;
assign addr[48082]= 2063024031;
assign addr[48083]= 1957443913;
assign addr[48084]= 1812196087;
assign addr[48085]= 1630224009;
assign addr[48086]= 1415215352;
assign addr[48087]= 1171527280;
assign addr[48088]= 904098143;
assign addr[48089]= 618347408;
assign addr[48090]= 320065829;
assign addr[48091]= 15298099;
assign addr[48092]= -289779648;
assign addr[48093]= -588984994;
assign addr[48094]= -876254528;
assign addr[48095]= -1145766716;
assign addr[48096]= -1392059879;
assign addr[48097]= -1610142873;
assign addr[48098]= -1795596234;
assign addr[48099]= -1944661739;
assign addr[48100]= -2054318569;
assign addr[48101]= -2122344521;
assign addr[48102]= -2147361045;
assign addr[48103]= -2128861181;
assign addr[48104]= -2067219829;
assign addr[48105]= -1963686155;
assign addr[48106]= -1820358275;
assign addr[48107]= -1640140734;
assign addr[48108]= -1426685652;
assign addr[48109]= -1184318708;
assign addr[48110]= -917951481;
assign addr[48111]= -632981917;
assign addr[48112]= -335184940;
assign addr[48113]= -30595422;
assign addr[48114]= 274614114;
assign addr[48115]= 574258580;
assign addr[48116]= 862265664;
assign addr[48117]= 1132798888;
assign addr[48118]= 1380375881;
assign addr[48119]= 1599979481;
assign addr[48120]= 1787159411;
assign addr[48121]= 1938122457;
assign addr[48122]= 2049809346;
assign addr[48123]= 2119956737;
assign addr[48124]= 2147143090;
assign addr[48125]= 2130817471;
assign addr[48126]= 2071310720;
assign addr[48127]= 1969828744;
assign addr[48128]= 1828428082;
assign addr[48129]= 1649974225;
assign addr[48130]= 1438083551;
assign addr[48131]= 1197050035;
assign addr[48132]= 931758235;
assign addr[48133]= 647584304;
assign addr[48134]= 350287041;
assign addr[48135]= 45891193;
assign addr[48136]= -259434643;
assign addr[48137]= -559503022;
assign addr[48138]= -848233042;
assign addr[48139]= -1119773573;
assign addr[48140]= -1368621831;
assign addr[48141]= -1589734894;
assign addr[48142]= -1778631892;
assign addr[48143]= -1931484818;
assign addr[48144]= -2045196100;
assign addr[48145]= -2117461370;
assign addr[48146]= -2146816171;
assign addr[48147]= -2132665626;
assign addr[48148]= -2075296495;
assign addr[48149]= -1975871368;
assign addr[48150]= -1836405100;
assign addr[48151]= -1659723983;
assign addr[48152]= -1449408469;
assign addr[48153]= -1209720613;
assign addr[48154]= -945517704;
assign addr[48155]= -662153826;
assign addr[48156]= -365371365;
assign addr[48157]= -61184634;
assign addr[48158]= 244242007;
assign addr[48159]= 544719071;
assign addr[48160]= 834157373;
assign addr[48161]= 1106691431;
assign addr[48162]= 1356798326;
assign addr[48163]= 1579409630;
assign addr[48164]= 1770014111;
assign addr[48165]= 1924749160;
assign addr[48166]= 2040479063;
assign addr[48167]= 2114858546;
assign addr[48168]= 2146380306;
assign addr[48169]= 2134405552;
assign addr[48170]= 2079176953;
assign addr[48171]= 1981813720;
assign addr[48172]= 1844288924;
assign addr[48173]= 1669389513;
assign addr[48174]= 1460659832;
assign addr[48175]= 1222329801;
assign addr[48176]= 959229189;
assign addr[48177]= 676689746;
assign addr[48178]= 380437148;
assign addr[48179]= 76474970;
assign addr[48180]= -229036977;
assign addr[48181]= -529907477;
assign addr[48182]= -820039373;
assign addr[48183]= -1093553126;
assign addr[48184]= -1344905966;
assign addr[48185]= -1569004214;
assign addr[48186]= -1761306505;
assign addr[48187]= -1917915825;
assign addr[48188]= -2035658475;
assign addr[48189]= -2112148396;
assign addr[48190]= -2145835515;
assign addr[48191]= -2136037160;
assign addr[48192]= -2082951896;
assign addr[48193]= -1987655498;
assign addr[48194]= -1852079154;
assign addr[48195]= -1678970324;
assign addr[48196]= -1471837070;
assign addr[48197]= -1234876957;
assign addr[48198]= -972891995;
assign addr[48199]= -691191324;
assign addr[48200]= -395483624;
assign addr[48201]= -91761426;
assign addr[48202]= 213820322;
assign addr[48203]= 515068990;
assign addr[48204]= 805879757;
assign addr[48205]= 1080359326;
assign addr[48206]= 1332945355;
assign addr[48207]= 1558519173;
assign addr[48208]= 1752509516;
assign addr[48209]= 1910985158;
assign addr[48210]= 2030734582;
assign addr[48211]= 2109331059;
assign addr[48212]= 2145181827;
assign addr[48213]= 2137560369;
assign addr[48214]= 2086621133;
assign addr[48215]= 1993396407;
assign addr[48216]= 1859775393;
assign addr[48217]= 1688465931;
assign addr[48218]= 1482939614;
assign addr[48219]= 1247361445;
assign addr[48220]= 986505429;
assign addr[48221]= 705657826;
assign addr[48222]= 410510029;
assign addr[48223]= 107043224;
assign addr[48224]= -198592817;
assign addr[48225]= -500204365;
assign addr[48226]= -791679244;
assign addr[48227]= -1067110699;
assign addr[48228]= -1320917099;
assign addr[48229]= -1547955041;
assign addr[48230]= -1743623590;
assign addr[48231]= -1903957513;
assign addr[48232]= -2025707632;
assign addr[48233]= -2106406677;
assign addr[48234]= -2144419275;
assign addr[48235]= -2138975100;
assign addr[48236]= -2090184478;
assign addr[48237]= -1999036154;
assign addr[48238]= -1867377253;
assign addr[48239]= -1697875851;
assign addr[48240]= -1493966902;
assign addr[48241]= -1259782632;
assign addr[48242]= -1000068799;
assign addr[48243]= -720088517;
assign addr[48244]= -425515602;
assign addr[48245]= -122319591;
assign addr[48246]= 183355234;
assign addr[48247]= 485314355;
assign addr[48248]= 777438554;
assign addr[48249]= 1053807919;
assign addr[48250]= 1308821808;
assign addr[48251]= 1537312353;
assign addr[48252]= 1734649179;
assign addr[48253]= 1896833245;
assign addr[48254]= 2020577882;
assign addr[48255]= 2103375398;
assign addr[48256]= 2143547897;
assign addr[48257]= 2140281282;
assign addr[48258]= 2093641749;
assign addr[48259]= 2004574453;
assign addr[48260]= 1874884346;
assign addr[48261]= 1707199606;
assign addr[48262]= 1504918373;
assign addr[48263]= 1272139887;
assign addr[48264]= 1013581418;
assign addr[48265]= 734482665;
assign addr[48266]= 440499581;
assign addr[48267]= 137589750;
assign addr[48268]= -168108346;
assign addr[48269]= -470399716;
assign addr[48270]= -763158411;
assign addr[48271]= -1040451659;
assign addr[48272]= -1296660098;
assign addr[48273]= -1526591649;
assign addr[48274]= -1725586737;
assign addr[48275]= -1889612716;
assign addr[48276]= -2015345591;
assign addr[48277]= -2100237377;
assign addr[48278]= -2142567738;
assign addr[48279]= -2141478848;
assign addr[48280]= -2096992772;
assign addr[48281]= -2010011024;
assign addr[48282]= -1882296293;
assign addr[48283]= -1716436725;
assign addr[48284]= -1515793473;
assign addr[48285]= -1284432584;
assign addr[48286]= -1027042599;
assign addr[48287]= -748839539;
assign addr[48288]= -455461206;
assign addr[48289]= -152852926;
assign addr[48290]= 152852926;
assign addr[48291]= 455461206;
assign addr[48292]= 748839539;
assign addr[48293]= 1027042599;
assign addr[48294]= 1284432584;
assign addr[48295]= 1515793473;
assign addr[48296]= 1716436725;
assign addr[48297]= 1882296293;
assign addr[48298]= 2010011024;
assign addr[48299]= 2096992772;
assign addr[48300]= 2141478848;
assign addr[48301]= 2142567738;
assign addr[48302]= 2100237377;
assign addr[48303]= 2015345591;
assign addr[48304]= 1889612716;
assign addr[48305]= 1725586737;
assign addr[48306]= 1526591649;
assign addr[48307]= 1296660098;
assign addr[48308]= 1040451659;
assign addr[48309]= 763158411;
assign addr[48310]= 470399716;
assign addr[48311]= 168108346;
assign addr[48312]= -137589750;
assign addr[48313]= -440499581;
assign addr[48314]= -734482665;
assign addr[48315]= -1013581418;
assign addr[48316]= -1272139887;
assign addr[48317]= -1504918373;
assign addr[48318]= -1707199606;
assign addr[48319]= -1874884346;
assign addr[48320]= -2004574453;
assign addr[48321]= -2093641749;
assign addr[48322]= -2140281282;
assign addr[48323]= -2143547897;
assign addr[48324]= -2103375398;
assign addr[48325]= -2020577882;
assign addr[48326]= -1896833245;
assign addr[48327]= -1734649179;
assign addr[48328]= -1537312353;
assign addr[48329]= -1308821808;
assign addr[48330]= -1053807919;
assign addr[48331]= -777438554;
assign addr[48332]= -485314355;
assign addr[48333]= -183355234;
assign addr[48334]= 122319591;
assign addr[48335]= 425515602;
assign addr[48336]= 720088517;
assign addr[48337]= 1000068799;
assign addr[48338]= 1259782632;
assign addr[48339]= 1493966902;
assign addr[48340]= 1697875851;
assign addr[48341]= 1867377253;
assign addr[48342]= 1999036154;
assign addr[48343]= 2090184478;
assign addr[48344]= 2138975100;
assign addr[48345]= 2144419275;
assign addr[48346]= 2106406677;
assign addr[48347]= 2025707632;
assign addr[48348]= 1903957513;
assign addr[48349]= 1743623590;
assign addr[48350]= 1547955041;
assign addr[48351]= 1320917099;
assign addr[48352]= 1067110699;
assign addr[48353]= 791679244;
assign addr[48354]= 500204365;
assign addr[48355]= 198592817;
assign addr[48356]= -107043224;
assign addr[48357]= -410510029;
assign addr[48358]= -705657826;
assign addr[48359]= -986505429;
assign addr[48360]= -1247361445;
assign addr[48361]= -1482939614;
assign addr[48362]= -1688465931;
assign addr[48363]= -1859775393;
assign addr[48364]= -1993396407;
assign addr[48365]= -2086621133;
assign addr[48366]= -2137560369;
assign addr[48367]= -2145181827;
assign addr[48368]= -2109331059;
assign addr[48369]= -2030734582;
assign addr[48370]= -1910985158;
assign addr[48371]= -1752509516;
assign addr[48372]= -1558519173;
assign addr[48373]= -1332945355;
assign addr[48374]= -1080359326;
assign addr[48375]= -805879757;
assign addr[48376]= -515068990;
assign addr[48377]= -213820322;
assign addr[48378]= 91761426;
assign addr[48379]= 395483624;
assign addr[48380]= 691191324;
assign addr[48381]= 972891995;
assign addr[48382]= 1234876957;
assign addr[48383]= 1471837070;
assign addr[48384]= 1678970324;
assign addr[48385]= 1852079154;
assign addr[48386]= 1987655498;
assign addr[48387]= 2082951896;
assign addr[48388]= 2136037160;
assign addr[48389]= 2145835515;
assign addr[48390]= 2112148396;
assign addr[48391]= 2035658475;
assign addr[48392]= 1917915825;
assign addr[48393]= 1761306505;
assign addr[48394]= 1569004214;
assign addr[48395]= 1344905966;
assign addr[48396]= 1093553126;
assign addr[48397]= 820039373;
assign addr[48398]= 529907477;
assign addr[48399]= 229036977;
assign addr[48400]= -76474970;
assign addr[48401]= -380437148;
assign addr[48402]= -676689746;
assign addr[48403]= -959229189;
assign addr[48404]= -1222329801;
assign addr[48405]= -1460659832;
assign addr[48406]= -1669389513;
assign addr[48407]= -1844288924;
assign addr[48408]= -1981813720;
assign addr[48409]= -2079176953;
assign addr[48410]= -2134405552;
assign addr[48411]= -2146380306;
assign addr[48412]= -2114858546;
assign addr[48413]= -2040479063;
assign addr[48414]= -1924749160;
assign addr[48415]= -1770014111;
assign addr[48416]= -1579409630;
assign addr[48417]= -1356798326;
assign addr[48418]= -1106691431;
assign addr[48419]= -834157373;
assign addr[48420]= -544719071;
assign addr[48421]= -244242007;
assign addr[48422]= 61184634;
assign addr[48423]= 365371365;
assign addr[48424]= 662153826;
assign addr[48425]= 945517704;
assign addr[48426]= 1209720613;
assign addr[48427]= 1449408469;
assign addr[48428]= 1659723983;
assign addr[48429]= 1836405100;
assign addr[48430]= 1975871368;
assign addr[48431]= 2075296495;
assign addr[48432]= 2132665626;
assign addr[48433]= 2146816171;
assign addr[48434]= 2117461370;
assign addr[48435]= 2045196100;
assign addr[48436]= 1931484818;
assign addr[48437]= 1778631892;
assign addr[48438]= 1589734894;
assign addr[48439]= 1368621831;
assign addr[48440]= 1119773573;
assign addr[48441]= 848233042;
assign addr[48442]= 559503022;
assign addr[48443]= 259434643;
assign addr[48444]= -45891193;
assign addr[48445]= -350287041;
assign addr[48446]= -647584304;
assign addr[48447]= -931758235;
assign addr[48448]= -1197050035;
assign addr[48449]= -1438083551;
assign addr[48450]= -1649974225;
assign addr[48451]= -1828428082;
assign addr[48452]= -1969828744;
assign addr[48453]= -2071310720;
assign addr[48454]= -2130817471;
assign addr[48455]= -2147143090;
assign addr[48456]= -2119956737;
assign addr[48457]= -2049809346;
assign addr[48458]= -1938122457;
assign addr[48459]= -1787159411;
assign addr[48460]= -1599979481;
assign addr[48461]= -1380375881;
assign addr[48462]= -1132798888;
assign addr[48463]= -862265664;
assign addr[48464]= -574258580;
assign addr[48465]= -274614114;
assign addr[48466]= 30595422;
assign addr[48467]= 335184940;
assign addr[48468]= 632981917;
assign addr[48469]= 917951481;
assign addr[48470]= 1184318708;
assign addr[48471]= 1426685652;
assign addr[48472]= 1640140734;
assign addr[48473]= 1820358275;
assign addr[48474]= 1963686155;
assign addr[48475]= 2067219829;
assign addr[48476]= 2128861181;
assign addr[48477]= 2147361045;
assign addr[48478]= 2122344521;
assign addr[48479]= 2054318569;
assign addr[48480]= 1944661739;
assign addr[48481]= 1795596234;
assign addr[48482]= 1610142873;
assign addr[48483]= 1392059879;
assign addr[48484]= 1145766716;
assign addr[48485]= 876254528;
assign addr[48486]= 588984994;
assign addr[48487]= 289779648;
assign addr[48488]= -15298099;
assign addr[48489]= -320065829;
assign addr[48490]= -618347408;
assign addr[48491]= -904098143;
assign addr[48492]= -1171527280;
assign addr[48493]= -1415215352;
assign addr[48494]= -1630224009;
assign addr[48495]= -1812196087;
assign addr[48496]= -1957443913;
assign addr[48497]= -2063024031;
assign addr[48498]= -2126796855;
assign addr[48499]= -2147470025;
assign addr[48500]= -2124624598;
assign addr[48501]= -2058723538;
assign addr[48502]= -1951102334;
assign addr[48503]= -1803941934;
assign addr[48504]= -1620224553;
assign addr[48505]= -1403673233;
assign addr[48506]= -1158676398;
assign addr[48507]= -890198924;
assign addr[48508]= -603681519;
assign addr[48509]= -304930476;
assign addr[48510]= 0;
assign addr[48511]= 304930476;
assign addr[48512]= 603681519;
assign addr[48513]= 890198924;
assign addr[48514]= 1158676398;
assign addr[48515]= 1403673233;
assign addr[48516]= 1620224553;
assign addr[48517]= 1803941934;
assign addr[48518]= 1951102334;
assign addr[48519]= 2058723538;
assign addr[48520]= 2124624598;
assign addr[48521]= 2147470025;
assign addr[48522]= 2126796855;
assign addr[48523]= 2063024031;
assign addr[48524]= 1957443913;
assign addr[48525]= 1812196087;
assign addr[48526]= 1630224009;
assign addr[48527]= 1415215352;
assign addr[48528]= 1171527280;
assign addr[48529]= 904098143;
assign addr[48530]= 618347408;
assign addr[48531]= 320065829;
assign addr[48532]= 15298099;
assign addr[48533]= -289779648;
assign addr[48534]= -588984994;
assign addr[48535]= -876254528;
assign addr[48536]= -1145766716;
assign addr[48537]= -1392059879;
assign addr[48538]= -1610142873;
assign addr[48539]= -1795596234;
assign addr[48540]= -1944661739;
assign addr[48541]= -2054318569;
assign addr[48542]= -2122344521;
assign addr[48543]= -2147361045;
assign addr[48544]= -2128861181;
assign addr[48545]= -2067219829;
assign addr[48546]= -1963686155;
assign addr[48547]= -1820358275;
assign addr[48548]= -1640140734;
assign addr[48549]= -1426685652;
assign addr[48550]= -1184318708;
assign addr[48551]= -917951481;
assign addr[48552]= -632981917;
assign addr[48553]= -335184940;
assign addr[48554]= -30595422;
assign addr[48555]= 274614114;
assign addr[48556]= 574258580;
assign addr[48557]= 862265664;
assign addr[48558]= 1132798888;
assign addr[48559]= 1380375881;
assign addr[48560]= 1599979481;
assign addr[48561]= 1787159411;
assign addr[48562]= 1938122457;
assign addr[48563]= 2049809346;
assign addr[48564]= 2119956737;
assign addr[48565]= 2147143090;
assign addr[48566]= 2130817471;
assign addr[48567]= 2071310720;
assign addr[48568]= 1969828744;
assign addr[48569]= 1828428082;
assign addr[48570]= 1649974225;
assign addr[48571]= 1438083551;
assign addr[48572]= 1197050035;
assign addr[48573]= 931758235;
assign addr[48574]= 647584304;
assign addr[48575]= 350287041;
assign addr[48576]= 45891193;
assign addr[48577]= -259434643;
assign addr[48578]= -559503022;
assign addr[48579]= -848233042;
assign addr[48580]= -1119773573;
assign addr[48581]= -1368621831;
assign addr[48582]= -1589734894;
assign addr[48583]= -1778631892;
assign addr[48584]= -1931484818;
assign addr[48585]= -2045196100;
assign addr[48586]= -2117461370;
assign addr[48587]= -2146816171;
assign addr[48588]= -2132665626;
assign addr[48589]= -2075296495;
assign addr[48590]= -1975871368;
assign addr[48591]= -1836405100;
assign addr[48592]= -1659723983;
assign addr[48593]= -1449408469;
assign addr[48594]= -1209720613;
assign addr[48595]= -945517704;
assign addr[48596]= -662153826;
assign addr[48597]= -365371365;
assign addr[48598]= -61184634;
assign addr[48599]= 244242007;
assign addr[48600]= 544719071;
assign addr[48601]= 834157373;
assign addr[48602]= 1106691431;
assign addr[48603]= 1356798326;
assign addr[48604]= 1579409630;
assign addr[48605]= 1770014111;
assign addr[48606]= 1924749160;
assign addr[48607]= 2040479063;
assign addr[48608]= 2114858546;
assign addr[48609]= 2146380306;
assign addr[48610]= 2134405552;
assign addr[48611]= 2079176953;
assign addr[48612]= 1981813720;
assign addr[48613]= 1844288924;
assign addr[48614]= 1669389513;
assign addr[48615]= 1460659832;
assign addr[48616]= 1222329801;
assign addr[48617]= 959229189;
assign addr[48618]= 676689746;
assign addr[48619]= 380437148;
assign addr[48620]= 76474970;
assign addr[48621]= -229036977;
assign addr[48622]= -529907477;
assign addr[48623]= -820039373;
assign addr[48624]= -1093553126;
assign addr[48625]= -1344905966;
assign addr[48626]= -1569004214;
assign addr[48627]= -1761306505;
assign addr[48628]= -1917915825;
assign addr[48629]= -2035658475;
assign addr[48630]= -2112148396;
assign addr[48631]= -2145835515;
assign addr[48632]= -2136037160;
assign addr[48633]= -2082951896;
assign addr[48634]= -1987655498;
assign addr[48635]= -1852079154;
assign addr[48636]= -1678970324;
assign addr[48637]= -1471837070;
assign addr[48638]= -1234876957;
assign addr[48639]= -972891995;
assign addr[48640]= -691191324;
assign addr[48641]= -395483624;
assign addr[48642]= -91761426;
assign addr[48643]= 213820322;
assign addr[48644]= 515068990;
assign addr[48645]= 805879757;
assign addr[48646]= 1080359326;
assign addr[48647]= 1332945355;
assign addr[48648]= 1558519173;
assign addr[48649]= 1752509516;
assign addr[48650]= 1910985158;
assign addr[48651]= 2030734582;
assign addr[48652]= 2109331059;
assign addr[48653]= 2145181827;
assign addr[48654]= 2137560369;
assign addr[48655]= 2086621133;
assign addr[48656]= 1993396407;
assign addr[48657]= 1859775393;
assign addr[48658]= 1688465931;
assign addr[48659]= 1482939614;
assign addr[48660]= 1247361445;
assign addr[48661]= 986505429;
assign addr[48662]= 705657826;
assign addr[48663]= 410510029;
assign addr[48664]= 107043224;
assign addr[48665]= -198592817;
assign addr[48666]= -500204365;
assign addr[48667]= -791679244;
assign addr[48668]= -1067110699;
assign addr[48669]= -1320917099;
assign addr[48670]= -1547955041;
assign addr[48671]= -1743623590;
assign addr[48672]= -1903957513;
assign addr[48673]= -2025707632;
assign addr[48674]= -2106406677;
assign addr[48675]= -2144419275;
assign addr[48676]= -2138975100;
assign addr[48677]= -2090184478;
assign addr[48678]= -1999036154;
assign addr[48679]= -1867377253;
assign addr[48680]= -1697875851;
assign addr[48681]= -1493966902;
assign addr[48682]= -1259782632;
assign addr[48683]= -1000068799;
assign addr[48684]= -720088517;
assign addr[48685]= -425515602;
assign addr[48686]= -122319591;
assign addr[48687]= 183355234;
assign addr[48688]= 485314355;
assign addr[48689]= 777438554;
assign addr[48690]= 1053807919;
assign addr[48691]= 1308821808;
assign addr[48692]= 1537312353;
assign addr[48693]= 1734649179;
assign addr[48694]= 1896833245;
assign addr[48695]= 2020577882;
assign addr[48696]= 2103375398;
assign addr[48697]= 2143547897;
assign addr[48698]= 2140281282;
assign addr[48699]= 2093641749;
assign addr[48700]= 2004574453;
assign addr[48701]= 1874884346;
assign addr[48702]= 1707199606;
assign addr[48703]= 1504918373;
assign addr[48704]= 1272139887;
assign addr[48705]= 1013581418;
assign addr[48706]= 734482665;
assign addr[48707]= 440499581;
assign addr[48708]= 137589750;
assign addr[48709]= -168108346;
assign addr[48710]= -470399716;
assign addr[48711]= -763158411;
assign addr[48712]= -1040451659;
assign addr[48713]= -1296660098;
assign addr[48714]= -1526591649;
assign addr[48715]= -1725586737;
assign addr[48716]= -1889612716;
assign addr[48717]= -2015345591;
assign addr[48718]= -2100237377;
assign addr[48719]= -2142567738;
assign addr[48720]= -2141478848;
assign addr[48721]= -2096992772;
assign addr[48722]= -2010011024;
assign addr[48723]= -1882296293;
assign addr[48724]= -1716436725;
assign addr[48725]= -1515793473;
assign addr[48726]= -1284432584;
assign addr[48727]= -1027042599;
assign addr[48728]= -748839539;
assign addr[48729]= -455461206;
assign addr[48730]= -152852926;
assign addr[48731]= 152852926;
assign addr[48732]= 455461206;
assign addr[48733]= 748839539;
assign addr[48734]= 1027042599;
assign addr[48735]= 1284432584;
assign addr[48736]= 1515793473;
assign addr[48737]= 1716436725;
assign addr[48738]= 1882296293;
assign addr[48739]= 2010011024;
assign addr[48740]= 2096992772;
assign addr[48741]= 2141478848;
assign addr[48742]= 2142567738;
assign addr[48743]= 2100237377;
assign addr[48744]= 2015345591;
assign addr[48745]= 1889612716;
assign addr[48746]= 1725586737;
assign addr[48747]= 1526591649;
assign addr[48748]= 1296660098;
assign addr[48749]= 1040451659;
assign addr[48750]= 763158411;
assign addr[48751]= 470399716;
assign addr[48752]= 168108346;
assign addr[48753]= -137589750;
assign addr[48754]= -440499581;
assign addr[48755]= -734482665;
assign addr[48756]= -1013581418;
assign addr[48757]= -1272139887;
assign addr[48758]= -1504918373;
assign addr[48759]= -1707199606;
assign addr[48760]= -1874884346;
assign addr[48761]= -2004574453;
assign addr[48762]= -2093641749;
assign addr[48763]= -2140281282;
assign addr[48764]= -2143547897;
assign addr[48765]= -2103375398;
assign addr[48766]= -2020577882;
assign addr[48767]= -1896833245;
assign addr[48768]= -1734649179;
assign addr[48769]= -1537312353;
assign addr[48770]= -1308821808;
assign addr[48771]= -1053807919;
assign addr[48772]= -777438554;
assign addr[48773]= -485314355;
assign addr[48774]= -183355234;
assign addr[48775]= 122319591;
assign addr[48776]= 425515602;
assign addr[48777]= 720088517;
assign addr[48778]= 1000068799;
assign addr[48779]= 1259782632;
assign addr[48780]= 1493966902;
assign addr[48781]= 1697875851;
assign addr[48782]= 1867377253;
assign addr[48783]= 1999036154;
assign addr[48784]= 2090184478;
assign addr[48785]= 2138975100;
assign addr[48786]= 2144419275;
assign addr[48787]= 2106406677;
assign addr[48788]= 2025707632;
assign addr[48789]= 1903957513;
assign addr[48790]= 1743623590;
assign addr[48791]= 1547955041;
assign addr[48792]= 1320917099;
assign addr[48793]= 1067110699;
assign addr[48794]= 791679244;
assign addr[48795]= 500204365;
assign addr[48796]= 198592817;
assign addr[48797]= -107043224;
assign addr[48798]= -410510029;
assign addr[48799]= -705657826;
assign addr[48800]= -986505429;
assign addr[48801]= -1247361445;
assign addr[48802]= -1482939614;
assign addr[48803]= -1688465931;
assign addr[48804]= -1859775393;
assign addr[48805]= -1993396407;
assign addr[48806]= -2086621133;
assign addr[48807]= -2137560369;
assign addr[48808]= -2145181827;
assign addr[48809]= -2109331059;
assign addr[48810]= -2030734582;
assign addr[48811]= -1910985158;
assign addr[48812]= -1752509516;
assign addr[48813]= -1558519173;
assign addr[48814]= -1332945355;
assign addr[48815]= -1080359326;
assign addr[48816]= -805879757;
assign addr[48817]= -515068990;
assign addr[48818]= -213820322;
assign addr[48819]= 91761426;
assign addr[48820]= 395483624;
assign addr[48821]= 691191324;
assign addr[48822]= 972891995;
assign addr[48823]= 1234876957;
assign addr[48824]= 1471837070;
assign addr[48825]= 1678970324;
assign addr[48826]= 1852079154;
assign addr[48827]= 1987655498;
assign addr[48828]= 2082951896;
assign addr[48829]= 2136037160;
assign addr[48830]= 2145835515;
assign addr[48831]= 2112148396;
assign addr[48832]= 2035658475;
assign addr[48833]= 1917915825;
assign addr[48834]= 1761306505;
assign addr[48835]= 1569004214;
assign addr[48836]= 1344905966;
assign addr[48837]= 1093553126;
assign addr[48838]= 820039373;
assign addr[48839]= 529907477;
assign addr[48840]= 229036977;
assign addr[48841]= -76474970;
assign addr[48842]= -380437148;
assign addr[48843]= -676689746;
assign addr[48844]= -959229189;
assign addr[48845]= -1222329801;
assign addr[48846]= -1460659832;
assign addr[48847]= -1669389513;
assign addr[48848]= -1844288924;
assign addr[48849]= -1981813720;
assign addr[48850]= -2079176953;
assign addr[48851]= -2134405552;
assign addr[48852]= -2146380306;
assign addr[48853]= -2114858546;
assign addr[48854]= -2040479063;
assign addr[48855]= -1924749160;
assign addr[48856]= -1770014111;
assign addr[48857]= -1579409630;
assign addr[48858]= -1356798326;
assign addr[48859]= -1106691431;
assign addr[48860]= -834157373;
assign addr[48861]= -544719071;
assign addr[48862]= -244242007;
assign addr[48863]= 61184634;
assign addr[48864]= 365371365;
assign addr[48865]= 662153826;
assign addr[48866]= 945517704;
assign addr[48867]= 1209720613;
assign addr[48868]= 1449408469;
assign addr[48869]= 1659723983;
assign addr[48870]= 1836405100;
assign addr[48871]= 1975871368;
assign addr[48872]= 2075296495;
assign addr[48873]= 2132665626;
assign addr[48874]= 2146816171;
assign addr[48875]= 2117461370;
assign addr[48876]= 2045196100;
assign addr[48877]= 1931484818;
assign addr[48878]= 1778631892;
assign addr[48879]= 1589734894;
assign addr[48880]= 1368621831;
assign addr[48881]= 1119773573;
assign addr[48882]= 848233042;
assign addr[48883]= 559503022;
assign addr[48884]= 259434643;
assign addr[48885]= -45891193;
assign addr[48886]= -350287041;
assign addr[48887]= -647584304;
assign addr[48888]= -931758235;
assign addr[48889]= -1197050035;
assign addr[48890]= -1438083551;
assign addr[48891]= -1649974225;
assign addr[48892]= -1828428082;
assign addr[48893]= -1969828744;
assign addr[48894]= -2071310720;
assign addr[48895]= -2130817471;
assign addr[48896]= -2147143090;
assign addr[48897]= -2119956737;
assign addr[48898]= -2049809346;
assign addr[48899]= -1938122457;
assign addr[48900]= -1787159411;
assign addr[48901]= -1599979481;
assign addr[48902]= -1380375881;
assign addr[48903]= -1132798888;
assign addr[48904]= -862265664;
assign addr[48905]= -574258580;
assign addr[48906]= -274614114;
assign addr[48907]= 30595422;
assign addr[48908]= 335184940;
assign addr[48909]= 632981917;
assign addr[48910]= 917951481;
assign addr[48911]= 1184318708;
assign addr[48912]= 1426685652;
assign addr[48913]= 1640140734;
assign addr[48914]= 1820358275;
assign addr[48915]= 1963686155;
assign addr[48916]= 2067219829;
assign addr[48917]= 2128861181;
assign addr[48918]= 2147361045;
assign addr[48919]= 2122344521;
assign addr[48920]= 2054318569;
assign addr[48921]= 1944661739;
assign addr[48922]= 1795596234;
assign addr[48923]= 1610142873;
assign addr[48924]= 1392059879;
assign addr[48925]= 1145766716;
assign addr[48926]= 876254528;
assign addr[48927]= 588984994;
assign addr[48928]= 289779648;
assign addr[48929]= -15298099;
assign addr[48930]= -320065829;
assign addr[48931]= -618347408;
assign addr[48932]= -904098143;
assign addr[48933]= -1171527280;
assign addr[48934]= -1415215352;
assign addr[48935]= -1630224009;
assign addr[48936]= -1812196087;
assign addr[48937]= -1957443913;
assign addr[48938]= -2063024031;
assign addr[48939]= -2126796855;
assign addr[48940]= -2147470025;
assign addr[48941]= -2124624598;
assign addr[48942]= -2058723538;
assign addr[48943]= -1951102334;
assign addr[48944]= -1803941934;
assign addr[48945]= -1620224553;
assign addr[48946]= -1403673233;
assign addr[48947]= -1158676398;
assign addr[48948]= -890198924;
assign addr[48949]= -603681519;
assign addr[48950]= -304930476;
assign addr[48951]= 0;
assign addr[48952]= 304930476;
assign addr[48953]= 603681519;
assign addr[48954]= 890198924;
assign addr[48955]= 1158676398;
assign addr[48956]= 1403673233;
assign addr[48957]= 1620224553;
assign addr[48958]= 1803941934;
assign addr[48959]= 1951102334;
assign addr[48960]= 2058723538;
assign addr[48961]= 2124624598;
assign addr[48962]= 2147470025;
assign addr[48963]= 2126796855;
assign addr[48964]= 2063024031;
assign addr[48965]= 1957443913;
assign addr[48966]= 1812196087;
assign addr[48967]= 1630224009;
assign addr[48968]= 1415215352;
assign addr[48969]= 1171527280;
assign addr[48970]= 904098143;
assign addr[48971]= 618347408;
assign addr[48972]= 320065829;
assign addr[48973]= 15298099;
assign addr[48974]= -289779648;
assign addr[48975]= -588984994;
assign addr[48976]= -876254528;
assign addr[48977]= -1145766716;
assign addr[48978]= -1392059879;
assign addr[48979]= -1610142873;
assign addr[48980]= -1795596234;
assign addr[48981]= -1944661739;
assign addr[48982]= -2054318569;
assign addr[48983]= -2122344521;
assign addr[48984]= -2147361045;
assign addr[48985]= -2128861181;
assign addr[48986]= -2067219829;
assign addr[48987]= -1963686155;
assign addr[48988]= -1820358275;
assign addr[48989]= -1640140734;
assign addr[48990]= -1426685652;
assign addr[48991]= -1184318708;
assign addr[48992]= -917951481;
assign addr[48993]= -632981917;
assign addr[48994]= -335184940;
assign addr[48995]= -30595422;
assign addr[48996]= 274614114;
assign addr[48997]= 574258580;
assign addr[48998]= 862265664;
assign addr[48999]= 1132798888;
assign addr[49000]= 1380375881;
assign addr[49001]= 1599979481;
assign addr[49002]= 1787159411;
assign addr[49003]= 1938122457;
assign addr[49004]= 2049809346;
assign addr[49005]= 2119956737;
assign addr[49006]= 2147143090;
assign addr[49007]= 2130817471;
assign addr[49008]= 2071310720;
assign addr[49009]= 1969828744;
assign addr[49010]= 1828428082;
assign addr[49011]= 1649974225;
assign addr[49012]= 1438083551;
assign addr[49013]= 1197050035;
assign addr[49014]= 931758235;
assign addr[49015]= 647584304;
assign addr[49016]= 350287041;
assign addr[49017]= 45891193;
assign addr[49018]= -259434643;
assign addr[49019]= -559503022;
assign addr[49020]= -848233042;
assign addr[49021]= -1119773573;
assign addr[49022]= -1368621831;
assign addr[49023]= -1589734894;
assign addr[49024]= -1778631892;
assign addr[49025]= -1931484818;
assign addr[49026]= -2045196100;
assign addr[49027]= -2117461370;
assign addr[49028]= -2146816171;
assign addr[49029]= -2132665626;
assign addr[49030]= -2075296495;
assign addr[49031]= -1975871368;
assign addr[49032]= -1836405100;
assign addr[49033]= -1659723983;
assign addr[49034]= -1449408469;
assign addr[49035]= -1209720613;
assign addr[49036]= -945517704;
assign addr[49037]= -662153826;
assign addr[49038]= -365371365;
assign addr[49039]= -61184634;
assign addr[49040]= 244242007;
assign addr[49041]= 544719071;
assign addr[49042]= 834157373;
assign addr[49043]= 1106691431;
assign addr[49044]= 1356798326;
assign addr[49045]= 1579409630;
assign addr[49046]= 1770014111;
assign addr[49047]= 1924749160;
assign addr[49048]= 2040479063;
assign addr[49049]= 2114858546;
assign addr[49050]= 2146380306;
assign addr[49051]= 2134405552;
assign addr[49052]= 2079176953;
assign addr[49053]= 1981813720;
assign addr[49054]= 1844288924;
assign addr[49055]= 1669389513;
assign addr[49056]= 1460659832;
assign addr[49057]= 1222329801;
assign addr[49058]= 959229189;
assign addr[49059]= 676689746;
assign addr[49060]= 380437148;
assign addr[49061]= 76474970;
assign addr[49062]= -229036977;
assign addr[49063]= -529907477;
assign addr[49064]= -820039373;
assign addr[49065]= -1093553126;
assign addr[49066]= -1344905966;
assign addr[49067]= -1569004214;
assign addr[49068]= -1761306505;
assign addr[49069]= -1917915825;
assign addr[49070]= -2035658475;
assign addr[49071]= -2112148396;
assign addr[49072]= -2145835515;
assign addr[49073]= -2136037160;
assign addr[49074]= -2082951896;
assign addr[49075]= -1987655498;
assign addr[49076]= -1852079154;
assign addr[49077]= -1678970324;
assign addr[49078]= -1471837070;
assign addr[49079]= -1234876957;
assign addr[49080]= -972891995;
assign addr[49081]= -691191324;
assign addr[49082]= -395483624;
assign addr[49083]= -91761426;
assign addr[49084]= 213820322;
assign addr[49085]= 515068990;
assign addr[49086]= 805879757;
assign addr[49087]= 1080359326;
assign addr[49088]= 1332945355;
assign addr[49089]= 1558519173;
assign addr[49090]= 1752509516;
assign addr[49091]= 1910985158;
assign addr[49092]= 2030734582;
assign addr[49093]= 2109331059;
assign addr[49094]= 2145181827;
assign addr[49095]= 2137560369;
assign addr[49096]= 2086621133;
assign addr[49097]= 1993396407;
assign addr[49098]= 1859775393;
assign addr[49099]= 1688465931;
assign addr[49100]= 1482939614;
assign addr[49101]= 1247361445;
assign addr[49102]= 986505429;
assign addr[49103]= 705657826;
assign addr[49104]= 410510029;
assign addr[49105]= 107043224;
assign addr[49106]= -198592817;
assign addr[49107]= -500204365;
assign addr[49108]= -791679244;
assign addr[49109]= -1067110699;
assign addr[49110]= -1320917099;
assign addr[49111]= -1547955041;
assign addr[49112]= -1743623590;
assign addr[49113]= -1903957513;
assign addr[49114]= -2025707632;
assign addr[49115]= -2106406677;
assign addr[49116]= -2144419275;
assign addr[49117]= -2138975100;
assign addr[49118]= -2090184478;
assign addr[49119]= -1999036154;
assign addr[49120]= -1867377253;
assign addr[49121]= -1697875851;
assign addr[49122]= -1493966902;
assign addr[49123]= -1259782632;
assign addr[49124]= -1000068799;
assign addr[49125]= -720088517;
assign addr[49126]= -425515602;
assign addr[49127]= -122319591;
assign addr[49128]= 183355234;
assign addr[49129]= 485314355;
assign addr[49130]= 777438554;
assign addr[49131]= 1053807919;
assign addr[49132]= 1308821808;
assign addr[49133]= 1537312353;
assign addr[49134]= 1734649179;
assign addr[49135]= 1896833245;
assign addr[49136]= 2020577882;
assign addr[49137]= 2103375398;
assign addr[49138]= 2143547897;
assign addr[49139]= 2140281282;
assign addr[49140]= 2093641749;
assign addr[49141]= 2004574453;
assign addr[49142]= 1874884346;
assign addr[49143]= 1707199606;
assign addr[49144]= 1504918373;
assign addr[49145]= 1272139887;
assign addr[49146]= 1013581418;
assign addr[49147]= 734482665;
assign addr[49148]= 440499581;
assign addr[49149]= 137589750;
assign addr[49150]= -168108346;
assign addr[49151]= -470399716;
assign addr[49152]= -763158411;
assign addr[49153]= -1040451659;
assign addr[49154]= -1296660098;
assign addr[49155]= -1526591649;
assign addr[49156]= -1725586737;
assign addr[49157]= -1889612716;
assign addr[49158]= -2015345591;
assign addr[49159]= -2100237377;
assign addr[49160]= -2142567738;
assign addr[49161]= -2141478848;
assign addr[49162]= -2096992772;
assign addr[49163]= -2010011024;
assign addr[49164]= -1882296293;
assign addr[49165]= -1716436725;
assign addr[49166]= -1515793473;
assign addr[49167]= -1284432584;
assign addr[49168]= -1027042599;
assign addr[49169]= -748839539;
assign addr[49170]= -455461206;
assign addr[49171]= -152852926;
assign addr[49172]= 152852926;
assign addr[49173]= 455461206;
assign addr[49174]= 748839539;
assign addr[49175]= 1027042599;
assign addr[49176]= 1284432584;
assign addr[49177]= 1515793473;
assign addr[49178]= 1716436725;
assign addr[49179]= 1882296293;
assign addr[49180]= 2010011024;
assign addr[49181]= 2096992772;
assign addr[49182]= 2141478848;
assign addr[49183]= 2142567738;
assign addr[49184]= 2100237377;
assign addr[49185]= 2015345591;
assign addr[49186]= 1889612716;
assign addr[49187]= 1725586737;
assign addr[49188]= 1526591649;
assign addr[49189]= 1296660098;
assign addr[49190]= 1040451659;
assign addr[49191]= 763158411;
assign addr[49192]= 470399716;
assign addr[49193]= 168108346;
assign addr[49194]= -137589750;
assign addr[49195]= -440499581;
assign addr[49196]= -734482665;
assign addr[49197]= -1013581418;
assign addr[49198]= -1272139887;
assign addr[49199]= -1504918373;
assign addr[49200]= -1707199606;
assign addr[49201]= -1874884346;
assign addr[49202]= -2004574453;
assign addr[49203]= -2093641749;
assign addr[49204]= -2140281282;
assign addr[49205]= -2143547897;
assign addr[49206]= -2103375398;
assign addr[49207]= -2020577882;
assign addr[49208]= -1896833245;
assign addr[49209]= -1734649179;
assign addr[49210]= -1537312353;
assign addr[49211]= -1308821808;
assign addr[49212]= -1053807919;
assign addr[49213]= -777438554;
assign addr[49214]= -485314355;
assign addr[49215]= -183355234;
assign addr[49216]= 122319591;
assign addr[49217]= 425515602;
assign addr[49218]= 720088517;
assign addr[49219]= 1000068799;
assign addr[49220]= 1259782632;
assign addr[49221]= 1493966902;
assign addr[49222]= 1697875851;
assign addr[49223]= 1867377253;
assign addr[49224]= 1999036154;
assign addr[49225]= 2090184478;
assign addr[49226]= 2138975100;
assign addr[49227]= 2144419275;
assign addr[49228]= 2106406677;
assign addr[49229]= 2025707632;
assign addr[49230]= 1903957513;
assign addr[49231]= 1743623590;
assign addr[49232]= 1547955041;
assign addr[49233]= 1320917099;
assign addr[49234]= 1067110699;
assign addr[49235]= 791679244;
assign addr[49236]= 500204365;
assign addr[49237]= 198592817;
assign addr[49238]= -107043224;
assign addr[49239]= -410510029;
assign addr[49240]= -705657826;
assign addr[49241]= -986505429;
assign addr[49242]= -1247361445;
assign addr[49243]= -1482939614;
assign addr[49244]= -1688465931;
assign addr[49245]= -1859775393;
assign addr[49246]= -1993396407;
assign addr[49247]= -2086621133;
assign addr[49248]= -2137560369;
assign addr[49249]= -2145181827;
assign addr[49250]= -2109331059;
assign addr[49251]= -2030734582;
assign addr[49252]= -1910985158;
assign addr[49253]= -1752509516;
assign addr[49254]= -1558519173;
assign addr[49255]= -1332945355;
assign addr[49256]= -1080359326;
assign addr[49257]= -805879757;
assign addr[49258]= -515068990;
assign addr[49259]= -213820322;
assign addr[49260]= 91761426;
assign addr[49261]= 395483624;
assign addr[49262]= 691191324;
assign addr[49263]= 972891995;
assign addr[49264]= 1234876957;
assign addr[49265]= 1471837070;
assign addr[49266]= 1678970324;
assign addr[49267]= 1852079154;
assign addr[49268]= 1987655498;
assign addr[49269]= 2082951896;
assign addr[49270]= 2136037160;
assign addr[49271]= 2145835515;
assign addr[49272]= 2112148396;
assign addr[49273]= 2035658475;
assign addr[49274]= 1917915825;
assign addr[49275]= 1761306505;
assign addr[49276]= 1569004214;
assign addr[49277]= 1344905966;
assign addr[49278]= 1093553126;
assign addr[49279]= 820039373;
assign addr[49280]= 529907477;
assign addr[49281]= 229036977;
assign addr[49282]= -76474970;
assign addr[49283]= -380437148;
assign addr[49284]= -676689746;
assign addr[49285]= -959229189;
assign addr[49286]= -1222329801;
assign addr[49287]= -1460659832;
assign addr[49288]= -1669389513;
assign addr[49289]= -1844288924;
assign addr[49290]= -1981813720;
assign addr[49291]= -2079176953;
assign addr[49292]= -2134405552;
assign addr[49293]= -2146380306;
assign addr[49294]= -2114858546;
assign addr[49295]= -2040479063;
assign addr[49296]= -1924749160;
assign addr[49297]= -1770014111;
assign addr[49298]= -1579409630;
assign addr[49299]= -1356798326;
assign addr[49300]= -1106691431;
assign addr[49301]= -834157373;
assign addr[49302]= -544719071;
assign addr[49303]= -244242007;
assign addr[49304]= 61184634;
assign addr[49305]= 365371365;
assign addr[49306]= 662153826;
assign addr[49307]= 945517704;
assign addr[49308]= 1209720613;
assign addr[49309]= 1449408469;
assign addr[49310]= 1659723983;
assign addr[49311]= 1836405100;
assign addr[49312]= 1975871368;
assign addr[49313]= 2075296495;
assign addr[49314]= 2132665626;
assign addr[49315]= 2146816171;
assign addr[49316]= 2117461370;
assign addr[49317]= 2045196100;
assign addr[49318]= 1931484818;
assign addr[49319]= 1778631892;
assign addr[49320]= 1589734894;
assign addr[49321]= 1368621831;
assign addr[49322]= 1119773573;
assign addr[49323]= 848233042;
assign addr[49324]= 559503022;
assign addr[49325]= 259434643;
assign addr[49326]= -45891193;
assign addr[49327]= -350287041;
assign addr[49328]= -647584304;
assign addr[49329]= -931758235;
assign addr[49330]= -1197050035;
assign addr[49331]= -1438083551;
assign addr[49332]= -1649974225;
assign addr[49333]= -1828428082;
assign addr[49334]= -1969828744;
assign addr[49335]= -2071310720;
assign addr[49336]= -2130817471;
assign addr[49337]= -2147143090;
assign addr[49338]= -2119956737;
assign addr[49339]= -2049809346;
assign addr[49340]= -1938122457;
assign addr[49341]= -1787159411;
assign addr[49342]= -1599979481;
assign addr[49343]= -1380375881;
assign addr[49344]= -1132798888;
assign addr[49345]= -862265664;
assign addr[49346]= -574258580;
assign addr[49347]= -274614114;
assign addr[49348]= 30595422;
assign addr[49349]= 335184940;
assign addr[49350]= 632981917;
assign addr[49351]= 917951481;
assign addr[49352]= 1184318708;
assign addr[49353]= 1426685652;
assign addr[49354]= 1640140734;
assign addr[49355]= 1820358275;
assign addr[49356]= 1963686155;
assign addr[49357]= 2067219829;
assign addr[49358]= 2128861181;
assign addr[49359]= 2147361045;
assign addr[49360]= 2122344521;
assign addr[49361]= 2054318569;
assign addr[49362]= 1944661739;
assign addr[49363]= 1795596234;
assign addr[49364]= 1610142873;
assign addr[49365]= 1392059879;
assign addr[49366]= 1145766716;
assign addr[49367]= 876254528;
assign addr[49368]= 588984994;
assign addr[49369]= 289779648;
assign addr[49370]= -15298099;
assign addr[49371]= -320065829;
assign addr[49372]= -618347408;
assign addr[49373]= -904098143;
assign addr[49374]= -1171527280;
assign addr[49375]= -1415215352;
assign addr[49376]= -1630224009;
assign addr[49377]= -1812196087;
assign addr[49378]= -1957443913;
assign addr[49379]= -2063024031;
assign addr[49380]= -2126796855;
assign addr[49381]= -2147470025;
assign addr[49382]= -2124624598;
assign addr[49383]= -2058723538;
assign addr[49384]= -1951102334;
assign addr[49385]= -1803941934;
assign addr[49386]= -1620224553;
assign addr[49387]= -1403673233;
assign addr[49388]= -1158676398;
assign addr[49389]= -890198924;
assign addr[49390]= -603681519;
assign addr[49391]= -304930476;
assign addr[49392]= 0;
assign addr[49393]= 304930476;
assign addr[49394]= 603681519;
assign addr[49395]= 890198924;
assign addr[49396]= 1158676398;
assign addr[49397]= 1403673233;
assign addr[49398]= 1620224553;
assign addr[49399]= 1803941934;
assign addr[49400]= 1951102334;
assign addr[49401]= 2058723538;
assign addr[49402]= 2124624598;
assign addr[49403]= 2147470025;
assign addr[49404]= 2126796855;
assign addr[49405]= 2063024031;
assign addr[49406]= 1957443913;
assign addr[49407]= 1812196087;
assign addr[49408]= 1630224009;
assign addr[49409]= 1415215352;
assign addr[49410]= 1171527280;
assign addr[49411]= 904098143;
assign addr[49412]= 618347408;
assign addr[49413]= 320065829;
assign addr[49414]= 15298099;
assign addr[49415]= -289779648;
assign addr[49416]= -588984994;
assign addr[49417]= -876254528;
assign addr[49418]= -1145766716;
assign addr[49419]= -1392059879;
assign addr[49420]= -1610142873;
assign addr[49421]= -1795596234;
assign addr[49422]= -1944661739;
assign addr[49423]= -2054318569;
assign addr[49424]= -2122344521;
assign addr[49425]= -2147361045;
assign addr[49426]= -2128861181;
assign addr[49427]= -2067219829;
assign addr[49428]= -1963686155;
assign addr[49429]= -1820358275;
assign addr[49430]= -1640140734;
assign addr[49431]= -1426685652;
assign addr[49432]= -1184318708;
assign addr[49433]= -917951481;
assign addr[49434]= -632981917;
assign addr[49435]= -335184940;
assign addr[49436]= -30595422;
assign addr[49437]= 274614114;
assign addr[49438]= 574258580;
assign addr[49439]= 862265664;
assign addr[49440]= 1132798888;
assign addr[49441]= 1380375881;
assign addr[49442]= 1599979481;
assign addr[49443]= 1787159411;
assign addr[49444]= 1938122457;
assign addr[49445]= 2049809346;
assign addr[49446]= 2119956737;
assign addr[49447]= 2147143090;
assign addr[49448]= 2130817471;
assign addr[49449]= 2071310720;
assign addr[49450]= 1969828744;
assign addr[49451]= 1828428082;
assign addr[49452]= 1649974225;
assign addr[49453]= 1438083551;
assign addr[49454]= 1197050035;
assign addr[49455]= 931758235;
assign addr[49456]= 647584304;
assign addr[49457]= 350287041;
assign addr[49458]= 45891193;
assign addr[49459]= -259434643;
assign addr[49460]= -559503022;
assign addr[49461]= -848233042;
assign addr[49462]= -1119773573;
assign addr[49463]= -1368621831;
assign addr[49464]= -1589734894;
assign addr[49465]= -1778631892;
assign addr[49466]= -1931484818;
assign addr[49467]= -2045196100;
assign addr[49468]= -2117461370;
assign addr[49469]= -2146816171;
assign addr[49470]= -2132665626;
assign addr[49471]= -2075296495;
assign addr[49472]= -1975871368;
assign addr[49473]= -1836405100;
assign addr[49474]= -1659723983;
assign addr[49475]= -1449408469;
assign addr[49476]= -1209720613;
assign addr[49477]= -945517704;
assign addr[49478]= -662153826;
assign addr[49479]= -365371365;
assign addr[49480]= -61184634;
assign addr[49481]= 244242007;
assign addr[49482]= 544719071;
assign addr[49483]= 834157373;
assign addr[49484]= 1106691431;
assign addr[49485]= 1356798326;
assign addr[49486]= 1579409630;
assign addr[49487]= 1770014111;
assign addr[49488]= 1924749160;
assign addr[49489]= 2040479063;
assign addr[49490]= 2114858546;
assign addr[49491]= 2146380306;
assign addr[49492]= 2134405552;
assign addr[49493]= 2079176953;
assign addr[49494]= 1981813720;
assign addr[49495]= 1844288924;
assign addr[49496]= 1669389513;
assign addr[49497]= 1460659832;
assign addr[49498]= 1222329801;
assign addr[49499]= 959229189;
assign addr[49500]= 676689746;
assign addr[49501]= 380437148;
assign addr[49502]= 76474970;
assign addr[49503]= -229036977;
assign addr[49504]= -529907477;
assign addr[49505]= -820039373;
assign addr[49506]= -1093553126;
assign addr[49507]= -1344905966;
assign addr[49508]= -1569004214;
assign addr[49509]= -1761306505;
assign addr[49510]= -1917915825;
assign addr[49511]= -2035658475;
assign addr[49512]= -2112148396;
assign addr[49513]= -2145835515;
assign addr[49514]= -2136037160;
assign addr[49515]= -2082951896;
assign addr[49516]= -1987655498;
assign addr[49517]= -1852079154;
assign addr[49518]= -1678970324;
assign addr[49519]= -1471837070;
assign addr[49520]= -1234876957;
assign addr[49521]= -972891995;
assign addr[49522]= -691191324;
assign addr[49523]= -395483624;
assign addr[49524]= -91761426;
assign addr[49525]= 213820322;
assign addr[49526]= 515068990;
assign addr[49527]= 805879757;
assign addr[49528]= 1080359326;
assign addr[49529]= 1332945355;
assign addr[49530]= 1558519173;
assign addr[49531]= 1752509516;
assign addr[49532]= 1910985158;
assign addr[49533]= 2030734582;
assign addr[49534]= 2109331059;
assign addr[49535]= 2145181827;
assign addr[49536]= 2137560369;
assign addr[49537]= 2086621133;
assign addr[49538]= 1993396407;
assign addr[49539]= 1859775393;
assign addr[49540]= 1688465931;
assign addr[49541]= 1482939614;
assign addr[49542]= 1247361445;
assign addr[49543]= 986505429;
assign addr[49544]= 705657826;
assign addr[49545]= 410510029;
assign addr[49546]= 107043224;
assign addr[49547]= -198592817;
assign addr[49548]= -500204365;
assign addr[49549]= -791679244;
assign addr[49550]= -1067110699;
assign addr[49551]= -1320917099;
assign addr[49552]= -1547955041;
assign addr[49553]= -1743623590;
assign addr[49554]= -1903957513;
assign addr[49555]= -2025707632;
assign addr[49556]= -2106406677;
assign addr[49557]= -2144419275;
assign addr[49558]= -2138975100;
assign addr[49559]= -2090184478;
assign addr[49560]= -1999036154;
assign addr[49561]= -1867377253;
assign addr[49562]= -1697875851;
assign addr[49563]= -1493966902;
assign addr[49564]= -1259782632;
assign addr[49565]= -1000068799;
assign addr[49566]= -720088517;
assign addr[49567]= -425515602;
assign addr[49568]= -122319591;
assign addr[49569]= 183355234;
assign addr[49570]= 485314355;
assign addr[49571]= 777438554;
assign addr[49572]= 1053807919;
assign addr[49573]= 1308821808;
assign addr[49574]= 1537312353;
assign addr[49575]= 1734649179;
assign addr[49576]= 1896833245;
assign addr[49577]= 2020577882;
assign addr[49578]= 2103375398;
assign addr[49579]= 2143547897;
assign addr[49580]= 2140281282;
assign addr[49581]= 2093641749;
assign addr[49582]= 2004574453;
assign addr[49583]= 1874884346;
assign addr[49584]= 1707199606;
assign addr[49585]= 1504918373;
assign addr[49586]= 1272139887;
assign addr[49587]= 1013581418;
assign addr[49588]= 734482665;
assign addr[49589]= 440499581;
assign addr[49590]= 137589750;
assign addr[49591]= -168108346;
assign addr[49592]= -470399716;
assign addr[49593]= -763158411;
assign addr[49594]= -1040451659;
assign addr[49595]= -1296660098;
assign addr[49596]= -1526591649;
assign addr[49597]= -1725586737;
assign addr[49598]= -1889612716;
assign addr[49599]= -2015345591;
assign addr[49600]= -2100237377;
assign addr[49601]= -2142567738;
assign addr[49602]= -2141478848;
assign addr[49603]= -2096992772;
assign addr[49604]= -2010011024;
assign addr[49605]= -1882296293;
assign addr[49606]= -1716436725;
assign addr[49607]= -1515793473;
assign addr[49608]= -1284432584;
assign addr[49609]= -1027042599;
assign addr[49610]= -748839539;
assign addr[49611]= -455461206;
assign addr[49612]= -152852926;
assign addr[49613]= 152852926;
assign addr[49614]= 455461206;
assign addr[49615]= 748839539;
assign addr[49616]= 1027042599;
assign addr[49617]= 1284432584;
assign addr[49618]= 1515793473;
assign addr[49619]= 1716436725;
assign addr[49620]= 1882296293;
assign addr[49621]= 2010011024;
assign addr[49622]= 2096992772;
assign addr[49623]= 2141478848;
assign addr[49624]= 2142567738;
assign addr[49625]= 2100237377;
assign addr[49626]= 2015345591;
assign addr[49627]= 1889612716;
assign addr[49628]= 1725586737;
assign addr[49629]= 1526591649;
assign addr[49630]= 1296660098;
assign addr[49631]= 1040451659;
assign addr[49632]= 763158411;
assign addr[49633]= 470399716;
assign addr[49634]= 168108346;
assign addr[49635]= -137589750;
assign addr[49636]= -440499581;
assign addr[49637]= -734482665;
assign addr[49638]= -1013581418;
assign addr[49639]= -1272139887;
assign addr[49640]= -1504918373;
assign addr[49641]= -1707199606;
assign addr[49642]= -1874884346;
assign addr[49643]= -2004574453;
assign addr[49644]= -2093641749;
assign addr[49645]= -2140281282;
assign addr[49646]= -2143547897;
assign addr[49647]= -2103375398;
assign addr[49648]= -2020577882;
assign addr[49649]= -1896833245;
assign addr[49650]= -1734649179;
assign addr[49651]= -1537312353;
assign addr[49652]= -1308821808;
assign addr[49653]= -1053807919;
assign addr[49654]= -777438554;
assign addr[49655]= -485314355;
assign addr[49656]= -183355234;
assign addr[49657]= 122319591;
assign addr[49658]= 425515602;
assign addr[49659]= 720088517;
assign addr[49660]= 1000068799;
assign addr[49661]= 1259782632;
assign addr[49662]= 1493966902;
assign addr[49663]= 1697875851;
assign addr[49664]= 1867377253;
assign addr[49665]= 1999036154;
assign addr[49666]= 2090184478;
assign addr[49667]= 2138975100;
assign addr[49668]= 2144419275;
assign addr[49669]= 2106406677;
assign addr[49670]= 2025707632;
assign addr[49671]= 1903957513;
assign addr[49672]= 1743623590;
assign addr[49673]= 1547955041;
assign addr[49674]= 1320917099;
assign addr[49675]= 1067110699;
assign addr[49676]= 791679244;
assign addr[49677]= 500204365;
assign addr[49678]= 198592817;
assign addr[49679]= -107043224;
assign addr[49680]= -410510029;
assign addr[49681]= -705657826;
assign addr[49682]= -986505429;
assign addr[49683]= -1247361445;
assign addr[49684]= -1482939614;
assign addr[49685]= -1688465931;
assign addr[49686]= -1859775393;
assign addr[49687]= -1993396407;
assign addr[49688]= -2086621133;
assign addr[49689]= -2137560369;
assign addr[49690]= -2145181827;
assign addr[49691]= -2109331059;
assign addr[49692]= -2030734582;
assign addr[49693]= -1910985158;
assign addr[49694]= -1752509516;
assign addr[49695]= -1558519173;
assign addr[49696]= -1332945355;
assign addr[49697]= -1080359326;
assign addr[49698]= -805879757;
assign addr[49699]= -515068990;
assign addr[49700]= -213820322;
assign addr[49701]= 91761426;
assign addr[49702]= 395483624;
assign addr[49703]= 691191324;
assign addr[49704]= 972891995;
assign addr[49705]= 1234876957;
assign addr[49706]= 1471837070;
assign addr[49707]= 1678970324;
assign addr[49708]= 1852079154;
assign addr[49709]= 1987655498;
assign addr[49710]= 2082951896;
assign addr[49711]= 2136037160;
assign addr[49712]= 2145835515;
assign addr[49713]= 2112148396;
assign addr[49714]= 2035658475;
assign addr[49715]= 1917915825;
assign addr[49716]= 1761306505;
assign addr[49717]= 1569004214;
assign addr[49718]= 1344905966;
assign addr[49719]= 1093553126;
assign addr[49720]= 820039373;
assign addr[49721]= 529907477;
assign addr[49722]= 229036977;
assign addr[49723]= -76474970;
assign addr[49724]= -380437148;
assign addr[49725]= -676689746;
assign addr[49726]= -959229189;
assign addr[49727]= -1222329801;
assign addr[49728]= -1460659832;
assign addr[49729]= -1669389513;
assign addr[49730]= -1844288924;
assign addr[49731]= -1981813720;
assign addr[49732]= -2079176953;
assign addr[49733]= -2134405552;
assign addr[49734]= -2146380306;
assign addr[49735]= -2114858546;
assign addr[49736]= -2040479063;
assign addr[49737]= -1924749160;
assign addr[49738]= -1770014111;
assign addr[49739]= -1579409630;
assign addr[49740]= -1356798326;
assign addr[49741]= -1106691431;
assign addr[49742]= -834157373;
assign addr[49743]= -544719071;
assign addr[49744]= -244242007;
assign addr[49745]= 61184634;
assign addr[49746]= 365371365;
assign addr[49747]= 662153826;
assign addr[49748]= 945517704;
assign addr[49749]= 1209720613;
assign addr[49750]= 1449408469;
assign addr[49751]= 1659723983;
assign addr[49752]= 1836405100;
assign addr[49753]= 1975871368;
assign addr[49754]= 2075296495;
assign addr[49755]= 2132665626;
assign addr[49756]= 2146816171;
assign addr[49757]= 2117461370;
assign addr[49758]= 2045196100;
assign addr[49759]= 1931484818;
assign addr[49760]= 1778631892;
assign addr[49761]= 1589734894;
assign addr[49762]= 1368621831;
assign addr[49763]= 1119773573;
assign addr[49764]= 848233042;
assign addr[49765]= 559503022;
assign addr[49766]= 259434643;
assign addr[49767]= -45891193;
assign addr[49768]= -350287041;
assign addr[49769]= -647584304;
assign addr[49770]= -931758235;
assign addr[49771]= -1197050035;
assign addr[49772]= -1438083551;
assign addr[49773]= -1649974225;
assign addr[49774]= -1828428082;
assign addr[49775]= -1969828744;
assign addr[49776]= -2071310720;
assign addr[49777]= -2130817471;
assign addr[49778]= -2147143090;
assign addr[49779]= -2119956737;
assign addr[49780]= -2049809346;
assign addr[49781]= -1938122457;
assign addr[49782]= -1787159411;
assign addr[49783]= -1599979481;
assign addr[49784]= -1380375881;
assign addr[49785]= -1132798888;
assign addr[49786]= -862265664;
assign addr[49787]= -574258580;
assign addr[49788]= -274614114;
assign addr[49789]= 30595422;
assign addr[49790]= 335184940;
assign addr[49791]= 632981917;
assign addr[49792]= 917951481;
assign addr[49793]= 1184318708;
assign addr[49794]= 1426685652;
assign addr[49795]= 1640140734;
assign addr[49796]= 1820358275;
assign addr[49797]= 1963686155;
assign addr[49798]= 2067219829;
assign addr[49799]= 2128861181;
assign addr[49800]= 2147361045;
assign addr[49801]= 2122344521;
assign addr[49802]= 2054318569;
assign addr[49803]= 1944661739;
assign addr[49804]= 1795596234;
assign addr[49805]= 1610142873;
assign addr[49806]= 1392059879;
assign addr[49807]= 1145766716;
assign addr[49808]= 876254528;
assign addr[49809]= 588984994;
assign addr[49810]= 289779648;
assign addr[49811]= -15298099;
assign addr[49812]= -320065829;
assign addr[49813]= -618347408;
assign addr[49814]= -904098143;
assign addr[49815]= -1171527280;
assign addr[49816]= -1415215352;
assign addr[49817]= -1630224009;
assign addr[49818]= -1812196087;
assign addr[49819]= -1957443913;
assign addr[49820]= -2063024031;
assign addr[49821]= -2126796855;
assign addr[49822]= -2147470025;
assign addr[49823]= -2124624598;
assign addr[49824]= -2058723538;
assign addr[49825]= -1951102334;
assign addr[49826]= -1803941934;
assign addr[49827]= -1620224553;
assign addr[49828]= -1403673233;
assign addr[49829]= -1158676398;
assign addr[49830]= -890198924;
assign addr[49831]= -603681519;
assign addr[49832]= -304930476;
assign addr[49833]= 0;
assign addr[49834]= 304930476;
assign addr[49835]= 603681519;
assign addr[49836]= 890198924;
assign addr[49837]= 1158676398;
assign addr[49838]= 1403673233;
assign addr[49839]= 1620224553;
assign addr[49840]= 1803941934;
assign addr[49841]= 1951102334;
assign addr[49842]= 2058723538;
assign addr[49843]= 2124624598;
assign addr[49844]= 2147470025;
assign addr[49845]= 2126796855;
assign addr[49846]= 2063024031;
assign addr[49847]= 1957443913;
assign addr[49848]= 1812196087;
assign addr[49849]= 1630224009;
assign addr[49850]= 1415215352;
assign addr[49851]= 1171527280;
assign addr[49852]= 904098143;
assign addr[49853]= 618347408;
assign addr[49854]= 320065829;
assign addr[49855]= 15298099;
assign addr[49856]= -289779648;
assign addr[49857]= -588984994;
assign addr[49858]= -876254528;
assign addr[49859]= -1145766716;
assign addr[49860]= -1392059879;
assign addr[49861]= -1610142873;
assign addr[49862]= -1795596234;
assign addr[49863]= -1944661739;
assign addr[49864]= -2054318569;
assign addr[49865]= -2122344521;
assign addr[49866]= -2147361045;
assign addr[49867]= -2128861181;
assign addr[49868]= -2067219829;
assign addr[49869]= -1963686155;
assign addr[49870]= -1820358275;
assign addr[49871]= -1640140734;
assign addr[49872]= -1426685652;
assign addr[49873]= -1184318708;
assign addr[49874]= -917951481;
assign addr[49875]= -632981917;
assign addr[49876]= -335184940;
assign addr[49877]= -30595422;
assign addr[49878]= 274614114;
assign addr[49879]= 574258580;
assign addr[49880]= 862265664;
assign addr[49881]= 1132798888;
assign addr[49882]= 1380375881;
assign addr[49883]= 1599979481;
assign addr[49884]= 1787159411;
assign addr[49885]= 1938122457;
assign addr[49886]= 2049809346;
assign addr[49887]= 2119956737;
assign addr[49888]= 2147143090;
assign addr[49889]= 2130817471;
assign addr[49890]= 2071310720;
assign addr[49891]= 1969828744;
assign addr[49892]= 1828428082;
assign addr[49893]= 1649974225;
assign addr[49894]= 1438083551;
assign addr[49895]= 1197050035;
assign addr[49896]= 931758235;
assign addr[49897]= 647584304;
assign addr[49898]= 350287041;
assign addr[49899]= 45891193;
assign addr[49900]= -259434643;
assign addr[49901]= -559503022;
assign addr[49902]= -848233042;
assign addr[49903]= -1119773573;
assign addr[49904]= -1368621831;
assign addr[49905]= -1589734894;
assign addr[49906]= -1778631892;
assign addr[49907]= -1931484818;
assign addr[49908]= -2045196100;
assign addr[49909]= -2117461370;
assign addr[49910]= -2146816171;
assign addr[49911]= -2132665626;
assign addr[49912]= -2075296495;
assign addr[49913]= -1975871368;
assign addr[49914]= -1836405100;
assign addr[49915]= -1659723983;
assign addr[49916]= -1449408469;
assign addr[49917]= -1209720613;
assign addr[49918]= -945517704;
assign addr[49919]= -662153826;
assign addr[49920]= -365371365;
assign addr[49921]= -61184634;
assign addr[49922]= 244242007;
assign addr[49923]= 544719071;
assign addr[49924]= 834157373;
assign addr[49925]= 1106691431;
assign addr[49926]= 1356798326;
assign addr[49927]= 1579409630;
assign addr[49928]= 1770014111;
assign addr[49929]= 1924749160;
assign addr[49930]= 2040479063;
assign addr[49931]= 2114858546;
assign addr[49932]= 2146380306;
assign addr[49933]= 2134405552;
assign addr[49934]= 2079176953;
assign addr[49935]= 1981813720;
assign addr[49936]= 1844288924;
assign addr[49937]= 1669389513;
assign addr[49938]= 1460659832;
assign addr[49939]= 1222329801;
assign addr[49940]= 959229189;
assign addr[49941]= 676689746;
assign addr[49942]= 380437148;
assign addr[49943]= 76474970;
assign addr[49944]= -229036977;
assign addr[49945]= -529907477;
assign addr[49946]= -820039373;
assign addr[49947]= -1093553126;
assign addr[49948]= -1344905966;
assign addr[49949]= -1569004214;
assign addr[49950]= -1761306505;
assign addr[49951]= -1917915825;
assign addr[49952]= -2035658475;
assign addr[49953]= -2112148396;
assign addr[49954]= -2145835515;
assign addr[49955]= -2136037160;
assign addr[49956]= -2082951896;
assign addr[49957]= -1987655498;
assign addr[49958]= -1852079154;
assign addr[49959]= -1678970324;
assign addr[49960]= -1471837070;
assign addr[49961]= -1234876957;
assign addr[49962]= -972891995;
assign addr[49963]= -691191324;
assign addr[49964]= -395483624;
assign addr[49965]= -91761426;
assign addr[49966]= 213820322;
assign addr[49967]= 515068990;
assign addr[49968]= 805879757;
assign addr[49969]= 1080359326;
assign addr[49970]= 1332945355;
assign addr[49971]= 1558519173;
assign addr[49972]= 1752509516;
assign addr[49973]= 1910985158;
assign addr[49974]= 2030734582;
assign addr[49975]= 2109331059;
assign addr[49976]= 2145181827;
assign addr[49977]= 2137560369;
assign addr[49978]= 2086621133;
assign addr[49979]= 1993396407;
assign addr[49980]= 1859775393;
assign addr[49981]= 1688465931;
assign addr[49982]= 1482939614;
assign addr[49983]= 1247361445;
assign addr[49984]= 986505429;
assign addr[49985]= 705657826;
assign addr[49986]= 410510029;
assign addr[49987]= 107043224;
assign addr[49988]= -198592817;
assign addr[49989]= -500204365;
assign addr[49990]= -791679244;
assign addr[49991]= -1067110699;
assign addr[49992]= -1320917099;
assign addr[49993]= -1547955041;
assign addr[49994]= -1743623590;
assign addr[49995]= -1903957513;
assign addr[49996]= -2025707632;
assign addr[49997]= -2106406677;
assign addr[49998]= -2144419275;
assign addr[49999]= -2138975100;
assign addr[50000]= -2090184478;
assign addr[50001]= -1999036154;
assign addr[50002]= -1867377253;
assign addr[50003]= -1697875851;
assign addr[50004]= -1493966902;
assign addr[50005]= -1259782632;
assign addr[50006]= -1000068799;
assign addr[50007]= -720088517;
assign addr[50008]= -425515602;
assign addr[50009]= -122319591;
assign addr[50010]= 183355234;
assign addr[50011]= 485314355;
assign addr[50012]= 777438554;
assign addr[50013]= 1053807919;
assign addr[50014]= 1308821808;
assign addr[50015]= 1537312353;
assign addr[50016]= 1734649179;
assign addr[50017]= 1896833245;
assign addr[50018]= 2020577882;
assign addr[50019]= 2103375398;
assign addr[50020]= 2143547897;
assign addr[50021]= 2140281282;
assign addr[50022]= 2093641749;
assign addr[50023]= 2004574453;
assign addr[50024]= 1874884346;
assign addr[50025]= 1707199606;
assign addr[50026]= 1504918373;
assign addr[50027]= 1272139887;
assign addr[50028]= 1013581418;
assign addr[50029]= 734482665;
assign addr[50030]= 440499581;
assign addr[50031]= 137589750;
assign addr[50032]= -168108346;
assign addr[50033]= -470399716;
assign addr[50034]= -763158411;
assign addr[50035]= -1040451659;
assign addr[50036]= -1296660098;
assign addr[50037]= -1526591649;
assign addr[50038]= -1725586737;
assign addr[50039]= -1889612716;
assign addr[50040]= -2015345591;
assign addr[50041]= -2100237377;
assign addr[50042]= -2142567738;
assign addr[50043]= -2141478848;
assign addr[50044]= -2096992772;
assign addr[50045]= -2010011024;
assign addr[50046]= -1882296293;
assign addr[50047]= -1716436725;
assign addr[50048]= -1515793473;
assign addr[50049]= -1284432584;
assign addr[50050]= -1027042599;
assign addr[50051]= -748839539;
assign addr[50052]= -455461206;
assign addr[50053]= -152852926;
assign addr[50054]= 152852926;
assign addr[50055]= 455461206;
assign addr[50056]= 748839539;
assign addr[50057]= 1027042599;
assign addr[50058]= 1284432584;
assign addr[50059]= 1515793473;
assign addr[50060]= 1716436725;
assign addr[50061]= 1882296293;
assign addr[50062]= 2010011024;
assign addr[50063]= 2096992772;
assign addr[50064]= 2141478848;
assign addr[50065]= 2142567738;
assign addr[50066]= 2100237377;
assign addr[50067]= 2015345591;
assign addr[50068]= 1889612716;
assign addr[50069]= 1725586737;
assign addr[50070]= 1526591649;
assign addr[50071]= 1296660098;
assign addr[50072]= 1040451659;
assign addr[50073]= 763158411;
assign addr[50074]= 470399716;
assign addr[50075]= 168108346;
assign addr[50076]= -137589750;
assign addr[50077]= -440499581;
assign addr[50078]= -734482665;
assign addr[50079]= -1013581418;
assign addr[50080]= -1272139887;
assign addr[50081]= -1504918373;
assign addr[50082]= -1707199606;
assign addr[50083]= -1874884346;
assign addr[50084]= -2004574453;
assign addr[50085]= -2093641749;
assign addr[50086]= -2140281282;
assign addr[50087]= -2143547897;
assign addr[50088]= -2103375398;
assign addr[50089]= -2020577882;
assign addr[50090]= -1896833245;
assign addr[50091]= -1734649179;
assign addr[50092]= -1537312353;
assign addr[50093]= -1308821808;
assign addr[50094]= -1053807919;
assign addr[50095]= -777438554;
assign addr[50096]= -485314355;
assign addr[50097]= -183355234;
assign addr[50098]= 122319591;
assign addr[50099]= 425515602;
assign addr[50100]= 720088517;
assign addr[50101]= 1000068799;
assign addr[50102]= 1259782632;
assign addr[50103]= 1493966902;
assign addr[50104]= 1697875851;
assign addr[50105]= 1867377253;
assign addr[50106]= 1999036154;
assign addr[50107]= 2090184478;
assign addr[50108]= 2138975100;
assign addr[50109]= 2144419275;
assign addr[50110]= 2106406677;
assign addr[50111]= 2025707632;
assign addr[50112]= 1903957513;
assign addr[50113]= 1743623590;
assign addr[50114]= 1547955041;
assign addr[50115]= 1320917099;
assign addr[50116]= 1067110699;
assign addr[50117]= 791679244;
assign addr[50118]= 500204365;
assign addr[50119]= 198592817;
assign addr[50120]= -107043224;
assign addr[50121]= -410510029;
assign addr[50122]= -705657826;
assign addr[50123]= -986505429;
assign addr[50124]= -1247361445;
assign addr[50125]= -1482939614;
assign addr[50126]= -1688465931;
assign addr[50127]= -1859775393;
assign addr[50128]= -1993396407;
assign addr[50129]= -2086621133;
assign addr[50130]= -2137560369;
assign addr[50131]= -2145181827;
assign addr[50132]= -2109331059;
assign addr[50133]= -2030734582;
assign addr[50134]= -1910985158;
assign addr[50135]= -1752509516;
assign addr[50136]= -1558519173;
assign addr[50137]= -1332945355;
assign addr[50138]= -1080359326;
assign addr[50139]= -805879757;
assign addr[50140]= -515068990;
assign addr[50141]= -213820322;
assign addr[50142]= 91761426;
assign addr[50143]= 395483624;
assign addr[50144]= 691191324;
assign addr[50145]= 972891995;
assign addr[50146]= 1234876957;
assign addr[50147]= 1471837070;
assign addr[50148]= 1678970324;
assign addr[50149]= 1852079154;
assign addr[50150]= 1987655498;
assign addr[50151]= 2082951896;
assign addr[50152]= 2136037160;
assign addr[50153]= 2145835515;
assign addr[50154]= 2112148396;
assign addr[50155]= 2035658475;
assign addr[50156]= 1917915825;
assign addr[50157]= 1761306505;
assign addr[50158]= 1569004214;
assign addr[50159]= 1344905966;
assign addr[50160]= 1093553126;
assign addr[50161]= 820039373;
assign addr[50162]= 529907477;
assign addr[50163]= 229036977;
assign addr[50164]= -76474970;
assign addr[50165]= -380437148;
assign addr[50166]= -676689746;
assign addr[50167]= -959229189;
assign addr[50168]= -1222329801;
assign addr[50169]= -1460659832;
assign addr[50170]= -1669389513;
assign addr[50171]= -1844288924;
assign addr[50172]= -1981813720;
assign addr[50173]= -2079176953;
assign addr[50174]= -2134405552;
assign addr[50175]= -2146380306;
assign addr[50176]= -2114858546;
assign addr[50177]= -2040479063;
assign addr[50178]= -1924749160;
assign addr[50179]= -1770014111;
assign addr[50180]= -1579409630;
assign addr[50181]= -1356798326;
assign addr[50182]= -1106691431;
assign addr[50183]= -834157373;
assign addr[50184]= -544719071;
assign addr[50185]= -244242007;
assign addr[50186]= 61184634;
assign addr[50187]= 365371365;
assign addr[50188]= 662153826;
assign addr[50189]= 945517704;
assign addr[50190]= 1209720613;
assign addr[50191]= 1449408469;
assign addr[50192]= 1659723983;
assign addr[50193]= 1836405100;
assign addr[50194]= 1975871368;
assign addr[50195]= 2075296495;
assign addr[50196]= 2132665626;
assign addr[50197]= 2146816171;
assign addr[50198]= 2117461370;
assign addr[50199]= 2045196100;
assign addr[50200]= 1931484818;
assign addr[50201]= 1778631892;
assign addr[50202]= 1589734894;
assign addr[50203]= 1368621831;
assign addr[50204]= 1119773573;
assign addr[50205]= 848233042;
assign addr[50206]= 559503022;
assign addr[50207]= 259434643;
assign addr[50208]= -45891193;
assign addr[50209]= -350287041;
assign addr[50210]= -647584304;
assign addr[50211]= -931758235;
assign addr[50212]= -1197050035;
assign addr[50213]= -1438083551;
assign addr[50214]= -1649974225;
assign addr[50215]= -1828428082;
assign addr[50216]= -1969828744;
assign addr[50217]= -2071310720;
assign addr[50218]= -2130817471;
assign addr[50219]= -2147143090;
assign addr[50220]= -2119956737;
assign addr[50221]= -2049809346;
assign addr[50222]= -1938122457;
assign addr[50223]= -1787159411;
assign addr[50224]= -1599979481;
assign addr[50225]= -1380375881;
assign addr[50226]= -1132798888;
assign addr[50227]= -862265664;
assign addr[50228]= -574258580;
assign addr[50229]= -274614114;
assign addr[50230]= 30595422;
assign addr[50231]= 335184940;
assign addr[50232]= 632981917;
assign addr[50233]= 917951481;
assign addr[50234]= 1184318708;
assign addr[50235]= 1426685652;
assign addr[50236]= 1640140734;
assign addr[50237]= 1820358275;
assign addr[50238]= 1963686155;
assign addr[50239]= 2067219829;
assign addr[50240]= 2128861181;
assign addr[50241]= 2147361045;
assign addr[50242]= 2122344521;
assign addr[50243]= 2054318569;
assign addr[50244]= 1944661739;
assign addr[50245]= 1795596234;
assign addr[50246]= 1610142873;
assign addr[50247]= 1392059879;
assign addr[50248]= 1145766716;
assign addr[50249]= 876254528;
assign addr[50250]= 588984994;
assign addr[50251]= 289779648;
assign addr[50252]= -15298099;
assign addr[50253]= -320065829;
assign addr[50254]= -618347408;
assign addr[50255]= -904098143;
assign addr[50256]= -1171527280;
assign addr[50257]= -1415215352;
assign addr[50258]= -1630224009;
assign addr[50259]= -1812196087;
assign addr[50260]= -1957443913;
assign addr[50261]= -2063024031;
assign addr[50262]= -2126796855;
assign addr[50263]= -2147470025;
assign addr[50264]= -2124624598;
assign addr[50265]= -2058723538;
assign addr[50266]= -1951102334;
assign addr[50267]= -1803941934;
assign addr[50268]= -1620224553;
assign addr[50269]= -1403673233;
assign addr[50270]= -1158676398;
assign addr[50271]= -890198924;
assign addr[50272]= -603681519;
assign addr[50273]= -304930476;
assign addr[50274]= 0;
assign addr[50275]= 304930476;
assign addr[50276]= 603681519;
assign addr[50277]= 890198924;
assign addr[50278]= 1158676398;
assign addr[50279]= 1403673233;
assign addr[50280]= 1620224553;
assign addr[50281]= 1803941934;
assign addr[50282]= 1951102334;
assign addr[50283]= 2058723538;
assign addr[50284]= 2124624598;
assign addr[50285]= 2147470025;
assign addr[50286]= 2126796855;
assign addr[50287]= 2063024031;
assign addr[50288]= 1957443913;
assign addr[50289]= 1812196087;
assign addr[50290]= 1630224009;
assign addr[50291]= 1415215352;
assign addr[50292]= 1171527280;
assign addr[50293]= 904098143;
assign addr[50294]= 618347408;
assign addr[50295]= 320065829;
assign addr[50296]= 15298099;
assign addr[50297]= -289779648;
assign addr[50298]= -588984994;
assign addr[50299]= -876254528;
assign addr[50300]= -1145766716;
assign addr[50301]= -1392059879;
assign addr[50302]= -1610142873;
assign addr[50303]= -1795596234;
assign addr[50304]= -1944661739;
assign addr[50305]= -2054318569;
assign addr[50306]= -2122344521;
assign addr[50307]= -2147361045;
assign addr[50308]= -2128861181;
assign addr[50309]= -2067219829;
assign addr[50310]= -1963686155;
assign addr[50311]= -1820358275;
assign addr[50312]= -1640140734;
assign addr[50313]= -1426685652;
assign addr[50314]= -1184318708;
assign addr[50315]= -917951481;
assign addr[50316]= -632981917;
assign addr[50317]= -335184940;
assign addr[50318]= -30595422;
assign addr[50319]= 274614114;
assign addr[50320]= 574258580;
assign addr[50321]= 862265664;
assign addr[50322]= 1132798888;
assign addr[50323]= 1380375881;
assign addr[50324]= 1599979481;
assign addr[50325]= 1787159411;
assign addr[50326]= 1938122457;
assign addr[50327]= 2049809346;
assign addr[50328]= 2119956737;
assign addr[50329]= 2147143090;
assign addr[50330]= 2130817471;
assign addr[50331]= 2071310720;
assign addr[50332]= 1969828744;
assign addr[50333]= 1828428082;
assign addr[50334]= 1649974225;
assign addr[50335]= 1438083551;
assign addr[50336]= 1197050035;
assign addr[50337]= 931758235;
assign addr[50338]= 647584304;
assign addr[50339]= 350287041;
assign addr[50340]= 45891193;
assign addr[50341]= -259434643;
assign addr[50342]= -559503022;
assign addr[50343]= -848233042;
assign addr[50344]= -1119773573;
assign addr[50345]= -1368621831;
assign addr[50346]= -1589734894;
assign addr[50347]= -1778631892;
assign addr[50348]= -1931484818;
assign addr[50349]= -2045196100;
assign addr[50350]= -2117461370;
assign addr[50351]= -2146816171;
assign addr[50352]= -2132665626;
assign addr[50353]= -2075296495;
assign addr[50354]= -1975871368;
assign addr[50355]= -1836405100;
assign addr[50356]= -1659723983;
assign addr[50357]= -1449408469;
assign addr[50358]= -1209720613;
assign addr[50359]= -945517704;
assign addr[50360]= -662153826;
assign addr[50361]= -365371365;
assign addr[50362]= -61184634;
assign addr[50363]= 244242007;
assign addr[50364]= 544719071;
assign addr[50365]= 834157373;
assign addr[50366]= 1106691431;
assign addr[50367]= 1356798326;
assign addr[50368]= 1579409630;
assign addr[50369]= 1770014111;
assign addr[50370]= 1924749160;
assign addr[50371]= 2040479063;
assign addr[50372]= 2114858546;
assign addr[50373]= 2146380306;
assign addr[50374]= 2134405552;
assign addr[50375]= 2079176953;
assign addr[50376]= 1981813720;
assign addr[50377]= 1844288924;
assign addr[50378]= 1669389513;
assign addr[50379]= 1460659832;
assign addr[50380]= 1222329801;
assign addr[50381]= 959229189;
assign addr[50382]= 676689746;
assign addr[50383]= 380437148;
assign addr[50384]= 76474970;
assign addr[50385]= -229036977;
assign addr[50386]= -529907477;
assign addr[50387]= -820039373;
assign addr[50388]= -1093553126;
assign addr[50389]= -1344905966;
assign addr[50390]= -1569004214;
assign addr[50391]= -1761306505;
assign addr[50392]= -1917915825;
assign addr[50393]= -2035658475;
assign addr[50394]= -2112148396;
assign addr[50395]= -2145835515;
assign addr[50396]= -2136037160;
assign addr[50397]= -2082951896;
assign addr[50398]= -1987655498;
assign addr[50399]= -1852079154;
assign addr[50400]= -1678970324;
assign addr[50401]= -1471837070;
assign addr[50402]= -1234876957;
assign addr[50403]= -972891995;
assign addr[50404]= -691191324;
assign addr[50405]= -395483624;
assign addr[50406]= -91761426;
assign addr[50407]= 213820322;
assign addr[50408]= 515068990;
assign addr[50409]= 805879757;
assign addr[50410]= 1080359326;
assign addr[50411]= 1332945355;
assign addr[50412]= 1558519173;
assign addr[50413]= 1752509516;
assign addr[50414]= 1910985158;
assign addr[50415]= 2030734582;
assign addr[50416]= 2109331059;
assign addr[50417]= 2145181827;
assign addr[50418]= 2137560369;
assign addr[50419]= 2086621133;
assign addr[50420]= 1993396407;
assign addr[50421]= 1859775393;
assign addr[50422]= 1688465931;
assign addr[50423]= 1482939614;
assign addr[50424]= 1247361445;
assign addr[50425]= 986505429;
assign addr[50426]= 705657826;
assign addr[50427]= 410510029;
assign addr[50428]= 107043224;
assign addr[50429]= -198592817;
assign addr[50430]= -500204365;
assign addr[50431]= -791679244;
assign addr[50432]= -1067110699;
assign addr[50433]= -1320917099;
assign addr[50434]= -1547955041;
assign addr[50435]= -1743623590;
assign addr[50436]= -1903957513;
assign addr[50437]= -2025707632;
assign addr[50438]= -2106406677;
assign addr[50439]= -2144419275;
assign addr[50440]= -2138975100;
assign addr[50441]= -2090184478;
assign addr[50442]= -1999036154;
assign addr[50443]= -1867377253;
assign addr[50444]= -1697875851;
assign addr[50445]= -1493966902;
assign addr[50446]= -1259782632;
assign addr[50447]= -1000068799;
assign addr[50448]= -720088517;
assign addr[50449]= -425515602;
assign addr[50450]= -122319591;
assign addr[50451]= 183355234;
assign addr[50452]= 485314355;
assign addr[50453]= 777438554;
assign addr[50454]= 1053807919;
assign addr[50455]= 1308821808;
assign addr[50456]= 1537312353;
assign addr[50457]= 1734649179;
assign addr[50458]= 1896833245;
assign addr[50459]= 2020577882;
assign addr[50460]= 2103375398;
assign addr[50461]= 2143547897;
assign addr[50462]= 2140281282;
assign addr[50463]= 2093641749;
assign addr[50464]= 2004574453;
assign addr[50465]= 1874884346;
assign addr[50466]= 1707199606;
assign addr[50467]= 1504918373;
assign addr[50468]= 1272139887;
assign addr[50469]= 1013581418;
assign addr[50470]= 734482665;
assign addr[50471]= 440499581;
assign addr[50472]= 137589750;
assign addr[50473]= -168108346;
assign addr[50474]= -470399716;
assign addr[50475]= -763158411;
assign addr[50476]= -1040451659;
assign addr[50477]= -1296660098;
assign addr[50478]= -1526591649;
assign addr[50479]= -1725586737;
assign addr[50480]= -1889612716;
assign addr[50481]= -2015345591;
assign addr[50482]= -2100237377;
assign addr[50483]= -2142567738;
assign addr[50484]= -2141478848;
assign addr[50485]= -2096992772;
assign addr[50486]= -2010011024;
assign addr[50487]= -1882296293;
assign addr[50488]= -1716436725;
assign addr[50489]= -1515793473;
assign addr[50490]= -1284432584;
assign addr[50491]= -1027042599;
assign addr[50492]= -748839539;
assign addr[50493]= -455461206;
assign addr[50494]= -152852926;
assign addr[50495]= 152852926;
assign addr[50496]= 455461206;
assign addr[50497]= 748839539;
assign addr[50498]= 1027042599;
assign addr[50499]= 1284432584;
assign addr[50500]= 1515793473;
assign addr[50501]= 1716436725;
assign addr[50502]= 1882296293;
assign addr[50503]= 2010011024;
assign addr[50504]= 2096992772;
assign addr[50505]= 2141478848;
assign addr[50506]= 2142567738;
assign addr[50507]= 2100237377;
assign addr[50508]= 2015345591;
assign addr[50509]= 1889612716;
assign addr[50510]= 1725586737;
assign addr[50511]= 1526591649;
assign addr[50512]= 1296660098;
assign addr[50513]= 1040451659;
assign addr[50514]= 763158411;
assign addr[50515]= 470399716;
assign addr[50516]= 168108346;
assign addr[50517]= -137589750;
assign addr[50518]= -440499581;
assign addr[50519]= -734482665;
assign addr[50520]= -1013581418;
assign addr[50521]= -1272139887;
assign addr[50522]= -1504918373;
assign addr[50523]= -1707199606;
assign addr[50524]= -1874884346;
assign addr[50525]= -2004574453;
assign addr[50526]= -2093641749;
assign addr[50527]= -2140281282;
assign addr[50528]= -2143547897;
assign addr[50529]= -2103375398;
assign addr[50530]= -2020577882;
assign addr[50531]= -1896833245;
assign addr[50532]= -1734649179;
assign addr[50533]= -1537312353;
assign addr[50534]= -1308821808;
assign addr[50535]= -1053807919;
assign addr[50536]= -777438554;
assign addr[50537]= -485314355;
assign addr[50538]= -183355234;
assign addr[50539]= 122319591;
assign addr[50540]= 425515602;
assign addr[50541]= 720088517;
assign addr[50542]= 1000068799;
assign addr[50543]= 1259782632;
assign addr[50544]= 1493966902;
assign addr[50545]= 1697875851;
assign addr[50546]= 1867377253;
assign addr[50547]= 1999036154;
assign addr[50548]= 2090184478;
assign addr[50549]= 2138975100;
assign addr[50550]= 2144419275;
assign addr[50551]= 2106406677;
assign addr[50552]= 2025707632;
assign addr[50553]= 1903957513;
assign addr[50554]= 1743623590;
assign addr[50555]= 1547955041;
assign addr[50556]= 1320917099;
assign addr[50557]= 1067110699;
assign addr[50558]= 791679244;
assign addr[50559]= 500204365;
assign addr[50560]= 198592817;
assign addr[50561]= -107043224;
assign addr[50562]= -410510029;
assign addr[50563]= -705657826;
assign addr[50564]= -986505429;
assign addr[50565]= -1247361445;
assign addr[50566]= -1482939614;
assign addr[50567]= -1688465931;
assign addr[50568]= -1859775393;
assign addr[50569]= -1993396407;
assign addr[50570]= -2086621133;
assign addr[50571]= -2137560369;
assign addr[50572]= -2145181827;
assign addr[50573]= -2109331059;
assign addr[50574]= -2030734582;
assign addr[50575]= -1910985158;
assign addr[50576]= -1752509516;
assign addr[50577]= -1558519173;
assign addr[50578]= -1332945355;
assign addr[50579]= -1080359326;
assign addr[50580]= -805879757;
assign addr[50581]= -515068990;
assign addr[50582]= -213820322;
assign addr[50583]= 91761426;
assign addr[50584]= 395483624;
assign addr[50585]= 691191324;
assign addr[50586]= 972891995;
assign addr[50587]= 1234876957;
assign addr[50588]= 1471837070;
assign addr[50589]= 1678970324;
assign addr[50590]= 1852079154;
assign addr[50591]= 1987655498;
assign addr[50592]= 2082951896;
assign addr[50593]= 2136037160;
assign addr[50594]= 2145835515;
assign addr[50595]= 2112148396;
assign addr[50596]= 2035658475;
assign addr[50597]= 1917915825;
assign addr[50598]= 1761306505;
assign addr[50599]= 1569004214;
assign addr[50600]= 1344905966;
assign addr[50601]= 1093553126;
assign addr[50602]= 820039373;
assign addr[50603]= 529907477;
assign addr[50604]= 229036977;
assign addr[50605]= -76474970;
assign addr[50606]= -380437148;
assign addr[50607]= -676689746;
assign addr[50608]= -959229189;
assign addr[50609]= -1222329801;
assign addr[50610]= -1460659832;
assign addr[50611]= -1669389513;
assign addr[50612]= -1844288924;
assign addr[50613]= -1981813720;
assign addr[50614]= -2079176953;
assign addr[50615]= -2134405552;
assign addr[50616]= -2146380306;
assign addr[50617]= -2114858546;
assign addr[50618]= -2040479063;
assign addr[50619]= -1924749160;
assign addr[50620]= -1770014111;
assign addr[50621]= -1579409630;
assign addr[50622]= -1356798326;
assign addr[50623]= -1106691431;
assign addr[50624]= -834157373;
assign addr[50625]= -544719071;
assign addr[50626]= -244242007;
assign addr[50627]= 61184634;
assign addr[50628]= 365371365;
assign addr[50629]= 662153826;
assign addr[50630]= 945517704;
assign addr[50631]= 1209720613;
assign addr[50632]= 1449408469;
assign addr[50633]= 1659723983;
assign addr[50634]= 1836405100;
assign addr[50635]= 1975871368;
assign addr[50636]= 2075296495;
assign addr[50637]= 2132665626;
assign addr[50638]= 2146816171;
assign addr[50639]= 2117461370;
assign addr[50640]= 2045196100;
assign addr[50641]= 1931484818;
assign addr[50642]= 1778631892;
assign addr[50643]= 1589734894;
assign addr[50644]= 1368621831;
assign addr[50645]= 1119773573;
assign addr[50646]= 848233042;
assign addr[50647]= 559503022;
assign addr[50648]= 259434643;
assign addr[50649]= -45891193;
assign addr[50650]= -350287041;
assign addr[50651]= -647584304;
assign addr[50652]= -931758235;
assign addr[50653]= -1197050035;
assign addr[50654]= -1438083551;
assign addr[50655]= -1649974225;
assign addr[50656]= -1828428082;
assign addr[50657]= -1969828744;
assign addr[50658]= -2071310720;
assign addr[50659]= -2130817471;
assign addr[50660]= -2147143090;
assign addr[50661]= -2119956737;
assign addr[50662]= -2049809346;
assign addr[50663]= -1938122457;
assign addr[50664]= -1787159411;
assign addr[50665]= -1599979481;
assign addr[50666]= -1380375881;
assign addr[50667]= -1132798888;
assign addr[50668]= -862265664;
assign addr[50669]= -574258580;
assign addr[50670]= -274614114;
assign addr[50671]= 30595422;
assign addr[50672]= 335184940;
assign addr[50673]= 632981917;
assign addr[50674]= 917951481;
assign addr[50675]= 1184318708;
assign addr[50676]= 1426685652;
assign addr[50677]= 1640140734;
assign addr[50678]= 1820358275;
assign addr[50679]= 1963686155;
assign addr[50680]= 2067219829;
assign addr[50681]= 2128861181;
assign addr[50682]= 2147361045;
assign addr[50683]= 2122344521;
assign addr[50684]= 2054318569;
assign addr[50685]= 1944661739;
assign addr[50686]= 1795596234;
assign addr[50687]= 1610142873;
assign addr[50688]= 1392059879;
assign addr[50689]= 1145766716;
assign addr[50690]= 876254528;
assign addr[50691]= 588984994;
assign addr[50692]= 289779648;
assign addr[50693]= -15298099;
assign addr[50694]= -320065829;
assign addr[50695]= -618347408;
assign addr[50696]= -904098143;
assign addr[50697]= -1171527280;
assign addr[50698]= -1415215352;
assign addr[50699]= -1630224009;
assign addr[50700]= -1812196087;
assign addr[50701]= -1957443913;
assign addr[50702]= -2063024031;
assign addr[50703]= -2126796855;
assign addr[50704]= -2147470025;
assign addr[50705]= -2124624598;
assign addr[50706]= -2058723538;
assign addr[50707]= -1951102334;
assign addr[50708]= -1803941934;
assign addr[50709]= -1620224553;
assign addr[50710]= -1403673233;
assign addr[50711]= -1158676398;
assign addr[50712]= -890198924;
assign addr[50713]= -603681519;
assign addr[50714]= -304930476;
assign addr[50715]= 0;
assign addr[50716]= 304930476;
assign addr[50717]= 603681519;
assign addr[50718]= 890198924;
assign addr[50719]= 1158676398;
assign addr[50720]= 1403673233;
assign addr[50721]= 1620224553;
assign addr[50722]= 1803941934;
assign addr[50723]= 1951102334;
assign addr[50724]= 2058723538;
assign addr[50725]= 2124624598;
assign addr[50726]= 2147470025;
assign addr[50727]= 2126796855;
assign addr[50728]= 2063024031;
assign addr[50729]= 1957443913;
assign addr[50730]= 1812196087;
assign addr[50731]= 1630224009;
assign addr[50732]= 1415215352;
assign addr[50733]= 1171527280;
assign addr[50734]= 904098143;
assign addr[50735]= 618347408;
assign addr[50736]= 320065829;
assign addr[50737]= 15298099;
assign addr[50738]= -289779648;
assign addr[50739]= -588984994;
assign addr[50740]= -876254528;
assign addr[50741]= -1145766716;
assign addr[50742]= -1392059879;
assign addr[50743]= -1610142873;
assign addr[50744]= -1795596234;
assign addr[50745]= -1944661739;
assign addr[50746]= -2054318569;
assign addr[50747]= -2122344521;
assign addr[50748]= -2147361045;
assign addr[50749]= -2128861181;
assign addr[50750]= -2067219829;
assign addr[50751]= -1963686155;
assign addr[50752]= -1820358275;
assign addr[50753]= -1640140734;
assign addr[50754]= -1426685652;
assign addr[50755]= -1184318708;
assign addr[50756]= -917951481;
assign addr[50757]= -632981917;
assign addr[50758]= -335184940;
assign addr[50759]= -30595422;
assign addr[50760]= 274614114;
assign addr[50761]= 574258580;
assign addr[50762]= 862265664;
assign addr[50763]= 1132798888;
assign addr[50764]= 1380375881;
assign addr[50765]= 1599979481;
assign addr[50766]= 1787159411;
assign addr[50767]= 1938122457;
assign addr[50768]= 2049809346;
assign addr[50769]= 2119956737;
assign addr[50770]= 2147143090;
assign addr[50771]= 2130817471;
assign addr[50772]= 2071310720;
assign addr[50773]= 1969828744;
assign addr[50774]= 1828428082;
assign addr[50775]= 1649974225;
assign addr[50776]= 1438083551;
assign addr[50777]= 1197050035;
assign addr[50778]= 931758235;
assign addr[50779]= 647584304;
assign addr[50780]= 350287041;
assign addr[50781]= 45891193;
assign addr[50782]= -259434643;
assign addr[50783]= -559503022;
assign addr[50784]= -848233042;
assign addr[50785]= -1119773573;
assign addr[50786]= -1368621831;
assign addr[50787]= -1589734894;
assign addr[50788]= -1778631892;
assign addr[50789]= -1931484818;
assign addr[50790]= -2045196100;
assign addr[50791]= -2117461370;
assign addr[50792]= -2146816171;
assign addr[50793]= -2132665626;
assign addr[50794]= -2075296495;
assign addr[50795]= -1975871368;
assign addr[50796]= -1836405100;
assign addr[50797]= -1659723983;
assign addr[50798]= -1449408469;
assign addr[50799]= -1209720613;
assign addr[50800]= -945517704;
assign addr[50801]= -662153826;
assign addr[50802]= -365371365;
assign addr[50803]= -61184634;
assign addr[50804]= 244242007;
assign addr[50805]= 544719071;
assign addr[50806]= 834157373;
assign addr[50807]= 1106691431;
assign addr[50808]= 1356798326;
assign addr[50809]= 1579409630;
assign addr[50810]= 1770014111;
assign addr[50811]= 1924749160;
assign addr[50812]= 2040479063;
assign addr[50813]= 2114858546;
assign addr[50814]= 2146380306;
assign addr[50815]= 2134405552;
assign addr[50816]= 2079176953;
assign addr[50817]= 1981813720;
assign addr[50818]= 1844288924;
assign addr[50819]= 1669389513;
assign addr[50820]= 1460659832;
assign addr[50821]= 1222329801;
assign addr[50822]= 959229189;
assign addr[50823]= 676689746;
assign addr[50824]= 380437148;
assign addr[50825]= 76474970;
assign addr[50826]= -229036977;
assign addr[50827]= -529907477;
assign addr[50828]= -820039373;
assign addr[50829]= -1093553126;
assign addr[50830]= -1344905966;
assign addr[50831]= -1569004214;
assign addr[50832]= -1761306505;
assign addr[50833]= -1917915825;
assign addr[50834]= -2035658475;
assign addr[50835]= -2112148396;
assign addr[50836]= -2145835515;
assign addr[50837]= -2136037160;
assign addr[50838]= -2082951896;
assign addr[50839]= -1987655498;
assign addr[50840]= -1852079154;
assign addr[50841]= -1678970324;
assign addr[50842]= -1471837070;
assign addr[50843]= -1234876957;
assign addr[50844]= -972891995;
assign addr[50845]= -691191324;
assign addr[50846]= -395483624;
assign addr[50847]= -91761426;
assign addr[50848]= 213820322;
assign addr[50849]= 515068990;
assign addr[50850]= 805879757;
assign addr[50851]= 1080359326;
assign addr[50852]= 1332945355;
assign addr[50853]= 1558519173;
assign addr[50854]= 1752509516;
assign addr[50855]= 1910985158;
assign addr[50856]= 2030734582;
assign addr[50857]= 2109331059;
assign addr[50858]= 2145181827;
assign addr[50859]= 2137560369;
assign addr[50860]= 2086621133;
assign addr[50861]= 1993396407;
assign addr[50862]= 1859775393;
assign addr[50863]= 1688465931;
assign addr[50864]= 1482939614;
assign addr[50865]= 1247361445;
assign addr[50866]= 986505429;
assign addr[50867]= 705657826;
assign addr[50868]= 410510029;
assign addr[50869]= 107043224;
assign addr[50870]= -198592817;
assign addr[50871]= -500204365;
assign addr[50872]= -791679244;
assign addr[50873]= -1067110699;
assign addr[50874]= -1320917099;
assign addr[50875]= -1547955041;
assign addr[50876]= -1743623590;
assign addr[50877]= -1903957513;
assign addr[50878]= -2025707632;
assign addr[50879]= -2106406677;
assign addr[50880]= -2144419275;
assign addr[50881]= -2138975100;
assign addr[50882]= -2090184478;
assign addr[50883]= -1999036154;
assign addr[50884]= -1867377253;
assign addr[50885]= -1697875851;
assign addr[50886]= -1493966902;
assign addr[50887]= -1259782632;
assign addr[50888]= -1000068799;
assign addr[50889]= -720088517;
assign addr[50890]= -425515602;
assign addr[50891]= -122319591;
assign addr[50892]= 183355234;
assign addr[50893]= 485314355;
assign addr[50894]= 777438554;
assign addr[50895]= 1053807919;
assign addr[50896]= 1308821808;
assign addr[50897]= 1537312353;
assign addr[50898]= 1734649179;
assign addr[50899]= 1896833245;
assign addr[50900]= 2020577882;
assign addr[50901]= 2103375398;
assign addr[50902]= 2143547897;
assign addr[50903]= 2140281282;
assign addr[50904]= 2093641749;
assign addr[50905]= 2004574453;
assign addr[50906]= 1874884346;
assign addr[50907]= 1707199606;
assign addr[50908]= 1504918373;
assign addr[50909]= 1272139887;
assign addr[50910]= 1013581418;
assign addr[50911]= 734482665;
assign addr[50912]= 440499581;
assign addr[50913]= 137589750;
assign addr[50914]= -168108346;
assign addr[50915]= -470399716;
assign addr[50916]= -763158411;
assign addr[50917]= -1040451659;
assign addr[50918]= -1296660098;
assign addr[50919]= -1526591649;
assign addr[50920]= -1725586737;
assign addr[50921]= -1889612716;
assign addr[50922]= -2015345591;
assign addr[50923]= -2100237377;
assign addr[50924]= -2142567738;
assign addr[50925]= -2141478848;
assign addr[50926]= -2096992772;
assign addr[50927]= -2010011024;
assign addr[50928]= -1882296293;
assign addr[50929]= -1716436725;
assign addr[50930]= -1515793473;
assign addr[50931]= -1284432584;
assign addr[50932]= -1027042599;
assign addr[50933]= -748839539;
assign addr[50934]= -455461206;
assign addr[50935]= -152852926;
assign addr[50936]= 152852926;
assign addr[50937]= 455461206;
assign addr[50938]= 748839539;
assign addr[50939]= 1027042599;
assign addr[50940]= 1284432584;
assign addr[50941]= 1515793473;
assign addr[50942]= 1716436725;
assign addr[50943]= 1882296293;
assign addr[50944]= 2010011024;
assign addr[50945]= 2096992772;
assign addr[50946]= 2141478848;
assign addr[50947]= 2142567738;
assign addr[50948]= 2100237377;
assign addr[50949]= 2015345591;
assign addr[50950]= 1889612716;
assign addr[50951]= 1725586737;
assign addr[50952]= 1526591649;
assign addr[50953]= 1296660098;
assign addr[50954]= 1040451659;
assign addr[50955]= 763158411;
assign addr[50956]= 470399716;
assign addr[50957]= 168108346;
assign addr[50958]= -137589750;
assign addr[50959]= -440499581;
assign addr[50960]= -734482665;
assign addr[50961]= -1013581418;
assign addr[50962]= -1272139887;
assign addr[50963]= -1504918373;
assign addr[50964]= -1707199606;
assign addr[50965]= -1874884346;
assign addr[50966]= -2004574453;
assign addr[50967]= -2093641749;
assign addr[50968]= -2140281282;
assign addr[50969]= -2143547897;
assign addr[50970]= -2103375398;
assign addr[50971]= -2020577882;
assign addr[50972]= -1896833245;
assign addr[50973]= -1734649179;
assign addr[50974]= -1537312353;
assign addr[50975]= -1308821808;
assign addr[50976]= -1053807919;
assign addr[50977]= -777438554;
assign addr[50978]= -485314355;
assign addr[50979]= -183355234;
assign addr[50980]= 122319591;
assign addr[50981]= 425515602;
assign addr[50982]= 720088517;
assign addr[50983]= 1000068799;
assign addr[50984]= 1259782632;
assign addr[50985]= 1493966902;
assign addr[50986]= 1697875851;
assign addr[50987]= 1867377253;
assign addr[50988]= 1999036154;
assign addr[50989]= 2090184478;
assign addr[50990]= 2138975100;
assign addr[50991]= 2144419275;
assign addr[50992]= 2106406677;
assign addr[50993]= 2025707632;
assign addr[50994]= 1903957513;
assign addr[50995]= 1743623590;
assign addr[50996]= 1547955041;
assign addr[50997]= 1320917099;
assign addr[50998]= 1067110699;
assign addr[50999]= 791679244;
assign addr[51000]= 500204365;
assign addr[51001]= 198592817;
assign addr[51002]= -107043224;
assign addr[51003]= -410510029;
assign addr[51004]= -705657826;
assign addr[51005]= -986505429;
assign addr[51006]= -1247361445;
assign addr[51007]= -1482939614;
assign addr[51008]= -1688465931;
assign addr[51009]= -1859775393;
assign addr[51010]= -1993396407;
assign addr[51011]= -2086621133;
assign addr[51012]= -2137560369;
assign addr[51013]= -2145181827;
assign addr[51014]= -2109331059;
assign addr[51015]= -2030734582;
assign addr[51016]= -1910985158;
assign addr[51017]= -1752509516;
assign addr[51018]= -1558519173;
assign addr[51019]= -1332945355;
assign addr[51020]= -1080359326;
assign addr[51021]= -805879757;
assign addr[51022]= -515068990;
assign addr[51023]= -213820322;
assign addr[51024]= 91761426;
assign addr[51025]= 395483624;
assign addr[51026]= 691191324;
assign addr[51027]= 972891995;
assign addr[51028]= 1234876957;
assign addr[51029]= 1471837070;
assign addr[51030]= 1678970324;
assign addr[51031]= 1852079154;
assign addr[51032]= 1987655498;
assign addr[51033]= 2082951896;
assign addr[51034]= 2136037160;
assign addr[51035]= 2145835515;
assign addr[51036]= 2112148396;
assign addr[51037]= 2035658475;
assign addr[51038]= 1917915825;
assign addr[51039]= 1761306505;
assign addr[51040]= 1569004214;
assign addr[51041]= 1344905966;
assign addr[51042]= 1093553126;
assign addr[51043]= 820039373;
assign addr[51044]= 529907477;
assign addr[51045]= 229036977;
assign addr[51046]= -76474970;
assign addr[51047]= -380437148;
assign addr[51048]= -676689746;
assign addr[51049]= -959229189;
assign addr[51050]= -1222329801;
assign addr[51051]= -1460659832;
assign addr[51052]= -1669389513;
assign addr[51053]= -1844288924;
assign addr[51054]= -1981813720;
assign addr[51055]= -2079176953;
assign addr[51056]= -2134405552;
assign addr[51057]= -2146380306;
assign addr[51058]= -2114858546;
assign addr[51059]= -2040479063;
assign addr[51060]= -1924749160;
assign addr[51061]= -1770014111;
assign addr[51062]= -1579409630;
assign addr[51063]= -1356798326;
assign addr[51064]= -1106691431;
assign addr[51065]= -834157373;
assign addr[51066]= -544719071;
assign addr[51067]= -244242007;
assign addr[51068]= 61184634;
assign addr[51069]= 365371365;
assign addr[51070]= 662153826;
assign addr[51071]= 945517704;
assign addr[51072]= 1209720613;
assign addr[51073]= 1449408469;
assign addr[51074]= 1659723983;
assign addr[51075]= 1836405100;
assign addr[51076]= 1975871368;
assign addr[51077]= 2075296495;
assign addr[51078]= 2132665626;
assign addr[51079]= 2146816171;
assign addr[51080]= 2117461370;
assign addr[51081]= 2045196100;
assign addr[51082]= 1931484818;
assign addr[51083]= 1778631892;
assign addr[51084]= 1589734894;
assign addr[51085]= 1368621831;
assign addr[51086]= 1119773573;
assign addr[51087]= 848233042;
assign addr[51088]= 559503022;
assign addr[51089]= 259434643;
assign addr[51090]= -45891193;
assign addr[51091]= -350287041;
assign addr[51092]= -647584304;
assign addr[51093]= -931758235;
assign addr[51094]= -1197050035;
assign addr[51095]= -1438083551;
assign addr[51096]= -1649974225;
assign addr[51097]= -1828428082;
assign addr[51098]= -1969828744;
assign addr[51099]= -2071310720;
assign addr[51100]= -2130817471;
assign addr[51101]= -2147143090;
assign addr[51102]= -2119956737;
assign addr[51103]= -2049809346;
assign addr[51104]= -1938122457;
assign addr[51105]= -1787159411;
assign addr[51106]= -1599979481;
assign addr[51107]= -1380375881;
assign addr[51108]= -1132798888;
assign addr[51109]= -862265664;
assign addr[51110]= -574258580;
assign addr[51111]= -274614114;
assign addr[51112]= 30595422;
assign addr[51113]= 335184940;
assign addr[51114]= 632981917;
assign addr[51115]= 917951481;
assign addr[51116]= 1184318708;
assign addr[51117]= 1426685652;
assign addr[51118]= 1640140734;
assign addr[51119]= 1820358275;
assign addr[51120]= 1963686155;
assign addr[51121]= 2067219829;
assign addr[51122]= 2128861181;
assign addr[51123]= 2147361045;
assign addr[51124]= 2122344521;
assign addr[51125]= 2054318569;
assign addr[51126]= 1944661739;
assign addr[51127]= 1795596234;
assign addr[51128]= 1610142873;
assign addr[51129]= 1392059879;
assign addr[51130]= 1145766716;
assign addr[51131]= 876254528;
assign addr[51132]= 588984994;
assign addr[51133]= 289779648;
assign addr[51134]= -15298099;
assign addr[51135]= -320065829;
assign addr[51136]= -618347408;
assign addr[51137]= -904098143;
assign addr[51138]= -1171527280;
assign addr[51139]= -1415215352;
assign addr[51140]= -1630224009;
assign addr[51141]= -1812196087;
assign addr[51142]= -1957443913;
assign addr[51143]= -2063024031;
assign addr[51144]= -2126796855;
assign addr[51145]= -2147470025;
assign addr[51146]= -2124624598;
assign addr[51147]= -2058723538;
assign addr[51148]= -1951102334;
assign addr[51149]= -1803941934;
assign addr[51150]= -1620224553;
assign addr[51151]= -1403673233;
assign addr[51152]= -1158676398;
assign addr[51153]= -890198924;
assign addr[51154]= -603681519;
assign addr[51155]= -304930476;
assign addr[51156]= 0;
assign addr[51157]= 304930476;
assign addr[51158]= 603681519;
assign addr[51159]= 890198924;
assign addr[51160]= 1158676398;
assign addr[51161]= 1403673233;
assign addr[51162]= 1620224553;
assign addr[51163]= 1803941934;
assign addr[51164]= 1951102334;
assign addr[51165]= 2058723538;
assign addr[51166]= 2124624598;
assign addr[51167]= 2147470025;
assign addr[51168]= 2126796855;
assign addr[51169]= 2063024031;
assign addr[51170]= 1957443913;
assign addr[51171]= 1812196087;
assign addr[51172]= 1630224009;
assign addr[51173]= 1415215352;
assign addr[51174]= 1171527280;
assign addr[51175]= 904098143;
assign addr[51176]= 618347408;
assign addr[51177]= 320065829;
assign addr[51178]= 15298099;
assign addr[51179]= -289779648;
assign addr[51180]= -588984994;
assign addr[51181]= -876254528;
assign addr[51182]= -1145766716;
assign addr[51183]= -1392059879;
assign addr[51184]= -1610142873;
assign addr[51185]= -1795596234;
assign addr[51186]= -1944661739;
assign addr[51187]= -2054318569;
assign addr[51188]= -2122344521;
assign addr[51189]= -2147361045;
assign addr[51190]= -2128861181;
assign addr[51191]= -2067219829;
assign addr[51192]= -1963686155;
assign addr[51193]= -1820358275;
assign addr[51194]= -1640140734;
assign addr[51195]= -1426685652;
assign addr[51196]= -1184318708;
assign addr[51197]= -917951481;
assign addr[51198]= -632981917;
assign addr[51199]= -335184940;
assign addr[51200]= -30595422;
assign addr[51201]= 274614114;
assign addr[51202]= 574258580;
assign addr[51203]= 862265664;
assign addr[51204]= 1132798888;
assign addr[51205]= 1380375881;
assign addr[51206]= 1599979481;
assign addr[51207]= 1787159411;
assign addr[51208]= 1938122457;
assign addr[51209]= 2049809346;
assign addr[51210]= 2119956737;
assign addr[51211]= 2147143090;
assign addr[51212]= 2130817471;
assign addr[51213]= 2071310720;
assign addr[51214]= 1969828744;
assign addr[51215]= 1828428082;
assign addr[51216]= 1649974225;
assign addr[51217]= 1438083551;
assign addr[51218]= 1197050035;
assign addr[51219]= 931758235;
assign addr[51220]= 647584304;
assign addr[51221]= 350287041;
assign addr[51222]= 45891193;
assign addr[51223]= -259434643;
assign addr[51224]= -559503022;
assign addr[51225]= -848233042;
assign addr[51226]= -1119773573;
assign addr[51227]= -1368621831;
assign addr[51228]= -1589734894;
assign addr[51229]= -1778631892;
assign addr[51230]= -1931484818;
assign addr[51231]= -2045196100;
assign addr[51232]= -2117461370;
assign addr[51233]= -2146816171;
assign addr[51234]= -2132665626;
assign addr[51235]= -2075296495;
assign addr[51236]= -1975871368;
assign addr[51237]= -1836405100;
assign addr[51238]= -1659723983;
assign addr[51239]= -1449408469;
assign addr[51240]= -1209720613;
assign addr[51241]= -945517704;
assign addr[51242]= -662153826;
assign addr[51243]= -365371365;
assign addr[51244]= -61184634;
assign addr[51245]= 244242007;
assign addr[51246]= 544719071;
assign addr[51247]= 834157373;
assign addr[51248]= 1106691431;
assign addr[51249]= 1356798326;
assign addr[51250]= 1579409630;
assign addr[51251]= 1770014111;
assign addr[51252]= 1924749160;
assign addr[51253]= 2040479063;
assign addr[51254]= 2114858546;
assign addr[51255]= 2146380306;
assign addr[51256]= 2134405552;
assign addr[51257]= 2079176953;
assign addr[51258]= 1981813720;
assign addr[51259]= 1844288924;
assign addr[51260]= 1669389513;
assign addr[51261]= 1460659832;
assign addr[51262]= 1222329801;
assign addr[51263]= 959229189;
assign addr[51264]= 676689746;
assign addr[51265]= 380437148;
assign addr[51266]= 76474970;
assign addr[51267]= -229036977;
assign addr[51268]= -529907477;
assign addr[51269]= -820039373;
assign addr[51270]= -1093553126;
assign addr[51271]= -1344905966;
assign addr[51272]= -1569004214;
assign addr[51273]= -1761306505;
assign addr[51274]= -1917915825;
assign addr[51275]= -2035658475;
assign addr[51276]= -2112148396;
assign addr[51277]= -2145835515;
assign addr[51278]= -2136037160;
assign addr[51279]= -2082951896;
assign addr[51280]= -1987655498;
assign addr[51281]= -1852079154;
assign addr[51282]= -1678970324;
assign addr[51283]= -1471837070;
assign addr[51284]= -1234876957;
assign addr[51285]= -972891995;
assign addr[51286]= -691191324;
assign addr[51287]= -395483624;
assign addr[51288]= -91761426;
assign addr[51289]= 213820322;
assign addr[51290]= 515068990;
assign addr[51291]= 805879757;
assign addr[51292]= 1080359326;
assign addr[51293]= 1332945355;
assign addr[51294]= 1558519173;
assign addr[51295]= 1752509516;
assign addr[51296]= 1910985158;
assign addr[51297]= 2030734582;
assign addr[51298]= 2109331059;
assign addr[51299]= 2145181827;
assign addr[51300]= 2137560369;
assign addr[51301]= 2086621133;
assign addr[51302]= 1993396407;
assign addr[51303]= 1859775393;
assign addr[51304]= 1688465931;
assign addr[51305]= 1482939614;
assign addr[51306]= 1247361445;
assign addr[51307]= 986505429;
assign addr[51308]= 705657826;
assign addr[51309]= 410510029;
assign addr[51310]= 107043224;
assign addr[51311]= -198592817;
assign addr[51312]= -500204365;
assign addr[51313]= -791679244;
assign addr[51314]= -1067110699;
assign addr[51315]= -1320917099;
assign addr[51316]= -1547955041;
assign addr[51317]= -1743623590;
assign addr[51318]= -1903957513;
assign addr[51319]= -2025707632;
assign addr[51320]= -2106406677;
assign addr[51321]= -2144419275;
assign addr[51322]= -2138975100;
assign addr[51323]= -2090184478;
assign addr[51324]= -1999036154;
assign addr[51325]= -1867377253;
assign addr[51326]= -1697875851;
assign addr[51327]= -1493966902;
assign addr[51328]= -1259782632;
assign addr[51329]= -1000068799;
assign addr[51330]= -720088517;
assign addr[51331]= -425515602;
assign addr[51332]= -122319591;
assign addr[51333]= 183355234;
assign addr[51334]= 485314355;
assign addr[51335]= 777438554;
assign addr[51336]= 1053807919;
assign addr[51337]= 1308821808;
assign addr[51338]= 1537312353;
assign addr[51339]= 1734649179;
assign addr[51340]= 1896833245;
assign addr[51341]= 2020577882;
assign addr[51342]= 2103375398;
assign addr[51343]= 2143547897;
assign addr[51344]= 2140281282;
assign addr[51345]= 2093641749;
assign addr[51346]= 2004574453;
assign addr[51347]= 1874884346;
assign addr[51348]= 1707199606;
assign addr[51349]= 1504918373;
assign addr[51350]= 1272139887;
assign addr[51351]= 1013581418;
assign addr[51352]= 734482665;
assign addr[51353]= 440499581;
assign addr[51354]= 137589750;
assign addr[51355]= -168108346;
assign addr[51356]= -470399716;
assign addr[51357]= -763158411;
assign addr[51358]= -1040451659;
assign addr[51359]= -1296660098;
assign addr[51360]= -1526591649;
assign addr[51361]= -1725586737;
assign addr[51362]= -1889612716;
assign addr[51363]= -2015345591;
assign addr[51364]= -2100237377;
assign addr[51365]= -2142567738;
assign addr[51366]= -2141478848;
assign addr[51367]= -2096992772;
assign addr[51368]= -2010011024;
assign addr[51369]= -1882296293;
assign addr[51370]= -1716436725;
assign addr[51371]= -1515793473;
assign addr[51372]= -1284432584;
assign addr[51373]= -1027042599;
assign addr[51374]= -748839539;
assign addr[51375]= -455461206;
assign addr[51376]= -152852926;
assign addr[51377]= 152852926;
assign addr[51378]= 455461206;
assign addr[51379]= 748839539;
assign addr[51380]= 1027042599;
assign addr[51381]= 1284432584;
assign addr[51382]= 1515793473;
assign addr[51383]= 1716436725;
assign addr[51384]= 1882296293;
assign addr[51385]= 2010011024;
assign addr[51386]= 2096992772;
assign addr[51387]= 2141478848;
assign addr[51388]= 2142567738;
assign addr[51389]= 2100237377;
assign addr[51390]= 2015345591;
assign addr[51391]= 1889612716;
assign addr[51392]= 1725586737;
assign addr[51393]= 1526591649;
assign addr[51394]= 1296660098;
assign addr[51395]= 1040451659;
assign addr[51396]= 763158411;
assign addr[51397]= 470399716;
assign addr[51398]= 168108346;
assign addr[51399]= -137589750;
assign addr[51400]= -440499581;
assign addr[51401]= -734482665;
assign addr[51402]= -1013581418;
assign addr[51403]= -1272139887;
assign addr[51404]= -1504918373;
assign addr[51405]= -1707199606;
assign addr[51406]= -1874884346;
assign addr[51407]= -2004574453;
assign addr[51408]= -2093641749;
assign addr[51409]= -2140281282;
assign addr[51410]= -2143547897;
assign addr[51411]= -2103375398;
assign addr[51412]= -2020577882;
assign addr[51413]= -1896833245;
assign addr[51414]= -1734649179;
assign addr[51415]= -1537312353;
assign addr[51416]= -1308821808;
assign addr[51417]= -1053807919;
assign addr[51418]= -777438554;
assign addr[51419]= -485314355;
assign addr[51420]= -183355234;
assign addr[51421]= 122319591;
assign addr[51422]= 425515602;
assign addr[51423]= 720088517;
assign addr[51424]= 1000068799;
assign addr[51425]= 1259782632;
assign addr[51426]= 1493966902;
assign addr[51427]= 1697875851;
assign addr[51428]= 1867377253;
assign addr[51429]= 1999036154;
assign addr[51430]= 2090184478;
assign addr[51431]= 2138975100;
assign addr[51432]= 2144419275;
assign addr[51433]= 2106406677;
assign addr[51434]= 2025707632;
assign addr[51435]= 1903957513;
assign addr[51436]= 1743623590;
assign addr[51437]= 1547955041;
assign addr[51438]= 1320917099;
assign addr[51439]= 1067110699;
assign addr[51440]= 791679244;
assign addr[51441]= 500204365;
assign addr[51442]= 198592817;
assign addr[51443]= -107043224;
assign addr[51444]= -410510029;
assign addr[51445]= -705657826;
assign addr[51446]= -986505429;
assign addr[51447]= -1247361445;
assign addr[51448]= -1482939614;
assign addr[51449]= -1688465931;
assign addr[51450]= -1859775393;
assign addr[51451]= -1993396407;
assign addr[51452]= -2086621133;
assign addr[51453]= -2137560369;
assign addr[51454]= -2145181827;
assign addr[51455]= -2109331059;
assign addr[51456]= -2030734582;
assign addr[51457]= -1910985158;
assign addr[51458]= -1752509516;
assign addr[51459]= -1558519173;
assign addr[51460]= -1332945355;
assign addr[51461]= -1080359326;
assign addr[51462]= -805879757;
assign addr[51463]= -515068990;
assign addr[51464]= -213820322;
assign addr[51465]= 91761426;
assign addr[51466]= 395483624;
assign addr[51467]= 691191324;
assign addr[51468]= 972891995;
assign addr[51469]= 1234876957;
assign addr[51470]= 1471837070;
assign addr[51471]= 1678970324;
assign addr[51472]= 1852079154;
assign addr[51473]= 1987655498;
assign addr[51474]= 2082951896;
assign addr[51475]= 2136037160;
assign addr[51476]= 2145835515;
assign addr[51477]= 2112148396;
assign addr[51478]= 2035658475;
assign addr[51479]= 1917915825;
assign addr[51480]= 1761306505;
assign addr[51481]= 1569004214;
assign addr[51482]= 1344905966;
assign addr[51483]= 1093553126;
assign addr[51484]= 820039373;
assign addr[51485]= 529907477;
assign addr[51486]= 229036977;
assign addr[51487]= -76474970;
assign addr[51488]= -380437148;
assign addr[51489]= -676689746;
assign addr[51490]= -959229189;
assign addr[51491]= -1222329801;
assign addr[51492]= -1460659832;
assign addr[51493]= -1669389513;
assign addr[51494]= -1844288924;
assign addr[51495]= -1981813720;
assign addr[51496]= -2079176953;
assign addr[51497]= -2134405552;
assign addr[51498]= -2146380306;
assign addr[51499]= -2114858546;
assign addr[51500]= -2040479063;
assign addr[51501]= -1924749160;
assign addr[51502]= -1770014111;
assign addr[51503]= -1579409630;
assign addr[51504]= -1356798326;
assign addr[51505]= -1106691431;
assign addr[51506]= -834157373;
assign addr[51507]= -544719071;
assign addr[51508]= -244242007;
assign addr[51509]= 61184634;
assign addr[51510]= 365371365;
assign addr[51511]= 662153826;
assign addr[51512]= 945517704;
assign addr[51513]= 1209720613;
assign addr[51514]= 1449408469;
assign addr[51515]= 1659723983;
assign addr[51516]= 1836405100;
assign addr[51517]= 1975871368;
assign addr[51518]= 2075296495;
assign addr[51519]= 2132665626;
assign addr[51520]= 2146816171;
assign addr[51521]= 2117461370;
assign addr[51522]= 2045196100;
assign addr[51523]= 1931484818;
assign addr[51524]= 1778631892;
assign addr[51525]= 1589734894;
assign addr[51526]= 1368621831;
assign addr[51527]= 1119773573;
assign addr[51528]= 848233042;
assign addr[51529]= 559503022;
assign addr[51530]= 259434643;
assign addr[51531]= -45891193;
assign addr[51532]= -350287041;
assign addr[51533]= -647584304;
assign addr[51534]= -931758235;
assign addr[51535]= -1197050035;
assign addr[51536]= -1438083551;
assign addr[51537]= -1649974225;
assign addr[51538]= -1828428082;
assign addr[51539]= -1969828744;
assign addr[51540]= -2071310720;
assign addr[51541]= -2130817471;
assign addr[51542]= -2147143090;
assign addr[51543]= -2119956737;
assign addr[51544]= -2049809346;
assign addr[51545]= -1938122457;
assign addr[51546]= -1787159411;
assign addr[51547]= -1599979481;
assign addr[51548]= -1380375881;
assign addr[51549]= -1132798888;
assign addr[51550]= -862265664;
assign addr[51551]= -574258580;
assign addr[51552]= -274614114;
assign addr[51553]= 30595422;
assign addr[51554]= 335184940;
assign addr[51555]= 632981917;
assign addr[51556]= 917951481;
assign addr[51557]= 1184318708;
assign addr[51558]= 1426685652;
assign addr[51559]= 1640140734;
assign addr[51560]= 1820358275;
assign addr[51561]= 1963686155;
assign addr[51562]= 2067219829;
assign addr[51563]= 2128861181;
assign addr[51564]= 2147361045;
assign addr[51565]= 2122344521;
assign addr[51566]= 2054318569;
assign addr[51567]= 1944661739;
assign addr[51568]= 1795596234;
assign addr[51569]= 1610142873;
assign addr[51570]= 1392059879;
assign addr[51571]= 1145766716;
assign addr[51572]= 876254528;
assign addr[51573]= 588984994;
assign addr[51574]= 289779648;
assign addr[51575]= -15298099;
assign addr[51576]= -320065829;
assign addr[51577]= -618347408;
assign addr[51578]= -904098143;
assign addr[51579]= -1171527280;
assign addr[51580]= -1415215352;
assign addr[51581]= -1630224009;
assign addr[51582]= -1812196087;
assign addr[51583]= -1957443913;
assign addr[51584]= -2063024031;
assign addr[51585]= -2126796855;
assign addr[51586]= -2147470025;
assign addr[51587]= -2124624598;
assign addr[51588]= -2058723538;
assign addr[51589]= -1951102334;
assign addr[51590]= -1803941934;
assign addr[51591]= -1620224553;
assign addr[51592]= -1403673233;
assign addr[51593]= -1158676398;
assign addr[51594]= -890198924;
assign addr[51595]= -603681519;
assign addr[51596]= -304930476;
assign addr[51597]= 0;
assign addr[51598]= 304930476;
assign addr[51599]= 603681519;
assign addr[51600]= 890198924;
assign addr[51601]= 1158676398;
assign addr[51602]= 1403673233;
assign addr[51603]= 1620224553;
assign addr[51604]= 1803941934;
assign addr[51605]= 1951102334;
assign addr[51606]= 2058723538;
assign addr[51607]= 2124624598;
assign addr[51608]= 2147470025;
assign addr[51609]= 2126796855;
assign addr[51610]= 2063024031;
assign addr[51611]= 1957443913;
assign addr[51612]= 1812196087;
assign addr[51613]= 1630224009;
assign addr[51614]= 1415215352;
assign addr[51615]= 1171527280;
assign addr[51616]= 904098143;
assign addr[51617]= 618347408;
assign addr[51618]= 320065829;
assign addr[51619]= 15298099;
assign addr[51620]= -289779648;
assign addr[51621]= -588984994;
assign addr[51622]= -876254528;
assign addr[51623]= -1145766716;
assign addr[51624]= -1392059879;
assign addr[51625]= -1610142873;
assign addr[51626]= -1795596234;
assign addr[51627]= -1944661739;
assign addr[51628]= -2054318569;
assign addr[51629]= -2122344521;
assign addr[51630]= -2147361045;
assign addr[51631]= -2128861181;
assign addr[51632]= -2067219829;
assign addr[51633]= -1963686155;
assign addr[51634]= -1820358275;
assign addr[51635]= -1640140734;
assign addr[51636]= -1426685652;
assign addr[51637]= -1184318708;
assign addr[51638]= -917951481;
assign addr[51639]= -632981917;
assign addr[51640]= -335184940;
assign addr[51641]= -30595422;
assign addr[51642]= 274614114;
assign addr[51643]= 574258580;
assign addr[51644]= 862265664;
assign addr[51645]= 1132798888;
assign addr[51646]= 1380375881;
assign addr[51647]= 1599979481;
assign addr[51648]= 1787159411;
assign addr[51649]= 1938122457;
assign addr[51650]= 2049809346;
assign addr[51651]= 2119956737;
assign addr[51652]= 2147143090;
assign addr[51653]= 2130817471;
assign addr[51654]= 2071310720;
assign addr[51655]= 1969828744;
assign addr[51656]= 1828428082;
assign addr[51657]= 1649974225;
assign addr[51658]= 1438083551;
assign addr[51659]= 1197050035;
assign addr[51660]= 931758235;
assign addr[51661]= 647584304;
assign addr[51662]= 350287041;
assign addr[51663]= 45891193;
assign addr[51664]= -259434643;
assign addr[51665]= -559503022;
assign addr[51666]= -848233042;
assign addr[51667]= -1119773573;
assign addr[51668]= -1368621831;
assign addr[51669]= -1589734894;
assign addr[51670]= -1778631892;
assign addr[51671]= -1931484818;
assign addr[51672]= -2045196100;
assign addr[51673]= -2117461370;
assign addr[51674]= -2146816171;
assign addr[51675]= -2132665626;
assign addr[51676]= -2075296495;
assign addr[51677]= -1975871368;
assign addr[51678]= -1836405100;
assign addr[51679]= -1659723983;
assign addr[51680]= -1449408469;
assign addr[51681]= -1209720613;
assign addr[51682]= -945517704;
assign addr[51683]= -662153826;
assign addr[51684]= -365371365;
assign addr[51685]= -61184634;
assign addr[51686]= 244242007;
assign addr[51687]= 544719071;
assign addr[51688]= 834157373;
assign addr[51689]= 1106691431;
assign addr[51690]= 1356798326;
assign addr[51691]= 1579409630;
assign addr[51692]= 1770014111;
assign addr[51693]= 1924749160;
assign addr[51694]= 2040479063;
assign addr[51695]= 2114858546;
assign addr[51696]= 2146380306;
assign addr[51697]= 2134405552;
assign addr[51698]= 2079176953;
assign addr[51699]= 1981813720;
assign addr[51700]= 1844288924;
assign addr[51701]= 1669389513;
assign addr[51702]= 1460659832;
assign addr[51703]= 1222329801;
assign addr[51704]= 959229189;
assign addr[51705]= 676689746;
assign addr[51706]= 380437148;
assign addr[51707]= 76474970;
assign addr[51708]= -229036977;
assign addr[51709]= -529907477;
assign addr[51710]= -820039373;
assign addr[51711]= -1093553126;
assign addr[51712]= -1344905966;
assign addr[51713]= -1569004214;
assign addr[51714]= -1761306505;
assign addr[51715]= -1917915825;
assign addr[51716]= -2035658475;
assign addr[51717]= -2112148396;
assign addr[51718]= -2145835515;
assign addr[51719]= -2136037160;
assign addr[51720]= -2082951896;
assign addr[51721]= -1987655498;
assign addr[51722]= -1852079154;
assign addr[51723]= -1678970324;
assign addr[51724]= -1471837070;
assign addr[51725]= -1234876957;
assign addr[51726]= -972891995;
assign addr[51727]= -691191324;
assign addr[51728]= -395483624;
assign addr[51729]= -91761426;
assign addr[51730]= 213820322;
assign addr[51731]= 515068990;
assign addr[51732]= 805879757;
assign addr[51733]= 1080359326;
assign addr[51734]= 1332945355;
assign addr[51735]= 1558519173;
assign addr[51736]= 1752509516;
assign addr[51737]= 1910985158;
assign addr[51738]= 2030734582;
assign addr[51739]= 2109331059;
assign addr[51740]= 2145181827;
assign addr[51741]= 2137560369;
assign addr[51742]= 2086621133;
assign addr[51743]= 1993396407;
assign addr[51744]= 1859775393;
assign addr[51745]= 1688465931;
assign addr[51746]= 1482939614;
assign addr[51747]= 1247361445;
assign addr[51748]= 986505429;
assign addr[51749]= 705657826;
assign addr[51750]= 410510029;
assign addr[51751]= 107043224;
assign addr[51752]= -198592817;
assign addr[51753]= -500204365;
assign addr[51754]= -791679244;
assign addr[51755]= -1067110699;
assign addr[51756]= -1320917099;
assign addr[51757]= -1547955041;
assign addr[51758]= -1743623590;
assign addr[51759]= -1903957513;
assign addr[51760]= -2025707632;
assign addr[51761]= -2106406677;
assign addr[51762]= -2144419275;
assign addr[51763]= -2138975100;
assign addr[51764]= -2090184478;
assign addr[51765]= -1999036154;
assign addr[51766]= -1867377253;
assign addr[51767]= -1697875851;
assign addr[51768]= -1493966902;
assign addr[51769]= -1259782632;
assign addr[51770]= -1000068799;
assign addr[51771]= -720088517;
assign addr[51772]= -425515602;
assign addr[51773]= -122319591;
assign addr[51774]= 183355234;
assign addr[51775]= 485314355;
assign addr[51776]= 777438554;
assign addr[51777]= 1053807919;
assign addr[51778]= 1308821808;
assign addr[51779]= 1537312353;
assign addr[51780]= 1734649179;
assign addr[51781]= 1896833245;
assign addr[51782]= 2020577882;
assign addr[51783]= 2103375398;
assign addr[51784]= 2143547897;
assign addr[51785]= 2140281282;
assign addr[51786]= 2093641749;
assign addr[51787]= 2004574453;
assign addr[51788]= 1874884346;
assign addr[51789]= 1707199606;
assign addr[51790]= 1504918373;
assign addr[51791]= 1272139887;
assign addr[51792]= 1013581418;
assign addr[51793]= 734482665;
assign addr[51794]= 440499581;
assign addr[51795]= 137589750;
assign addr[51796]= -168108346;
assign addr[51797]= -470399716;
assign addr[51798]= -763158411;
assign addr[51799]= -1040451659;
assign addr[51800]= -1296660098;
assign addr[51801]= -1526591649;
assign addr[51802]= -1725586737;
assign addr[51803]= -1889612716;
assign addr[51804]= -2015345591;
assign addr[51805]= -2100237377;
assign addr[51806]= -2142567738;
assign addr[51807]= -2141478848;
assign addr[51808]= -2096992772;
assign addr[51809]= -2010011024;
assign addr[51810]= -1882296293;
assign addr[51811]= -1716436725;
assign addr[51812]= -1515793473;
assign addr[51813]= -1284432584;
assign addr[51814]= -1027042599;
assign addr[51815]= -748839539;
assign addr[51816]= -455461206;
assign addr[51817]= -152852926;
assign addr[51818]= 152852926;
assign addr[51819]= 455461206;
assign addr[51820]= 748839539;
assign addr[51821]= 1027042599;
assign addr[51822]= 1284432584;
assign addr[51823]= 1515793473;
assign addr[51824]= 1716436725;
assign addr[51825]= 1882296293;
assign addr[51826]= 2010011024;
assign addr[51827]= 2096992772;
assign addr[51828]= 2141478848;
assign addr[51829]= 2142567738;
assign addr[51830]= 2100237377;
assign addr[51831]= 2015345591;
assign addr[51832]= 1889612716;
assign addr[51833]= 1725586737;
assign addr[51834]= 1526591649;
assign addr[51835]= 1296660098;
assign addr[51836]= 1040451659;
assign addr[51837]= 763158411;
assign addr[51838]= 470399716;
assign addr[51839]= 168108346;
assign addr[51840]= -137589750;
assign addr[51841]= -440499581;
assign addr[51842]= -734482665;
assign addr[51843]= -1013581418;
assign addr[51844]= -1272139887;
assign addr[51845]= -1504918373;
assign addr[51846]= -1707199606;
assign addr[51847]= -1874884346;
assign addr[51848]= -2004574453;
assign addr[51849]= -2093641749;
assign addr[51850]= -2140281282;
assign addr[51851]= -2143547897;
assign addr[51852]= -2103375398;
assign addr[51853]= -2020577882;
assign addr[51854]= -1896833245;
assign addr[51855]= -1734649179;
assign addr[51856]= -1537312353;
assign addr[51857]= -1308821808;
assign addr[51858]= -1053807919;
assign addr[51859]= -777438554;
assign addr[51860]= -485314355;
assign addr[51861]= -183355234;
assign addr[51862]= 122319591;
assign addr[51863]= 425515602;
assign addr[51864]= 720088517;
assign addr[51865]= 1000068799;
assign addr[51866]= 1259782632;
assign addr[51867]= 1493966902;
assign addr[51868]= 1697875851;
assign addr[51869]= 1867377253;
assign addr[51870]= 1999036154;
assign addr[51871]= 2090184478;
assign addr[51872]= 2138975100;
assign addr[51873]= 2144419275;
assign addr[51874]= 2106406677;
assign addr[51875]= 2025707632;
assign addr[51876]= 1903957513;
assign addr[51877]= 1743623590;
assign addr[51878]= 1547955041;
assign addr[51879]= 1320917099;
assign addr[51880]= 1067110699;
assign addr[51881]= 791679244;
assign addr[51882]= 500204365;
assign addr[51883]= 198592817;
assign addr[51884]= -107043224;
assign addr[51885]= -410510029;
assign addr[51886]= -705657826;
assign addr[51887]= -986505429;
assign addr[51888]= -1247361445;
assign addr[51889]= -1482939614;
assign addr[51890]= -1688465931;
assign addr[51891]= -1859775393;
assign addr[51892]= -1993396407;
assign addr[51893]= -2086621133;
assign addr[51894]= -2137560369;
assign addr[51895]= -2145181827;
assign addr[51896]= -2109331059;
assign addr[51897]= -2030734582;
assign addr[51898]= -1910985158;
assign addr[51899]= -1752509516;
assign addr[51900]= -1558519173;
assign addr[51901]= -1332945355;
assign addr[51902]= -1080359326;
assign addr[51903]= -805879757;
assign addr[51904]= -515068990;
assign addr[51905]= -213820322;
assign addr[51906]= 91761426;
assign addr[51907]= 395483624;
assign addr[51908]= 691191324;
assign addr[51909]= 972891995;
assign addr[51910]= 1234876957;
assign addr[51911]= 1471837070;
assign addr[51912]= 1678970324;
assign addr[51913]= 1852079154;
assign addr[51914]= 1987655498;
assign addr[51915]= 2082951896;
assign addr[51916]= 2136037160;
assign addr[51917]= 2145835515;
assign addr[51918]= 2112148396;
assign addr[51919]= 2035658475;
assign addr[51920]= 1917915825;
assign addr[51921]= 1761306505;
assign addr[51922]= 1569004214;
assign addr[51923]= 1344905966;
assign addr[51924]= 1093553126;
assign addr[51925]= 820039373;
assign addr[51926]= 529907477;
assign addr[51927]= 229036977;
assign addr[51928]= -76474970;
assign addr[51929]= -380437148;
assign addr[51930]= -676689746;
assign addr[51931]= -959229189;
assign addr[51932]= -1222329801;
assign addr[51933]= -1460659832;
assign addr[51934]= -1669389513;
assign addr[51935]= -1844288924;
assign addr[51936]= -1981813720;
assign addr[51937]= -2079176953;
assign addr[51938]= -2134405552;
assign addr[51939]= -2146380306;
assign addr[51940]= -2114858546;
assign addr[51941]= -2040479063;
assign addr[51942]= -1924749160;
assign addr[51943]= -1770014111;
assign addr[51944]= -1579409630;
assign addr[51945]= -1356798326;
assign addr[51946]= -1106691431;
assign addr[51947]= -834157373;
assign addr[51948]= -544719071;
assign addr[51949]= -244242007;
assign addr[51950]= 61184634;
assign addr[51951]= 365371365;
assign addr[51952]= 662153826;
assign addr[51953]= 945517704;
assign addr[51954]= 1209720613;
assign addr[51955]= 1449408469;
assign addr[51956]= 1659723983;
assign addr[51957]= 1836405100;
assign addr[51958]= 1975871368;
assign addr[51959]= 2075296495;
assign addr[51960]= 2132665626;
assign addr[51961]= 2146816171;
assign addr[51962]= 2117461370;
assign addr[51963]= 2045196100;
assign addr[51964]= 1931484818;
assign addr[51965]= 1778631892;
assign addr[51966]= 1589734894;
assign addr[51967]= 1368621831;
assign addr[51968]= 1119773573;
assign addr[51969]= 848233042;
assign addr[51970]= 559503022;
assign addr[51971]= 259434643;
assign addr[51972]= -45891193;
assign addr[51973]= -350287041;
assign addr[51974]= -647584304;
assign addr[51975]= -931758235;
assign addr[51976]= -1197050035;
assign addr[51977]= -1438083551;
assign addr[51978]= -1649974225;
assign addr[51979]= -1828428082;
assign addr[51980]= -1969828744;
assign addr[51981]= -2071310720;
assign addr[51982]= -2130817471;
assign addr[51983]= -2147143090;
assign addr[51984]= -2119956737;
assign addr[51985]= -2049809346;
assign addr[51986]= -1938122457;
assign addr[51987]= -1787159411;
assign addr[51988]= -1599979481;
assign addr[51989]= -1380375881;
assign addr[51990]= -1132798888;
assign addr[51991]= -862265664;
assign addr[51992]= -574258580;
assign addr[51993]= -274614114;
assign addr[51994]= 30595422;
assign addr[51995]= 335184940;
assign addr[51996]= 632981917;
assign addr[51997]= 917951481;
assign addr[51998]= 1184318708;
assign addr[51999]= 1426685652;
assign addr[52000]= 1640140734;
assign addr[52001]= 1820358275;
assign addr[52002]= 1963686155;
assign addr[52003]= 2067219829;
assign addr[52004]= 2128861181;
assign addr[52005]= 2147361045;
assign addr[52006]= 2122344521;
assign addr[52007]= 2054318569;
assign addr[52008]= 1944661739;
assign addr[52009]= 1795596234;
assign addr[52010]= 1610142873;
assign addr[52011]= 1392059879;
assign addr[52012]= 1145766716;
assign addr[52013]= 876254528;
assign addr[52014]= 588984994;
assign addr[52015]= 289779648;
assign addr[52016]= -15298099;
assign addr[52017]= -320065829;
assign addr[52018]= -618347408;
assign addr[52019]= -904098143;
assign addr[52020]= -1171527280;
assign addr[52021]= -1415215352;
assign addr[52022]= -1630224009;
assign addr[52023]= -1812196087;
assign addr[52024]= -1957443913;
assign addr[52025]= -2063024031;
assign addr[52026]= -2126796855;
assign addr[52027]= -2147470025;
assign addr[52028]= -2124624598;
assign addr[52029]= -2058723538;
assign addr[52030]= -1951102334;
assign addr[52031]= -1803941934;
assign addr[52032]= -1620224553;
assign addr[52033]= -1403673233;
assign addr[52034]= -1158676398;
assign addr[52035]= -890198924;
assign addr[52036]= -603681519;
assign addr[52037]= -304930476;
assign addr[52038]= 0;
assign addr[52039]= 304930476;
assign addr[52040]= 603681519;
assign addr[52041]= 890198924;
assign addr[52042]= 1158676398;
assign addr[52043]= 1403673233;
assign addr[52044]= 1620224553;
assign addr[52045]= 1803941934;
assign addr[52046]= 1951102334;
assign addr[52047]= 2058723538;
assign addr[52048]= 2124624598;
assign addr[52049]= 2147470025;
assign addr[52050]= 2126796855;
assign addr[52051]= 2063024031;
assign addr[52052]= 1957443913;
assign addr[52053]= 1812196087;
assign addr[52054]= 1630224009;
assign addr[52055]= 1415215352;
assign addr[52056]= 1171527280;
assign addr[52057]= 904098143;
assign addr[52058]= 618347408;
assign addr[52059]= 320065829;
assign addr[52060]= 15298099;
assign addr[52061]= -289779648;
assign addr[52062]= -588984994;
assign addr[52063]= -876254528;
assign addr[52064]= -1145766716;
assign addr[52065]= -1392059879;
assign addr[52066]= -1610142873;
assign addr[52067]= -1795596234;
assign addr[52068]= -1944661739;
assign addr[52069]= -2054318569;
assign addr[52070]= -2122344521;
assign addr[52071]= -2147361045;
assign addr[52072]= -2128861181;
assign addr[52073]= -2067219829;
assign addr[52074]= -1963686155;
assign addr[52075]= -1820358275;
assign addr[52076]= -1640140734;
assign addr[52077]= -1426685652;
assign addr[52078]= -1184318708;
assign addr[52079]= -917951481;
assign addr[52080]= -632981917;
assign addr[52081]= -335184940;
assign addr[52082]= -30595422;
assign addr[52083]= 274614114;
assign addr[52084]= 574258580;
assign addr[52085]= 862265664;
assign addr[52086]= 1132798888;
assign addr[52087]= 1380375881;
assign addr[52088]= 1599979481;
assign addr[52089]= 1787159411;
assign addr[52090]= 1938122457;
assign addr[52091]= 2049809346;
assign addr[52092]= 2119956737;
assign addr[52093]= 2147143090;
assign addr[52094]= 2130817471;
assign addr[52095]= 2071310720;
assign addr[52096]= 1969828744;
assign addr[52097]= 1828428082;
assign addr[52098]= 1649974225;
assign addr[52099]= 1438083551;
assign addr[52100]= 1197050035;
assign addr[52101]= 931758235;
assign addr[52102]= 647584304;
assign addr[52103]= 350287041;
assign addr[52104]= 45891193;
assign addr[52105]= -259434643;
assign addr[52106]= -559503022;
assign addr[52107]= -848233042;
assign addr[52108]= -1119773573;
assign addr[52109]= -1368621831;
assign addr[52110]= -1589734894;
assign addr[52111]= -1778631892;
assign addr[52112]= -1931484818;
assign addr[52113]= -2045196100;
assign addr[52114]= -2117461370;
assign addr[52115]= -2146816171;
assign addr[52116]= -2132665626;
assign addr[52117]= -2075296495;
assign addr[52118]= -1975871368;
assign addr[52119]= -1836405100;
assign addr[52120]= -1659723983;
assign addr[52121]= -1449408469;
assign addr[52122]= -1209720613;
assign addr[52123]= -945517704;
assign addr[52124]= -662153826;
assign addr[52125]= -365371365;
assign addr[52126]= -61184634;
assign addr[52127]= 244242007;
assign addr[52128]= 544719071;
assign addr[52129]= 834157373;
assign addr[52130]= 1106691431;
assign addr[52131]= 1356798326;
assign addr[52132]= 1579409630;
assign addr[52133]= 1770014111;
assign addr[52134]= 1924749160;
assign addr[52135]= 2040479063;
assign addr[52136]= 2114858546;
assign addr[52137]= 2146380306;
assign addr[52138]= 2134405552;
assign addr[52139]= 2079176953;
assign addr[52140]= 1981813720;
assign addr[52141]= 1844288924;
assign addr[52142]= 1669389513;
assign addr[52143]= 1460659832;
assign addr[52144]= 1222329801;
assign addr[52145]= 959229189;
assign addr[52146]= 676689746;
assign addr[52147]= 380437148;
assign addr[52148]= 76474970;
assign addr[52149]= -229036977;
assign addr[52150]= -529907477;
assign addr[52151]= -820039373;
assign addr[52152]= -1093553126;
assign addr[52153]= -1344905966;
assign addr[52154]= -1569004214;
assign addr[52155]= -1761306505;
assign addr[52156]= -1917915825;
assign addr[52157]= -2035658475;
assign addr[52158]= -2112148396;
assign addr[52159]= -2145835515;
assign addr[52160]= -2136037160;
assign addr[52161]= -2082951896;
assign addr[52162]= -1987655498;
assign addr[52163]= -1852079154;
assign addr[52164]= -1678970324;
assign addr[52165]= -1471837070;
assign addr[52166]= -1234876957;
assign addr[52167]= -972891995;
assign addr[52168]= -691191324;
assign addr[52169]= -395483624;
assign addr[52170]= -91761426;
assign addr[52171]= 213820322;
assign addr[52172]= 515068990;
assign addr[52173]= 805879757;
assign addr[52174]= 1080359326;
assign addr[52175]= 1332945355;
assign addr[52176]= 1558519173;
assign addr[52177]= 1752509516;
assign addr[52178]= 1910985158;
assign addr[52179]= 2030734582;
assign addr[52180]= 2109331059;
assign addr[52181]= 2145181827;
assign addr[52182]= 2137560369;
assign addr[52183]= 2086621133;
assign addr[52184]= 1993396407;
assign addr[52185]= 1859775393;
assign addr[52186]= 1688465931;
assign addr[52187]= 1482939614;
assign addr[52188]= 1247361445;
assign addr[52189]= 986505429;
assign addr[52190]= 705657826;
assign addr[52191]= 410510029;
assign addr[52192]= 107043224;
assign addr[52193]= -198592817;
assign addr[52194]= -500204365;
assign addr[52195]= -791679244;
assign addr[52196]= -1067110699;
assign addr[52197]= -1320917099;
assign addr[52198]= -1547955041;
assign addr[52199]= -1743623590;
assign addr[52200]= -1903957513;
assign addr[52201]= -2025707632;
assign addr[52202]= -2106406677;
assign addr[52203]= -2144419275;
assign addr[52204]= -2138975100;
assign addr[52205]= -2090184478;
assign addr[52206]= -1999036154;
assign addr[52207]= -1867377253;
assign addr[52208]= -1697875851;
assign addr[52209]= -1493966902;
assign addr[52210]= -1259782632;
assign addr[52211]= -1000068799;
assign addr[52212]= -720088517;
assign addr[52213]= -425515602;
assign addr[52214]= -122319591;
assign addr[52215]= 183355234;
assign addr[52216]= 485314355;
assign addr[52217]= 777438554;
assign addr[52218]= 1053807919;
assign addr[52219]= 1308821808;
assign addr[52220]= 1537312353;
assign addr[52221]= 1734649179;
assign addr[52222]= 1896833245;
assign addr[52223]= 2020577882;
assign addr[52224]= 2103375398;
assign addr[52225]= 2143547897;
assign addr[52226]= 2140281282;
assign addr[52227]= 2093641749;
assign addr[52228]= 2004574453;
assign addr[52229]= 1874884346;
assign addr[52230]= 1707199606;
assign addr[52231]= 1504918373;
assign addr[52232]= 1272139887;
assign addr[52233]= 1013581418;
assign addr[52234]= 734482665;
assign addr[52235]= 440499581;
assign addr[52236]= 137589750;
assign addr[52237]= -168108346;
assign addr[52238]= -470399716;
assign addr[52239]= -763158411;
assign addr[52240]= -1040451659;
assign addr[52241]= -1296660098;
assign addr[52242]= -1526591649;
assign addr[52243]= -1725586737;
assign addr[52244]= -1889612716;
assign addr[52245]= -2015345591;
assign addr[52246]= -2100237377;
assign addr[52247]= -2142567738;
assign addr[52248]= -2141478848;
assign addr[52249]= -2096992772;
assign addr[52250]= -2010011024;
assign addr[52251]= -1882296293;
assign addr[52252]= -1716436725;
assign addr[52253]= -1515793473;
assign addr[52254]= -1284432584;
assign addr[52255]= -1027042599;
assign addr[52256]= -748839539;
assign addr[52257]= -455461206;
assign addr[52258]= -152852926;
assign addr[52259]= 152852926;
assign addr[52260]= 455461206;
assign addr[52261]= 748839539;
assign addr[52262]= 1027042599;
assign addr[52263]= 1284432584;
assign addr[52264]= 1515793473;
assign addr[52265]= 1716436725;
assign addr[52266]= 1882296293;
assign addr[52267]= 2010011024;
assign addr[52268]= 2096992772;
assign addr[52269]= 2141478848;
assign addr[52270]= 2142567738;
assign addr[52271]= 2100237377;
assign addr[52272]= 2015345591;
assign addr[52273]= 1889612716;
assign addr[52274]= 1725586737;
assign addr[52275]= 1526591649;
assign addr[52276]= 1296660098;
assign addr[52277]= 1040451659;
assign addr[52278]= 763158411;
assign addr[52279]= 470399716;
assign addr[52280]= 168108346;
assign addr[52281]= -137589750;
assign addr[52282]= -440499581;
assign addr[52283]= -734482665;
assign addr[52284]= -1013581418;
assign addr[52285]= -1272139887;
assign addr[52286]= -1504918373;
assign addr[52287]= -1707199606;
assign addr[52288]= -1874884346;
assign addr[52289]= -2004574453;
assign addr[52290]= -2093641749;
assign addr[52291]= -2140281282;
assign addr[52292]= -2143547897;
assign addr[52293]= -2103375398;
assign addr[52294]= -2020577882;
assign addr[52295]= -1896833245;
assign addr[52296]= -1734649179;
assign addr[52297]= -1537312353;
assign addr[52298]= -1308821808;
assign addr[52299]= -1053807919;
assign addr[52300]= -777438554;
assign addr[52301]= -485314355;
assign addr[52302]= -183355234;
assign addr[52303]= 122319591;
assign addr[52304]= 425515602;
assign addr[52305]= 720088517;
assign addr[52306]= 1000068799;
assign addr[52307]= 1259782632;
assign addr[52308]= 1493966902;
assign addr[52309]= 1697875851;
assign addr[52310]= 1867377253;
assign addr[52311]= 1999036154;
assign addr[52312]= 2090184478;
assign addr[52313]= 2138975100;
assign addr[52314]= 2144419275;
assign addr[52315]= 2106406677;
assign addr[52316]= 2025707632;
assign addr[52317]= 1903957513;
assign addr[52318]= 1743623590;
assign addr[52319]= 1547955041;
assign addr[52320]= 1320917099;
assign addr[52321]= 1067110699;
assign addr[52322]= 791679244;
assign addr[52323]= 500204365;
assign addr[52324]= 198592817;
assign addr[52325]= -107043224;
assign addr[52326]= -410510029;
assign addr[52327]= -705657826;
assign addr[52328]= -986505429;
assign addr[52329]= -1247361445;
assign addr[52330]= -1482939614;
assign addr[52331]= -1688465931;
assign addr[52332]= -1859775393;
assign addr[52333]= -1993396407;
assign addr[52334]= -2086621133;
assign addr[52335]= -2137560369;
assign addr[52336]= -2145181827;
assign addr[52337]= -2109331059;
assign addr[52338]= -2030734582;
assign addr[52339]= -1910985158;
assign addr[52340]= -1752509516;
assign addr[52341]= -1558519173;
assign addr[52342]= -1332945355;
assign addr[52343]= -1080359326;
assign addr[52344]= -805879757;
assign addr[52345]= -515068990;
assign addr[52346]= -213820322;
assign addr[52347]= 91761426;
assign addr[52348]= 395483624;
assign addr[52349]= 691191324;
assign addr[52350]= 972891995;
assign addr[52351]= 1234876957;
assign addr[52352]= 1471837070;
assign addr[52353]= 1678970324;
assign addr[52354]= 1852079154;
assign addr[52355]= 1987655498;
assign addr[52356]= 2082951896;
assign addr[52357]= 2136037160;
assign addr[52358]= 2145835515;
assign addr[52359]= 2112148396;
assign addr[52360]= 2035658475;
assign addr[52361]= 1917915825;
assign addr[52362]= 1761306505;
assign addr[52363]= 1569004214;
assign addr[52364]= 1344905966;
assign addr[52365]= 1093553126;
assign addr[52366]= 820039373;
assign addr[52367]= 529907477;
assign addr[52368]= 229036977;
assign addr[52369]= -76474970;
assign addr[52370]= -380437148;
assign addr[52371]= -676689746;
assign addr[52372]= -959229189;
assign addr[52373]= -1222329801;
assign addr[52374]= -1460659832;
assign addr[52375]= -1669389513;
assign addr[52376]= -1844288924;
assign addr[52377]= -1981813720;
assign addr[52378]= -2079176953;
assign addr[52379]= -2134405552;
assign addr[52380]= -2146380306;
assign addr[52381]= -2114858546;
assign addr[52382]= -2040479063;
assign addr[52383]= -1924749160;
assign addr[52384]= -1770014111;
assign addr[52385]= -1579409630;
assign addr[52386]= -1356798326;
assign addr[52387]= -1106691431;
assign addr[52388]= -834157373;
assign addr[52389]= -544719071;
assign addr[52390]= -244242007;
assign addr[52391]= 61184634;
assign addr[52392]= 365371365;
assign addr[52393]= 662153826;
assign addr[52394]= 945517704;
assign addr[52395]= 1209720613;
assign addr[52396]= 1449408469;
assign addr[52397]= 1659723983;
assign addr[52398]= 1836405100;
assign addr[52399]= 1975871368;
assign addr[52400]= 2075296495;
assign addr[52401]= 2132665626;
assign addr[52402]= 2146816171;
assign addr[52403]= 2117461370;
assign addr[52404]= 2045196100;
assign addr[52405]= 1931484818;
assign addr[52406]= 1778631892;
assign addr[52407]= 1589734894;
assign addr[52408]= 1368621831;
assign addr[52409]= 1119773573;
assign addr[52410]= 848233042;
assign addr[52411]= 559503022;
assign addr[52412]= 259434643;
assign addr[52413]= -45891193;
assign addr[52414]= -350287041;
assign addr[52415]= -647584304;
assign addr[52416]= -931758235;
assign addr[52417]= -1197050035;
assign addr[52418]= -1438083551;
assign addr[52419]= -1649974225;
assign addr[52420]= -1828428082;
assign addr[52421]= -1969828744;
assign addr[52422]= -2071310720;
assign addr[52423]= -2130817471;
assign addr[52424]= -2147143090;
assign addr[52425]= -2119956737;
assign addr[52426]= -2049809346;
assign addr[52427]= -1938122457;
assign addr[52428]= -1787159411;
assign addr[52429]= -1599979481;
assign addr[52430]= -1380375881;
assign addr[52431]= -1132798888;
assign addr[52432]= -862265664;
assign addr[52433]= -574258580;
assign addr[52434]= -274614114;
assign addr[52435]= 30595422;
assign addr[52436]= 335184940;
assign addr[52437]= 632981917;
assign addr[52438]= 917951481;
assign addr[52439]= 1184318708;
assign addr[52440]= 1426685652;
assign addr[52441]= 1640140734;
assign addr[52442]= 1820358275;
assign addr[52443]= 1963686155;
assign addr[52444]= 2067219829;
assign addr[52445]= 2128861181;
assign addr[52446]= 2147361045;
assign addr[52447]= 2122344521;
assign addr[52448]= 2054318569;
assign addr[52449]= 1944661739;
assign addr[52450]= 1795596234;
assign addr[52451]= 1610142873;
assign addr[52452]= 1392059879;
assign addr[52453]= 1145766716;
assign addr[52454]= 876254528;
assign addr[52455]= 588984994;
assign addr[52456]= 289779648;
assign addr[52457]= -15298099;
assign addr[52458]= -320065829;
assign addr[52459]= -618347408;
assign addr[52460]= -904098143;
assign addr[52461]= -1171527280;
assign addr[52462]= -1415215352;
assign addr[52463]= -1630224009;
assign addr[52464]= -1812196087;
assign addr[52465]= -1957443913;
assign addr[52466]= -2063024031;
assign addr[52467]= -2126796855;
assign addr[52468]= -2147470025;
assign addr[52469]= -2124624598;
assign addr[52470]= -2058723538;
assign addr[52471]= -1951102334;
assign addr[52472]= -1803941934;
assign addr[52473]= -1620224553;
assign addr[52474]= -1403673233;
assign addr[52475]= -1158676398;
assign addr[52476]= -890198924;
assign addr[52477]= -603681519;
assign addr[52478]= -304930476;
assign addr[52479]= 0;
assign addr[52480]= 304930476;
assign addr[52481]= 603681519;
assign addr[52482]= 890198924;
assign addr[52483]= 1158676398;
assign addr[52484]= 1403673233;
assign addr[52485]= 1620224553;
assign addr[52486]= 1803941934;
assign addr[52487]= 1951102334;
assign addr[52488]= 2058723538;
assign addr[52489]= 2124624598;
assign addr[52490]= 2147470025;
assign addr[52491]= 2126796855;
assign addr[52492]= 2063024031;
assign addr[52493]= 1957443913;
assign addr[52494]= 1812196087;
assign addr[52495]= 1630224009;
assign addr[52496]= 1415215352;
assign addr[52497]= 1171527280;
assign addr[52498]= 904098143;
assign addr[52499]= 618347408;
assign addr[52500]= 320065829;
assign addr[52501]= 15298099;
assign addr[52502]= -289779648;
assign addr[52503]= -588984994;
assign addr[52504]= -876254528;
assign addr[52505]= -1145766716;
assign addr[52506]= -1392059879;
assign addr[52507]= -1610142873;
assign addr[52508]= -1795596234;
assign addr[52509]= -1944661739;
assign addr[52510]= -2054318569;
assign addr[52511]= -2122344521;
assign addr[52512]= -2147361045;
assign addr[52513]= -2128861181;
assign addr[52514]= -2067219829;
assign addr[52515]= -1963686155;
assign addr[52516]= -1820358275;
assign addr[52517]= -1640140734;
assign addr[52518]= -1426685652;
assign addr[52519]= -1184318708;
assign addr[52520]= -917951481;
assign addr[52521]= -632981917;
assign addr[52522]= -335184940;
assign addr[52523]= -30595422;
assign addr[52524]= 274614114;
assign addr[52525]= 574258580;
assign addr[52526]= 862265664;
assign addr[52527]= 1132798888;
assign addr[52528]= 1380375881;
assign addr[52529]= 1599979481;
assign addr[52530]= 1787159411;
assign addr[52531]= 1938122457;
assign addr[52532]= 2049809346;
assign addr[52533]= 2119956737;
assign addr[52534]= 2147143090;
assign addr[52535]= 2130817471;
assign addr[52536]= 2071310720;
assign addr[52537]= 1969828744;
assign addr[52538]= 1828428082;
assign addr[52539]= 1649974225;
assign addr[52540]= 1438083551;
assign addr[52541]= 1197050035;
assign addr[52542]= 931758235;
assign addr[52543]= 647584304;
assign addr[52544]= 350287041;
assign addr[52545]= 45891193;
assign addr[52546]= -259434643;
assign addr[52547]= -559503022;
assign addr[52548]= -848233042;
assign addr[52549]= -1119773573;
assign addr[52550]= -1368621831;
assign addr[52551]= -1589734894;
assign addr[52552]= -1778631892;
assign addr[52553]= -1931484818;
assign addr[52554]= -2045196100;
assign addr[52555]= -2117461370;
assign addr[52556]= -2146816171;
assign addr[52557]= -2132665626;
assign addr[52558]= -2075296495;
assign addr[52559]= -1975871368;
assign addr[52560]= -1836405100;
assign addr[52561]= -1659723983;
assign addr[52562]= -1449408469;
assign addr[52563]= -1209720613;
assign addr[52564]= -945517704;
assign addr[52565]= -662153826;
assign addr[52566]= -365371365;
assign addr[52567]= -61184634;
assign addr[52568]= 244242007;
assign addr[52569]= 544719071;
assign addr[52570]= 834157373;
assign addr[52571]= 1106691431;
assign addr[52572]= 1356798326;
assign addr[52573]= 1579409630;
assign addr[52574]= 1770014111;
assign addr[52575]= 1924749160;
assign addr[52576]= 2040479063;
assign addr[52577]= 2114858546;
assign addr[52578]= 2146380306;
assign addr[52579]= 2134405552;
assign addr[52580]= 2079176953;
assign addr[52581]= 1981813720;
assign addr[52582]= 1844288924;
assign addr[52583]= 1669389513;
assign addr[52584]= 1460659832;
assign addr[52585]= 1222329801;
assign addr[52586]= 959229189;
assign addr[52587]= 676689746;
assign addr[52588]= 380437148;
assign addr[52589]= 76474970;
assign addr[52590]= -229036977;
assign addr[52591]= -529907477;
assign addr[52592]= -820039373;
assign addr[52593]= -1093553126;
assign addr[52594]= -1344905966;
assign addr[52595]= -1569004214;
assign addr[52596]= -1761306505;
assign addr[52597]= -1917915825;
assign addr[52598]= -2035658475;
assign addr[52599]= -2112148396;
assign addr[52600]= -2145835515;
assign addr[52601]= -2136037160;
assign addr[52602]= -2082951896;
assign addr[52603]= -1987655498;
assign addr[52604]= -1852079154;
assign addr[52605]= -1678970324;
assign addr[52606]= -1471837070;
assign addr[52607]= -1234876957;
assign addr[52608]= -972891995;
assign addr[52609]= -691191324;
assign addr[52610]= -395483624;
assign addr[52611]= -91761426;
assign addr[52612]= 213820322;
assign addr[52613]= 515068990;
assign addr[52614]= 805879757;
assign addr[52615]= 1080359326;
assign addr[52616]= 1332945355;
assign addr[52617]= 1558519173;
assign addr[52618]= 1752509516;
assign addr[52619]= 1910985158;
assign addr[52620]= 2030734582;
assign addr[52621]= 2109331059;
assign addr[52622]= 2145181827;
assign addr[52623]= 2137560369;
assign addr[52624]= 2086621133;
assign addr[52625]= 1993396407;
assign addr[52626]= 1859775393;
assign addr[52627]= 1688465931;
assign addr[52628]= 1482939614;
assign addr[52629]= 1247361445;
assign addr[52630]= 986505429;
assign addr[52631]= 705657826;
assign addr[52632]= 410510029;
assign addr[52633]= 107043224;
assign addr[52634]= -198592817;
assign addr[52635]= -500204365;
assign addr[52636]= -791679244;
assign addr[52637]= -1067110699;
assign addr[52638]= -1320917099;
assign addr[52639]= -1547955041;
assign addr[52640]= -1743623590;
assign addr[52641]= -1903957513;
assign addr[52642]= -2025707632;
assign addr[52643]= -2106406677;
assign addr[52644]= -2144419275;
assign addr[52645]= -2138975100;
assign addr[52646]= -2090184478;
assign addr[52647]= -1999036154;
assign addr[52648]= -1867377253;
assign addr[52649]= -1697875851;
assign addr[52650]= -1493966902;
assign addr[52651]= -1259782632;
assign addr[52652]= -1000068799;
assign addr[52653]= -720088517;
assign addr[52654]= -425515602;
assign addr[52655]= -122319591;
assign addr[52656]= 183355234;
assign addr[52657]= 485314355;
assign addr[52658]= 777438554;
assign addr[52659]= 1053807919;
assign addr[52660]= 1308821808;
assign addr[52661]= 1537312353;
assign addr[52662]= 1734649179;
assign addr[52663]= 1896833245;
assign addr[52664]= 2020577882;
assign addr[52665]= 2103375398;
assign addr[52666]= 2143547897;
assign addr[52667]= 2140281282;
assign addr[52668]= 2093641749;
assign addr[52669]= 2004574453;
assign addr[52670]= 1874884346;
assign addr[52671]= 1707199606;
assign addr[52672]= 1504918373;
assign addr[52673]= 1272139887;
assign addr[52674]= 1013581418;
assign addr[52675]= 734482665;
assign addr[52676]= 440499581;
assign addr[52677]= 137589750;
assign addr[52678]= -168108346;
assign addr[52679]= -470399716;
assign addr[52680]= -763158411;
assign addr[52681]= -1040451659;
assign addr[52682]= -1296660098;
assign addr[52683]= -1526591649;
assign addr[52684]= -1725586737;
assign addr[52685]= -1889612716;
assign addr[52686]= -2015345591;
assign addr[52687]= -2100237377;
assign addr[52688]= -2142567738;
assign addr[52689]= -2141478848;
assign addr[52690]= -2096992772;
assign addr[52691]= -2010011024;
assign addr[52692]= -1882296293;
assign addr[52693]= -1716436725;
assign addr[52694]= -1515793473;
assign addr[52695]= -1284432584;
assign addr[52696]= -1027042599;
assign addr[52697]= -748839539;
assign addr[52698]= -455461206;
assign addr[52699]= -152852926;
assign addr[52700]= 152852926;
assign addr[52701]= 455461206;
assign addr[52702]= 748839539;
assign addr[52703]= 1027042599;
assign addr[52704]= 1284432584;
assign addr[52705]= 1515793473;
assign addr[52706]= 1716436725;
assign addr[52707]= 1882296293;
assign addr[52708]= 2010011024;
assign addr[52709]= 2096992772;
assign addr[52710]= 2141478848;
assign addr[52711]= 2142567738;
assign addr[52712]= 2100237377;
assign addr[52713]= 2015345591;
assign addr[52714]= 1889612716;
assign addr[52715]= 1725586737;
assign addr[52716]= 1526591649;
assign addr[52717]= 1296660098;
assign addr[52718]= 1040451659;
assign addr[52719]= 763158411;
assign addr[52720]= 470399716;
assign addr[52721]= 168108346;
assign addr[52722]= -137589750;
assign addr[52723]= -440499581;
assign addr[52724]= -734482665;
assign addr[52725]= -1013581418;
assign addr[52726]= -1272139887;
assign addr[52727]= -1504918373;
assign addr[52728]= -1707199606;
assign addr[52729]= -1874884346;
assign addr[52730]= -2004574453;
assign addr[52731]= -2093641749;
assign addr[52732]= -2140281282;
assign addr[52733]= -2143547897;
assign addr[52734]= -2103375398;
assign addr[52735]= -2020577882;
assign addr[52736]= -1896833245;
assign addr[52737]= -1734649179;
assign addr[52738]= -1537312353;
assign addr[52739]= -1308821808;
assign addr[52740]= -1053807919;
assign addr[52741]= -777438554;
assign addr[52742]= -485314355;
assign addr[52743]= -183355234;
assign addr[52744]= 122319591;
assign addr[52745]= 425515602;
assign addr[52746]= 720088517;
assign addr[52747]= 1000068799;
assign addr[52748]= 1259782632;
assign addr[52749]= 1493966902;
assign addr[52750]= 1697875851;
assign addr[52751]= 1867377253;
assign addr[52752]= 1999036154;
assign addr[52753]= 2090184478;
assign addr[52754]= 2138975100;
assign addr[52755]= 2144419275;
assign addr[52756]= 2106406677;
assign addr[52757]= 2025707632;
assign addr[52758]= 1903957513;
assign addr[52759]= 1743623590;
assign addr[52760]= 1547955041;
assign addr[52761]= 1320917099;
assign addr[52762]= 1067110699;
assign addr[52763]= 791679244;
assign addr[52764]= 500204365;
assign addr[52765]= 198592817;
assign addr[52766]= -107043224;
assign addr[52767]= -410510029;
assign addr[52768]= -705657826;
assign addr[52769]= -986505429;
assign addr[52770]= -1247361445;
assign addr[52771]= -1482939614;
assign addr[52772]= -1688465931;
assign addr[52773]= -1859775393;
assign addr[52774]= -1993396407;
assign addr[52775]= -2086621133;
assign addr[52776]= -2137560369;
assign addr[52777]= -2145181827;
assign addr[52778]= -2109331059;
assign addr[52779]= -2030734582;
assign addr[52780]= -1910985158;
assign addr[52781]= -1752509516;
assign addr[52782]= -1558519173;
assign addr[52783]= -1332945355;
assign addr[52784]= -1080359326;
assign addr[52785]= -805879757;
assign addr[52786]= -515068990;
assign addr[52787]= -213820322;
assign addr[52788]= 91761426;
assign addr[52789]= 395483624;
assign addr[52790]= 691191324;
assign addr[52791]= 972891995;
assign addr[52792]= 1234876957;
assign addr[52793]= 1471837070;
assign addr[52794]= 1678970324;
assign addr[52795]= 1852079154;
assign addr[52796]= 1987655498;
assign addr[52797]= 2082951896;
assign addr[52798]= 2136037160;
assign addr[52799]= 2145835515;
assign addr[52800]= 2112148396;
assign addr[52801]= 2035658475;
assign addr[52802]= 1917915825;
assign addr[52803]= 1761306505;
assign addr[52804]= 1569004214;
assign addr[52805]= 1344905966;
assign addr[52806]= 1093553126;
assign addr[52807]= 820039373;
assign addr[52808]= 529907477;
assign addr[52809]= 229036977;
assign addr[52810]= -76474970;
assign addr[52811]= -380437148;
assign addr[52812]= -676689746;
assign addr[52813]= -959229189;
assign addr[52814]= -1222329801;
assign addr[52815]= -1460659832;
assign addr[52816]= -1669389513;
assign addr[52817]= -1844288924;
assign addr[52818]= -1981813720;
assign addr[52819]= -2079176953;
assign addr[52820]= -2134405552;
assign addr[52821]= -2146380306;
assign addr[52822]= -2114858546;
assign addr[52823]= -2040479063;
assign addr[52824]= -1924749160;
assign addr[52825]= -1770014111;
assign addr[52826]= -1579409630;
assign addr[52827]= -1356798326;
assign addr[52828]= -1106691431;
assign addr[52829]= -834157373;
assign addr[52830]= -544719071;
assign addr[52831]= -244242007;
assign addr[52832]= 61184634;
assign addr[52833]= 365371365;
assign addr[52834]= 662153826;
assign addr[52835]= 945517704;
assign addr[52836]= 1209720613;
assign addr[52837]= 1449408469;
assign addr[52838]= 1659723983;
assign addr[52839]= 1836405100;
assign addr[52840]= 1975871368;
assign addr[52841]= 2075296495;
assign addr[52842]= 2132665626;
assign addr[52843]= 2146816171;
assign addr[52844]= 2117461370;
assign addr[52845]= 2045196100;
assign addr[52846]= 1931484818;
assign addr[52847]= 1778631892;
assign addr[52848]= 1589734894;
assign addr[52849]= 1368621831;
assign addr[52850]= 1119773573;
assign addr[52851]= 848233042;
assign addr[52852]= 559503022;
assign addr[52853]= 259434643;
assign addr[52854]= -45891193;
assign addr[52855]= -350287041;
assign addr[52856]= -647584304;
assign addr[52857]= -931758235;
assign addr[52858]= -1197050035;
assign addr[52859]= -1438083551;
assign addr[52860]= -1649974225;
assign addr[52861]= -1828428082;
assign addr[52862]= -1969828744;
assign addr[52863]= -2071310720;
assign addr[52864]= -2130817471;
assign addr[52865]= -2147143090;
assign addr[52866]= -2119956737;
assign addr[52867]= -2049809346;
assign addr[52868]= -1938122457;
assign addr[52869]= -1787159411;
assign addr[52870]= -1599979481;
assign addr[52871]= -1380375881;
assign addr[52872]= -1132798888;
assign addr[52873]= -862265664;
assign addr[52874]= -574258580;
assign addr[52875]= -274614114;
assign addr[52876]= 30595422;
assign addr[52877]= 335184940;
assign addr[52878]= 632981917;
assign addr[52879]= 917951481;
assign addr[52880]= 1184318708;
assign addr[52881]= 1426685652;
assign addr[52882]= 1640140734;
assign addr[52883]= 1820358275;
assign addr[52884]= 1963686155;
assign addr[52885]= 2067219829;
assign addr[52886]= 2128861181;
assign addr[52887]= 2147361045;
assign addr[52888]= 2122344521;
assign addr[52889]= 2054318569;
assign addr[52890]= 1944661739;
assign addr[52891]= 1795596234;
assign addr[52892]= 1610142873;
assign addr[52893]= 1392059879;
assign addr[52894]= 1145766716;
assign addr[52895]= 876254528;
assign addr[52896]= 588984994;
assign addr[52897]= 289779648;
assign addr[52898]= -15298099;
assign addr[52899]= -320065829;
assign addr[52900]= -618347408;
assign addr[52901]= -904098143;
assign addr[52902]= -1171527280;
assign addr[52903]= -1415215352;
assign addr[52904]= -1630224009;
assign addr[52905]= -1812196087;
assign addr[52906]= -1957443913;
assign addr[52907]= -2063024031;
assign addr[52908]= -2126796855;
assign addr[52909]= -2147470025;
assign addr[52910]= -2124624598;
assign addr[52911]= -2058723538;
assign addr[52912]= -1951102334;
assign addr[52913]= -1803941934;
assign addr[52914]= -1620224553;
assign addr[52915]= -1403673233;
assign addr[52916]= -1158676398;
assign addr[52917]= -890198924;
assign addr[52918]= -603681519;
assign addr[52919]= -304930476;
assign addr[52920]= 0;
assign addr[52921]= 304930476;
assign addr[52922]= 603681519;
assign addr[52923]= 890198924;
assign addr[52924]= 1158676398;
assign addr[52925]= 1403673233;
assign addr[52926]= 1620224553;
assign addr[52927]= 1803941934;
assign addr[52928]= 1951102334;
assign addr[52929]= 2058723538;
assign addr[52930]= 2124624598;
assign addr[52931]= 2147470025;
assign addr[52932]= 2126796855;
assign addr[52933]= 2063024031;
assign addr[52934]= 1957443913;
assign addr[52935]= 1812196087;
assign addr[52936]= 1630224009;
assign addr[52937]= 1415215352;
assign addr[52938]= 1171527280;
assign addr[52939]= 904098143;
assign addr[52940]= 618347408;
assign addr[52941]= 320065829;
assign addr[52942]= 15298099;
assign addr[52943]= -289779648;
assign addr[52944]= -588984994;
assign addr[52945]= -876254528;
assign addr[52946]= -1145766716;
assign addr[52947]= -1392059879;
assign addr[52948]= -1610142873;
assign addr[52949]= -1795596234;
assign addr[52950]= -1944661739;
assign addr[52951]= -2054318569;
assign addr[52952]= -2122344521;
assign addr[52953]= -2147361045;
assign addr[52954]= -2128861181;
assign addr[52955]= -2067219829;
assign addr[52956]= -1963686155;
assign addr[52957]= -1820358275;
assign addr[52958]= -1640140734;
assign addr[52959]= -1426685652;
assign addr[52960]= -1184318708;
assign addr[52961]= -917951481;
assign addr[52962]= -632981917;
assign addr[52963]= -335184940;
assign addr[52964]= -30595422;
assign addr[52965]= 274614114;
assign addr[52966]= 574258580;
assign addr[52967]= 862265664;
assign addr[52968]= 1132798888;
assign addr[52969]= 1380375881;
assign addr[52970]= 1599979481;
assign addr[52971]= 1787159411;
assign addr[52972]= 1938122457;
assign addr[52973]= 2049809346;
assign addr[52974]= 2119956737;
assign addr[52975]= 2147143090;
assign addr[52976]= 2130817471;
assign addr[52977]= 2071310720;
assign addr[52978]= 1969828744;
assign addr[52979]= 1828428082;
assign addr[52980]= 1649974225;
assign addr[52981]= 1438083551;
assign addr[52982]= 1197050035;
assign addr[52983]= 931758235;
assign addr[52984]= 647584304;
assign addr[52985]= 350287041;
assign addr[52986]= 45891193;
assign addr[52987]= -259434643;
assign addr[52988]= -559503022;
assign addr[52989]= -848233042;
assign addr[52990]= -1119773573;
assign addr[52991]= -1368621831;
assign addr[52992]= -1589734894;
assign addr[52993]= -1778631892;
assign addr[52994]= -1931484818;
assign addr[52995]= -2045196100;
assign addr[52996]= -2117461370;
assign addr[52997]= -2146816171;
assign addr[52998]= -2132665626;
assign addr[52999]= -2075296495;
assign addr[53000]= -1975871368;
assign addr[53001]= -1836405100;
assign addr[53002]= -1659723983;
assign addr[53003]= -1449408469;
assign addr[53004]= -1209720613;
assign addr[53005]= -945517704;
assign addr[53006]= -662153826;
assign addr[53007]= -365371365;
assign addr[53008]= -61184634;
assign addr[53009]= 244242007;
assign addr[53010]= 544719071;
assign addr[53011]= 834157373;
assign addr[53012]= 1106691431;
assign addr[53013]= 1356798326;
assign addr[53014]= 1579409630;
assign addr[53015]= 1770014111;
assign addr[53016]= 1924749160;
assign addr[53017]= 2040479063;
assign addr[53018]= 2114858546;
assign addr[53019]= 2146380306;
assign addr[53020]= 2134405552;
assign addr[53021]= 2079176953;
assign addr[53022]= 1981813720;
assign addr[53023]= 1844288924;
assign addr[53024]= 1669389513;
assign addr[53025]= 1460659832;
assign addr[53026]= 1222329801;
assign addr[53027]= 959229189;
assign addr[53028]= 676689746;
assign addr[53029]= 380437148;
assign addr[53030]= 76474970;
assign addr[53031]= -229036977;
assign addr[53032]= -529907477;
assign addr[53033]= -820039373;
assign addr[53034]= -1093553126;
assign addr[53035]= -1344905966;
assign addr[53036]= -1569004214;
assign addr[53037]= -1761306505;
assign addr[53038]= -1917915825;
assign addr[53039]= -2035658475;
assign addr[53040]= -2112148396;
assign addr[53041]= -2145835515;
assign addr[53042]= -2136037160;
assign addr[53043]= -2082951896;
assign addr[53044]= -1987655498;
assign addr[53045]= -1852079154;
assign addr[53046]= -1678970324;
assign addr[53047]= -1471837070;
assign addr[53048]= -1234876957;
assign addr[53049]= -972891995;
assign addr[53050]= -691191324;
assign addr[53051]= -395483624;
assign addr[53052]= -91761426;
assign addr[53053]= 213820322;
assign addr[53054]= 515068990;
assign addr[53055]= 805879757;
assign addr[53056]= 1080359326;
assign addr[53057]= 1332945355;
assign addr[53058]= 1558519173;
assign addr[53059]= 1752509516;
assign addr[53060]= 1910985158;
assign addr[53061]= 2030734582;
assign addr[53062]= 2109331059;
assign addr[53063]= 2145181827;
assign addr[53064]= 2137560369;
assign addr[53065]= 2086621133;
assign addr[53066]= 1993396407;
assign addr[53067]= 1859775393;
assign addr[53068]= 1688465931;
assign addr[53069]= 1482939614;
assign addr[53070]= 1247361445;
assign addr[53071]= 986505429;
assign addr[53072]= 705657826;
assign addr[53073]= 410510029;
assign addr[53074]= 107043224;
assign addr[53075]= -198592817;
assign addr[53076]= -500204365;
assign addr[53077]= -791679244;
assign addr[53078]= -1067110699;
assign addr[53079]= -1320917099;
assign addr[53080]= -1547955041;
assign addr[53081]= -1743623590;
assign addr[53082]= -1903957513;
assign addr[53083]= -2025707632;
assign addr[53084]= -2106406677;
assign addr[53085]= -2144419275;
assign addr[53086]= -2138975100;
assign addr[53087]= -2090184478;
assign addr[53088]= -1999036154;
assign addr[53089]= -1867377253;
assign addr[53090]= -1697875851;
assign addr[53091]= -1493966902;
assign addr[53092]= -1259782632;
assign addr[53093]= -1000068799;
assign addr[53094]= -720088517;
assign addr[53095]= -425515602;
assign addr[53096]= -122319591;
assign addr[53097]= 183355234;
assign addr[53098]= 485314355;
assign addr[53099]= 777438554;
assign addr[53100]= 1053807919;
assign addr[53101]= 1308821808;
assign addr[53102]= 1537312353;
assign addr[53103]= 1734649179;
assign addr[53104]= 1896833245;
assign addr[53105]= 2020577882;
assign addr[53106]= 2103375398;
assign addr[53107]= 2143547897;
assign addr[53108]= 2140281282;
assign addr[53109]= 2093641749;
assign addr[53110]= 2004574453;
assign addr[53111]= 1874884346;
assign addr[53112]= 1707199606;
assign addr[53113]= 1504918373;
assign addr[53114]= 1272139887;
assign addr[53115]= 1013581418;
assign addr[53116]= 734482665;
assign addr[53117]= 440499581;
assign addr[53118]= 137589750;
assign addr[53119]= -168108346;
assign addr[53120]= -470399716;
assign addr[53121]= -763158411;
assign addr[53122]= -1040451659;
assign addr[53123]= -1296660098;
assign addr[53124]= -1526591649;
assign addr[53125]= -1725586737;
assign addr[53126]= -1889612716;
assign addr[53127]= -2015345591;
assign addr[53128]= -2100237377;
assign addr[53129]= -2142567738;
assign addr[53130]= -2141478848;
assign addr[53131]= -2096992772;
assign addr[53132]= -2010011024;
assign addr[53133]= -1882296293;
assign addr[53134]= -1716436725;
assign addr[53135]= -1515793473;
assign addr[53136]= -1284432584;
assign addr[53137]= -1027042599;
assign addr[53138]= -748839539;
assign addr[53139]= -455461206;
assign addr[53140]= -152852926;
assign addr[53141]= 152852926;
assign addr[53142]= 455461206;
assign addr[53143]= 748839539;
assign addr[53144]= 1027042599;
assign addr[53145]= 1284432584;
assign addr[53146]= 1515793473;
assign addr[53147]= 1716436725;
assign addr[53148]= 1882296293;
assign addr[53149]= 2010011024;
assign addr[53150]= 2096992772;
assign addr[53151]= 2141478848;
assign addr[53152]= 2142567738;
assign addr[53153]= 2100237377;
assign addr[53154]= 2015345591;
assign addr[53155]= 1889612716;
assign addr[53156]= 1725586737;
assign addr[53157]= 1526591649;
assign addr[53158]= 1296660098;
assign addr[53159]= 1040451659;
assign addr[53160]= 763158411;
assign addr[53161]= 470399716;
assign addr[53162]= 168108346;
assign addr[53163]= -137589750;
assign addr[53164]= -440499581;
assign addr[53165]= -734482665;
assign addr[53166]= -1013581418;
assign addr[53167]= -1272139887;
assign addr[53168]= -1504918373;
assign addr[53169]= -1707199606;
assign addr[53170]= -1874884346;
assign addr[53171]= -2004574453;
assign addr[53172]= -2093641749;
assign addr[53173]= -2140281282;
assign addr[53174]= -2143547897;
assign addr[53175]= -2103375398;
assign addr[53176]= -2020577882;
assign addr[53177]= -1896833245;
assign addr[53178]= -1734649179;
assign addr[53179]= -1537312353;
assign addr[53180]= -1308821808;
assign addr[53181]= -1053807919;
assign addr[53182]= -777438554;
assign addr[53183]= -485314355;
assign addr[53184]= -183355234;
assign addr[53185]= 122319591;
assign addr[53186]= 425515602;
assign addr[53187]= 720088517;
assign addr[53188]= 1000068799;
assign addr[53189]= 1259782632;
assign addr[53190]= 1493966902;
assign addr[53191]= 1697875851;
assign addr[53192]= 1867377253;
assign addr[53193]= 1999036154;
assign addr[53194]= 2090184478;
assign addr[53195]= 2138975100;
assign addr[53196]= 2144419275;
assign addr[53197]= 2106406677;
assign addr[53198]= 2025707632;
assign addr[53199]= 1903957513;
assign addr[53200]= 1743623590;
assign addr[53201]= 1547955041;
assign addr[53202]= 1320917099;
assign addr[53203]= 1067110699;
assign addr[53204]= 791679244;
assign addr[53205]= 500204365;
assign addr[53206]= 198592817;
assign addr[53207]= -107043224;
assign addr[53208]= -410510029;
assign addr[53209]= -705657826;
assign addr[53210]= -986505429;
assign addr[53211]= -1247361445;
assign addr[53212]= -1482939614;
assign addr[53213]= -1688465931;
assign addr[53214]= -1859775393;
assign addr[53215]= -1993396407;
assign addr[53216]= -2086621133;
assign addr[53217]= -2137560369;
assign addr[53218]= -2145181827;
assign addr[53219]= -2109331059;
assign addr[53220]= -2030734582;
assign addr[53221]= -1910985158;
assign addr[53222]= -1752509516;
assign addr[53223]= -1558519173;
assign addr[53224]= -1332945355;
assign addr[53225]= -1080359326;
assign addr[53226]= -805879757;
assign addr[53227]= -515068990;
assign addr[53228]= -213820322;
assign addr[53229]= 91761426;
assign addr[53230]= 395483624;
assign addr[53231]= 691191324;
assign addr[53232]= 972891995;
assign addr[53233]= 1234876957;
assign addr[53234]= 1471837070;
assign addr[53235]= 1678970324;
assign addr[53236]= 1852079154;
assign addr[53237]= 1987655498;
assign addr[53238]= 2082951896;
assign addr[53239]= 2136037160;
assign addr[53240]= 2145835515;
assign addr[53241]= 2112148396;
assign addr[53242]= 2035658475;
assign addr[53243]= 1917915825;
assign addr[53244]= 1761306505;
assign addr[53245]= 1569004214;
assign addr[53246]= 1344905966;
assign addr[53247]= 1093553126;
assign addr[53248]= 820039373;
assign addr[53249]= 529907477;
assign addr[53250]= 229036977;
assign addr[53251]= -76474970;
assign addr[53252]= -380437148;
assign addr[53253]= -676689746;
assign addr[53254]= -959229189;
assign addr[53255]= -1222329801;
assign addr[53256]= -1460659832;
assign addr[53257]= -1669389513;
assign addr[53258]= -1844288924;
assign addr[53259]= -1981813720;
assign addr[53260]= -2079176953;
assign addr[53261]= -2134405552;
assign addr[53262]= -2146380306;
assign addr[53263]= -2114858546;
assign addr[53264]= -2040479063;
assign addr[53265]= -1924749160;
assign addr[53266]= -1770014111;
assign addr[53267]= -1579409630;
assign addr[53268]= -1356798326;
assign addr[53269]= -1106691431;
assign addr[53270]= -834157373;
assign addr[53271]= -544719071;
assign addr[53272]= -244242007;
assign addr[53273]= 61184634;
assign addr[53274]= 365371365;
assign addr[53275]= 662153826;
assign addr[53276]= 945517704;
assign addr[53277]= 1209720613;
assign addr[53278]= 1449408469;
assign addr[53279]= 1659723983;
assign addr[53280]= 1836405100;
assign addr[53281]= 1975871368;
assign addr[53282]= 2075296495;
assign addr[53283]= 2132665626;
assign addr[53284]= 2146816171;
assign addr[53285]= 2117461370;
assign addr[53286]= 2045196100;
assign addr[53287]= 1931484818;
assign addr[53288]= 1778631892;
assign addr[53289]= 1589734894;
assign addr[53290]= 1368621831;
assign addr[53291]= 1119773573;
assign addr[53292]= 848233042;
assign addr[53293]= 559503022;
assign addr[53294]= 259434643;
assign addr[53295]= -45891193;
assign addr[53296]= -350287041;
assign addr[53297]= -647584304;
assign addr[53298]= -931758235;
assign addr[53299]= -1197050035;
assign addr[53300]= -1438083551;
assign addr[53301]= -1649974225;
assign addr[53302]= -1828428082;
assign addr[53303]= -1969828744;
assign addr[53304]= -2071310720;
assign addr[53305]= -2130817471;
assign addr[53306]= -2147143090;
assign addr[53307]= -2119956737;
assign addr[53308]= -2049809346;
assign addr[53309]= -1938122457;
assign addr[53310]= -1787159411;
assign addr[53311]= -1599979481;
assign addr[53312]= -1380375881;
assign addr[53313]= -1132798888;
assign addr[53314]= -862265664;
assign addr[53315]= -574258580;
assign addr[53316]= -274614114;
assign addr[53317]= 30595422;
assign addr[53318]= 335184940;
assign addr[53319]= 632981917;
assign addr[53320]= 917951481;
assign addr[53321]= 1184318708;
assign addr[53322]= 1426685652;
assign addr[53323]= 1640140734;
assign addr[53324]= 1820358275;
assign addr[53325]= 1963686155;
assign addr[53326]= 2067219829;
assign addr[53327]= 2128861181;
assign addr[53328]= 2147361045;
assign addr[53329]= 2122344521;
assign addr[53330]= 2054318569;
assign addr[53331]= 1944661739;
assign addr[53332]= 1795596234;
assign addr[53333]= 1610142873;
assign addr[53334]= 1392059879;
assign addr[53335]= 1145766716;
assign addr[53336]= 876254528;
assign addr[53337]= 588984994;
assign addr[53338]= 289779648;
assign addr[53339]= -15298099;
assign addr[53340]= -320065829;
assign addr[53341]= -618347408;
assign addr[53342]= -904098143;
assign addr[53343]= -1171527280;
assign addr[53344]= -1415215352;
assign addr[53345]= -1630224009;
assign addr[53346]= -1812196087;
assign addr[53347]= -1957443913;
assign addr[53348]= -2063024031;
assign addr[53349]= -2126796855;
assign addr[53350]= -2147470025;
assign addr[53351]= -2124624598;
assign addr[53352]= -2058723538;
assign addr[53353]= -1951102334;
assign addr[53354]= -1803941934;
assign addr[53355]= -1620224553;
assign addr[53356]= -1403673233;
assign addr[53357]= -1158676398;
assign addr[53358]= -890198924;
assign addr[53359]= -603681519;
assign addr[53360]= -304930476;
assign addr[53361]= 0;
assign addr[53362]= 304930476;
assign addr[53363]= 603681519;
assign addr[53364]= 890198924;
assign addr[53365]= 1158676398;
assign addr[53366]= 1403673233;
assign addr[53367]= 1620224553;
assign addr[53368]= 1803941934;
assign addr[53369]= 1951102334;
assign addr[53370]= 2058723538;
assign addr[53371]= 2124624598;
assign addr[53372]= 2147470025;
assign addr[53373]= 2126796855;
assign addr[53374]= 2063024031;
assign addr[53375]= 1957443913;
assign addr[53376]= 1812196087;
assign addr[53377]= 1630224009;
assign addr[53378]= 1415215352;
assign addr[53379]= 1171527280;
assign addr[53380]= 904098143;
assign addr[53381]= 618347408;
assign addr[53382]= 320065829;
assign addr[53383]= 15298099;
assign addr[53384]= -289779648;
assign addr[53385]= -588984994;
assign addr[53386]= -876254528;
assign addr[53387]= -1145766716;
assign addr[53388]= -1392059879;
assign addr[53389]= -1610142873;
assign addr[53390]= -1795596234;
assign addr[53391]= -1944661739;
assign addr[53392]= -2054318569;
assign addr[53393]= -2122344521;
assign addr[53394]= -2147361045;
assign addr[53395]= -2128861181;
assign addr[53396]= -2067219829;
assign addr[53397]= -1963686155;
assign addr[53398]= -1820358275;
assign addr[53399]= -1640140734;
assign addr[53400]= -1426685652;
assign addr[53401]= -1184318708;
assign addr[53402]= -917951481;
assign addr[53403]= -632981917;
assign addr[53404]= -335184940;
assign addr[53405]= -30595422;
assign addr[53406]= 274614114;
assign addr[53407]= 574258580;
assign addr[53408]= 862265664;
assign addr[53409]= 1132798888;
assign addr[53410]= 1380375881;
assign addr[53411]= 1599979481;
assign addr[53412]= 1787159411;
assign addr[53413]= 1938122457;
assign addr[53414]= 2049809346;
assign addr[53415]= 2119956737;
assign addr[53416]= 2147143090;
assign addr[53417]= 2130817471;
assign addr[53418]= 2071310720;
assign addr[53419]= 1969828744;
assign addr[53420]= 1828428082;
assign addr[53421]= 1649974225;
assign addr[53422]= 1438083551;
assign addr[53423]= 1197050035;
assign addr[53424]= 931758235;
assign addr[53425]= 647584304;
assign addr[53426]= 350287041;
assign addr[53427]= 45891193;
assign addr[53428]= -259434643;
assign addr[53429]= -559503022;
assign addr[53430]= -848233042;
assign addr[53431]= -1119773573;
assign addr[53432]= -1368621831;
assign addr[53433]= -1589734894;
assign addr[53434]= -1778631892;
assign addr[53435]= -1931484818;
assign addr[53436]= -2045196100;
assign addr[53437]= -2117461370;
assign addr[53438]= -2146816171;
assign addr[53439]= -2132665626;
assign addr[53440]= -2075296495;
assign addr[53441]= -1975871368;
assign addr[53442]= -1836405100;
assign addr[53443]= -1659723983;
assign addr[53444]= -1449408469;
assign addr[53445]= -1209720613;
assign addr[53446]= -945517704;
assign addr[53447]= -662153826;
assign addr[53448]= -365371365;
assign addr[53449]= -61184634;
assign addr[53450]= 244242007;
assign addr[53451]= 544719071;
assign addr[53452]= 834157373;
assign addr[53453]= 1106691431;
assign addr[53454]= 1356798326;
assign addr[53455]= 1579409630;
assign addr[53456]= 1770014111;
assign addr[53457]= 1924749160;
assign addr[53458]= 2040479063;
assign addr[53459]= 2114858546;
assign addr[53460]= 2146380306;
assign addr[53461]= 2134405552;
assign addr[53462]= 2079176953;
assign addr[53463]= 1981813720;
assign addr[53464]= 1844288924;
assign addr[53465]= 1669389513;
assign addr[53466]= 1460659832;
assign addr[53467]= 1222329801;
assign addr[53468]= 959229189;
assign addr[53469]= 676689746;
assign addr[53470]= 380437148;
assign addr[53471]= 76474970;
assign addr[53472]= -229036977;
assign addr[53473]= -529907477;
assign addr[53474]= -820039373;
assign addr[53475]= -1093553126;
assign addr[53476]= -1344905966;
assign addr[53477]= -1569004214;
assign addr[53478]= -1761306505;
assign addr[53479]= -1917915825;
assign addr[53480]= -2035658475;
assign addr[53481]= -2112148396;
assign addr[53482]= -2145835515;
assign addr[53483]= -2136037160;
assign addr[53484]= -2082951896;
assign addr[53485]= -1987655498;
assign addr[53486]= -1852079154;
assign addr[53487]= -1678970324;
assign addr[53488]= -1471837070;
assign addr[53489]= -1234876957;
assign addr[53490]= -972891995;
assign addr[53491]= -691191324;
assign addr[53492]= -395483624;
assign addr[53493]= -91761426;
assign addr[53494]= 213820322;
assign addr[53495]= 515068990;
assign addr[53496]= 805879757;
assign addr[53497]= 1080359326;
assign addr[53498]= 1332945355;
assign addr[53499]= 1558519173;
assign addr[53500]= 1752509516;
assign addr[53501]= 1910985158;
assign addr[53502]= 2030734582;
assign addr[53503]= 2109331059;
assign addr[53504]= 2145181827;
assign addr[53505]= 2137560369;
assign addr[53506]= 2086621133;
assign addr[53507]= 1993396407;
assign addr[53508]= 1859775393;
assign addr[53509]= 1688465931;
assign addr[53510]= 1482939614;
assign addr[53511]= 1247361445;
assign addr[53512]= 986505429;
assign addr[53513]= 705657826;
assign addr[53514]= 410510029;
assign addr[53515]= 107043224;
assign addr[53516]= -198592817;
assign addr[53517]= -500204365;
assign addr[53518]= -791679244;
assign addr[53519]= -1067110699;
assign addr[53520]= -1320917099;
assign addr[53521]= -1547955041;
assign addr[53522]= -1743623590;
assign addr[53523]= -1903957513;
assign addr[53524]= -2025707632;
assign addr[53525]= -2106406677;
assign addr[53526]= -2144419275;
assign addr[53527]= -2138975100;
assign addr[53528]= -2090184478;
assign addr[53529]= -1999036154;
assign addr[53530]= -1867377253;
assign addr[53531]= -1697875851;
assign addr[53532]= -1493966902;
assign addr[53533]= -1259782632;
assign addr[53534]= -1000068799;
assign addr[53535]= -720088517;
assign addr[53536]= -425515602;
assign addr[53537]= -122319591;
assign addr[53538]= 183355234;
assign addr[53539]= 485314355;
assign addr[53540]= 777438554;
assign addr[53541]= 1053807919;
assign addr[53542]= 1308821808;
assign addr[53543]= 1537312353;
assign addr[53544]= 1734649179;
assign addr[53545]= 1896833245;
assign addr[53546]= 2020577882;
assign addr[53547]= 2103375398;
assign addr[53548]= 2143547897;
assign addr[53549]= 2140281282;
assign addr[53550]= 2093641749;
assign addr[53551]= 2004574453;
assign addr[53552]= 1874884346;
assign addr[53553]= 1707199606;
assign addr[53554]= 1504918373;
assign addr[53555]= 1272139887;
assign addr[53556]= 1013581418;
assign addr[53557]= 734482665;
assign addr[53558]= 440499581;
assign addr[53559]= 137589750;
assign addr[53560]= -168108346;
assign addr[53561]= -470399716;
assign addr[53562]= -763158411;
assign addr[53563]= -1040451659;
assign addr[53564]= -1296660098;
assign addr[53565]= -1526591649;
assign addr[53566]= -1725586737;
assign addr[53567]= -1889612716;
assign addr[53568]= -2015345591;
assign addr[53569]= -2100237377;
assign addr[53570]= -2142567738;
assign addr[53571]= -2141478848;
assign addr[53572]= -2096992772;
assign addr[53573]= -2010011024;
assign addr[53574]= -1882296293;
assign addr[53575]= -1716436725;
assign addr[53576]= -1515793473;
assign addr[53577]= -1284432584;
assign addr[53578]= -1027042599;
assign addr[53579]= -748839539;
assign addr[53580]= -455461206;
assign addr[53581]= -152852926;
assign addr[53582]= 152852926;
assign addr[53583]= 455461206;
assign addr[53584]= 748839539;
assign addr[53585]= 1027042599;
assign addr[53586]= 1284432584;
assign addr[53587]= 1515793473;
assign addr[53588]= 1716436725;
assign addr[53589]= 1882296293;
assign addr[53590]= 2010011024;
assign addr[53591]= 2096992772;
assign addr[53592]= 2141478848;
assign addr[53593]= 2142567738;
assign addr[53594]= 2100237377;
assign addr[53595]= 2015345591;
assign addr[53596]= 1889612716;
assign addr[53597]= 1725586737;
assign addr[53598]= 1526591649;
assign addr[53599]= 1296660098;
assign addr[53600]= 1040451659;
assign addr[53601]= 763158411;
assign addr[53602]= 470399716;
assign addr[53603]= 168108346;
assign addr[53604]= -137589750;
assign addr[53605]= -440499581;
assign addr[53606]= -734482665;
assign addr[53607]= -1013581418;
assign addr[53608]= -1272139887;
assign addr[53609]= -1504918373;
assign addr[53610]= -1707199606;
assign addr[53611]= -1874884346;
assign addr[53612]= -2004574453;
assign addr[53613]= -2093641749;
assign addr[53614]= -2140281282;
assign addr[53615]= -2143547897;
assign addr[53616]= -2103375398;
assign addr[53617]= -2020577882;
assign addr[53618]= -1896833245;
assign addr[53619]= -1734649179;
assign addr[53620]= -1537312353;
assign addr[53621]= -1308821808;
assign addr[53622]= -1053807919;
assign addr[53623]= -777438554;
assign addr[53624]= -485314355;
assign addr[53625]= -183355234;
assign addr[53626]= 122319591;
assign addr[53627]= 425515602;
assign addr[53628]= 720088517;
assign addr[53629]= 1000068799;
assign addr[53630]= 1259782632;
assign addr[53631]= 1493966902;
assign addr[53632]= 1697875851;
assign addr[53633]= 1867377253;
assign addr[53634]= 1999036154;
assign addr[53635]= 2090184478;
assign addr[53636]= 2138975100;
assign addr[53637]= 2144419275;
assign addr[53638]= 2106406677;
assign addr[53639]= 2025707632;
assign addr[53640]= 1903957513;
assign addr[53641]= 1743623590;
assign addr[53642]= 1547955041;
assign addr[53643]= 1320917099;
assign addr[53644]= 1067110699;
assign addr[53645]= 791679244;
assign addr[53646]= 500204365;
assign addr[53647]= 198592817;
assign addr[53648]= -107043224;
assign addr[53649]= -410510029;
assign addr[53650]= -705657826;
assign addr[53651]= -986505429;
assign addr[53652]= -1247361445;
assign addr[53653]= -1482939614;
assign addr[53654]= -1688465931;
assign addr[53655]= -1859775393;
assign addr[53656]= -1993396407;
assign addr[53657]= -2086621133;
assign addr[53658]= -2137560369;
assign addr[53659]= -2145181827;
assign addr[53660]= -2109331059;
assign addr[53661]= -2030734582;
assign addr[53662]= -1910985158;
assign addr[53663]= -1752509516;
assign addr[53664]= -1558519173;
assign addr[53665]= -1332945355;
assign addr[53666]= -1080359326;
assign addr[53667]= -805879757;
assign addr[53668]= -515068990;
assign addr[53669]= -213820322;
assign addr[53670]= 91761426;
assign addr[53671]= 395483624;
assign addr[53672]= 691191324;
assign addr[53673]= 972891995;
assign addr[53674]= 1234876957;
assign addr[53675]= 1471837070;
assign addr[53676]= 1678970324;
assign addr[53677]= 1852079154;
assign addr[53678]= 1987655498;
assign addr[53679]= 2082951896;
assign addr[53680]= 2136037160;
assign addr[53681]= 2145835515;
assign addr[53682]= 2112148396;
assign addr[53683]= 2035658475;
assign addr[53684]= 1917915825;
assign addr[53685]= 1761306505;
assign addr[53686]= 1569004214;
assign addr[53687]= 1344905966;
assign addr[53688]= 1093553126;
assign addr[53689]= 820039373;
assign addr[53690]= 529907477;
assign addr[53691]= 229036977;
assign addr[53692]= -76474970;
assign addr[53693]= -380437148;
assign addr[53694]= -676689746;
assign addr[53695]= -959229189;
assign addr[53696]= -1222329801;
assign addr[53697]= -1460659832;
assign addr[53698]= -1669389513;
assign addr[53699]= -1844288924;
assign addr[53700]= -1981813720;
assign addr[53701]= -2079176953;
assign addr[53702]= -2134405552;
assign addr[53703]= -2146380306;
assign addr[53704]= -2114858546;
assign addr[53705]= -2040479063;
assign addr[53706]= -1924749160;
assign addr[53707]= -1770014111;
assign addr[53708]= -1579409630;
assign addr[53709]= -1356798326;
assign addr[53710]= -1106691431;
assign addr[53711]= -834157373;
assign addr[53712]= -544719071;
assign addr[53713]= -244242007;
assign addr[53714]= 61184634;
assign addr[53715]= 365371365;
assign addr[53716]= 662153826;
assign addr[53717]= 945517704;
assign addr[53718]= 1209720613;
assign addr[53719]= 1449408469;
assign addr[53720]= 1659723983;
assign addr[53721]= 1836405100;
assign addr[53722]= 1975871368;
assign addr[53723]= 2075296495;
assign addr[53724]= 2132665626;
assign addr[53725]= 2146816171;
assign addr[53726]= 2117461370;
assign addr[53727]= 2045196100;
assign addr[53728]= 1931484818;
assign addr[53729]= 1778631892;
assign addr[53730]= 1589734894;
assign addr[53731]= 1368621831;
assign addr[53732]= 1119773573;
assign addr[53733]= 848233042;
assign addr[53734]= 559503022;
assign addr[53735]= 259434643;
assign addr[53736]= -45891193;
assign addr[53737]= -350287041;
assign addr[53738]= -647584304;
assign addr[53739]= -931758235;
assign addr[53740]= -1197050035;
assign addr[53741]= -1438083551;
assign addr[53742]= -1649974225;
assign addr[53743]= -1828428082;
assign addr[53744]= -1969828744;
assign addr[53745]= -2071310720;
assign addr[53746]= -2130817471;
assign addr[53747]= -2147143090;
assign addr[53748]= -2119956737;
assign addr[53749]= -2049809346;
assign addr[53750]= -1938122457;
assign addr[53751]= -1787159411;
assign addr[53752]= -1599979481;
assign addr[53753]= -1380375881;
assign addr[53754]= -1132798888;
assign addr[53755]= -862265664;
assign addr[53756]= -574258580;
assign addr[53757]= -274614114;
assign addr[53758]= 30595422;
assign addr[53759]= 335184940;
assign addr[53760]= 632981917;
assign addr[53761]= 917951481;
assign addr[53762]= 1184318708;
assign addr[53763]= 1426685652;
assign addr[53764]= 1640140734;
assign addr[53765]= 1820358275;
assign addr[53766]= 1963686155;
assign addr[53767]= 2067219829;
assign addr[53768]= 2128861181;
assign addr[53769]= 2147361045;
assign addr[53770]= 2122344521;
assign addr[53771]= 2054318569;
assign addr[53772]= 1944661739;
assign addr[53773]= 1795596234;
assign addr[53774]= 1610142873;
assign addr[53775]= 1392059879;
assign addr[53776]= 1145766716;
assign addr[53777]= 876254528;
assign addr[53778]= 588984994;
assign addr[53779]= 289779648;
assign addr[53780]= -15298099;
assign addr[53781]= -320065829;
assign addr[53782]= -618347408;
assign addr[53783]= -904098143;
assign addr[53784]= -1171527280;
assign addr[53785]= -1415215352;
assign addr[53786]= -1630224009;
assign addr[53787]= -1812196087;
assign addr[53788]= -1957443913;
assign addr[53789]= -2063024031;
assign addr[53790]= -2126796855;
assign addr[53791]= -2147470025;
assign addr[53792]= -2124624598;
assign addr[53793]= -2058723538;
assign addr[53794]= -1951102334;
assign addr[53795]= -1803941934;
assign addr[53796]= -1620224553;
assign addr[53797]= -1403673233;
assign addr[53798]= -1158676398;
assign addr[53799]= -890198924;
assign addr[53800]= -603681519;
assign addr[53801]= -304930476;
assign addr[53802]= 0;
assign addr[53803]= 304930476;
assign addr[53804]= 603681519;
assign addr[53805]= 890198924;
assign addr[53806]= 1158676398;
assign addr[53807]= 1403673233;
assign addr[53808]= 1620224553;
assign addr[53809]= 1803941934;
assign addr[53810]= 1951102334;
assign addr[53811]= 2058723538;
assign addr[53812]= 2124624598;
assign addr[53813]= 2147470025;
assign addr[53814]= 2126796855;
assign addr[53815]= 2063024031;
assign addr[53816]= 1957443913;
assign addr[53817]= 1812196087;
assign addr[53818]= 1630224009;
assign addr[53819]= 1415215352;
assign addr[53820]= 1171527280;
assign addr[53821]= 904098143;
assign addr[53822]= 618347408;
assign addr[53823]= 320065829;
assign addr[53824]= 15298099;
assign addr[53825]= -289779648;
assign addr[53826]= -588984994;
assign addr[53827]= -876254528;
assign addr[53828]= -1145766716;
assign addr[53829]= -1392059879;
assign addr[53830]= -1610142873;
assign addr[53831]= -1795596234;
assign addr[53832]= -1944661739;
assign addr[53833]= -2054318569;
assign addr[53834]= -2122344521;
assign addr[53835]= -2147361045;
assign addr[53836]= -2128861181;
assign addr[53837]= -2067219829;
assign addr[53838]= -1963686155;
assign addr[53839]= -1820358275;
assign addr[53840]= -1640140734;
assign addr[53841]= -1426685652;
assign addr[53842]= -1184318708;
assign addr[53843]= -917951481;
assign addr[53844]= -632981917;
assign addr[53845]= -335184940;
assign addr[53846]= -30595422;
assign addr[53847]= 274614114;
assign addr[53848]= 574258580;
assign addr[53849]= 862265664;
assign addr[53850]= 1132798888;
assign addr[53851]= 1380375881;
assign addr[53852]= 1599979481;
assign addr[53853]= 1787159411;
assign addr[53854]= 1938122457;
assign addr[53855]= 2049809346;
assign addr[53856]= 2119956737;
assign addr[53857]= 2147143090;
assign addr[53858]= 2130817471;
assign addr[53859]= 2071310720;
assign addr[53860]= 1969828744;
assign addr[53861]= 1828428082;
assign addr[53862]= 1649974225;
assign addr[53863]= 1438083551;
assign addr[53864]= 1197050035;
assign addr[53865]= 931758235;
assign addr[53866]= 647584304;
assign addr[53867]= 350287041;
assign addr[53868]= 45891193;
assign addr[53869]= -259434643;
assign addr[53870]= -559503022;
assign addr[53871]= -848233042;
assign addr[53872]= -1119773573;
assign addr[53873]= -1368621831;
assign addr[53874]= -1589734894;
assign addr[53875]= -1778631892;
assign addr[53876]= -1931484818;
assign addr[53877]= -2045196100;
assign addr[53878]= -2117461370;
assign addr[53879]= -2146816171;
assign addr[53880]= -2132665626;
assign addr[53881]= -2075296495;
assign addr[53882]= -1975871368;
assign addr[53883]= -1836405100;
assign addr[53884]= -1659723983;
assign addr[53885]= -1449408469;
assign addr[53886]= -1209720613;
assign addr[53887]= -945517704;
assign addr[53888]= -662153826;
assign addr[53889]= -365371365;
assign addr[53890]= -61184634;
assign addr[53891]= 244242007;
assign addr[53892]= 544719071;
assign addr[53893]= 834157373;
assign addr[53894]= 1106691431;
assign addr[53895]= 1356798326;
assign addr[53896]= 1579409630;
assign addr[53897]= 1770014111;
assign addr[53898]= 1924749160;
assign addr[53899]= 2040479063;
assign addr[53900]= 2114858546;
assign addr[53901]= 2146380306;
assign addr[53902]= 2134405552;
assign addr[53903]= 2079176953;
assign addr[53904]= 1981813720;
assign addr[53905]= 1844288924;
assign addr[53906]= 1669389513;
assign addr[53907]= 1460659832;
assign addr[53908]= 1222329801;
assign addr[53909]= 959229189;
assign addr[53910]= 676689746;
assign addr[53911]= 380437148;
assign addr[53912]= 76474970;
assign addr[53913]= -229036977;
assign addr[53914]= -529907477;
assign addr[53915]= -820039373;
assign addr[53916]= -1093553126;
assign addr[53917]= -1344905966;
assign addr[53918]= -1569004214;
assign addr[53919]= -1761306505;
assign addr[53920]= -1917915825;
assign addr[53921]= -2035658475;
assign addr[53922]= -2112148396;
assign addr[53923]= -2145835515;
assign addr[53924]= -2136037160;
assign addr[53925]= -2082951896;
assign addr[53926]= -1987655498;
assign addr[53927]= -1852079154;
assign addr[53928]= -1678970324;
assign addr[53929]= -1471837070;
assign addr[53930]= -1234876957;
assign addr[53931]= -972891995;
assign addr[53932]= -691191324;
assign addr[53933]= -395483624;
assign addr[53934]= -91761426;
assign addr[53935]= 213820322;
assign addr[53936]= 515068990;
assign addr[53937]= 805879757;
assign addr[53938]= 1080359326;
assign addr[53939]= 1332945355;
assign addr[53940]= 1558519173;
assign addr[53941]= 1752509516;
assign addr[53942]= 1910985158;
assign addr[53943]= 2030734582;
assign addr[53944]= 2109331059;
assign addr[53945]= 2145181827;
assign addr[53946]= 2137560369;
assign addr[53947]= 2086621133;
assign addr[53948]= 1993396407;
assign addr[53949]= 1859775393;
assign addr[53950]= 1688465931;
assign addr[53951]= 1482939614;
assign addr[53952]= 1247361445;
assign addr[53953]= 986505429;
assign addr[53954]= 705657826;
assign addr[53955]= 410510029;
assign addr[53956]= 107043224;
assign addr[53957]= -198592817;
assign addr[53958]= -500204365;
assign addr[53959]= -791679244;
assign addr[53960]= -1067110699;
assign addr[53961]= -1320917099;
assign addr[53962]= -1547955041;
assign addr[53963]= -1743623590;
assign addr[53964]= -1903957513;
assign addr[53965]= -2025707632;
assign addr[53966]= -2106406677;
assign addr[53967]= -2144419275;
assign addr[53968]= -2138975100;
assign addr[53969]= -2090184478;
assign addr[53970]= -1999036154;
assign addr[53971]= -1867377253;
assign addr[53972]= -1697875851;
assign addr[53973]= -1493966902;
assign addr[53974]= -1259782632;
assign addr[53975]= -1000068799;
assign addr[53976]= -720088517;
assign addr[53977]= -425515602;
assign addr[53978]= -122319591;
assign addr[53979]= 183355234;
assign addr[53980]= 485314355;
assign addr[53981]= 777438554;
assign addr[53982]= 1053807919;
assign addr[53983]= 1308821808;
assign addr[53984]= 1537312353;
assign addr[53985]= 1734649179;
assign addr[53986]= 1896833245;
assign addr[53987]= 2020577882;
assign addr[53988]= 2103375398;
assign addr[53989]= 2143547897;
assign addr[53990]= 2140281282;
assign addr[53991]= 2093641749;
assign addr[53992]= 2004574453;
assign addr[53993]= 1874884346;
assign addr[53994]= 1707199606;
assign addr[53995]= 1504918373;
assign addr[53996]= 1272139887;
assign addr[53997]= 1013581418;
assign addr[53998]= 734482665;
assign addr[53999]= 440499581;
assign addr[54000]= 137589750;
assign addr[54001]= -168108346;
assign addr[54002]= -470399716;
assign addr[54003]= -763158411;
assign addr[54004]= -1040451659;
assign addr[54005]= -1296660098;
assign addr[54006]= -1526591649;
assign addr[54007]= -1725586737;
assign addr[54008]= -1889612716;
assign addr[54009]= -2015345591;
assign addr[54010]= -2100237377;
assign addr[54011]= -2142567738;
assign addr[54012]= -2141478848;
assign addr[54013]= -2096992772;
assign addr[54014]= -2010011024;
assign addr[54015]= -1882296293;
assign addr[54016]= -1716436725;
assign addr[54017]= -1515793473;
assign addr[54018]= -1284432584;
assign addr[54019]= -1027042599;
assign addr[54020]= -748839539;
assign addr[54021]= -455461206;
assign addr[54022]= -152852926;
assign addr[54023]= 152852926;
assign addr[54024]= 455461206;
assign addr[54025]= 748839539;
assign addr[54026]= 1027042599;
assign addr[54027]= 1284432584;
assign addr[54028]= 1515793473;
assign addr[54029]= 1716436725;
assign addr[54030]= 1882296293;
assign addr[54031]= 2010011024;
assign addr[54032]= 2096992772;
assign addr[54033]= 2141478848;
assign addr[54034]= 2142567738;
assign addr[54035]= 2100237377;
assign addr[54036]= 2015345591;
assign addr[54037]= 1889612716;
assign addr[54038]= 1725586737;
assign addr[54039]= 1526591649;
assign addr[54040]= 1296660098;
assign addr[54041]= 1040451659;
assign addr[54042]= 763158411;
assign addr[54043]= 470399716;
assign addr[54044]= 168108346;
assign addr[54045]= -137589750;
assign addr[54046]= -440499581;
assign addr[54047]= -734482665;
assign addr[54048]= -1013581418;
assign addr[54049]= -1272139887;
assign addr[54050]= -1504918373;
assign addr[54051]= -1707199606;
assign addr[54052]= -1874884346;
assign addr[54053]= -2004574453;
assign addr[54054]= -2093641749;
assign addr[54055]= -2140281282;
assign addr[54056]= -2143547897;
assign addr[54057]= -2103375398;
assign addr[54058]= -2020577882;
assign addr[54059]= -1896833245;
assign addr[54060]= -1734649179;
assign addr[54061]= -1537312353;
assign addr[54062]= -1308821808;
assign addr[54063]= -1053807919;
assign addr[54064]= -777438554;
assign addr[54065]= -485314355;
assign addr[54066]= -183355234;
assign addr[54067]= 122319591;
assign addr[54068]= 425515602;
assign addr[54069]= 720088517;
assign addr[54070]= 1000068799;
assign addr[54071]= 1259782632;
assign addr[54072]= 1493966902;
assign addr[54073]= 1697875851;
assign addr[54074]= 1867377253;
assign addr[54075]= 1999036154;
assign addr[54076]= 2090184478;
assign addr[54077]= 2138975100;
assign addr[54078]= 2144419275;
assign addr[54079]= 2106406677;
assign addr[54080]= 2025707632;
assign addr[54081]= 1903957513;
assign addr[54082]= 1743623590;
assign addr[54083]= 1547955041;
assign addr[54084]= 1320917099;
assign addr[54085]= 1067110699;
assign addr[54086]= 791679244;
assign addr[54087]= 500204365;
assign addr[54088]= 198592817;
assign addr[54089]= -107043224;
assign addr[54090]= -410510029;
assign addr[54091]= -705657826;
assign addr[54092]= -986505429;
assign addr[54093]= -1247361445;
assign addr[54094]= -1482939614;
assign addr[54095]= -1688465931;
assign addr[54096]= -1859775393;
assign addr[54097]= -1993396407;
assign addr[54098]= -2086621133;
assign addr[54099]= -2137560369;
assign addr[54100]= -2145181827;
assign addr[54101]= -2109331059;
assign addr[54102]= -2030734582;
assign addr[54103]= -1910985158;
assign addr[54104]= -1752509516;
assign addr[54105]= -1558519173;
assign addr[54106]= -1332945355;
assign addr[54107]= -1080359326;
assign addr[54108]= -805879757;
assign addr[54109]= -515068990;
assign addr[54110]= -213820322;
assign addr[54111]= 91761426;
assign addr[54112]= 395483624;
assign addr[54113]= 691191324;
assign addr[54114]= 972891995;
assign addr[54115]= 1234876957;
assign addr[54116]= 1471837070;
assign addr[54117]= 1678970324;
assign addr[54118]= 1852079154;
assign addr[54119]= 1987655498;
assign addr[54120]= 2082951896;
assign addr[54121]= 2136037160;
assign addr[54122]= 2145835515;
assign addr[54123]= 2112148396;
assign addr[54124]= 2035658475;
assign addr[54125]= 1917915825;
assign addr[54126]= 1761306505;
assign addr[54127]= 1569004214;
assign addr[54128]= 1344905966;
assign addr[54129]= 1093553126;
assign addr[54130]= 820039373;
assign addr[54131]= 529907477;
assign addr[54132]= 229036977;
assign addr[54133]= -76474970;
assign addr[54134]= -380437148;
assign addr[54135]= -676689746;
assign addr[54136]= -959229189;
assign addr[54137]= -1222329801;
assign addr[54138]= -1460659832;
assign addr[54139]= -1669389513;
assign addr[54140]= -1844288924;
assign addr[54141]= -1981813720;
assign addr[54142]= -2079176953;
assign addr[54143]= -2134405552;
assign addr[54144]= -2146380306;
assign addr[54145]= -2114858546;
assign addr[54146]= -2040479063;
assign addr[54147]= -1924749160;
assign addr[54148]= -1770014111;
assign addr[54149]= -1579409630;
assign addr[54150]= -1356798326;
assign addr[54151]= -1106691431;
assign addr[54152]= -834157373;
assign addr[54153]= -544719071;
assign addr[54154]= -244242007;
assign addr[54155]= 61184634;
assign addr[54156]= 365371365;
assign addr[54157]= 662153826;
assign addr[54158]= 945517704;
assign addr[54159]= 1209720613;
assign addr[54160]= 1449408469;
assign addr[54161]= 1659723983;
assign addr[54162]= 1836405100;
assign addr[54163]= 1975871368;
assign addr[54164]= 2075296495;
assign addr[54165]= 2132665626;
assign addr[54166]= 2146816171;
assign addr[54167]= 2117461370;
assign addr[54168]= 2045196100;
assign addr[54169]= 1931484818;
assign addr[54170]= 1778631892;
assign addr[54171]= 1589734894;
assign addr[54172]= 1368621831;
assign addr[54173]= 1119773573;
assign addr[54174]= 848233042;
assign addr[54175]= 559503022;
assign addr[54176]= 259434643;
assign addr[54177]= -45891193;
assign addr[54178]= -350287041;
assign addr[54179]= -647584304;
assign addr[54180]= -931758235;
assign addr[54181]= -1197050035;
assign addr[54182]= -1438083551;
assign addr[54183]= -1649974225;
assign addr[54184]= -1828428082;
assign addr[54185]= -1969828744;
assign addr[54186]= -2071310720;
assign addr[54187]= -2130817471;
assign addr[54188]= -2147143090;
assign addr[54189]= -2119956737;
assign addr[54190]= -2049809346;
assign addr[54191]= -1938122457;
assign addr[54192]= -1787159411;
assign addr[54193]= -1599979481;
assign addr[54194]= -1380375881;
assign addr[54195]= -1132798888;
assign addr[54196]= -862265664;
assign addr[54197]= -574258580;
assign addr[54198]= -274614114;
assign addr[54199]= 30595422;
assign addr[54200]= 335184940;
assign addr[54201]= 632981917;
assign addr[54202]= 917951481;
assign addr[54203]= 1184318708;
assign addr[54204]= 1426685652;
assign addr[54205]= 1640140734;
assign addr[54206]= 1820358275;
assign addr[54207]= 1963686155;
assign addr[54208]= 2067219829;
assign addr[54209]= 2128861181;
assign addr[54210]= 2147361045;
assign addr[54211]= 2122344521;
assign addr[54212]= 2054318569;
assign addr[54213]= 1944661739;
assign addr[54214]= 1795596234;
assign addr[54215]= 1610142873;
assign addr[54216]= 1392059879;
assign addr[54217]= 1145766716;
assign addr[54218]= 876254528;
assign addr[54219]= 588984994;
assign addr[54220]= 289779648;
assign addr[54221]= -15298099;
assign addr[54222]= -320065829;
assign addr[54223]= -618347408;
assign addr[54224]= -904098143;
assign addr[54225]= -1171527280;
assign addr[54226]= -1415215352;
assign addr[54227]= -1630224009;
assign addr[54228]= -1812196087;
assign addr[54229]= -1957443913;
assign addr[54230]= -2063024031;
assign addr[54231]= -2126796855;
assign addr[54232]= -2147470025;
assign addr[54233]= -2124624598;
assign addr[54234]= -2058723538;
assign addr[54235]= -1951102334;
assign addr[54236]= -1803941934;
assign addr[54237]= -1620224553;
assign addr[54238]= -1403673233;
assign addr[54239]= -1158676398;
assign addr[54240]= -890198924;
assign addr[54241]= -603681519;
assign addr[54242]= -304930476;
assign addr[54243]= 0;
assign addr[54244]= 304930476;
assign addr[54245]= 603681519;
assign addr[54246]= 890198924;
assign addr[54247]= 1158676398;
assign addr[54248]= 1403673233;
assign addr[54249]= 1620224553;
assign addr[54250]= 1803941934;
assign addr[54251]= 1951102334;
assign addr[54252]= 2058723538;
assign addr[54253]= 2124624598;
assign addr[54254]= 2147470025;
assign addr[54255]= 2126796855;
assign addr[54256]= 2063024031;
assign addr[54257]= 1957443913;
assign addr[54258]= 1812196087;
assign addr[54259]= 1630224009;
assign addr[54260]= 1415215352;
assign addr[54261]= 1171527280;
assign addr[54262]= 904098143;
assign addr[54263]= 618347408;
assign addr[54264]= 320065829;
assign addr[54265]= 15298099;
assign addr[54266]= -289779648;
assign addr[54267]= -588984994;
assign addr[54268]= -876254528;
assign addr[54269]= -1145766716;
assign addr[54270]= -1392059879;
assign addr[54271]= -1610142873;
assign addr[54272]= -1795596234;
assign addr[54273]= -1944661739;
assign addr[54274]= -2054318569;
assign addr[54275]= -2122344521;
assign addr[54276]= -2147361045;
assign addr[54277]= -2128861181;
assign addr[54278]= -2067219829;
assign addr[54279]= -1963686155;
assign addr[54280]= -1820358275;
assign addr[54281]= -1640140734;
assign addr[54282]= -1426685652;
assign addr[54283]= -1184318708;
assign addr[54284]= -917951481;
assign addr[54285]= -632981917;
assign addr[54286]= -335184940;
assign addr[54287]= -30595422;
assign addr[54288]= 274614114;
assign addr[54289]= 574258580;
assign addr[54290]= 862265664;
assign addr[54291]= 1132798888;
assign addr[54292]= 1380375881;
assign addr[54293]= 1599979481;
assign addr[54294]= 1787159411;
assign addr[54295]= 1938122457;
assign addr[54296]= 2049809346;
assign addr[54297]= 2119956737;
assign addr[54298]= 2147143090;
assign addr[54299]= 2130817471;
assign addr[54300]= 2071310720;
assign addr[54301]= 1969828744;
assign addr[54302]= 1828428082;
assign addr[54303]= 1649974225;
assign addr[54304]= 1438083551;
assign addr[54305]= 1197050035;
assign addr[54306]= 931758235;
assign addr[54307]= 647584304;
assign addr[54308]= 350287041;
assign addr[54309]= 45891193;
assign addr[54310]= -259434643;
assign addr[54311]= -559503022;
assign addr[54312]= -848233042;
assign addr[54313]= -1119773573;
assign addr[54314]= -1368621831;
assign addr[54315]= -1589734894;
assign addr[54316]= -1778631892;
assign addr[54317]= -1931484818;
assign addr[54318]= -2045196100;
assign addr[54319]= -2117461370;
assign addr[54320]= -2146816171;
assign addr[54321]= -2132665626;
assign addr[54322]= -2075296495;
assign addr[54323]= -1975871368;
assign addr[54324]= -1836405100;
assign addr[54325]= -1659723983;
assign addr[54326]= -1449408469;
assign addr[54327]= -1209720613;
assign addr[54328]= -945517704;
assign addr[54329]= -662153826;
assign addr[54330]= -365371365;
assign addr[54331]= -61184634;
assign addr[54332]= 244242007;
assign addr[54333]= 544719071;
assign addr[54334]= 834157373;
assign addr[54335]= 1106691431;
assign addr[54336]= 1356798326;
assign addr[54337]= 1579409630;
assign addr[54338]= 1770014111;
assign addr[54339]= 1924749160;
assign addr[54340]= 2040479063;
assign addr[54341]= 2114858546;
assign addr[54342]= 2146380306;
assign addr[54343]= 2134405552;
assign addr[54344]= 2079176953;
assign addr[54345]= 1981813720;
assign addr[54346]= 1844288924;
assign addr[54347]= 1669389513;
assign addr[54348]= 1460659832;
assign addr[54349]= 1222329801;
assign addr[54350]= 959229189;
assign addr[54351]= 676689746;
assign addr[54352]= 380437148;
assign addr[54353]= 76474970;
assign addr[54354]= -229036977;
assign addr[54355]= -529907477;
assign addr[54356]= -820039373;
assign addr[54357]= -1093553126;
assign addr[54358]= -1344905966;
assign addr[54359]= -1569004214;
assign addr[54360]= -1761306505;
assign addr[54361]= -1917915825;
assign addr[54362]= -2035658475;
assign addr[54363]= -2112148396;
assign addr[54364]= -2145835515;
assign addr[54365]= -2136037160;
assign addr[54366]= -2082951896;
assign addr[54367]= -1987655498;
assign addr[54368]= -1852079154;
assign addr[54369]= -1678970324;
assign addr[54370]= -1471837070;
assign addr[54371]= -1234876957;
assign addr[54372]= -972891995;
assign addr[54373]= -691191324;
assign addr[54374]= -395483624;
assign addr[54375]= -91761426;
assign addr[54376]= 213820322;
assign addr[54377]= 515068990;
assign addr[54378]= 805879757;
assign addr[54379]= 1080359326;
assign addr[54380]= 1332945355;
assign addr[54381]= 1558519173;
assign addr[54382]= 1752509516;
assign addr[54383]= 1910985158;
assign addr[54384]= 2030734582;
assign addr[54385]= 2109331059;
assign addr[54386]= 2145181827;
assign addr[54387]= 2137560369;
assign addr[54388]= 2086621133;
assign addr[54389]= 1993396407;
assign addr[54390]= 1859775393;
assign addr[54391]= 1688465931;
assign addr[54392]= 1482939614;
assign addr[54393]= 1247361445;
assign addr[54394]= 986505429;
assign addr[54395]= 705657826;
assign addr[54396]= 410510029;
assign addr[54397]= 107043224;
assign addr[54398]= -198592817;
assign addr[54399]= -500204365;
assign addr[54400]= -791679244;
assign addr[54401]= -1067110699;
assign addr[54402]= -1320917099;
assign addr[54403]= -1547955041;
assign addr[54404]= -1743623590;
assign addr[54405]= -1903957513;
assign addr[54406]= -2025707632;
assign addr[54407]= -2106406677;
assign addr[54408]= -2144419275;
assign addr[54409]= -2138975100;
assign addr[54410]= -2090184478;
assign addr[54411]= -1999036154;
assign addr[54412]= -1867377253;
assign addr[54413]= -1697875851;
assign addr[54414]= -1493966902;
assign addr[54415]= -1259782632;
assign addr[54416]= -1000068799;
assign addr[54417]= -720088517;
assign addr[54418]= -425515602;
assign addr[54419]= -122319591;
assign addr[54420]= 183355234;
assign addr[54421]= 485314355;
assign addr[54422]= 777438554;
assign addr[54423]= 1053807919;
assign addr[54424]= 1308821808;
assign addr[54425]= 1537312353;
assign addr[54426]= 1734649179;
assign addr[54427]= 1896833245;
assign addr[54428]= 2020577882;
assign addr[54429]= 2103375398;
assign addr[54430]= 2143547897;
assign addr[54431]= 2140281282;
assign addr[54432]= 2093641749;
assign addr[54433]= 2004574453;
assign addr[54434]= 1874884346;
assign addr[54435]= 1707199606;
assign addr[54436]= 1504918373;
assign addr[54437]= 1272139887;
assign addr[54438]= 1013581418;
assign addr[54439]= 734482665;
assign addr[54440]= 440499581;
assign addr[54441]= 137589750;
assign addr[54442]= -168108346;
assign addr[54443]= -470399716;
assign addr[54444]= -763158411;
assign addr[54445]= -1040451659;
assign addr[54446]= -1296660098;
assign addr[54447]= -1526591649;
assign addr[54448]= -1725586737;
assign addr[54449]= -1889612716;
assign addr[54450]= -2015345591;
assign addr[54451]= -2100237377;
assign addr[54452]= -2142567738;
assign addr[54453]= -2141478848;
assign addr[54454]= -2096992772;
assign addr[54455]= -2010011024;
assign addr[54456]= -1882296293;
assign addr[54457]= -1716436725;
assign addr[54458]= -1515793473;
assign addr[54459]= -1284432584;
assign addr[54460]= -1027042599;
assign addr[54461]= -748839539;
assign addr[54462]= -455461206;
assign addr[54463]= -152852926;
assign addr[54464]= 152852926;
assign addr[54465]= 455461206;
assign addr[54466]= 748839539;
assign addr[54467]= 1027042599;
assign addr[54468]= 1284432584;
assign addr[54469]= 1515793473;
assign addr[54470]= 1716436725;
assign addr[54471]= 1882296293;
assign addr[54472]= 2010011024;
assign addr[54473]= 2096992772;
assign addr[54474]= 2141478848;
assign addr[54475]= 2142567738;
assign addr[54476]= 2100237377;
assign addr[54477]= 2015345591;
assign addr[54478]= 1889612716;
assign addr[54479]= 1725586737;
assign addr[54480]= 1526591649;
assign addr[54481]= 1296660098;
assign addr[54482]= 1040451659;
assign addr[54483]= 763158411;
assign addr[54484]= 470399716;
assign addr[54485]= 168108346;
assign addr[54486]= -137589750;
assign addr[54487]= -440499581;
assign addr[54488]= -734482665;
assign addr[54489]= -1013581418;
assign addr[54490]= -1272139887;
assign addr[54491]= -1504918373;
assign addr[54492]= -1707199606;
assign addr[54493]= -1874884346;
assign addr[54494]= -2004574453;
assign addr[54495]= -2093641749;
assign addr[54496]= -2140281282;
assign addr[54497]= -2143547897;
assign addr[54498]= -2103375398;
assign addr[54499]= -2020577882;
assign addr[54500]= -1896833245;
assign addr[54501]= -1734649179;
assign addr[54502]= -1537312353;
assign addr[54503]= -1308821808;
assign addr[54504]= -1053807919;
assign addr[54505]= -777438554;
assign addr[54506]= -485314355;
assign addr[54507]= -183355234;
assign addr[54508]= 122319591;
assign addr[54509]= 425515602;
assign addr[54510]= 720088517;
assign addr[54511]= 1000068799;
assign addr[54512]= 1259782632;
assign addr[54513]= 1493966902;
assign addr[54514]= 1697875851;
assign addr[54515]= 1867377253;
assign addr[54516]= 1999036154;
assign addr[54517]= 2090184478;
assign addr[54518]= 2138975100;
assign addr[54519]= 2144419275;
assign addr[54520]= 2106406677;
assign addr[54521]= 2025707632;
assign addr[54522]= 1903957513;
assign addr[54523]= 1743623590;
assign addr[54524]= 1547955041;
assign addr[54525]= 1320917099;
assign addr[54526]= 1067110699;
assign addr[54527]= 791679244;
assign addr[54528]= 500204365;
assign addr[54529]= 198592817;
assign addr[54530]= -107043224;
assign addr[54531]= -410510029;
assign addr[54532]= -705657826;
assign addr[54533]= -986505429;
assign addr[54534]= -1247361445;
assign addr[54535]= -1482939614;
assign addr[54536]= -1688465931;
assign addr[54537]= -1859775393;
assign addr[54538]= -1993396407;
assign addr[54539]= -2086621133;
assign addr[54540]= -2137560369;
assign addr[54541]= -2145181827;
assign addr[54542]= -2109331059;
assign addr[54543]= -2030734582;
assign addr[54544]= -1910985158;
assign addr[54545]= -1752509516;
assign addr[54546]= -1558519173;
assign addr[54547]= -1332945355;
assign addr[54548]= -1080359326;
assign addr[54549]= -805879757;
assign addr[54550]= -515068990;
assign addr[54551]= -213820322;
assign addr[54552]= 91761426;
assign addr[54553]= 395483624;
assign addr[54554]= 691191324;
assign addr[54555]= 972891995;
assign addr[54556]= 1234876957;
assign addr[54557]= 1471837070;
assign addr[54558]= 1678970324;
assign addr[54559]= 1852079154;
assign addr[54560]= 1987655498;
assign addr[54561]= 2082951896;
assign addr[54562]= 2136037160;
assign addr[54563]= 2145835515;
assign addr[54564]= 2112148396;
assign addr[54565]= 2035658475;
assign addr[54566]= 1917915825;
assign addr[54567]= 1761306505;
assign addr[54568]= 1569004214;
assign addr[54569]= 1344905966;
assign addr[54570]= 1093553126;
assign addr[54571]= 820039373;
assign addr[54572]= 529907477;
assign addr[54573]= 229036977;
assign addr[54574]= -76474970;
assign addr[54575]= -380437148;
assign addr[54576]= -676689746;
assign addr[54577]= -959229189;
assign addr[54578]= -1222329801;
assign addr[54579]= -1460659832;
assign addr[54580]= -1669389513;
assign addr[54581]= -1844288924;
assign addr[54582]= -1981813720;
assign addr[54583]= -2079176953;
assign addr[54584]= -2134405552;
assign addr[54585]= -2146380306;
assign addr[54586]= -2114858546;
assign addr[54587]= -2040479063;
assign addr[54588]= -1924749160;
assign addr[54589]= -1770014111;
assign addr[54590]= -1579409630;
assign addr[54591]= -1356798326;
assign addr[54592]= -1106691431;
assign addr[54593]= -834157373;
assign addr[54594]= -544719071;
assign addr[54595]= -244242007;
assign addr[54596]= 61184634;
assign addr[54597]= 365371365;
assign addr[54598]= 662153826;
assign addr[54599]= 945517704;
assign addr[54600]= 1209720613;
assign addr[54601]= 1449408469;
assign addr[54602]= 1659723983;
assign addr[54603]= 1836405100;
assign addr[54604]= 1975871368;
assign addr[54605]= 2075296495;
assign addr[54606]= 2132665626;
assign addr[54607]= 2146816171;
assign addr[54608]= 2117461370;
assign addr[54609]= 2045196100;
assign addr[54610]= 1931484818;
assign addr[54611]= 1778631892;
assign addr[54612]= 1589734894;
assign addr[54613]= 1368621831;
assign addr[54614]= 1119773573;
assign addr[54615]= 848233042;
assign addr[54616]= 559503022;
assign addr[54617]= 259434643;
assign addr[54618]= -45891193;
assign addr[54619]= -350287041;
assign addr[54620]= -647584304;
assign addr[54621]= -931758235;
assign addr[54622]= -1197050035;
assign addr[54623]= -1438083551;
assign addr[54624]= -1649974225;
assign addr[54625]= -1828428082;
assign addr[54626]= -1969828744;
assign addr[54627]= -2071310720;
assign addr[54628]= -2130817471;
assign addr[54629]= -2147143090;
assign addr[54630]= -2119956737;
assign addr[54631]= -2049809346;
assign addr[54632]= -1938122457;
assign addr[54633]= -1787159411;
assign addr[54634]= -1599979481;
assign addr[54635]= -1380375881;
assign addr[54636]= -1132798888;
assign addr[54637]= -862265664;
assign addr[54638]= -574258580;
assign addr[54639]= -274614114;
assign addr[54640]= 30595422;
assign addr[54641]= 335184940;
assign addr[54642]= 632981917;
assign addr[54643]= 917951481;
assign addr[54644]= 1184318708;
assign addr[54645]= 1426685652;
assign addr[54646]= 1640140734;
assign addr[54647]= 1820358275;
assign addr[54648]= 1963686155;
assign addr[54649]= 2067219829;
assign addr[54650]= 2128861181;
assign addr[54651]= 2147361045;
assign addr[54652]= 2122344521;
assign addr[54653]= 2054318569;
assign addr[54654]= 1944661739;
assign addr[54655]= 1795596234;
assign addr[54656]= 1610142873;
assign addr[54657]= 1392059879;
assign addr[54658]= 1145766716;
assign addr[54659]= 876254528;
assign addr[54660]= 588984994;
assign addr[54661]= 289779648;
assign addr[54662]= -15298099;
assign addr[54663]= -320065829;
assign addr[54664]= -618347408;
assign addr[54665]= -904098143;
assign addr[54666]= -1171527280;
assign addr[54667]= -1415215352;
assign addr[54668]= -1630224009;
assign addr[54669]= -1812196087;
assign addr[54670]= -1957443913;
assign addr[54671]= -2063024031;
assign addr[54672]= -2126796855;
assign addr[54673]= -2147470025;
assign addr[54674]= -2124624598;
assign addr[54675]= -2058723538;
assign addr[54676]= -1951102334;
assign addr[54677]= -1803941934;
assign addr[54678]= -1620224553;
assign addr[54679]= -1403673233;
assign addr[54680]= -1158676398;
assign addr[54681]= -890198924;
assign addr[54682]= -603681519;
assign addr[54683]= -304930476;
assign addr[54684]= 0;
assign addr[54685]= 304930476;
assign addr[54686]= 603681519;
assign addr[54687]= 890198924;
assign addr[54688]= 1158676398;
assign addr[54689]= 1403673233;
assign addr[54690]= 1620224553;
assign addr[54691]= 1803941934;
assign addr[54692]= 1951102334;
assign addr[54693]= 2058723538;
assign addr[54694]= 2124624598;
assign addr[54695]= 2147470025;
assign addr[54696]= 2126796855;
assign addr[54697]= 2063024031;
assign addr[54698]= 1957443913;
assign addr[54699]= 1812196087;
assign addr[54700]= 1630224009;
assign addr[54701]= 1415215352;
assign addr[54702]= 1171527280;
assign addr[54703]= 904098143;
assign addr[54704]= 618347408;
assign addr[54705]= 320065829;
assign addr[54706]= 15298099;
assign addr[54707]= -289779648;
assign addr[54708]= -588984994;
assign addr[54709]= -876254528;
assign addr[54710]= -1145766716;
assign addr[54711]= -1392059879;
assign addr[54712]= -1610142873;
assign addr[54713]= -1795596234;
assign addr[54714]= -1944661739;
assign addr[54715]= -2054318569;
assign addr[54716]= -2122344521;
assign addr[54717]= -2147361045;
assign addr[54718]= -2128861181;
assign addr[54719]= -2067219829;
assign addr[54720]= -1963686155;
assign addr[54721]= -1820358275;
assign addr[54722]= -1640140734;
assign addr[54723]= -1426685652;
assign addr[54724]= -1184318708;
assign addr[54725]= -917951481;
assign addr[54726]= -632981917;
assign addr[54727]= -335184940;
assign addr[54728]= -30595422;
assign addr[54729]= 274614114;
assign addr[54730]= 574258580;
assign addr[54731]= 862265664;
assign addr[54732]= 1132798888;
assign addr[54733]= 1380375881;
assign addr[54734]= 1599979481;
assign addr[54735]= 1787159411;
assign addr[54736]= 1938122457;
assign addr[54737]= 2049809346;
assign addr[54738]= 2119956737;
assign addr[54739]= 2147143090;
assign addr[54740]= 2130817471;
assign addr[54741]= 2071310720;
assign addr[54742]= 1969828744;
assign addr[54743]= 1828428082;
assign addr[54744]= 1649974225;
assign addr[54745]= 1438083551;
assign addr[54746]= 1197050035;
assign addr[54747]= 931758235;
assign addr[54748]= 647584304;
assign addr[54749]= 350287041;
assign addr[54750]= 45891193;
assign addr[54751]= -259434643;
assign addr[54752]= -559503022;
assign addr[54753]= -848233042;
assign addr[54754]= -1119773573;
assign addr[54755]= -1368621831;
assign addr[54756]= -1589734894;
assign addr[54757]= -1778631892;
assign addr[54758]= -1931484818;
assign addr[54759]= -2045196100;
assign addr[54760]= -2117461370;
assign addr[54761]= -2146816171;
assign addr[54762]= -2132665626;
assign addr[54763]= -2075296495;
assign addr[54764]= -1975871368;
assign addr[54765]= -1836405100;
assign addr[54766]= -1659723983;
assign addr[54767]= -1449408469;
assign addr[54768]= -1209720613;
assign addr[54769]= -945517704;
assign addr[54770]= -662153826;
assign addr[54771]= -365371365;
assign addr[54772]= -61184634;
assign addr[54773]= 244242007;
assign addr[54774]= 544719071;
assign addr[54775]= 834157373;
assign addr[54776]= 1106691431;
assign addr[54777]= 1356798326;
assign addr[54778]= 1579409630;
assign addr[54779]= 1770014111;
assign addr[54780]= 1924749160;
assign addr[54781]= 2040479063;
assign addr[54782]= 2114858546;
assign addr[54783]= 2146380306;
assign addr[54784]= 2134405552;
assign addr[54785]= 2079176953;
assign addr[54786]= 1981813720;
assign addr[54787]= 1844288924;
assign addr[54788]= 1669389513;
assign addr[54789]= 1460659832;
assign addr[54790]= 1222329801;
assign addr[54791]= 959229189;
assign addr[54792]= 676689746;
assign addr[54793]= 380437148;
assign addr[54794]= 76474970;
assign addr[54795]= -229036977;
assign addr[54796]= -529907477;
assign addr[54797]= -820039373;
assign addr[54798]= -1093553126;
assign addr[54799]= -1344905966;
assign addr[54800]= -1569004214;
assign addr[54801]= -1761306505;
assign addr[54802]= -1917915825;
assign addr[54803]= -2035658475;
assign addr[54804]= -2112148396;
assign addr[54805]= -2145835515;
assign addr[54806]= -2136037160;
assign addr[54807]= -2082951896;
assign addr[54808]= -1987655498;
assign addr[54809]= -1852079154;
assign addr[54810]= -1678970324;
assign addr[54811]= -1471837070;
assign addr[54812]= -1234876957;
assign addr[54813]= -972891995;
assign addr[54814]= -691191324;
assign addr[54815]= -395483624;
assign addr[54816]= -91761426;
assign addr[54817]= 213820322;
assign addr[54818]= 515068990;
assign addr[54819]= 805879757;
assign addr[54820]= 1080359326;
assign addr[54821]= 1332945355;
assign addr[54822]= 1558519173;
assign addr[54823]= 1752509516;
assign addr[54824]= 1910985158;
assign addr[54825]= 2030734582;
assign addr[54826]= 2109331059;
assign addr[54827]= 2145181827;
assign addr[54828]= 2137560369;
assign addr[54829]= 2086621133;
assign addr[54830]= 1993396407;
assign addr[54831]= 1859775393;
assign addr[54832]= 1688465931;
assign addr[54833]= 1482939614;
assign addr[54834]= 1247361445;
assign addr[54835]= 986505429;
assign addr[54836]= 705657826;
assign addr[54837]= 410510029;
assign addr[54838]= 107043224;
assign addr[54839]= -198592817;
assign addr[54840]= -500204365;
assign addr[54841]= -791679244;
assign addr[54842]= -1067110699;
assign addr[54843]= -1320917099;
assign addr[54844]= -1547955041;
assign addr[54845]= -1743623590;
assign addr[54846]= -1903957513;
assign addr[54847]= -2025707632;
assign addr[54848]= -2106406677;
assign addr[54849]= -2144419275;
assign addr[54850]= -2138975100;
assign addr[54851]= -2090184478;
assign addr[54852]= -1999036154;
assign addr[54853]= -1867377253;
assign addr[54854]= -1697875851;
assign addr[54855]= -1493966902;
assign addr[54856]= -1259782632;
assign addr[54857]= -1000068799;
assign addr[54858]= -720088517;
assign addr[54859]= -425515602;
assign addr[54860]= -122319591;
assign addr[54861]= 183355234;
assign addr[54862]= 485314355;
assign addr[54863]= 777438554;
assign addr[54864]= 1053807919;
assign addr[54865]= 1308821808;
assign addr[54866]= 1537312353;
assign addr[54867]= 1734649179;
assign addr[54868]= 1896833245;
assign addr[54869]= 2020577882;
assign addr[54870]= 2103375398;
assign addr[54871]= 2143547897;
assign addr[54872]= 2140281282;
assign addr[54873]= 2093641749;
assign addr[54874]= 2004574453;
assign addr[54875]= 1874884346;
assign addr[54876]= 1707199606;
assign addr[54877]= 1504918373;
assign addr[54878]= 1272139887;
assign addr[54879]= 1013581418;
assign addr[54880]= 734482665;
assign addr[54881]= 440499581;
assign addr[54882]= 137589750;
assign addr[54883]= -168108346;
assign addr[54884]= -470399716;
assign addr[54885]= -763158411;
assign addr[54886]= -1040451659;
assign addr[54887]= -1296660098;
assign addr[54888]= -1526591649;
assign addr[54889]= -1725586737;
assign addr[54890]= -1889612716;
assign addr[54891]= -2015345591;
assign addr[54892]= -2100237377;
assign addr[54893]= -2142567738;
assign addr[54894]= -2141478848;
assign addr[54895]= -2096992772;
assign addr[54896]= -2010011024;
assign addr[54897]= -1882296293;
assign addr[54898]= -1716436725;
assign addr[54899]= -1515793473;
assign addr[54900]= -1284432584;
assign addr[54901]= -1027042599;
assign addr[54902]= -748839539;
assign addr[54903]= -455461206;
assign addr[54904]= -152852926;
assign addr[54905]= 152852926;
assign addr[54906]= 455461206;
assign addr[54907]= 748839539;
assign addr[54908]= 1027042599;
assign addr[54909]= 1284432584;
assign addr[54910]= 1515793473;
assign addr[54911]= 1716436725;
assign addr[54912]= 1882296293;
assign addr[54913]= 2010011024;
assign addr[54914]= 2096992772;
assign addr[54915]= 2141478848;
assign addr[54916]= 2142567738;
assign addr[54917]= 2100237377;
assign addr[54918]= 2015345591;
assign addr[54919]= 1889612716;
assign addr[54920]= 1725586737;
assign addr[54921]= 1526591649;
assign addr[54922]= 1296660098;
assign addr[54923]= 1040451659;
assign addr[54924]= 763158411;
assign addr[54925]= 470399716;
assign addr[54926]= 168108346;
assign addr[54927]= -137589750;
assign addr[54928]= -440499581;
assign addr[54929]= -734482665;
assign addr[54930]= -1013581418;
assign addr[54931]= -1272139887;
assign addr[54932]= -1504918373;
assign addr[54933]= -1707199606;
assign addr[54934]= -1874884346;
assign addr[54935]= -2004574453;
assign addr[54936]= -2093641749;
assign addr[54937]= -2140281282;
assign addr[54938]= -2143547897;
assign addr[54939]= -2103375398;
assign addr[54940]= -2020577882;
assign addr[54941]= -1896833245;
assign addr[54942]= -1734649179;
assign addr[54943]= -1537312353;
assign addr[54944]= -1308821808;
assign addr[54945]= -1053807919;
assign addr[54946]= -777438554;
assign addr[54947]= -485314355;
assign addr[54948]= -183355234;
assign addr[54949]= 122319591;
assign addr[54950]= 425515602;
assign addr[54951]= 720088517;
assign addr[54952]= 1000068799;
assign addr[54953]= 1259782632;
assign addr[54954]= 1493966902;
assign addr[54955]= 1697875851;
assign addr[54956]= 1867377253;
assign addr[54957]= 1999036154;
assign addr[54958]= 2090184478;
assign addr[54959]= 2138975100;
assign addr[54960]= 2144419275;
assign addr[54961]= 2106406677;
assign addr[54962]= 2025707632;
assign addr[54963]= 1903957513;
assign addr[54964]= 1743623590;
assign addr[54965]= 1547955041;
assign addr[54966]= 1320917099;
assign addr[54967]= 1067110699;
assign addr[54968]= 791679244;
assign addr[54969]= 500204365;
assign addr[54970]= 198592817;
assign addr[54971]= -107043224;
assign addr[54972]= -410510029;
assign addr[54973]= -705657826;
assign addr[54974]= -986505429;
assign addr[54975]= -1247361445;
assign addr[54976]= -1482939614;
assign addr[54977]= -1688465931;
assign addr[54978]= -1859775393;
assign addr[54979]= -1993396407;
assign addr[54980]= -2086621133;
assign addr[54981]= -2137560369;
assign addr[54982]= -2145181827;
assign addr[54983]= -2109331059;
assign addr[54984]= -2030734582;
assign addr[54985]= -1910985158;
assign addr[54986]= -1752509516;
assign addr[54987]= -1558519173;
assign addr[54988]= -1332945355;
assign addr[54989]= -1080359326;
assign addr[54990]= -805879757;
assign addr[54991]= -515068990;
assign addr[54992]= -213820322;
assign addr[54993]= 91761426;
assign addr[54994]= 395483624;
assign addr[54995]= 691191324;
assign addr[54996]= 972891995;
assign addr[54997]= 1234876957;
assign addr[54998]= 1471837070;
assign addr[54999]= 1678970324;
assign addr[55000]= 1852079154;
assign addr[55001]= 1987655498;
assign addr[55002]= 2082951896;
assign addr[55003]= 2136037160;
assign addr[55004]= 2145835515;
assign addr[55005]= 2112148396;
assign addr[55006]= 2035658475;
assign addr[55007]= 1917915825;
assign addr[55008]= 1761306505;
assign addr[55009]= 1569004214;
assign addr[55010]= 1344905966;
assign addr[55011]= 1093553126;
assign addr[55012]= 820039373;
assign addr[55013]= 529907477;
assign addr[55014]= 229036977;
assign addr[55015]= -76474970;
assign addr[55016]= -380437148;
assign addr[55017]= -676689746;
assign addr[55018]= -959229189;
assign addr[55019]= -1222329801;
assign addr[55020]= -1460659832;
assign addr[55021]= -1669389513;
assign addr[55022]= -1844288924;
assign addr[55023]= -1981813720;
assign addr[55024]= -2079176953;
assign addr[55025]= -2134405552;
assign addr[55026]= -2146380306;
assign addr[55027]= -2114858546;
assign addr[55028]= -2040479063;
assign addr[55029]= -1924749160;
assign addr[55030]= -1770014111;
assign addr[55031]= -1579409630;
assign addr[55032]= -1356798326;
assign addr[55033]= -1106691431;
assign addr[55034]= -834157373;
assign addr[55035]= -544719071;
assign addr[55036]= -244242007;
assign addr[55037]= 61184634;
assign addr[55038]= 365371365;
assign addr[55039]= 662153826;
assign addr[55040]= 945517704;
assign addr[55041]= 1209720613;
assign addr[55042]= 1449408469;
assign addr[55043]= 1659723983;
assign addr[55044]= 1836405100;
assign addr[55045]= 1975871368;
assign addr[55046]= 2075296495;
assign addr[55047]= 2132665626;
assign addr[55048]= 2146816171;
assign addr[55049]= 2117461370;
assign addr[55050]= 2045196100;
assign addr[55051]= 1931484818;
assign addr[55052]= 1778631892;
assign addr[55053]= 1589734894;
assign addr[55054]= 1368621831;
assign addr[55055]= 1119773573;
assign addr[55056]= 848233042;
assign addr[55057]= 559503022;
assign addr[55058]= 259434643;
assign addr[55059]= -45891193;
assign addr[55060]= -350287041;
assign addr[55061]= -647584304;
assign addr[55062]= -931758235;
assign addr[55063]= -1197050035;
assign addr[55064]= -1438083551;
assign addr[55065]= -1649974225;
assign addr[55066]= -1828428082;
assign addr[55067]= -1969828744;
assign addr[55068]= -2071310720;
assign addr[55069]= -2130817471;
assign addr[55070]= -2147143090;
assign addr[55071]= -2119956737;
assign addr[55072]= -2049809346;
assign addr[55073]= -1938122457;
assign addr[55074]= -1787159411;
assign addr[55075]= -1599979481;
assign addr[55076]= -1380375881;
assign addr[55077]= -1132798888;
assign addr[55078]= -862265664;
assign addr[55079]= -574258580;
assign addr[55080]= -274614114;
assign addr[55081]= 30595422;
assign addr[55082]= 335184940;
assign addr[55083]= 632981917;
assign addr[55084]= 917951481;
assign addr[55085]= 1184318708;
assign addr[55086]= 1426685652;
assign addr[55087]= 1640140734;
assign addr[55088]= 1820358275;
assign addr[55089]= 1963686155;
assign addr[55090]= 2067219829;
assign addr[55091]= 2128861181;
assign addr[55092]= 2147361045;
assign addr[55093]= 2122344521;
assign addr[55094]= 2054318569;
assign addr[55095]= 1944661739;
assign addr[55096]= 1795596234;
assign addr[55097]= 1610142873;
assign addr[55098]= 1392059879;
assign addr[55099]= 1145766716;
assign addr[55100]= 876254528;
assign addr[55101]= 588984994;
assign addr[55102]= 289779648;
assign addr[55103]= -15298099;
assign addr[55104]= -320065829;
assign addr[55105]= -618347408;
assign addr[55106]= -904098143;
assign addr[55107]= -1171527280;
assign addr[55108]= -1415215352;
assign addr[55109]= -1630224009;
assign addr[55110]= -1812196087;
assign addr[55111]= -1957443913;
assign addr[55112]= -2063024031;
assign addr[55113]= -2126796855;
assign addr[55114]= -2147470025;
assign addr[55115]= -2124624598;
assign addr[55116]= -2058723538;
assign addr[55117]= -1951102334;
assign addr[55118]= -1803941934;
assign addr[55119]= -1620224553;
assign addr[55120]= -1403673233;
assign addr[55121]= -1158676398;
assign addr[55122]= -890198924;
assign addr[55123]= -603681519;
assign addr[55124]= -304930476;
assign addr[55125]= 0;
assign addr[55126]= 304930476;
assign addr[55127]= 603681519;
assign addr[55128]= 890198924;
assign addr[55129]= 1158676398;
assign addr[55130]= 1403673233;
assign addr[55131]= 1620224553;
assign addr[55132]= 1803941934;
assign addr[55133]= 1951102334;
assign addr[55134]= 2058723538;
assign addr[55135]= 2124624598;
assign addr[55136]= 2147470025;
assign addr[55137]= 2126796855;
assign addr[55138]= 2063024031;
assign addr[55139]= 1957443913;
assign addr[55140]= 1812196087;
assign addr[55141]= 1630224009;
assign addr[55142]= 1415215352;
assign addr[55143]= 1171527280;
assign addr[55144]= 904098143;
assign addr[55145]= 618347408;
assign addr[55146]= 320065829;
assign addr[55147]= 15298099;
assign addr[55148]= -289779648;
assign addr[55149]= -588984994;
assign addr[55150]= -876254528;
assign addr[55151]= -1145766716;
assign addr[55152]= -1392059879;
assign addr[55153]= -1610142873;
assign addr[55154]= -1795596234;
assign addr[55155]= -1944661739;
assign addr[55156]= -2054318569;
assign addr[55157]= -2122344521;
assign addr[55158]= -2147361045;
assign addr[55159]= -2128861181;
assign addr[55160]= -2067219829;
assign addr[55161]= -1963686155;
assign addr[55162]= -1820358275;
assign addr[55163]= -1640140734;
assign addr[55164]= -1426685652;
assign addr[55165]= -1184318708;
assign addr[55166]= -917951481;
assign addr[55167]= -632981917;
assign addr[55168]= -335184940;
assign addr[55169]= -30595422;
assign addr[55170]= 274614114;
assign addr[55171]= 574258580;
assign addr[55172]= 862265664;
assign addr[55173]= 1132798888;
assign addr[55174]= 1380375881;
assign addr[55175]= 1599979481;
assign addr[55176]= 1787159411;
assign addr[55177]= 1938122457;
assign addr[55178]= 2049809346;
assign addr[55179]= 2119956737;
assign addr[55180]= 2147143090;
assign addr[55181]= 2130817471;
assign addr[55182]= 2071310720;
assign addr[55183]= 1969828744;
assign addr[55184]= 1828428082;
assign addr[55185]= 1649974225;
assign addr[55186]= 1438083551;
assign addr[55187]= 1197050035;
assign addr[55188]= 931758235;
assign addr[55189]= 647584304;
assign addr[55190]= 350287041;
assign addr[55191]= 45891193;
assign addr[55192]= -259434643;
assign addr[55193]= -559503022;
assign addr[55194]= -848233042;
assign addr[55195]= -1119773573;
assign addr[55196]= -1368621831;
assign addr[55197]= -1589734894;
assign addr[55198]= -1778631892;
assign addr[55199]= -1931484818;
assign addr[55200]= -2045196100;
assign addr[55201]= -2117461370;
assign addr[55202]= -2146816171;
assign addr[55203]= -2132665626;
assign addr[55204]= -2075296495;
assign addr[55205]= -1975871368;
assign addr[55206]= -1836405100;
assign addr[55207]= -1659723983;
assign addr[55208]= -1449408469;
assign addr[55209]= -1209720613;
assign addr[55210]= -945517704;
assign addr[55211]= -662153826;
assign addr[55212]= -365371365;
assign addr[55213]= -61184634;
assign addr[55214]= 244242007;
assign addr[55215]= 544719071;
assign addr[55216]= 834157373;
assign addr[55217]= 1106691431;
assign addr[55218]= 1356798326;
assign addr[55219]= 1579409630;
assign addr[55220]= 1770014111;
assign addr[55221]= 1924749160;
assign addr[55222]= 2040479063;
assign addr[55223]= 2114858546;
assign addr[55224]= 2146380306;
assign addr[55225]= 2134405552;
assign addr[55226]= 2079176953;
assign addr[55227]= 1981813720;
assign addr[55228]= 1844288924;
assign addr[55229]= 1669389513;
assign addr[55230]= 1460659832;
assign addr[55231]= 1222329801;
assign addr[55232]= 959229189;
assign addr[55233]= 676689746;
assign addr[55234]= 380437148;
assign addr[55235]= 76474970;
assign addr[55236]= -229036977;
assign addr[55237]= -529907477;
assign addr[55238]= -820039373;
assign addr[55239]= -1093553126;
assign addr[55240]= -1344905966;
assign addr[55241]= -1569004214;
assign addr[55242]= -1761306505;
assign addr[55243]= -1917915825;
assign addr[55244]= -2035658475;
assign addr[55245]= -2112148396;
assign addr[55246]= -2145835515;
assign addr[55247]= -2136037160;
assign addr[55248]= -2082951896;
assign addr[55249]= -1987655498;
assign addr[55250]= -1852079154;
assign addr[55251]= -1678970324;
assign addr[55252]= -1471837070;
assign addr[55253]= -1234876957;
assign addr[55254]= -972891995;
assign addr[55255]= -691191324;
assign addr[55256]= -395483624;
assign addr[55257]= -91761426;
assign addr[55258]= 213820322;
assign addr[55259]= 515068990;
assign addr[55260]= 805879757;
assign addr[55261]= 1080359326;
assign addr[55262]= 1332945355;
assign addr[55263]= 1558519173;
assign addr[55264]= 1752509516;
assign addr[55265]= 1910985158;
assign addr[55266]= 2030734582;
assign addr[55267]= 2109331059;
assign addr[55268]= 2145181827;
assign addr[55269]= 2137560369;
assign addr[55270]= 2086621133;
assign addr[55271]= 1993396407;
assign addr[55272]= 1859775393;
assign addr[55273]= 1688465931;
assign addr[55274]= 1482939614;
assign addr[55275]= 1247361445;
assign addr[55276]= 986505429;
assign addr[55277]= 705657826;
assign addr[55278]= 410510029;
assign addr[55279]= 107043224;
assign addr[55280]= -198592817;
assign addr[55281]= -500204365;
assign addr[55282]= -791679244;
assign addr[55283]= -1067110699;
assign addr[55284]= -1320917099;
assign addr[55285]= -1547955041;
assign addr[55286]= -1743623590;
assign addr[55287]= -1903957513;
assign addr[55288]= -2025707632;
assign addr[55289]= -2106406677;
assign addr[55290]= -2144419275;
assign addr[55291]= -2138975100;
assign addr[55292]= -2090184478;
assign addr[55293]= -1999036154;
assign addr[55294]= -1867377253;
assign addr[55295]= -1697875851;
assign addr[55296]= -1493966902;
assign addr[55297]= -1259782632;
assign addr[55298]= -1000068799;
assign addr[55299]= -720088517;
assign addr[55300]= -425515602;
assign addr[55301]= -122319591;
assign addr[55302]= 183355234;
assign addr[55303]= 485314355;
assign addr[55304]= 777438554;
assign addr[55305]= 1053807919;
assign addr[55306]= 1308821808;
assign addr[55307]= 1537312353;
assign addr[55308]= 1734649179;
assign addr[55309]= 1896833245;
assign addr[55310]= 2020577882;
assign addr[55311]= 2103375398;
assign addr[55312]= 2143547897;
assign addr[55313]= 2140281282;
assign addr[55314]= 2093641749;
assign addr[55315]= 2004574453;
assign addr[55316]= 1874884346;
assign addr[55317]= 1707199606;
assign addr[55318]= 1504918373;
assign addr[55319]= 1272139887;
assign addr[55320]= 1013581418;
assign addr[55321]= 734482665;
assign addr[55322]= 440499581;
assign addr[55323]= 137589750;
assign addr[55324]= -168108346;
assign addr[55325]= -470399716;
assign addr[55326]= -763158411;
assign addr[55327]= -1040451659;
assign addr[55328]= -1296660098;
assign addr[55329]= -1526591649;
assign addr[55330]= -1725586737;
assign addr[55331]= -1889612716;
assign addr[55332]= -2015345591;
assign addr[55333]= -2100237377;
assign addr[55334]= -2142567738;
assign addr[55335]= -2141478848;
assign addr[55336]= -2096992772;
assign addr[55337]= -2010011024;
assign addr[55338]= -1882296293;
assign addr[55339]= -1716436725;
assign addr[55340]= -1515793473;
assign addr[55341]= -1284432584;
assign addr[55342]= -1027042599;
assign addr[55343]= -748839539;
assign addr[55344]= -455461206;
assign addr[55345]= -152852926;
assign addr[55346]= 152852926;
assign addr[55347]= 455461206;
assign addr[55348]= 748839539;
assign addr[55349]= 1027042599;
assign addr[55350]= 1284432584;
assign addr[55351]= 1515793473;
assign addr[55352]= 1716436725;
assign addr[55353]= 1882296293;
assign addr[55354]= 2010011024;
assign addr[55355]= 2096992772;
assign addr[55356]= 2141478848;
assign addr[55357]= 2142567738;
assign addr[55358]= 2100237377;
assign addr[55359]= 2015345591;
assign addr[55360]= 1889612716;
assign addr[55361]= 1725586737;
assign addr[55362]= 1526591649;
assign addr[55363]= 1296660098;
assign addr[55364]= 1040451659;
assign addr[55365]= 763158411;
assign addr[55366]= 470399716;
assign addr[55367]= 168108346;
assign addr[55368]= -137589750;
assign addr[55369]= -440499581;
assign addr[55370]= -734482665;
assign addr[55371]= -1013581418;
assign addr[55372]= -1272139887;
assign addr[55373]= -1504918373;
assign addr[55374]= -1707199606;
assign addr[55375]= -1874884346;
assign addr[55376]= -2004574453;
assign addr[55377]= -2093641749;
assign addr[55378]= -2140281282;
assign addr[55379]= -2143547897;
assign addr[55380]= -2103375398;
assign addr[55381]= -2020577882;
assign addr[55382]= -1896833245;
assign addr[55383]= -1734649179;
assign addr[55384]= -1537312353;
assign addr[55385]= -1308821808;
assign addr[55386]= -1053807919;
assign addr[55387]= -777438554;
assign addr[55388]= -485314355;
assign addr[55389]= -183355234;
assign addr[55390]= 122319591;
assign addr[55391]= 425515602;
assign addr[55392]= 720088517;
assign addr[55393]= 1000068799;
assign addr[55394]= 1259782632;
assign addr[55395]= 1493966902;
assign addr[55396]= 1697875851;
assign addr[55397]= 1867377253;
assign addr[55398]= 1999036154;
assign addr[55399]= 2090184478;
assign addr[55400]= 2138975100;
assign addr[55401]= 2144419275;
assign addr[55402]= 2106406677;
assign addr[55403]= 2025707632;
assign addr[55404]= 1903957513;
assign addr[55405]= 1743623590;
assign addr[55406]= 1547955041;
assign addr[55407]= 1320917099;
assign addr[55408]= 1067110699;
assign addr[55409]= 791679244;
assign addr[55410]= 500204365;
assign addr[55411]= 198592817;
assign addr[55412]= -107043224;
assign addr[55413]= -410510029;
assign addr[55414]= -705657826;
assign addr[55415]= -986505429;
assign addr[55416]= -1247361445;
assign addr[55417]= -1482939614;
assign addr[55418]= -1688465931;
assign addr[55419]= -1859775393;
assign addr[55420]= -1993396407;
assign addr[55421]= -2086621133;
assign addr[55422]= -2137560369;
assign addr[55423]= -2145181827;
assign addr[55424]= -2109331059;
assign addr[55425]= -2030734582;
assign addr[55426]= -1910985158;
assign addr[55427]= -1752509516;
assign addr[55428]= -1558519173;
assign addr[55429]= -1332945355;
assign addr[55430]= -1080359326;
assign addr[55431]= -805879757;
assign addr[55432]= -515068990;
assign addr[55433]= -213820322;
assign addr[55434]= 91761426;
assign addr[55435]= 395483624;
assign addr[55436]= 691191324;
assign addr[55437]= 972891995;
assign addr[55438]= 1234876957;
assign addr[55439]= 1471837070;
assign addr[55440]= 1678970324;
assign addr[55441]= 1852079154;
assign addr[55442]= 1987655498;
assign addr[55443]= 2082951896;
assign addr[55444]= 2136037160;
assign addr[55445]= 2145835515;
assign addr[55446]= 2112148396;
assign addr[55447]= 2035658475;
assign addr[55448]= 1917915825;
assign addr[55449]= 1761306505;
assign addr[55450]= 1569004214;
assign addr[55451]= 1344905966;
assign addr[55452]= 1093553126;
assign addr[55453]= 820039373;
assign addr[55454]= 529907477;
assign addr[55455]= 229036977;
assign addr[55456]= -76474970;
assign addr[55457]= -380437148;
assign addr[55458]= -676689746;
assign addr[55459]= -959229189;
assign addr[55460]= -1222329801;
assign addr[55461]= -1460659832;
assign addr[55462]= -1669389513;
assign addr[55463]= -1844288924;
assign addr[55464]= -1981813720;
assign addr[55465]= -2079176953;
assign addr[55466]= -2134405552;
assign addr[55467]= -2146380306;
assign addr[55468]= -2114858546;
assign addr[55469]= -2040479063;
assign addr[55470]= -1924749160;
assign addr[55471]= -1770014111;
assign addr[55472]= -1579409630;
assign addr[55473]= -1356798326;
assign addr[55474]= -1106691431;
assign addr[55475]= -834157373;
assign addr[55476]= -544719071;
assign addr[55477]= -244242007;
assign addr[55478]= 61184634;
assign addr[55479]= 365371365;
assign addr[55480]= 662153826;
assign addr[55481]= 945517704;
assign addr[55482]= 1209720613;
assign addr[55483]= 1449408469;
assign addr[55484]= 1659723983;
assign addr[55485]= 1836405100;
assign addr[55486]= 1975871368;
assign addr[55487]= 2075296495;
assign addr[55488]= 2132665626;
assign addr[55489]= 2146816171;
assign addr[55490]= 2117461370;
assign addr[55491]= 2045196100;
assign addr[55492]= 1931484818;
assign addr[55493]= 1778631892;
assign addr[55494]= 1589734894;
assign addr[55495]= 1368621831;
assign addr[55496]= 1119773573;
assign addr[55497]= 848233042;
assign addr[55498]= 559503022;
assign addr[55499]= 259434643;
assign addr[55500]= -45891193;
assign addr[55501]= -350287041;
assign addr[55502]= -647584304;
assign addr[55503]= -931758235;
assign addr[55504]= -1197050035;
assign addr[55505]= -1438083551;
assign addr[55506]= -1649974225;
assign addr[55507]= -1828428082;
assign addr[55508]= -1969828744;
assign addr[55509]= -2071310720;
assign addr[55510]= -2130817471;
assign addr[55511]= -2147143090;
assign addr[55512]= -2119956737;
assign addr[55513]= -2049809346;
assign addr[55514]= -1938122457;
assign addr[55515]= -1787159411;
assign addr[55516]= -1599979481;
assign addr[55517]= -1380375881;
assign addr[55518]= -1132798888;
assign addr[55519]= -862265664;
assign addr[55520]= -574258580;
assign addr[55521]= -274614114;
assign addr[55522]= 30595422;
assign addr[55523]= 335184940;
assign addr[55524]= 632981917;
assign addr[55525]= 917951481;
assign addr[55526]= 1184318708;
assign addr[55527]= 1426685652;
assign addr[55528]= 1640140734;
assign addr[55529]= 1820358275;
assign addr[55530]= 1963686155;
assign addr[55531]= 2067219829;
assign addr[55532]= 2128861181;
assign addr[55533]= 2147361045;
assign addr[55534]= 2122344521;
assign addr[55535]= 2054318569;
assign addr[55536]= 1944661739;
assign addr[55537]= 1795596234;
assign addr[55538]= 1610142873;
assign addr[55539]= 1392059879;
assign addr[55540]= 1145766716;
assign addr[55541]= 876254528;
assign addr[55542]= 588984994;
assign addr[55543]= 289779648;
assign addr[55544]= -15298099;
assign addr[55545]= -320065829;
assign addr[55546]= -618347408;
assign addr[55547]= -904098143;
assign addr[55548]= -1171527280;
assign addr[55549]= -1415215352;
assign addr[55550]= -1630224009;
assign addr[55551]= -1812196087;
assign addr[55552]= -1957443913;
assign addr[55553]= -2063024031;
assign addr[55554]= -2126796855;
assign addr[55555]= -2147470025;
assign addr[55556]= -2124624598;
assign addr[55557]= -2058723538;
assign addr[55558]= -1951102334;
assign addr[55559]= -1803941934;
assign addr[55560]= -1620224553;
assign addr[55561]= -1403673233;
assign addr[55562]= -1158676398;
assign addr[55563]= -890198924;
assign addr[55564]= -603681519;
assign addr[55565]= -304930476;
assign addr[55566]= 0;
assign addr[55567]= 304930476;
assign addr[55568]= 603681519;
assign addr[55569]= 890198924;
assign addr[55570]= 1158676398;
assign addr[55571]= 1403673233;
assign addr[55572]= 1620224553;
assign addr[55573]= 1803941934;
assign addr[55574]= 1951102334;
assign addr[55575]= 2058723538;
assign addr[55576]= 2124624598;
assign addr[55577]= 2147470025;
assign addr[55578]= 2126796855;
assign addr[55579]= 2063024031;
assign addr[55580]= 1957443913;
assign addr[55581]= 1812196087;
assign addr[55582]= 1630224009;
assign addr[55583]= 1415215352;
assign addr[55584]= 1171527280;
assign addr[55585]= 904098143;
assign addr[55586]= 618347408;
assign addr[55587]= 320065829;
assign addr[55588]= 15298099;
assign addr[55589]= -289779648;
assign addr[55590]= -588984994;
assign addr[55591]= -876254528;
assign addr[55592]= -1145766716;
assign addr[55593]= -1392059879;
assign addr[55594]= -1610142873;
assign addr[55595]= -1795596234;
assign addr[55596]= -1944661739;
assign addr[55597]= -2054318569;
assign addr[55598]= -2122344521;
assign addr[55599]= -2147361045;
assign addr[55600]= -2128861181;
assign addr[55601]= -2067219829;
assign addr[55602]= -1963686155;
assign addr[55603]= -1820358275;
assign addr[55604]= -1640140734;
assign addr[55605]= -1426685652;
assign addr[55606]= -1184318708;
assign addr[55607]= -917951481;
assign addr[55608]= -632981917;
assign addr[55609]= -335184940;
assign addr[55610]= -30595422;
assign addr[55611]= 274614114;
assign addr[55612]= 574258580;
assign addr[55613]= 862265664;
assign addr[55614]= 1132798888;
assign addr[55615]= 1380375881;
assign addr[55616]= 1599979481;
assign addr[55617]= 1787159411;
assign addr[55618]= 1938122457;
assign addr[55619]= 2049809346;
assign addr[55620]= 2119956737;
assign addr[55621]= 2147143090;
assign addr[55622]= 2130817471;
assign addr[55623]= 2071310720;
assign addr[55624]= 1969828744;
assign addr[55625]= 1828428082;
assign addr[55626]= 1649974225;
assign addr[55627]= 1438083551;
assign addr[55628]= 1197050035;
assign addr[55629]= 931758235;
assign addr[55630]= 647584304;
assign addr[55631]= 350287041;
assign addr[55632]= 45891193;
assign addr[55633]= -259434643;
assign addr[55634]= -559503022;
assign addr[55635]= -848233042;
assign addr[55636]= -1119773573;
assign addr[55637]= -1368621831;
assign addr[55638]= -1589734894;
assign addr[55639]= -1778631892;
assign addr[55640]= -1931484818;
assign addr[55641]= -2045196100;
assign addr[55642]= -2117461370;
assign addr[55643]= -2146816171;
assign addr[55644]= -2132665626;
assign addr[55645]= -2075296495;
assign addr[55646]= -1975871368;
assign addr[55647]= -1836405100;
assign addr[55648]= -1659723983;
assign addr[55649]= -1449408469;
assign addr[55650]= -1209720613;
assign addr[55651]= -945517704;
assign addr[55652]= -662153826;
assign addr[55653]= -365371365;
assign addr[55654]= -61184634;
assign addr[55655]= 244242007;
assign addr[55656]= 544719071;
assign addr[55657]= 834157373;
assign addr[55658]= 1106691431;
assign addr[55659]= 1356798326;
assign addr[55660]= 1579409630;
assign addr[55661]= 1770014111;
assign addr[55662]= 1924749160;
assign addr[55663]= 2040479063;
assign addr[55664]= 2114858546;
assign addr[55665]= 2146380306;
assign addr[55666]= 2134405552;
assign addr[55667]= 2079176953;
assign addr[55668]= 1981813720;
assign addr[55669]= 1844288924;
assign addr[55670]= 1669389513;
assign addr[55671]= 1460659832;
assign addr[55672]= 1222329801;
assign addr[55673]= 959229189;
assign addr[55674]= 676689746;
assign addr[55675]= 380437148;
assign addr[55676]= 76474970;
assign addr[55677]= -229036977;
assign addr[55678]= -529907477;
assign addr[55679]= -820039373;
assign addr[55680]= -1093553126;
assign addr[55681]= -1344905966;
assign addr[55682]= -1569004214;
assign addr[55683]= -1761306505;
assign addr[55684]= -1917915825;
assign addr[55685]= -2035658475;
assign addr[55686]= -2112148396;
assign addr[55687]= -2145835515;
assign addr[55688]= -2136037160;
assign addr[55689]= -2082951896;
assign addr[55690]= -1987655498;
assign addr[55691]= -1852079154;
assign addr[55692]= -1678970324;
assign addr[55693]= -1471837070;
assign addr[55694]= -1234876957;
assign addr[55695]= -972891995;
assign addr[55696]= -691191324;
assign addr[55697]= -395483624;
assign addr[55698]= -91761426;
assign addr[55699]= 213820322;
assign addr[55700]= 515068990;
assign addr[55701]= 805879757;
assign addr[55702]= 1080359326;
assign addr[55703]= 1332945355;
assign addr[55704]= 1558519173;
assign addr[55705]= 1752509516;
assign addr[55706]= 1910985158;
assign addr[55707]= 2030734582;
assign addr[55708]= 2109331059;
assign addr[55709]= 2145181827;
assign addr[55710]= 2137560369;
assign addr[55711]= 2086621133;
assign addr[55712]= 1993396407;
assign addr[55713]= 1859775393;
assign addr[55714]= 1688465931;
assign addr[55715]= 1482939614;
assign addr[55716]= 1247361445;
assign addr[55717]= 986505429;
assign addr[55718]= 705657826;
assign addr[55719]= 410510029;
assign addr[55720]= 107043224;
assign addr[55721]= -198592817;
assign addr[55722]= -500204365;
assign addr[55723]= -791679244;
assign addr[55724]= -1067110699;
assign addr[55725]= -1320917099;
assign addr[55726]= -1547955041;
assign addr[55727]= -1743623590;
assign addr[55728]= -1903957513;
assign addr[55729]= -2025707632;
assign addr[55730]= -2106406677;
assign addr[55731]= -2144419275;
assign addr[55732]= -2138975100;
assign addr[55733]= -2090184478;
assign addr[55734]= -1999036154;
assign addr[55735]= -1867377253;
assign addr[55736]= -1697875851;
assign addr[55737]= -1493966902;
assign addr[55738]= -1259782632;
assign addr[55739]= -1000068799;
assign addr[55740]= -720088517;
assign addr[55741]= -425515602;
assign addr[55742]= -122319591;
assign addr[55743]= 183355234;
assign addr[55744]= 485314355;
assign addr[55745]= 777438554;
assign addr[55746]= 1053807919;
assign addr[55747]= 1308821808;
assign addr[55748]= 1537312353;
assign addr[55749]= 1734649179;
assign addr[55750]= 1896833245;
assign addr[55751]= 2020577882;
assign addr[55752]= 2103375398;
assign addr[55753]= 2143547897;
assign addr[55754]= 2140281282;
assign addr[55755]= 2093641749;
assign addr[55756]= 2004574453;
assign addr[55757]= 1874884346;
assign addr[55758]= 1707199606;
assign addr[55759]= 1504918373;
assign addr[55760]= 1272139887;
assign addr[55761]= 1013581418;
assign addr[55762]= 734482665;
assign addr[55763]= 440499581;
assign addr[55764]= 137589750;
assign addr[55765]= -168108346;
assign addr[55766]= -470399716;
assign addr[55767]= -763158411;
assign addr[55768]= -1040451659;
assign addr[55769]= -1296660098;
assign addr[55770]= -1526591649;
assign addr[55771]= -1725586737;
assign addr[55772]= -1889612716;
assign addr[55773]= -2015345591;
assign addr[55774]= -2100237377;
assign addr[55775]= -2142567738;
assign addr[55776]= -2141478848;
assign addr[55777]= -2096992772;
assign addr[55778]= -2010011024;
assign addr[55779]= -1882296293;
assign addr[55780]= -1716436725;
assign addr[55781]= -1515793473;
assign addr[55782]= -1284432584;
assign addr[55783]= -1027042599;
assign addr[55784]= -748839539;
assign addr[55785]= -455461206;
assign addr[55786]= -152852926;
assign addr[55787]= 152852926;
assign addr[55788]= 455461206;
assign addr[55789]= 748839539;
assign addr[55790]= 1027042599;
assign addr[55791]= 1284432584;
assign addr[55792]= 1515793473;
assign addr[55793]= 1716436725;
assign addr[55794]= 1882296293;
assign addr[55795]= 2010011024;
assign addr[55796]= 2096992772;
assign addr[55797]= 2141478848;
assign addr[55798]= 2142567738;
assign addr[55799]= 2100237377;
assign addr[55800]= 2015345591;
assign addr[55801]= 1889612716;
assign addr[55802]= 1725586737;
assign addr[55803]= 1526591649;
assign addr[55804]= 1296660098;
assign addr[55805]= 1040451659;
assign addr[55806]= 763158411;
assign addr[55807]= 470399716;
assign addr[55808]= 168108346;
assign addr[55809]= -137589750;
assign addr[55810]= -440499581;
assign addr[55811]= -734482665;
assign addr[55812]= -1013581418;
assign addr[55813]= -1272139887;
assign addr[55814]= -1504918373;
assign addr[55815]= -1707199606;
assign addr[55816]= -1874884346;
assign addr[55817]= -2004574453;
assign addr[55818]= -2093641749;
assign addr[55819]= -2140281282;
assign addr[55820]= -2143547897;
assign addr[55821]= -2103375398;
assign addr[55822]= -2020577882;
assign addr[55823]= -1896833245;
assign addr[55824]= -1734649179;
assign addr[55825]= -1537312353;
assign addr[55826]= -1308821808;
assign addr[55827]= -1053807919;
assign addr[55828]= -777438554;
assign addr[55829]= -485314355;
assign addr[55830]= -183355234;
assign addr[55831]= 122319591;
assign addr[55832]= 425515602;
assign addr[55833]= 720088517;
assign addr[55834]= 1000068799;
assign addr[55835]= 1259782632;
assign addr[55836]= 1493966902;
assign addr[55837]= 1697875851;
assign addr[55838]= 1867377253;
assign addr[55839]= 1999036154;
assign addr[55840]= 2090184478;
assign addr[55841]= 2138975100;
assign addr[55842]= 2144419275;
assign addr[55843]= 2106406677;
assign addr[55844]= 2025707632;
assign addr[55845]= 1903957513;
assign addr[55846]= 1743623590;
assign addr[55847]= 1547955041;
assign addr[55848]= 1320917099;
assign addr[55849]= 1067110699;
assign addr[55850]= 791679244;
assign addr[55851]= 500204365;
assign addr[55852]= 198592817;
assign addr[55853]= -107043224;
assign addr[55854]= -410510029;
assign addr[55855]= -705657826;
assign addr[55856]= -986505429;
assign addr[55857]= -1247361445;
assign addr[55858]= -1482939614;
assign addr[55859]= -1688465931;
assign addr[55860]= -1859775393;
assign addr[55861]= -1993396407;
assign addr[55862]= -2086621133;
assign addr[55863]= -2137560369;
assign addr[55864]= -2145181827;
assign addr[55865]= -2109331059;
assign addr[55866]= -2030734582;
assign addr[55867]= -1910985158;
assign addr[55868]= -1752509516;
assign addr[55869]= -1558519173;
assign addr[55870]= -1332945355;
assign addr[55871]= -1080359326;
assign addr[55872]= -805879757;
assign addr[55873]= -515068990;
assign addr[55874]= -213820322;
assign addr[55875]= 91761426;
assign addr[55876]= 395483624;
assign addr[55877]= 691191324;
assign addr[55878]= 972891995;
assign addr[55879]= 1234876957;
assign addr[55880]= 1471837070;
assign addr[55881]= 1678970324;
assign addr[55882]= 1852079154;
assign addr[55883]= 1987655498;
assign addr[55884]= 2082951896;
assign addr[55885]= 2136037160;
assign addr[55886]= 2145835515;
assign addr[55887]= 2112148396;
assign addr[55888]= 2035658475;
assign addr[55889]= 1917915825;
assign addr[55890]= 1761306505;
assign addr[55891]= 1569004214;
assign addr[55892]= 1344905966;
assign addr[55893]= 1093553126;
assign addr[55894]= 820039373;
assign addr[55895]= 529907477;
assign addr[55896]= 229036977;
assign addr[55897]= -76474970;
assign addr[55898]= -380437148;
assign addr[55899]= -676689746;
assign addr[55900]= -959229189;
assign addr[55901]= -1222329801;
assign addr[55902]= -1460659832;
assign addr[55903]= -1669389513;
assign addr[55904]= -1844288924;
assign addr[55905]= -1981813720;
assign addr[55906]= -2079176953;
assign addr[55907]= -2134405552;
assign addr[55908]= -2146380306;
assign addr[55909]= -2114858546;
assign addr[55910]= -2040479063;
assign addr[55911]= -1924749160;
assign addr[55912]= -1770014111;
assign addr[55913]= -1579409630;
assign addr[55914]= -1356798326;
assign addr[55915]= -1106691431;
assign addr[55916]= -834157373;
assign addr[55917]= -544719071;
assign addr[55918]= -244242007;
assign addr[55919]= 61184634;
assign addr[55920]= 365371365;
assign addr[55921]= 662153826;
assign addr[55922]= 945517704;
assign addr[55923]= 1209720613;
assign addr[55924]= 1449408469;
assign addr[55925]= 1659723983;
assign addr[55926]= 1836405100;
assign addr[55927]= 1975871368;
assign addr[55928]= 2075296495;
assign addr[55929]= 2132665626;
assign addr[55930]= 2146816171;
assign addr[55931]= 2117461370;
assign addr[55932]= 2045196100;
assign addr[55933]= 1931484818;
assign addr[55934]= 1778631892;
assign addr[55935]= 1589734894;
assign addr[55936]= 1368621831;
assign addr[55937]= 1119773573;
assign addr[55938]= 848233042;
assign addr[55939]= 559503022;
assign addr[55940]= 259434643;
assign addr[55941]= -45891193;
assign addr[55942]= -350287041;
assign addr[55943]= -647584304;
assign addr[55944]= -931758235;
assign addr[55945]= -1197050035;
assign addr[55946]= -1438083551;
assign addr[55947]= -1649974225;
assign addr[55948]= -1828428082;
assign addr[55949]= -1969828744;
assign addr[55950]= -2071310720;
assign addr[55951]= -2130817471;
assign addr[55952]= -2147143090;
assign addr[55953]= -2119956737;
assign addr[55954]= -2049809346;
assign addr[55955]= -1938122457;
assign addr[55956]= -1787159411;
assign addr[55957]= -1599979481;
assign addr[55958]= -1380375881;
assign addr[55959]= -1132798888;
assign addr[55960]= -862265664;
assign addr[55961]= -574258580;
assign addr[55962]= -274614114;
assign addr[55963]= 30595422;
assign addr[55964]= 335184940;
assign addr[55965]= 632981917;
assign addr[55966]= 917951481;
assign addr[55967]= 1184318708;
assign addr[55968]= 1426685652;
assign addr[55969]= 1640140734;
assign addr[55970]= 1820358275;
assign addr[55971]= 1963686155;
assign addr[55972]= 2067219829;
assign addr[55973]= 2128861181;
assign addr[55974]= 2147361045;
assign addr[55975]= 2122344521;
assign addr[55976]= 2054318569;
assign addr[55977]= 1944661739;
assign addr[55978]= 1795596234;
assign addr[55979]= 1610142873;
assign addr[55980]= 1392059879;
assign addr[55981]= 1145766716;
assign addr[55982]= 876254528;
assign addr[55983]= 588984994;
assign addr[55984]= 289779648;
assign addr[55985]= -15298099;
assign addr[55986]= -320065829;
assign addr[55987]= -618347408;
assign addr[55988]= -904098143;
assign addr[55989]= -1171527280;
assign addr[55990]= -1415215352;
assign addr[55991]= -1630224009;
assign addr[55992]= -1812196087;
assign addr[55993]= -1957443913;
assign addr[55994]= -2063024031;
assign addr[55995]= -2126796855;
assign addr[55996]= -2147470025;
assign addr[55997]= -2124624598;
assign addr[55998]= -2058723538;
assign addr[55999]= -1951102334;
assign addr[56000]= -1803941934;
assign addr[56001]= -1620224553;
assign addr[56002]= -1403673233;
assign addr[56003]= -1158676398;
assign addr[56004]= -890198924;
assign addr[56005]= -603681519;
assign addr[56006]= -304930476;
assign addr[56007]= 0;
assign addr[56008]= 304930476;
assign addr[56009]= 603681519;
assign addr[56010]= 890198924;
assign addr[56011]= 1158676398;
assign addr[56012]= 1403673233;
assign addr[56013]= 1620224553;
assign addr[56014]= 1803941934;
assign addr[56015]= 1951102334;
assign addr[56016]= 2058723538;
assign addr[56017]= 2124624598;
assign addr[56018]= 2147470025;
assign addr[56019]= 2126796855;
assign addr[56020]= 2063024031;
assign addr[56021]= 1957443913;
assign addr[56022]= 1812196087;
assign addr[56023]= 1630224009;
assign addr[56024]= 1415215352;
assign addr[56025]= 1171527280;
assign addr[56026]= 904098143;
assign addr[56027]= 618347408;
assign addr[56028]= 320065829;
assign addr[56029]= 15298099;
assign addr[56030]= -289779648;
assign addr[56031]= -588984994;
assign addr[56032]= -876254528;
assign addr[56033]= -1145766716;
assign addr[56034]= -1392059879;
assign addr[56035]= -1610142873;
assign addr[56036]= -1795596234;
assign addr[56037]= -1944661739;
assign addr[56038]= -2054318569;
assign addr[56039]= -2122344521;
assign addr[56040]= -2147361045;
assign addr[56041]= -2128861181;
assign addr[56042]= -2067219829;
assign addr[56043]= -1963686155;
assign addr[56044]= -1820358275;
assign addr[56045]= -1640140734;
assign addr[56046]= -1426685652;
assign addr[56047]= -1184318708;
assign addr[56048]= -917951481;
assign addr[56049]= -632981917;
assign addr[56050]= -335184940;
assign addr[56051]= -30595422;
assign addr[56052]= 274614114;
assign addr[56053]= 574258580;
assign addr[56054]= 862265664;
assign addr[56055]= 1132798888;
assign addr[56056]= 1380375881;
assign addr[56057]= 1599979481;
assign addr[56058]= 1787159411;
assign addr[56059]= 1938122457;
assign addr[56060]= 2049809346;
assign addr[56061]= 2119956737;
assign addr[56062]= 2147143090;
assign addr[56063]= 2130817471;
assign addr[56064]= 2071310720;
assign addr[56065]= 1969828744;
assign addr[56066]= 1828428082;
assign addr[56067]= 1649974225;
assign addr[56068]= 1438083551;
assign addr[56069]= 1197050035;
assign addr[56070]= 931758235;
assign addr[56071]= 647584304;
assign addr[56072]= 350287041;
assign addr[56073]= 45891193;
assign addr[56074]= -259434643;
assign addr[56075]= -559503022;
assign addr[56076]= -848233042;
assign addr[56077]= -1119773573;
assign addr[56078]= -1368621831;
assign addr[56079]= -1589734894;
assign addr[56080]= -1778631892;
assign addr[56081]= -1931484818;
assign addr[56082]= -2045196100;
assign addr[56083]= -2117461370;
assign addr[56084]= -2146816171;
assign addr[56085]= -2132665626;
assign addr[56086]= -2075296495;
assign addr[56087]= -1975871368;
assign addr[56088]= -1836405100;
assign addr[56089]= -1659723983;
assign addr[56090]= -1449408469;
assign addr[56091]= -1209720613;
assign addr[56092]= -945517704;
assign addr[56093]= -662153826;
assign addr[56094]= -365371365;
assign addr[56095]= -61184634;
assign addr[56096]= 244242007;
assign addr[56097]= 544719071;
assign addr[56098]= 834157373;
assign addr[56099]= 1106691431;
assign addr[56100]= 1356798326;
assign addr[56101]= 1579409630;
assign addr[56102]= 1770014111;
assign addr[56103]= 1924749160;
assign addr[56104]= 2040479063;
assign addr[56105]= 2114858546;
assign addr[56106]= 2146380306;
assign addr[56107]= 2134405552;
assign addr[56108]= 2079176953;
assign addr[56109]= 1981813720;
assign addr[56110]= 1844288924;
assign addr[56111]= 1669389513;
assign addr[56112]= 1460659832;
assign addr[56113]= 1222329801;
assign addr[56114]= 959229189;
assign addr[56115]= 676689746;
assign addr[56116]= 380437148;
assign addr[56117]= 76474970;
assign addr[56118]= -229036977;
assign addr[56119]= -529907477;
assign addr[56120]= -820039373;
assign addr[56121]= -1093553126;
assign addr[56122]= -1344905966;
assign addr[56123]= -1569004214;
assign addr[56124]= -1761306505;
assign addr[56125]= -1917915825;
assign addr[56126]= -2035658475;
assign addr[56127]= -2112148396;
assign addr[56128]= -2145835515;
assign addr[56129]= -2136037160;
assign addr[56130]= -2082951896;
assign addr[56131]= -1987655498;
assign addr[56132]= -1852079154;
assign addr[56133]= -1678970324;
assign addr[56134]= -1471837070;
assign addr[56135]= -1234876957;
assign addr[56136]= -972891995;
assign addr[56137]= -691191324;
assign addr[56138]= -395483624;
assign addr[56139]= -91761426;
assign addr[56140]= 213820322;
assign addr[56141]= 515068990;
assign addr[56142]= 805879757;
assign addr[56143]= 1080359326;
assign addr[56144]= 1332945355;
assign addr[56145]= 1558519173;
assign addr[56146]= 1752509516;
assign addr[56147]= 1910985158;
assign addr[56148]= 2030734582;
assign addr[56149]= 2109331059;
assign addr[56150]= 2145181827;
assign addr[56151]= 2137560369;
assign addr[56152]= 2086621133;
assign addr[56153]= 1993396407;
assign addr[56154]= 1859775393;
assign addr[56155]= 1688465931;
assign addr[56156]= 1482939614;
assign addr[56157]= 1247361445;
assign addr[56158]= 986505429;
assign addr[56159]= 705657826;
assign addr[56160]= 410510029;
assign addr[56161]= 107043224;
assign addr[56162]= -198592817;
assign addr[56163]= -500204365;
assign addr[56164]= -791679244;
assign addr[56165]= -1067110699;
assign addr[56166]= -1320917099;
assign addr[56167]= -1547955041;
assign addr[56168]= -1743623590;
assign addr[56169]= -1903957513;
assign addr[56170]= -2025707632;
assign addr[56171]= -2106406677;
assign addr[56172]= -2144419275;
assign addr[56173]= -2138975100;
assign addr[56174]= -2090184478;
assign addr[56175]= -1999036154;
assign addr[56176]= -1867377253;
assign addr[56177]= -1697875851;
assign addr[56178]= -1493966902;
assign addr[56179]= -1259782632;
assign addr[56180]= -1000068799;
assign addr[56181]= -720088517;
assign addr[56182]= -425515602;
assign addr[56183]= -122319591;
assign addr[56184]= 183355234;
assign addr[56185]= 485314355;
assign addr[56186]= 777438554;
assign addr[56187]= 1053807919;
assign addr[56188]= 1308821808;
assign addr[56189]= 1537312353;
assign addr[56190]= 1734649179;
assign addr[56191]= 1896833245;
assign addr[56192]= 2020577882;
assign addr[56193]= 2103375398;
assign addr[56194]= 2143547897;
assign addr[56195]= 2140281282;
assign addr[56196]= 2093641749;
assign addr[56197]= 2004574453;
assign addr[56198]= 1874884346;
assign addr[56199]= 1707199606;
assign addr[56200]= 1504918373;
assign addr[56201]= 1272139887;
assign addr[56202]= 1013581418;
assign addr[56203]= 734482665;
assign addr[56204]= 440499581;
assign addr[56205]= 137589750;
assign addr[56206]= -168108346;
assign addr[56207]= -470399716;
assign addr[56208]= -763158411;
assign addr[56209]= -1040451659;
assign addr[56210]= -1296660098;
assign addr[56211]= -1526591649;
assign addr[56212]= -1725586737;
assign addr[56213]= -1889612716;
assign addr[56214]= -2015345591;
assign addr[56215]= -2100237377;
assign addr[56216]= -2142567738;
assign addr[56217]= -2141478848;
assign addr[56218]= -2096992772;
assign addr[56219]= -2010011024;
assign addr[56220]= -1882296293;
assign addr[56221]= -1716436725;
assign addr[56222]= -1515793473;
assign addr[56223]= -1284432584;
assign addr[56224]= -1027042599;
assign addr[56225]= -748839539;
assign addr[56226]= -455461206;
assign addr[56227]= -152852926;
assign addr[56228]= 152852926;
assign addr[56229]= 455461206;
assign addr[56230]= 748839539;
assign addr[56231]= 1027042599;
assign addr[56232]= 1284432584;
assign addr[56233]= 1515793473;
assign addr[56234]= 1716436725;
assign addr[56235]= 1882296293;
assign addr[56236]= 2010011024;
assign addr[56237]= 2096992772;
assign addr[56238]= 2141478848;
assign addr[56239]= 2142567738;
assign addr[56240]= 2100237377;
assign addr[56241]= 2015345591;
assign addr[56242]= 1889612716;
assign addr[56243]= 1725586737;
assign addr[56244]= 1526591649;
assign addr[56245]= 1296660098;
assign addr[56246]= 1040451659;
assign addr[56247]= 763158411;
assign addr[56248]= 470399716;
assign addr[56249]= 168108346;
assign addr[56250]= -137589750;
assign addr[56251]= -440499581;
assign addr[56252]= -734482665;
assign addr[56253]= -1013581418;
assign addr[56254]= -1272139887;
assign addr[56255]= -1504918373;
assign addr[56256]= -1707199606;
assign addr[56257]= -1874884346;
assign addr[56258]= -2004574453;
assign addr[56259]= -2093641749;
assign addr[56260]= -2140281282;
assign addr[56261]= -2143547897;
assign addr[56262]= -2103375398;
assign addr[56263]= -2020577882;
assign addr[56264]= -1896833245;
assign addr[56265]= -1734649179;
assign addr[56266]= -1537312353;
assign addr[56267]= -1308821808;
assign addr[56268]= -1053807919;
assign addr[56269]= -777438554;
assign addr[56270]= -485314355;
assign addr[56271]= -183355234;
assign addr[56272]= 122319591;
assign addr[56273]= 425515602;
assign addr[56274]= 720088517;
assign addr[56275]= 1000068799;
assign addr[56276]= 1259782632;
assign addr[56277]= 1493966902;
assign addr[56278]= 1697875851;
assign addr[56279]= 1867377253;
assign addr[56280]= 1999036154;
assign addr[56281]= 2090184478;
assign addr[56282]= 2138975100;
assign addr[56283]= 2144419275;
assign addr[56284]= 2106406677;
assign addr[56285]= 2025707632;
assign addr[56286]= 1903957513;
assign addr[56287]= 1743623590;
assign addr[56288]= 1547955041;
assign addr[56289]= 1320917099;
assign addr[56290]= 1067110699;
assign addr[56291]= 791679244;
assign addr[56292]= 500204365;
assign addr[56293]= 198592817;
assign addr[56294]= -107043224;
assign addr[56295]= -410510029;
assign addr[56296]= -705657826;
assign addr[56297]= -986505429;
assign addr[56298]= -1247361445;
assign addr[56299]= -1482939614;
assign addr[56300]= -1688465931;
assign addr[56301]= -1859775393;
assign addr[56302]= -1993396407;
assign addr[56303]= -2086621133;
assign addr[56304]= -2137560369;
assign addr[56305]= -2145181827;
assign addr[56306]= -2109331059;
assign addr[56307]= -2030734582;
assign addr[56308]= -1910985158;
assign addr[56309]= -1752509516;
assign addr[56310]= -1558519173;
assign addr[56311]= -1332945355;
assign addr[56312]= -1080359326;
assign addr[56313]= -805879757;
assign addr[56314]= -515068990;
assign addr[56315]= -213820322;
assign addr[56316]= 91761426;
assign addr[56317]= 395483624;
assign addr[56318]= 691191324;
assign addr[56319]= 972891995;
assign addr[56320]= 1234876957;
assign addr[56321]= 1471837070;
assign addr[56322]= 1678970324;
assign addr[56323]= 1852079154;
assign addr[56324]= 1987655498;
assign addr[56325]= 2082951896;
assign addr[56326]= 2136037160;
assign addr[56327]= 2145835515;
assign addr[56328]= 2112148396;
assign addr[56329]= 2035658475;
assign addr[56330]= 1917915825;
assign addr[56331]= 1761306505;
assign addr[56332]= 1569004214;
assign addr[56333]= 1344905966;
assign addr[56334]= 1093553126;
assign addr[56335]= 820039373;
assign addr[56336]= 529907477;
assign addr[56337]= 229036977;
assign addr[56338]= -76474970;
assign addr[56339]= -380437148;
assign addr[56340]= -676689746;
assign addr[56341]= -959229189;
assign addr[56342]= -1222329801;
assign addr[56343]= -1460659832;
assign addr[56344]= -1669389513;
assign addr[56345]= -1844288924;
assign addr[56346]= -1981813720;
assign addr[56347]= -2079176953;
assign addr[56348]= -2134405552;
assign addr[56349]= -2146380306;
assign addr[56350]= -2114858546;
assign addr[56351]= -2040479063;
assign addr[56352]= -1924749160;
assign addr[56353]= -1770014111;
assign addr[56354]= -1579409630;
assign addr[56355]= -1356798326;
assign addr[56356]= -1106691431;
assign addr[56357]= -834157373;
assign addr[56358]= -544719071;
assign addr[56359]= -244242007;
assign addr[56360]= 61184634;
assign addr[56361]= 365371365;
assign addr[56362]= 662153826;
assign addr[56363]= 945517704;
assign addr[56364]= 1209720613;
assign addr[56365]= 1449408469;
assign addr[56366]= 1659723983;
assign addr[56367]= 1836405100;
assign addr[56368]= 1975871368;
assign addr[56369]= 2075296495;
assign addr[56370]= 2132665626;
assign addr[56371]= 2146816171;
assign addr[56372]= 2117461370;
assign addr[56373]= 2045196100;
assign addr[56374]= 1931484818;
assign addr[56375]= 1778631892;
assign addr[56376]= 1589734894;
assign addr[56377]= 1368621831;
assign addr[56378]= 1119773573;
assign addr[56379]= 848233042;
assign addr[56380]= 559503022;
assign addr[56381]= 259434643;
assign addr[56382]= -45891193;
assign addr[56383]= -350287041;
assign addr[56384]= -647584304;
assign addr[56385]= -931758235;
assign addr[56386]= -1197050035;
assign addr[56387]= -1438083551;
assign addr[56388]= -1649974225;
assign addr[56389]= -1828428082;
assign addr[56390]= -1969828744;
assign addr[56391]= -2071310720;
assign addr[56392]= -2130817471;
assign addr[56393]= -2147143090;
assign addr[56394]= -2119956737;
assign addr[56395]= -2049809346;
assign addr[56396]= -1938122457;
assign addr[56397]= -1787159411;
assign addr[56398]= -1599979481;
assign addr[56399]= -1380375881;
assign addr[56400]= -1132798888;
assign addr[56401]= -862265664;
assign addr[56402]= -574258580;
assign addr[56403]= -274614114;
assign addr[56404]= 30595422;
assign addr[56405]= 335184940;
assign addr[56406]= 632981917;
assign addr[56407]= 917951481;
assign addr[56408]= 1184318708;
assign addr[56409]= 1426685652;
assign addr[56410]= 1640140734;
assign addr[56411]= 1820358275;
assign addr[56412]= 1963686155;
assign addr[56413]= 2067219829;
assign addr[56414]= 2128861181;
assign addr[56415]= 2147361045;
assign addr[56416]= 2122344521;
assign addr[56417]= 2054318569;
assign addr[56418]= 1944661739;
assign addr[56419]= 1795596234;
assign addr[56420]= 1610142873;
assign addr[56421]= 1392059879;
assign addr[56422]= 1145766716;
assign addr[56423]= 876254528;
assign addr[56424]= 588984994;
assign addr[56425]= 289779648;
assign addr[56426]= -15298099;
assign addr[56427]= -320065829;
assign addr[56428]= -618347408;
assign addr[56429]= -904098143;
assign addr[56430]= -1171527280;
assign addr[56431]= -1415215352;
assign addr[56432]= -1630224009;
assign addr[56433]= -1812196087;
assign addr[56434]= -1957443913;
assign addr[56435]= -2063024031;
assign addr[56436]= -2126796855;
assign addr[56437]= -2147470025;
assign addr[56438]= -2124624598;
assign addr[56439]= -2058723538;
assign addr[56440]= -1951102334;
assign addr[56441]= -1803941934;
assign addr[56442]= -1620224553;
assign addr[56443]= -1403673233;
assign addr[56444]= -1158676398;
assign addr[56445]= -890198924;
assign addr[56446]= -603681519;
assign addr[56447]= -304930476;
assign addr[56448]= 0;
assign addr[56449]= 304930476;
assign addr[56450]= 603681519;
assign addr[56451]= 890198924;
assign addr[56452]= 1158676398;
assign addr[56453]= 1403673233;
assign addr[56454]= 1620224553;
assign addr[56455]= 1803941934;
assign addr[56456]= 1951102334;
assign addr[56457]= 2058723538;
assign addr[56458]= 2124624598;
assign addr[56459]= 2147470025;
assign addr[56460]= 2126796855;
assign addr[56461]= 2063024031;
assign addr[56462]= 1957443913;
assign addr[56463]= 1812196087;
assign addr[56464]= 1630224009;
assign addr[56465]= 1415215352;
assign addr[56466]= 1171527280;
assign addr[56467]= 904098143;
assign addr[56468]= 618347408;
assign addr[56469]= 320065829;
assign addr[56470]= 15298099;
assign addr[56471]= -289779648;
assign addr[56472]= -588984994;
assign addr[56473]= -876254528;
assign addr[56474]= -1145766716;
assign addr[56475]= -1392059879;
assign addr[56476]= -1610142873;
assign addr[56477]= -1795596234;
assign addr[56478]= -1944661739;
assign addr[56479]= -2054318569;
assign addr[56480]= -2122344521;
assign addr[56481]= -2147361045;
assign addr[56482]= -2128861181;
assign addr[56483]= -2067219829;
assign addr[56484]= -1963686155;
assign addr[56485]= -1820358275;
assign addr[56486]= -1640140734;
assign addr[56487]= -1426685652;
assign addr[56488]= -1184318708;
assign addr[56489]= -917951481;
assign addr[56490]= -632981917;
assign addr[56491]= -335184940;
assign addr[56492]= -30595422;
assign addr[56493]= 274614114;
assign addr[56494]= 574258580;
assign addr[56495]= 862265664;
assign addr[56496]= 1132798888;
assign addr[56497]= 1380375881;
assign addr[56498]= 1599979481;
assign addr[56499]= 1787159411;
assign addr[56500]= 1938122457;
assign addr[56501]= 2049809346;
assign addr[56502]= 2119956737;
assign addr[56503]= 2147143090;
assign addr[56504]= 2130817471;
assign addr[56505]= 2071310720;
assign addr[56506]= 1969828744;
assign addr[56507]= 1828428082;
assign addr[56508]= 1649974225;
assign addr[56509]= 1438083551;
assign addr[56510]= 1197050035;
assign addr[56511]= 931758235;
assign addr[56512]= 647584304;
assign addr[56513]= 350287041;
assign addr[56514]= 45891193;
assign addr[56515]= -259434643;
assign addr[56516]= -559503022;
assign addr[56517]= -848233042;
assign addr[56518]= -1119773573;
assign addr[56519]= -1368621831;
assign addr[56520]= -1589734894;
assign addr[56521]= -1778631892;
assign addr[56522]= -1931484818;
assign addr[56523]= -2045196100;
assign addr[56524]= -2117461370;
assign addr[56525]= -2146816171;
assign addr[56526]= -2132665626;
assign addr[56527]= -2075296495;
assign addr[56528]= -1975871368;
assign addr[56529]= -1836405100;
assign addr[56530]= -1659723983;
assign addr[56531]= -1449408469;
assign addr[56532]= -1209720613;
assign addr[56533]= -945517704;
assign addr[56534]= -662153826;
assign addr[56535]= -365371365;
assign addr[56536]= -61184634;
assign addr[56537]= 244242007;
assign addr[56538]= 544719071;
assign addr[56539]= 834157373;
assign addr[56540]= 1106691431;
assign addr[56541]= 1356798326;
assign addr[56542]= 1579409630;
assign addr[56543]= 1770014111;
assign addr[56544]= 1924749160;
assign addr[56545]= 2040479063;
assign addr[56546]= 2114858546;
assign addr[56547]= 2146380306;
assign addr[56548]= 2134405552;
assign addr[56549]= 2079176953;
assign addr[56550]= 1981813720;
assign addr[56551]= 1844288924;
assign addr[56552]= 1669389513;
assign addr[56553]= 1460659832;
assign addr[56554]= 1222329801;
assign addr[56555]= 959229189;
assign addr[56556]= 676689746;
assign addr[56557]= 380437148;
assign addr[56558]= 76474970;
assign addr[56559]= -229036977;
assign addr[56560]= -529907477;
assign addr[56561]= -820039373;
assign addr[56562]= -1093553126;
assign addr[56563]= -1344905966;
assign addr[56564]= -1569004214;
assign addr[56565]= -1761306505;
assign addr[56566]= -1917915825;
assign addr[56567]= -2035658475;
assign addr[56568]= -2112148396;
assign addr[56569]= -2145835515;
assign addr[56570]= -2136037160;
assign addr[56571]= -2082951896;
assign addr[56572]= -1987655498;
assign addr[56573]= -1852079154;
assign addr[56574]= -1678970324;
assign addr[56575]= -1471837070;
assign addr[56576]= -1234876957;
assign addr[56577]= -972891995;
assign addr[56578]= -691191324;
assign addr[56579]= -395483624;
assign addr[56580]= -91761426;
assign addr[56581]= 213820322;
assign addr[56582]= 515068990;
assign addr[56583]= 805879757;
assign addr[56584]= 1080359326;
assign addr[56585]= 1332945355;
assign addr[56586]= 1558519173;
assign addr[56587]= 1752509516;
assign addr[56588]= 1910985158;
assign addr[56589]= 2030734582;
assign addr[56590]= 2109331059;
assign addr[56591]= 2145181827;
assign addr[56592]= 2137560369;
assign addr[56593]= 2086621133;
assign addr[56594]= 1993396407;
assign addr[56595]= 1859775393;
assign addr[56596]= 1688465931;
assign addr[56597]= 1482939614;
assign addr[56598]= 1247361445;
assign addr[56599]= 986505429;
assign addr[56600]= 705657826;
assign addr[56601]= 410510029;
assign addr[56602]= 107043224;
assign addr[56603]= -198592817;
assign addr[56604]= -500204365;
assign addr[56605]= -791679244;
assign addr[56606]= -1067110699;
assign addr[56607]= -1320917099;
assign addr[56608]= -1547955041;
assign addr[56609]= -1743623590;
assign addr[56610]= -1903957513;
assign addr[56611]= -2025707632;
assign addr[56612]= -2106406677;
assign addr[56613]= -2144419275;
assign addr[56614]= -2138975100;
assign addr[56615]= -2090184478;
assign addr[56616]= -1999036154;
assign addr[56617]= -1867377253;
assign addr[56618]= -1697875851;
assign addr[56619]= -1493966902;
assign addr[56620]= -1259782632;
assign addr[56621]= -1000068799;
assign addr[56622]= -720088517;
assign addr[56623]= -425515602;
assign addr[56624]= -122319591;
assign addr[56625]= 183355234;
assign addr[56626]= 485314355;
assign addr[56627]= 777438554;
assign addr[56628]= 1053807919;
assign addr[56629]= 1308821808;
assign addr[56630]= 1537312353;
assign addr[56631]= 1734649179;
assign addr[56632]= 1896833245;
assign addr[56633]= 2020577882;
assign addr[56634]= 2103375398;
assign addr[56635]= 2143547897;
assign addr[56636]= 2140281282;
assign addr[56637]= 2093641749;
assign addr[56638]= 2004574453;
assign addr[56639]= 1874884346;
assign addr[56640]= 1707199606;
assign addr[56641]= 1504918373;
assign addr[56642]= 1272139887;
assign addr[56643]= 1013581418;
assign addr[56644]= 734482665;
assign addr[56645]= 440499581;
assign addr[56646]= 137589750;
assign addr[56647]= -168108346;
assign addr[56648]= -470399716;
assign addr[56649]= -763158411;
assign addr[56650]= -1040451659;
assign addr[56651]= -1296660098;
assign addr[56652]= -1526591649;
assign addr[56653]= -1725586737;
assign addr[56654]= -1889612716;
assign addr[56655]= -2015345591;
assign addr[56656]= -2100237377;
assign addr[56657]= -2142567738;
assign addr[56658]= -2141478848;
assign addr[56659]= -2096992772;
assign addr[56660]= -2010011024;
assign addr[56661]= -1882296293;
assign addr[56662]= -1716436725;
assign addr[56663]= -1515793473;
assign addr[56664]= -1284432584;
assign addr[56665]= -1027042599;
assign addr[56666]= -748839539;
assign addr[56667]= -455461206;
assign addr[56668]= -152852926;
assign addr[56669]= 152852926;
assign addr[56670]= 455461206;
assign addr[56671]= 748839539;
assign addr[56672]= 1027042599;
assign addr[56673]= 1284432584;
assign addr[56674]= 1515793473;
assign addr[56675]= 1716436725;
assign addr[56676]= 1882296293;
assign addr[56677]= 2010011024;
assign addr[56678]= 2096992772;
assign addr[56679]= 2141478848;
assign addr[56680]= 2142567738;
assign addr[56681]= 2100237377;
assign addr[56682]= 2015345591;
assign addr[56683]= 1889612716;
assign addr[56684]= 1725586737;
assign addr[56685]= 1526591649;
assign addr[56686]= 1296660098;
assign addr[56687]= 1040451659;
assign addr[56688]= 763158411;
assign addr[56689]= 470399716;
assign addr[56690]= 168108346;
assign addr[56691]= -137589750;
assign addr[56692]= -440499581;
assign addr[56693]= -734482665;
assign addr[56694]= -1013581418;
assign addr[56695]= -1272139887;
assign addr[56696]= -1504918373;
assign addr[56697]= -1707199606;
assign addr[56698]= -1874884346;
assign addr[56699]= -2004574453;
assign addr[56700]= -2093641749;
assign addr[56701]= -2140281282;
assign addr[56702]= -2143547897;
assign addr[56703]= -2103375398;
assign addr[56704]= -2020577882;
assign addr[56705]= -1896833245;
assign addr[56706]= -1734649179;
assign addr[56707]= -1537312353;
assign addr[56708]= -1308821808;
assign addr[56709]= -1053807919;
assign addr[56710]= -777438554;
assign addr[56711]= -485314355;
assign addr[56712]= -183355234;
assign addr[56713]= 122319591;
assign addr[56714]= 425515602;
assign addr[56715]= 720088517;
assign addr[56716]= 1000068799;
assign addr[56717]= 1259782632;
assign addr[56718]= 1493966902;
assign addr[56719]= 1697875851;
assign addr[56720]= 1867377253;
assign addr[56721]= 1999036154;
assign addr[56722]= 2090184478;
assign addr[56723]= 2138975100;
assign addr[56724]= 2144419275;
assign addr[56725]= 2106406677;
assign addr[56726]= 2025707632;
assign addr[56727]= 1903957513;
assign addr[56728]= 1743623590;
assign addr[56729]= 1547955041;
assign addr[56730]= 1320917099;
assign addr[56731]= 1067110699;
assign addr[56732]= 791679244;
assign addr[56733]= 500204365;
assign addr[56734]= 198592817;
assign addr[56735]= -107043224;
assign addr[56736]= -410510029;
assign addr[56737]= -705657826;
assign addr[56738]= -986505429;
assign addr[56739]= -1247361445;
assign addr[56740]= -1482939614;
assign addr[56741]= -1688465931;
assign addr[56742]= -1859775393;
assign addr[56743]= -1993396407;
assign addr[56744]= -2086621133;
assign addr[56745]= -2137560369;
assign addr[56746]= -2145181827;
assign addr[56747]= -2109331059;
assign addr[56748]= -2030734582;
assign addr[56749]= -1910985158;
assign addr[56750]= -1752509516;
assign addr[56751]= -1558519173;
assign addr[56752]= -1332945355;
assign addr[56753]= -1080359326;
assign addr[56754]= -805879757;
assign addr[56755]= -515068990;
assign addr[56756]= -213820322;
assign addr[56757]= 91761426;
assign addr[56758]= 395483624;
assign addr[56759]= 691191324;
assign addr[56760]= 972891995;
assign addr[56761]= 1234876957;
assign addr[56762]= 1471837070;
assign addr[56763]= 1678970324;
assign addr[56764]= 1852079154;
assign addr[56765]= 1987655498;
assign addr[56766]= 2082951896;
assign addr[56767]= 2136037160;
assign addr[56768]= 2145835515;
assign addr[56769]= 2112148396;
assign addr[56770]= 2035658475;
assign addr[56771]= 1917915825;
assign addr[56772]= 1761306505;
assign addr[56773]= 1569004214;
assign addr[56774]= 1344905966;
assign addr[56775]= 1093553126;
assign addr[56776]= 820039373;
assign addr[56777]= 529907477;
assign addr[56778]= 229036977;
assign addr[56779]= -76474970;
assign addr[56780]= -380437148;
assign addr[56781]= -676689746;
assign addr[56782]= -959229189;
assign addr[56783]= -1222329801;
assign addr[56784]= -1460659832;
assign addr[56785]= -1669389513;
assign addr[56786]= -1844288924;
assign addr[56787]= -1981813720;
assign addr[56788]= -2079176953;
assign addr[56789]= -2134405552;
assign addr[56790]= -2146380306;
assign addr[56791]= -2114858546;
assign addr[56792]= -2040479063;
assign addr[56793]= -1924749160;
assign addr[56794]= -1770014111;
assign addr[56795]= -1579409630;
assign addr[56796]= -1356798326;
assign addr[56797]= -1106691431;
assign addr[56798]= -834157373;
assign addr[56799]= -544719071;
assign addr[56800]= -244242007;
assign addr[56801]= 61184634;
assign addr[56802]= 365371365;
assign addr[56803]= 662153826;
assign addr[56804]= 945517704;
assign addr[56805]= 1209720613;
assign addr[56806]= 1449408469;
assign addr[56807]= 1659723983;
assign addr[56808]= 1836405100;
assign addr[56809]= 1975871368;
assign addr[56810]= 2075296495;
assign addr[56811]= 2132665626;
assign addr[56812]= 2146816171;
assign addr[56813]= 2117461370;
assign addr[56814]= 2045196100;
assign addr[56815]= 1931484818;
assign addr[56816]= 1778631892;
assign addr[56817]= 1589734894;
assign addr[56818]= 1368621831;
assign addr[56819]= 1119773573;
assign addr[56820]= 848233042;
assign addr[56821]= 559503022;
assign addr[56822]= 259434643;
assign addr[56823]= -45891193;
assign addr[56824]= -350287041;
assign addr[56825]= -647584304;
assign addr[56826]= -931758235;
assign addr[56827]= -1197050035;
assign addr[56828]= -1438083551;
assign addr[56829]= -1649974225;
assign addr[56830]= -1828428082;
assign addr[56831]= -1969828744;
assign addr[56832]= -2071310720;
assign addr[56833]= -2130817471;
assign addr[56834]= -2147143090;
assign addr[56835]= -2119956737;
assign addr[56836]= -2049809346;
assign addr[56837]= -1938122457;
assign addr[56838]= -1787159411;
assign addr[56839]= -1599979481;
assign addr[56840]= -1380375881;
assign addr[56841]= -1132798888;
assign addr[56842]= -862265664;
assign addr[56843]= -574258580;
assign addr[56844]= -274614114;
assign addr[56845]= 30595422;
assign addr[56846]= 335184940;
assign addr[56847]= 632981917;
assign addr[56848]= 917951481;
assign addr[56849]= 1184318708;
assign addr[56850]= 1426685652;
assign addr[56851]= 1640140734;
assign addr[56852]= 1820358275;
assign addr[56853]= 1963686155;
assign addr[56854]= 2067219829;
assign addr[56855]= 2128861181;
assign addr[56856]= 2147361045;
assign addr[56857]= 2122344521;
assign addr[56858]= 2054318569;
assign addr[56859]= 1944661739;
assign addr[56860]= 1795596234;
assign addr[56861]= 1610142873;
assign addr[56862]= 1392059879;
assign addr[56863]= 1145766716;
assign addr[56864]= 876254528;
assign addr[56865]= 588984994;
assign addr[56866]= 289779648;
assign addr[56867]= -15298099;
assign addr[56868]= -320065829;
assign addr[56869]= -618347408;
assign addr[56870]= -904098143;
assign addr[56871]= -1171527280;
assign addr[56872]= -1415215352;
assign addr[56873]= -1630224009;
assign addr[56874]= -1812196087;
assign addr[56875]= -1957443913;
assign addr[56876]= -2063024031;
assign addr[56877]= -2126796855;
assign addr[56878]= -2147470025;
assign addr[56879]= -2124624598;
assign addr[56880]= -2058723538;
assign addr[56881]= -1951102334;
assign addr[56882]= -1803941934;
assign addr[56883]= -1620224553;
assign addr[56884]= -1403673233;
assign addr[56885]= -1158676398;
assign addr[56886]= -890198924;
assign addr[56887]= -603681519;
assign addr[56888]= -304930476;
assign addr[56889]= 0;
assign addr[56890]= 304930476;
assign addr[56891]= 603681519;
assign addr[56892]= 890198924;
assign addr[56893]= 1158676398;
assign addr[56894]= 1403673233;
assign addr[56895]= 1620224553;
assign addr[56896]= 1803941934;
assign addr[56897]= 1951102334;
assign addr[56898]= 2058723538;
assign addr[56899]= 2124624598;
assign addr[56900]= 2147470025;
assign addr[56901]= 2126796855;
assign addr[56902]= 2063024031;
assign addr[56903]= 1957443913;
assign addr[56904]= 1812196087;
assign addr[56905]= 1630224009;
assign addr[56906]= 1415215352;
assign addr[56907]= 1171527280;
assign addr[56908]= 904098143;
assign addr[56909]= 618347408;
assign addr[56910]= 320065829;
assign addr[56911]= 15298099;
assign addr[56912]= -289779648;
assign addr[56913]= -588984994;
assign addr[56914]= -876254528;
assign addr[56915]= -1145766716;
assign addr[56916]= -1392059879;
assign addr[56917]= -1610142873;
assign addr[56918]= -1795596234;
assign addr[56919]= -1944661739;
assign addr[56920]= -2054318569;
assign addr[56921]= -2122344521;
assign addr[56922]= -2147361045;
assign addr[56923]= -2128861181;
assign addr[56924]= -2067219829;
assign addr[56925]= -1963686155;
assign addr[56926]= -1820358275;
assign addr[56927]= -1640140734;
assign addr[56928]= -1426685652;
assign addr[56929]= -1184318708;
assign addr[56930]= -917951481;
assign addr[56931]= -632981917;
assign addr[56932]= -335184940;
assign addr[56933]= -30595422;
assign addr[56934]= 274614114;
assign addr[56935]= 574258580;
assign addr[56936]= 862265664;
assign addr[56937]= 1132798888;
assign addr[56938]= 1380375881;
assign addr[56939]= 1599979481;
assign addr[56940]= 1787159411;
assign addr[56941]= 1938122457;
assign addr[56942]= 2049809346;
assign addr[56943]= 2119956737;
assign addr[56944]= 2147143090;
assign addr[56945]= 2130817471;
assign addr[56946]= 2071310720;
assign addr[56947]= 1969828744;
assign addr[56948]= 1828428082;
assign addr[56949]= 1649974225;
assign addr[56950]= 1438083551;
assign addr[56951]= 1197050035;
assign addr[56952]= 931758235;
assign addr[56953]= 647584304;
assign addr[56954]= 350287041;
assign addr[56955]= 45891193;
assign addr[56956]= -259434643;
assign addr[56957]= -559503022;
assign addr[56958]= -848233042;
assign addr[56959]= -1119773573;
assign addr[56960]= -1368621831;
assign addr[56961]= -1589734894;
assign addr[56962]= -1778631892;
assign addr[56963]= -1931484818;
assign addr[56964]= -2045196100;
assign addr[56965]= -2117461370;
assign addr[56966]= -2146816171;
assign addr[56967]= -2132665626;
assign addr[56968]= -2075296495;
assign addr[56969]= -1975871368;
assign addr[56970]= -1836405100;
assign addr[56971]= -1659723983;
assign addr[56972]= -1449408469;
assign addr[56973]= -1209720613;
assign addr[56974]= -945517704;
assign addr[56975]= -662153826;
assign addr[56976]= -365371365;
assign addr[56977]= -61184634;
assign addr[56978]= 244242007;
assign addr[56979]= 544719071;
assign addr[56980]= 834157373;
assign addr[56981]= 1106691431;
assign addr[56982]= 1356798326;
assign addr[56983]= 1579409630;
assign addr[56984]= 1770014111;
assign addr[56985]= 1924749160;
assign addr[56986]= 2040479063;
assign addr[56987]= 2114858546;
assign addr[56988]= 2146380306;
assign addr[56989]= 2134405552;
assign addr[56990]= 2079176953;
assign addr[56991]= 1981813720;
assign addr[56992]= 1844288924;
assign addr[56993]= 1669389513;
assign addr[56994]= 1460659832;
assign addr[56995]= 1222329801;
assign addr[56996]= 959229189;
assign addr[56997]= 676689746;
assign addr[56998]= 380437148;
assign addr[56999]= 76474970;
assign addr[57000]= -229036977;
assign addr[57001]= -529907477;
assign addr[57002]= -820039373;
assign addr[57003]= -1093553126;
assign addr[57004]= -1344905966;
assign addr[57005]= -1569004214;
assign addr[57006]= -1761306505;
assign addr[57007]= -1917915825;
assign addr[57008]= -2035658475;
assign addr[57009]= -2112148396;
assign addr[57010]= -2145835515;
assign addr[57011]= -2136037160;
assign addr[57012]= -2082951896;
assign addr[57013]= -1987655498;
assign addr[57014]= -1852079154;
assign addr[57015]= -1678970324;
assign addr[57016]= -1471837070;
assign addr[57017]= -1234876957;
assign addr[57018]= -972891995;
assign addr[57019]= -691191324;
assign addr[57020]= -395483624;
assign addr[57021]= -91761426;
assign addr[57022]= 213820322;
assign addr[57023]= 515068990;
assign addr[57024]= 805879757;
assign addr[57025]= 1080359326;
assign addr[57026]= 1332945355;
assign addr[57027]= 1558519173;
assign addr[57028]= 1752509516;
assign addr[57029]= 1910985158;
assign addr[57030]= 2030734582;
assign addr[57031]= 2109331059;
assign addr[57032]= 2145181827;
assign addr[57033]= 2137560369;
assign addr[57034]= 2086621133;
assign addr[57035]= 1993396407;
assign addr[57036]= 1859775393;
assign addr[57037]= 1688465931;
assign addr[57038]= 1482939614;
assign addr[57039]= 1247361445;
assign addr[57040]= 986505429;
assign addr[57041]= 705657826;
assign addr[57042]= 410510029;
assign addr[57043]= 107043224;
assign addr[57044]= -198592817;
assign addr[57045]= -500204365;
assign addr[57046]= -791679244;
assign addr[57047]= -1067110699;
assign addr[57048]= -1320917099;
assign addr[57049]= -1547955041;
assign addr[57050]= -1743623590;
assign addr[57051]= -1903957513;
assign addr[57052]= -2025707632;
assign addr[57053]= -2106406677;
assign addr[57054]= -2144419275;
assign addr[57055]= -2138975100;
assign addr[57056]= -2090184478;
assign addr[57057]= -1999036154;
assign addr[57058]= -1867377253;
assign addr[57059]= -1697875851;
assign addr[57060]= -1493966902;
assign addr[57061]= -1259782632;
assign addr[57062]= -1000068799;
assign addr[57063]= -720088517;
assign addr[57064]= -425515602;
assign addr[57065]= -122319591;
assign addr[57066]= 183355234;
assign addr[57067]= 485314355;
assign addr[57068]= 777438554;
assign addr[57069]= 1053807919;
assign addr[57070]= 1308821808;
assign addr[57071]= 1537312353;
assign addr[57072]= 1734649179;
assign addr[57073]= 1896833245;
assign addr[57074]= 2020577882;
assign addr[57075]= 2103375398;
assign addr[57076]= 2143547897;
assign addr[57077]= 2140281282;
assign addr[57078]= 2093641749;
assign addr[57079]= 2004574453;
assign addr[57080]= 1874884346;
assign addr[57081]= 1707199606;
assign addr[57082]= 1504918373;
assign addr[57083]= 1272139887;
assign addr[57084]= 1013581418;
assign addr[57085]= 734482665;
assign addr[57086]= 440499581;
assign addr[57087]= 137589750;
assign addr[57088]= -168108346;
assign addr[57089]= -470399716;
assign addr[57090]= -763158411;
assign addr[57091]= -1040451659;
assign addr[57092]= -1296660098;
assign addr[57093]= -1526591649;
assign addr[57094]= -1725586737;
assign addr[57095]= -1889612716;
assign addr[57096]= -2015345591;
assign addr[57097]= -2100237377;
assign addr[57098]= -2142567738;
assign addr[57099]= -2141478848;
assign addr[57100]= -2096992772;
assign addr[57101]= -2010011024;
assign addr[57102]= -1882296293;
assign addr[57103]= -1716436725;
assign addr[57104]= -1515793473;
assign addr[57105]= -1284432584;
assign addr[57106]= -1027042599;
assign addr[57107]= -748839539;
assign addr[57108]= -455461206;
assign addr[57109]= -152852926;
assign addr[57110]= 152852926;
assign addr[57111]= 455461206;
assign addr[57112]= 748839539;
assign addr[57113]= 1027042599;
assign addr[57114]= 1284432584;
assign addr[57115]= 1515793473;
assign addr[57116]= 1716436725;
assign addr[57117]= 1882296293;
assign addr[57118]= 2010011024;
assign addr[57119]= 2096992772;
assign addr[57120]= 2141478848;
assign addr[57121]= 2142567738;
assign addr[57122]= 2100237377;
assign addr[57123]= 2015345591;
assign addr[57124]= 1889612716;
assign addr[57125]= 1725586737;
assign addr[57126]= 1526591649;
assign addr[57127]= 1296660098;
assign addr[57128]= 1040451659;
assign addr[57129]= 763158411;
assign addr[57130]= 470399716;
assign addr[57131]= 168108346;
assign addr[57132]= -137589750;
assign addr[57133]= -440499581;
assign addr[57134]= -734482665;
assign addr[57135]= -1013581418;
assign addr[57136]= -1272139887;
assign addr[57137]= -1504918373;
assign addr[57138]= -1707199606;
assign addr[57139]= -1874884346;
assign addr[57140]= -2004574453;
assign addr[57141]= -2093641749;
assign addr[57142]= -2140281282;
assign addr[57143]= -2143547897;
assign addr[57144]= -2103375398;
assign addr[57145]= -2020577882;
assign addr[57146]= -1896833245;
assign addr[57147]= -1734649179;
assign addr[57148]= -1537312353;
assign addr[57149]= -1308821808;
assign addr[57150]= -1053807919;
assign addr[57151]= -777438554;
assign addr[57152]= -485314355;
assign addr[57153]= -183355234;
assign addr[57154]= 122319591;
assign addr[57155]= 425515602;
assign addr[57156]= 720088517;
assign addr[57157]= 1000068799;
assign addr[57158]= 1259782632;
assign addr[57159]= 1493966902;
assign addr[57160]= 1697875851;
assign addr[57161]= 1867377253;
assign addr[57162]= 1999036154;
assign addr[57163]= 2090184478;
assign addr[57164]= 2138975100;
assign addr[57165]= 2144419275;
assign addr[57166]= 2106406677;
assign addr[57167]= 2025707632;
assign addr[57168]= 1903957513;
assign addr[57169]= 1743623590;
assign addr[57170]= 1547955041;
assign addr[57171]= 1320917099;
assign addr[57172]= 1067110699;
assign addr[57173]= 791679244;
assign addr[57174]= 500204365;
assign addr[57175]= 198592817;
assign addr[57176]= -107043224;
assign addr[57177]= -410510029;
assign addr[57178]= -705657826;
assign addr[57179]= -986505429;
assign addr[57180]= -1247361445;
assign addr[57181]= -1482939614;
assign addr[57182]= -1688465931;
assign addr[57183]= -1859775393;
assign addr[57184]= -1993396407;
assign addr[57185]= -2086621133;
assign addr[57186]= -2137560369;
assign addr[57187]= -2145181827;
assign addr[57188]= -2109331059;
assign addr[57189]= -2030734582;
assign addr[57190]= -1910985158;
assign addr[57191]= -1752509516;
assign addr[57192]= -1558519173;
assign addr[57193]= -1332945355;
assign addr[57194]= -1080359326;
assign addr[57195]= -805879757;
assign addr[57196]= -515068990;
assign addr[57197]= -213820322;
assign addr[57198]= 91761426;
assign addr[57199]= 395483624;
assign addr[57200]= 691191324;
assign addr[57201]= 972891995;
assign addr[57202]= 1234876957;
assign addr[57203]= 1471837070;
assign addr[57204]= 1678970324;
assign addr[57205]= 1852079154;
assign addr[57206]= 1987655498;
assign addr[57207]= 2082951896;
assign addr[57208]= 2136037160;
assign addr[57209]= 2145835515;
assign addr[57210]= 2112148396;
assign addr[57211]= 2035658475;
assign addr[57212]= 1917915825;
assign addr[57213]= 1761306505;
assign addr[57214]= 1569004214;
assign addr[57215]= 1344905966;
assign addr[57216]= 1093553126;
assign addr[57217]= 820039373;
assign addr[57218]= 529907477;
assign addr[57219]= 229036977;
assign addr[57220]= -76474970;
assign addr[57221]= -380437148;
assign addr[57222]= -676689746;
assign addr[57223]= -959229189;
assign addr[57224]= -1222329801;
assign addr[57225]= -1460659832;
assign addr[57226]= -1669389513;
assign addr[57227]= -1844288924;
assign addr[57228]= -1981813720;
assign addr[57229]= -2079176953;
assign addr[57230]= -2134405552;
assign addr[57231]= -2146380306;
assign addr[57232]= -2114858546;
assign addr[57233]= -2040479063;
assign addr[57234]= -1924749160;
assign addr[57235]= -1770014111;
assign addr[57236]= -1579409630;
assign addr[57237]= -1356798326;
assign addr[57238]= -1106691431;
assign addr[57239]= -834157373;
assign addr[57240]= -544719071;
assign addr[57241]= -244242007;
assign addr[57242]= 61184634;
assign addr[57243]= 365371365;
assign addr[57244]= 662153826;
assign addr[57245]= 945517704;
assign addr[57246]= 1209720613;
assign addr[57247]= 1449408469;
assign addr[57248]= 1659723983;
assign addr[57249]= 1836405100;
assign addr[57250]= 1975871368;
assign addr[57251]= 2075296495;
assign addr[57252]= 2132665626;
assign addr[57253]= 2146816171;
assign addr[57254]= 2117461370;
assign addr[57255]= 2045196100;
assign addr[57256]= 1931484818;
assign addr[57257]= 1778631892;
assign addr[57258]= 1589734894;
assign addr[57259]= 1368621831;
assign addr[57260]= 1119773573;
assign addr[57261]= 848233042;
assign addr[57262]= 559503022;
assign addr[57263]= 259434643;
assign addr[57264]= -45891193;
assign addr[57265]= -350287041;
assign addr[57266]= -647584304;
assign addr[57267]= -931758235;
assign addr[57268]= -1197050035;
assign addr[57269]= -1438083551;
assign addr[57270]= -1649974225;
assign addr[57271]= -1828428082;
assign addr[57272]= -1969828744;
assign addr[57273]= -2071310720;
assign addr[57274]= -2130817471;
assign addr[57275]= -2147143090;
assign addr[57276]= -2119956737;
assign addr[57277]= -2049809346;
assign addr[57278]= -1938122457;
assign addr[57279]= -1787159411;
assign addr[57280]= -1599979481;
assign addr[57281]= -1380375881;
assign addr[57282]= -1132798888;
assign addr[57283]= -862265664;
assign addr[57284]= -574258580;
assign addr[57285]= -274614114;
assign addr[57286]= 30595422;
assign addr[57287]= 335184940;
assign addr[57288]= 632981917;
assign addr[57289]= 917951481;
assign addr[57290]= 1184318708;
assign addr[57291]= 1426685652;
assign addr[57292]= 1640140734;
assign addr[57293]= 1820358275;
assign addr[57294]= 1963686155;
assign addr[57295]= 2067219829;
assign addr[57296]= 2128861181;
assign addr[57297]= 2147361045;
assign addr[57298]= 2122344521;
assign addr[57299]= 2054318569;
assign addr[57300]= 1944661739;
assign addr[57301]= 1795596234;
assign addr[57302]= 1610142873;
assign addr[57303]= 1392059879;
assign addr[57304]= 1145766716;
assign addr[57305]= 876254528;
assign addr[57306]= 588984994;
assign addr[57307]= 289779648;
assign addr[57308]= -15298099;
assign addr[57309]= -320065829;
assign addr[57310]= -618347408;
assign addr[57311]= -904098143;
assign addr[57312]= -1171527280;
assign addr[57313]= -1415215352;
assign addr[57314]= -1630224009;
assign addr[57315]= -1812196087;
assign addr[57316]= -1957443913;
assign addr[57317]= -2063024031;
assign addr[57318]= -2126796855;
assign addr[57319]= -2147470025;
assign addr[57320]= -2124624598;
assign addr[57321]= -2058723538;
assign addr[57322]= -1951102334;
assign addr[57323]= -1803941934;
assign addr[57324]= -1620224553;
assign addr[57325]= -1403673233;
assign addr[57326]= -1158676398;
assign addr[57327]= -890198924;
assign addr[57328]= -603681519;
assign addr[57329]= -304930476;
assign addr[57330]= 0;
assign addr[57331]= 304930476;
assign addr[57332]= 603681519;
assign addr[57333]= 890198924;
assign addr[57334]= 1158676398;
assign addr[57335]= 1403673233;
assign addr[57336]= 1620224553;
assign addr[57337]= 1803941934;
assign addr[57338]= 1951102334;
assign addr[57339]= 2058723538;
assign addr[57340]= 2124624598;
assign addr[57341]= 2147470025;
assign addr[57342]= 2126796855;
assign addr[57343]= 2063024031;
assign addr[57344]= 1957443913;
assign addr[57345]= 1812196087;
assign addr[57346]= 1630224009;
assign addr[57347]= 1415215352;
assign addr[57348]= 1171527280;
assign addr[57349]= 904098143;
assign addr[57350]= 618347408;
assign addr[57351]= 320065829;
assign addr[57352]= 15298099;
assign addr[57353]= -289779648;
assign addr[57354]= -588984994;
assign addr[57355]= -876254528;
assign addr[57356]= -1145766716;
assign addr[57357]= -1392059879;
assign addr[57358]= -1610142873;
assign addr[57359]= -1795596234;
assign addr[57360]= -1944661739;
assign addr[57361]= -2054318569;
assign addr[57362]= -2122344521;
assign addr[57363]= -2147361045;
assign addr[57364]= -2128861181;
assign addr[57365]= -2067219829;
assign addr[57366]= -1963686155;
assign addr[57367]= -1820358275;
assign addr[57368]= -1640140734;
assign addr[57369]= -1426685652;
assign addr[57370]= -1184318708;
assign addr[57371]= -917951481;
assign addr[57372]= -632981917;
assign addr[57373]= -335184940;
assign addr[57374]= -30595422;
assign addr[57375]= 274614114;
assign addr[57376]= 574258580;
assign addr[57377]= 862265664;
assign addr[57378]= 1132798888;
assign addr[57379]= 1380375881;
assign addr[57380]= 1599979481;
assign addr[57381]= 1787159411;
assign addr[57382]= 1938122457;
assign addr[57383]= 2049809346;
assign addr[57384]= 2119956737;
assign addr[57385]= 2147143090;
assign addr[57386]= 2130817471;
assign addr[57387]= 2071310720;
assign addr[57388]= 1969828744;
assign addr[57389]= 1828428082;
assign addr[57390]= 1649974225;
assign addr[57391]= 1438083551;
assign addr[57392]= 1197050035;
assign addr[57393]= 931758235;
assign addr[57394]= 647584304;
assign addr[57395]= 350287041;
assign addr[57396]= 45891193;
assign addr[57397]= -259434643;
assign addr[57398]= -559503022;
assign addr[57399]= -848233042;
assign addr[57400]= -1119773573;
assign addr[57401]= -1368621831;
assign addr[57402]= -1589734894;
assign addr[57403]= -1778631892;
assign addr[57404]= -1931484818;
assign addr[57405]= -2045196100;
assign addr[57406]= -2117461370;
assign addr[57407]= -2146816171;
assign addr[57408]= -2132665626;
assign addr[57409]= -2075296495;
assign addr[57410]= -1975871368;
assign addr[57411]= -1836405100;
assign addr[57412]= -1659723983;
assign addr[57413]= -1449408469;
assign addr[57414]= -1209720613;
assign addr[57415]= -945517704;
assign addr[57416]= -662153826;
assign addr[57417]= -365371365;
assign addr[57418]= -61184634;
assign addr[57419]= 244242007;
assign addr[57420]= 544719071;
assign addr[57421]= 834157373;
assign addr[57422]= 1106691431;
assign addr[57423]= 1356798326;
assign addr[57424]= 1579409630;
assign addr[57425]= 1770014111;
assign addr[57426]= 1924749160;
assign addr[57427]= 2040479063;
assign addr[57428]= 2114858546;
assign addr[57429]= 2146380306;
assign addr[57430]= 2134405552;
assign addr[57431]= 2079176953;
assign addr[57432]= 1981813720;
assign addr[57433]= 1844288924;
assign addr[57434]= 1669389513;
assign addr[57435]= 1460659832;
assign addr[57436]= 1222329801;
assign addr[57437]= 959229189;
assign addr[57438]= 676689746;
assign addr[57439]= 380437148;
assign addr[57440]= 76474970;
assign addr[57441]= -229036977;
assign addr[57442]= -529907477;
assign addr[57443]= -820039373;
assign addr[57444]= -1093553126;
assign addr[57445]= -1344905966;
assign addr[57446]= -1569004214;
assign addr[57447]= -1761306505;
assign addr[57448]= -1917915825;
assign addr[57449]= -2035658475;
assign addr[57450]= -2112148396;
assign addr[57451]= -2145835515;
assign addr[57452]= -2136037160;
assign addr[57453]= -2082951896;
assign addr[57454]= -1987655498;
assign addr[57455]= -1852079154;
assign addr[57456]= -1678970324;
assign addr[57457]= -1471837070;
assign addr[57458]= -1234876957;
assign addr[57459]= -972891995;
assign addr[57460]= -691191324;
assign addr[57461]= -395483624;
assign addr[57462]= -91761426;
assign addr[57463]= 213820322;
assign addr[57464]= 515068990;
assign addr[57465]= 805879757;
assign addr[57466]= 1080359326;
assign addr[57467]= 1332945355;
assign addr[57468]= 1558519173;
assign addr[57469]= 1752509516;
assign addr[57470]= 1910985158;
assign addr[57471]= 2030734582;
assign addr[57472]= 2109331059;
assign addr[57473]= 2145181827;
assign addr[57474]= 2137560369;
assign addr[57475]= 2086621133;
assign addr[57476]= 1993396407;
assign addr[57477]= 1859775393;
assign addr[57478]= 1688465931;
assign addr[57479]= 1482939614;
assign addr[57480]= 1247361445;
assign addr[57481]= 986505429;
assign addr[57482]= 705657826;
assign addr[57483]= 410510029;
assign addr[57484]= 107043224;
assign addr[57485]= -198592817;
assign addr[57486]= -500204365;
assign addr[57487]= -791679244;
assign addr[57488]= -1067110699;
assign addr[57489]= -1320917099;
assign addr[57490]= -1547955041;
assign addr[57491]= -1743623590;
assign addr[57492]= -1903957513;
assign addr[57493]= -2025707632;
assign addr[57494]= -2106406677;
assign addr[57495]= -2144419275;
assign addr[57496]= -2138975100;
assign addr[57497]= -2090184478;
assign addr[57498]= -1999036154;
assign addr[57499]= -1867377253;
assign addr[57500]= -1697875851;
assign addr[57501]= -1493966902;
assign addr[57502]= -1259782632;
assign addr[57503]= -1000068799;
assign addr[57504]= -720088517;
assign addr[57505]= -425515602;
assign addr[57506]= -122319591;
assign addr[57507]= 183355234;
assign addr[57508]= 485314355;
assign addr[57509]= 777438554;
assign addr[57510]= 1053807919;
assign addr[57511]= 1308821808;
assign addr[57512]= 1537312353;
assign addr[57513]= 1734649179;
assign addr[57514]= 1896833245;
assign addr[57515]= 2020577882;
assign addr[57516]= 2103375398;
assign addr[57517]= 2143547897;
assign addr[57518]= 2140281282;
assign addr[57519]= 2093641749;
assign addr[57520]= 2004574453;
assign addr[57521]= 1874884346;
assign addr[57522]= 1707199606;
assign addr[57523]= 1504918373;
assign addr[57524]= 1272139887;
assign addr[57525]= 1013581418;
assign addr[57526]= 734482665;
assign addr[57527]= 440499581;
assign addr[57528]= 137589750;
assign addr[57529]= -168108346;
assign addr[57530]= -470399716;
assign addr[57531]= -763158411;
assign addr[57532]= -1040451659;
assign addr[57533]= -1296660098;
assign addr[57534]= -1526591649;
assign addr[57535]= -1725586737;
assign addr[57536]= -1889612716;
assign addr[57537]= -2015345591;
assign addr[57538]= -2100237377;
assign addr[57539]= -2142567738;
assign addr[57540]= -2141478848;
assign addr[57541]= -2096992772;
assign addr[57542]= -2010011024;
assign addr[57543]= -1882296293;
assign addr[57544]= -1716436725;
assign addr[57545]= -1515793473;
assign addr[57546]= -1284432584;
assign addr[57547]= -1027042599;
assign addr[57548]= -748839539;
assign addr[57549]= -455461206;
assign addr[57550]= -152852926;
assign addr[57551]= 152852926;
assign addr[57552]= 455461206;
assign addr[57553]= 748839539;
assign addr[57554]= 1027042599;
assign addr[57555]= 1284432584;
assign addr[57556]= 1515793473;
assign addr[57557]= 1716436725;
assign addr[57558]= 1882296293;
assign addr[57559]= 2010011024;
assign addr[57560]= 2096992772;
assign addr[57561]= 2141478848;
assign addr[57562]= 2142567738;
assign addr[57563]= 2100237377;
assign addr[57564]= 2015345591;
assign addr[57565]= 1889612716;
assign addr[57566]= 1725586737;
assign addr[57567]= 1526591649;
assign addr[57568]= 1296660098;
assign addr[57569]= 1040451659;
assign addr[57570]= 763158411;
assign addr[57571]= 470399716;
assign addr[57572]= 168108346;
assign addr[57573]= -137589750;
assign addr[57574]= -440499581;
assign addr[57575]= -734482665;
assign addr[57576]= -1013581418;
assign addr[57577]= -1272139887;
assign addr[57578]= -1504918373;
assign addr[57579]= -1707199606;
assign addr[57580]= -1874884346;
assign addr[57581]= -2004574453;
assign addr[57582]= -2093641749;
assign addr[57583]= -2140281282;
assign addr[57584]= -2143547897;
assign addr[57585]= -2103375398;
assign addr[57586]= -2020577882;
assign addr[57587]= -1896833245;
assign addr[57588]= -1734649179;
assign addr[57589]= -1537312353;
assign addr[57590]= -1308821808;
assign addr[57591]= -1053807919;
assign addr[57592]= -777438554;
assign addr[57593]= -485314355;
assign addr[57594]= -183355234;
assign addr[57595]= 122319591;
assign addr[57596]= 425515602;
assign addr[57597]= 720088517;
assign addr[57598]= 1000068799;
assign addr[57599]= 1259782632;
assign addr[57600]= 1493966902;
assign addr[57601]= 1697875851;
assign addr[57602]= 1867377253;
assign addr[57603]= 1999036154;
assign addr[57604]= 2090184478;
assign addr[57605]= 2138975100;
assign addr[57606]= 2144419275;
assign addr[57607]= 2106406677;
assign addr[57608]= 2025707632;
assign addr[57609]= 1903957513;
assign addr[57610]= 1743623590;
assign addr[57611]= 1547955041;
assign addr[57612]= 1320917099;
assign addr[57613]= 1067110699;
assign addr[57614]= 791679244;
assign addr[57615]= 500204365;
assign addr[57616]= 198592817;
assign addr[57617]= -107043224;
assign addr[57618]= -410510029;
assign addr[57619]= -705657826;
assign addr[57620]= -986505429;
assign addr[57621]= -1247361445;
assign addr[57622]= -1482939614;
assign addr[57623]= -1688465931;
assign addr[57624]= -1859775393;
assign addr[57625]= -1993396407;
assign addr[57626]= -2086621133;
assign addr[57627]= -2137560369;
assign addr[57628]= -2145181827;
assign addr[57629]= -2109331059;
assign addr[57630]= -2030734582;
assign addr[57631]= -1910985158;
assign addr[57632]= -1752509516;
assign addr[57633]= -1558519173;
assign addr[57634]= -1332945355;
assign addr[57635]= -1080359326;
assign addr[57636]= -805879757;
assign addr[57637]= -515068990;
assign addr[57638]= -213820322;
assign addr[57639]= 91761426;
assign addr[57640]= 395483624;
assign addr[57641]= 691191324;
assign addr[57642]= 972891995;
assign addr[57643]= 1234876957;
assign addr[57644]= 1471837070;
assign addr[57645]= 1678970324;
assign addr[57646]= 1852079154;
assign addr[57647]= 1987655498;
assign addr[57648]= 2082951896;
assign addr[57649]= 2136037160;
assign addr[57650]= 2145835515;
assign addr[57651]= 2112148396;
assign addr[57652]= 2035658475;
assign addr[57653]= 1917915825;
assign addr[57654]= 1761306505;
assign addr[57655]= 1569004214;
assign addr[57656]= 1344905966;
assign addr[57657]= 1093553126;
assign addr[57658]= 820039373;
assign addr[57659]= 529907477;
assign addr[57660]= 229036977;
assign addr[57661]= -76474970;
assign addr[57662]= -380437148;
assign addr[57663]= -676689746;
assign addr[57664]= -959229189;
assign addr[57665]= -1222329801;
assign addr[57666]= -1460659832;
assign addr[57667]= -1669389513;
assign addr[57668]= -1844288924;
assign addr[57669]= -1981813720;
assign addr[57670]= -2079176953;
assign addr[57671]= -2134405552;
assign addr[57672]= -2146380306;
assign addr[57673]= -2114858546;
assign addr[57674]= -2040479063;
assign addr[57675]= -1924749160;
assign addr[57676]= -1770014111;
assign addr[57677]= -1579409630;
assign addr[57678]= -1356798326;
assign addr[57679]= -1106691431;
assign addr[57680]= -834157373;
assign addr[57681]= -544719071;
assign addr[57682]= -244242007;
assign addr[57683]= 61184634;
assign addr[57684]= 365371365;
assign addr[57685]= 662153826;
assign addr[57686]= 945517704;
assign addr[57687]= 1209720613;
assign addr[57688]= 1449408469;
assign addr[57689]= 1659723983;
assign addr[57690]= 1836405100;
assign addr[57691]= 1975871368;
assign addr[57692]= 2075296495;
assign addr[57693]= 2132665626;
assign addr[57694]= 2146816171;
assign addr[57695]= 2117461370;
assign addr[57696]= 2045196100;
assign addr[57697]= 1931484818;
assign addr[57698]= 1778631892;
assign addr[57699]= 1589734894;
assign addr[57700]= 1368621831;
assign addr[57701]= 1119773573;
assign addr[57702]= 848233042;
assign addr[57703]= 559503022;
assign addr[57704]= 259434643;
assign addr[57705]= -45891193;
assign addr[57706]= -350287041;
assign addr[57707]= -647584304;
assign addr[57708]= -931758235;
assign addr[57709]= -1197050035;
assign addr[57710]= -1438083551;
assign addr[57711]= -1649974225;
assign addr[57712]= -1828428082;
assign addr[57713]= -1969828744;
assign addr[57714]= -2071310720;
assign addr[57715]= -2130817471;
assign addr[57716]= -2147143090;
assign addr[57717]= -2119956737;
assign addr[57718]= -2049809346;
assign addr[57719]= -1938122457;
assign addr[57720]= -1787159411;
assign addr[57721]= -1599979481;
assign addr[57722]= -1380375881;
assign addr[57723]= -1132798888;
assign addr[57724]= -862265664;
assign addr[57725]= -574258580;
assign addr[57726]= -274614114;
assign addr[57727]= 30595422;
assign addr[57728]= 335184940;
assign addr[57729]= 632981917;
assign addr[57730]= 917951481;
assign addr[57731]= 1184318708;
assign addr[57732]= 1426685652;
assign addr[57733]= 1640140734;
assign addr[57734]= 1820358275;
assign addr[57735]= 1963686155;
assign addr[57736]= 2067219829;
assign addr[57737]= 2128861181;
assign addr[57738]= 2147361045;
assign addr[57739]= 2122344521;
assign addr[57740]= 2054318569;
assign addr[57741]= 1944661739;
assign addr[57742]= 1795596234;
assign addr[57743]= 1610142873;
assign addr[57744]= 1392059879;
assign addr[57745]= 1145766716;
assign addr[57746]= 876254528;
assign addr[57747]= 588984994;
assign addr[57748]= 289779648;
assign addr[57749]= -15298099;
assign addr[57750]= -320065829;
assign addr[57751]= -618347408;
assign addr[57752]= -904098143;
assign addr[57753]= -1171527280;
assign addr[57754]= -1415215352;
assign addr[57755]= -1630224009;
assign addr[57756]= -1812196087;
assign addr[57757]= -1957443913;
assign addr[57758]= -2063024031;
assign addr[57759]= -2126796855;
assign addr[57760]= -2147470025;
assign addr[57761]= -2124624598;
assign addr[57762]= -2058723538;
assign addr[57763]= -1951102334;
assign addr[57764]= -1803941934;
assign addr[57765]= -1620224553;
assign addr[57766]= -1403673233;
assign addr[57767]= -1158676398;
assign addr[57768]= -890198924;
assign addr[57769]= -603681519;
assign addr[57770]= -304930476;
assign addr[57771]= 0;
assign addr[57772]= 304930476;
assign addr[57773]= 603681519;
assign addr[57774]= 890198924;
assign addr[57775]= 1158676398;
assign addr[57776]= 1403673233;
assign addr[57777]= 1620224553;
assign addr[57778]= 1803941934;
assign addr[57779]= 1951102334;
assign addr[57780]= 2058723538;
assign addr[57781]= 2124624598;
assign addr[57782]= 2147470025;
assign addr[57783]= 2126796855;
assign addr[57784]= 2063024031;
assign addr[57785]= 1957443913;
assign addr[57786]= 1812196087;
assign addr[57787]= 1630224009;
assign addr[57788]= 1415215352;
assign addr[57789]= 1171527280;
assign addr[57790]= 904098143;
assign addr[57791]= 618347408;
assign addr[57792]= 320065829;
assign addr[57793]= 15298099;
assign addr[57794]= -289779648;
assign addr[57795]= -588984994;
assign addr[57796]= -876254528;
assign addr[57797]= -1145766716;
assign addr[57798]= -1392059879;
assign addr[57799]= -1610142873;
assign addr[57800]= -1795596234;
assign addr[57801]= -1944661739;
assign addr[57802]= -2054318569;
assign addr[57803]= -2122344521;
assign addr[57804]= -2147361045;
assign addr[57805]= -2128861181;
assign addr[57806]= -2067219829;
assign addr[57807]= -1963686155;
assign addr[57808]= -1820358275;
assign addr[57809]= -1640140734;
assign addr[57810]= -1426685652;
assign addr[57811]= -1184318708;
assign addr[57812]= -917951481;
assign addr[57813]= -632981917;
assign addr[57814]= -335184940;
assign addr[57815]= -30595422;
assign addr[57816]= 274614114;
assign addr[57817]= 574258580;
assign addr[57818]= 862265664;
assign addr[57819]= 1132798888;
assign addr[57820]= 1380375881;
assign addr[57821]= 1599979481;
assign addr[57822]= 1787159411;
assign addr[57823]= 1938122457;
assign addr[57824]= 2049809346;
assign addr[57825]= 2119956737;
assign addr[57826]= 2147143090;
assign addr[57827]= 2130817471;
assign addr[57828]= 2071310720;
assign addr[57829]= 1969828744;
assign addr[57830]= 1828428082;
assign addr[57831]= 1649974225;
assign addr[57832]= 1438083551;
assign addr[57833]= 1197050035;
assign addr[57834]= 931758235;
assign addr[57835]= 647584304;
assign addr[57836]= 350287041;
assign addr[57837]= 45891193;
assign addr[57838]= -259434643;
assign addr[57839]= -559503022;
assign addr[57840]= -848233042;
assign addr[57841]= -1119773573;
assign addr[57842]= -1368621831;
assign addr[57843]= -1589734894;
assign addr[57844]= -1778631892;
assign addr[57845]= -1931484818;
assign addr[57846]= -2045196100;
assign addr[57847]= -2117461370;
assign addr[57848]= -2146816171;
assign addr[57849]= -2132665626;
assign addr[57850]= -2075296495;
assign addr[57851]= -1975871368;
assign addr[57852]= -1836405100;
assign addr[57853]= -1659723983;
assign addr[57854]= -1449408469;
assign addr[57855]= -1209720613;
assign addr[57856]= -945517704;
assign addr[57857]= -662153826;
assign addr[57858]= -365371365;
assign addr[57859]= -61184634;
assign addr[57860]= 244242007;
assign addr[57861]= 544719071;
assign addr[57862]= 834157373;
assign addr[57863]= 1106691431;
assign addr[57864]= 1356798326;
assign addr[57865]= 1579409630;
assign addr[57866]= 1770014111;
assign addr[57867]= 1924749160;
assign addr[57868]= 2040479063;
assign addr[57869]= 2114858546;
assign addr[57870]= 2146380306;
assign addr[57871]= 2134405552;
assign addr[57872]= 2079176953;
assign addr[57873]= 1981813720;
assign addr[57874]= 1844288924;
assign addr[57875]= 1669389513;
assign addr[57876]= 1460659832;
assign addr[57877]= 1222329801;
assign addr[57878]= 959229189;
assign addr[57879]= 676689746;
assign addr[57880]= 380437148;
assign addr[57881]= 76474970;
assign addr[57882]= -229036977;
assign addr[57883]= -529907477;
assign addr[57884]= -820039373;
assign addr[57885]= -1093553126;
assign addr[57886]= -1344905966;
assign addr[57887]= -1569004214;
assign addr[57888]= -1761306505;
assign addr[57889]= -1917915825;
assign addr[57890]= -2035658475;
assign addr[57891]= -2112148396;
assign addr[57892]= -2145835515;
assign addr[57893]= -2136037160;
assign addr[57894]= -2082951896;
assign addr[57895]= -1987655498;
assign addr[57896]= -1852079154;
assign addr[57897]= -1678970324;
assign addr[57898]= -1471837070;
assign addr[57899]= -1234876957;
assign addr[57900]= -972891995;
assign addr[57901]= -691191324;
assign addr[57902]= -395483624;
assign addr[57903]= -91761426;
assign addr[57904]= 213820322;
assign addr[57905]= 515068990;
assign addr[57906]= 805879757;
assign addr[57907]= 1080359326;
assign addr[57908]= 1332945355;
assign addr[57909]= 1558519173;
assign addr[57910]= 1752509516;
assign addr[57911]= 1910985158;
assign addr[57912]= 2030734582;
assign addr[57913]= 2109331059;
assign addr[57914]= 2145181827;
assign addr[57915]= 2137560369;
assign addr[57916]= 2086621133;
assign addr[57917]= 1993396407;
assign addr[57918]= 1859775393;
assign addr[57919]= 1688465931;
assign addr[57920]= 1482939614;
assign addr[57921]= 1247361445;
assign addr[57922]= 986505429;
assign addr[57923]= 705657826;
assign addr[57924]= 410510029;
assign addr[57925]= 107043224;
assign addr[57926]= -198592817;
assign addr[57927]= -500204365;
assign addr[57928]= -791679244;
assign addr[57929]= -1067110699;
assign addr[57930]= -1320917099;
assign addr[57931]= -1547955041;
assign addr[57932]= -1743623590;
assign addr[57933]= -1903957513;
assign addr[57934]= -2025707632;
assign addr[57935]= -2106406677;
assign addr[57936]= -2144419275;
assign addr[57937]= -2138975100;
assign addr[57938]= -2090184478;
assign addr[57939]= -1999036154;
assign addr[57940]= -1867377253;
assign addr[57941]= -1697875851;
assign addr[57942]= -1493966902;
assign addr[57943]= -1259782632;
assign addr[57944]= -1000068799;
assign addr[57945]= -720088517;
assign addr[57946]= -425515602;
assign addr[57947]= -122319591;
assign addr[57948]= 183355234;
assign addr[57949]= 485314355;
assign addr[57950]= 777438554;
assign addr[57951]= 1053807919;
assign addr[57952]= 1308821808;
assign addr[57953]= 1537312353;
assign addr[57954]= 1734649179;
assign addr[57955]= 1896833245;
assign addr[57956]= 2020577882;
assign addr[57957]= 2103375398;
assign addr[57958]= 2143547897;
assign addr[57959]= 2140281282;
assign addr[57960]= 2093641749;
assign addr[57961]= 2004574453;
assign addr[57962]= 1874884346;
assign addr[57963]= 1707199606;
assign addr[57964]= 1504918373;
assign addr[57965]= 1272139887;
assign addr[57966]= 1013581418;
assign addr[57967]= 734482665;
assign addr[57968]= 440499581;
assign addr[57969]= 137589750;
assign addr[57970]= -168108346;
assign addr[57971]= -470399716;
assign addr[57972]= -763158411;
assign addr[57973]= -1040451659;
assign addr[57974]= -1296660098;
assign addr[57975]= -1526591649;
assign addr[57976]= -1725586737;
assign addr[57977]= -1889612716;
assign addr[57978]= -2015345591;
assign addr[57979]= -2100237377;
assign addr[57980]= -2142567738;
assign addr[57981]= -2141478848;
assign addr[57982]= -2096992772;
assign addr[57983]= -2010011024;
assign addr[57984]= -1882296293;
assign addr[57985]= -1716436725;
assign addr[57986]= -1515793473;
assign addr[57987]= -1284432584;
assign addr[57988]= -1027042599;
assign addr[57989]= -748839539;
assign addr[57990]= -455461206;
assign addr[57991]= -152852926;
assign addr[57992]= 152852926;
assign addr[57993]= 455461206;
assign addr[57994]= 748839539;
assign addr[57995]= 1027042599;
assign addr[57996]= 1284432584;
assign addr[57997]= 1515793473;
assign addr[57998]= 1716436725;
assign addr[57999]= 1882296293;
assign addr[58000]= 2010011024;
assign addr[58001]= 2096992772;
assign addr[58002]= 2141478848;
assign addr[58003]= 2142567738;
assign addr[58004]= 2100237377;
assign addr[58005]= 2015345591;
assign addr[58006]= 1889612716;
assign addr[58007]= 1725586737;
assign addr[58008]= 1526591649;
assign addr[58009]= 1296660098;
assign addr[58010]= 1040451659;
assign addr[58011]= 763158411;
assign addr[58012]= 470399716;
assign addr[58013]= 168108346;
assign addr[58014]= -137589750;
assign addr[58015]= -440499581;
assign addr[58016]= -734482665;
assign addr[58017]= -1013581418;
assign addr[58018]= -1272139887;
assign addr[58019]= -1504918373;
assign addr[58020]= -1707199606;
assign addr[58021]= -1874884346;
assign addr[58022]= -2004574453;
assign addr[58023]= -2093641749;
assign addr[58024]= -2140281282;
assign addr[58025]= -2143547897;
assign addr[58026]= -2103375398;
assign addr[58027]= -2020577882;
assign addr[58028]= -1896833245;
assign addr[58029]= -1734649179;
assign addr[58030]= -1537312353;
assign addr[58031]= -1308821808;
assign addr[58032]= -1053807919;
assign addr[58033]= -777438554;
assign addr[58034]= -485314355;
assign addr[58035]= -183355234;
assign addr[58036]= 122319591;
assign addr[58037]= 425515602;
assign addr[58038]= 720088517;
assign addr[58039]= 1000068799;
assign addr[58040]= 1259782632;
assign addr[58041]= 1493966902;
assign addr[58042]= 1697875851;
assign addr[58043]= 1867377253;
assign addr[58044]= 1999036154;
assign addr[58045]= 2090184478;
assign addr[58046]= 2138975100;
assign addr[58047]= 2144419275;
assign addr[58048]= 2106406677;
assign addr[58049]= 2025707632;
assign addr[58050]= 1903957513;
assign addr[58051]= 1743623590;
assign addr[58052]= 1547955041;
assign addr[58053]= 1320917099;
assign addr[58054]= 1067110699;
assign addr[58055]= 791679244;
assign addr[58056]= 500204365;
assign addr[58057]= 198592817;
assign addr[58058]= -107043224;
assign addr[58059]= -410510029;
assign addr[58060]= -705657826;
assign addr[58061]= -986505429;
assign addr[58062]= -1247361445;
assign addr[58063]= -1482939614;
assign addr[58064]= -1688465931;
assign addr[58065]= -1859775393;
assign addr[58066]= -1993396407;
assign addr[58067]= -2086621133;
assign addr[58068]= -2137560369;
assign addr[58069]= -2145181827;
assign addr[58070]= -2109331059;
assign addr[58071]= -2030734582;
assign addr[58072]= -1910985158;
assign addr[58073]= -1752509516;
assign addr[58074]= -1558519173;
assign addr[58075]= -1332945355;
assign addr[58076]= -1080359326;
assign addr[58077]= -805879757;
assign addr[58078]= -515068990;
assign addr[58079]= -213820322;
assign addr[58080]= 91761426;
assign addr[58081]= 395483624;
assign addr[58082]= 691191324;
assign addr[58083]= 972891995;
assign addr[58084]= 1234876957;
assign addr[58085]= 1471837070;
assign addr[58086]= 1678970324;
assign addr[58087]= 1852079154;
assign addr[58088]= 1987655498;
assign addr[58089]= 2082951896;
assign addr[58090]= 2136037160;
assign addr[58091]= 2145835515;
assign addr[58092]= 2112148396;
assign addr[58093]= 2035658475;
assign addr[58094]= 1917915825;
assign addr[58095]= 1761306505;
assign addr[58096]= 1569004214;
assign addr[58097]= 1344905966;
assign addr[58098]= 1093553126;
assign addr[58099]= 820039373;
assign addr[58100]= 529907477;
assign addr[58101]= 229036977;
assign addr[58102]= -76474970;
assign addr[58103]= -380437148;
assign addr[58104]= -676689746;
assign addr[58105]= -959229189;
assign addr[58106]= -1222329801;
assign addr[58107]= -1460659832;
assign addr[58108]= -1669389513;
assign addr[58109]= -1844288924;
assign addr[58110]= -1981813720;
assign addr[58111]= -2079176953;
assign addr[58112]= -2134405552;
assign addr[58113]= -2146380306;
assign addr[58114]= -2114858546;
assign addr[58115]= -2040479063;
assign addr[58116]= -1924749160;
assign addr[58117]= -1770014111;
assign addr[58118]= -1579409630;
assign addr[58119]= -1356798326;
assign addr[58120]= -1106691431;
assign addr[58121]= -834157373;
assign addr[58122]= -544719071;
assign addr[58123]= -244242007;
assign addr[58124]= 61184634;
assign addr[58125]= 365371365;
assign addr[58126]= 662153826;
assign addr[58127]= 945517704;
assign addr[58128]= 1209720613;
assign addr[58129]= 1449408469;
assign addr[58130]= 1659723983;
assign addr[58131]= 1836405100;
assign addr[58132]= 1975871368;
assign addr[58133]= 2075296495;
assign addr[58134]= 2132665626;
assign addr[58135]= 2146816171;
assign addr[58136]= 2117461370;
assign addr[58137]= 2045196100;
assign addr[58138]= 1931484818;
assign addr[58139]= 1778631892;
assign addr[58140]= 1589734894;
assign addr[58141]= 1368621831;
assign addr[58142]= 1119773573;
assign addr[58143]= 848233042;
assign addr[58144]= 559503022;
assign addr[58145]= 259434643;
assign addr[58146]= -45891193;
assign addr[58147]= -350287041;
assign addr[58148]= -647584304;
assign addr[58149]= -931758235;
assign addr[58150]= -1197050035;
assign addr[58151]= -1438083551;
assign addr[58152]= -1649974225;
assign addr[58153]= -1828428082;
assign addr[58154]= -1969828744;
assign addr[58155]= -2071310720;
assign addr[58156]= -2130817471;
assign addr[58157]= -2147143090;
assign addr[58158]= -2119956737;
assign addr[58159]= -2049809346;
assign addr[58160]= -1938122457;
assign addr[58161]= -1787159411;
assign addr[58162]= -1599979481;
assign addr[58163]= -1380375881;
assign addr[58164]= -1132798888;
assign addr[58165]= -862265664;
assign addr[58166]= -574258580;
assign addr[58167]= -274614114;
assign addr[58168]= 30595422;
assign addr[58169]= 335184940;
assign addr[58170]= 632981917;
assign addr[58171]= 917951481;
assign addr[58172]= 1184318708;
assign addr[58173]= 1426685652;
assign addr[58174]= 1640140734;
assign addr[58175]= 1820358275;
assign addr[58176]= 1963686155;
assign addr[58177]= 2067219829;
assign addr[58178]= 2128861181;
assign addr[58179]= 2147361045;
assign addr[58180]= 2122344521;
assign addr[58181]= 2054318569;
assign addr[58182]= 1944661739;
assign addr[58183]= 1795596234;
assign addr[58184]= 1610142873;
assign addr[58185]= 1392059879;
assign addr[58186]= 1145766716;
assign addr[58187]= 876254528;
assign addr[58188]= 588984994;
assign addr[58189]= 289779648;
assign addr[58190]= -15298099;
assign addr[58191]= -320065829;
assign addr[58192]= -618347408;
assign addr[58193]= -904098143;
assign addr[58194]= -1171527280;
assign addr[58195]= -1415215352;
assign addr[58196]= -1630224009;
assign addr[58197]= -1812196087;
assign addr[58198]= -1957443913;
assign addr[58199]= -2063024031;
assign addr[58200]= -2126796855;
assign addr[58201]= -2147470025;
assign addr[58202]= -2124624598;
assign addr[58203]= -2058723538;
assign addr[58204]= -1951102334;
assign addr[58205]= -1803941934;
assign addr[58206]= -1620224553;
assign addr[58207]= -1403673233;
assign addr[58208]= -1158676398;
assign addr[58209]= -890198924;
assign addr[58210]= -603681519;
assign addr[58211]= -304930476;
assign addr[58212]= 0;
assign addr[58213]= 304930476;
assign addr[58214]= 603681519;
assign addr[58215]= 890198924;
assign addr[58216]= 1158676398;
assign addr[58217]= 1403673233;
assign addr[58218]= 1620224553;
assign addr[58219]= 1803941934;
assign addr[58220]= 1951102334;
assign addr[58221]= 2058723538;
assign addr[58222]= 2124624598;
assign addr[58223]= 2147470025;
assign addr[58224]= 2126796855;
assign addr[58225]= 2063024031;
assign addr[58226]= 1957443913;
assign addr[58227]= 1812196087;
assign addr[58228]= 1630224009;
assign addr[58229]= 1415215352;
assign addr[58230]= 1171527280;
assign addr[58231]= 904098143;
assign addr[58232]= 618347408;
assign addr[58233]= 320065829;
assign addr[58234]= 15298099;
assign addr[58235]= -289779648;
assign addr[58236]= -588984994;
assign addr[58237]= -876254528;
assign addr[58238]= -1145766716;
assign addr[58239]= -1392059879;
assign addr[58240]= -1610142873;
assign addr[58241]= -1795596234;
assign addr[58242]= -1944661739;
assign addr[58243]= -2054318569;
assign addr[58244]= -2122344521;
assign addr[58245]= -2147361045;
assign addr[58246]= -2128861181;
assign addr[58247]= -2067219829;
assign addr[58248]= -1963686155;
assign addr[58249]= -1820358275;
assign addr[58250]= -1640140734;
assign addr[58251]= -1426685652;
assign addr[58252]= -1184318708;
assign addr[58253]= -917951481;
assign addr[58254]= -632981917;
assign addr[58255]= -335184940;
assign addr[58256]= -30595422;
assign addr[58257]= 274614114;
assign addr[58258]= 574258580;
assign addr[58259]= 862265664;
assign addr[58260]= 1132798888;
assign addr[58261]= 1380375881;
assign addr[58262]= 1599979481;
assign addr[58263]= 1787159411;
assign addr[58264]= 1938122457;
assign addr[58265]= 2049809346;
assign addr[58266]= 2119956737;
assign addr[58267]= 2147143090;
assign addr[58268]= 2130817471;
assign addr[58269]= 2071310720;
assign addr[58270]= 1969828744;
assign addr[58271]= 1828428082;
assign addr[58272]= 1649974225;
assign addr[58273]= 1438083551;
assign addr[58274]= 1197050035;
assign addr[58275]= 931758235;
assign addr[58276]= 647584304;
assign addr[58277]= 350287041;
assign addr[58278]= 45891193;
assign addr[58279]= -259434643;
assign addr[58280]= -559503022;
assign addr[58281]= -848233042;
assign addr[58282]= -1119773573;
assign addr[58283]= -1368621831;
assign addr[58284]= -1589734894;
assign addr[58285]= -1778631892;
assign addr[58286]= -1931484818;
assign addr[58287]= -2045196100;
assign addr[58288]= -2117461370;
assign addr[58289]= -2146816171;
assign addr[58290]= -2132665626;
assign addr[58291]= -2075296495;
assign addr[58292]= -1975871368;
assign addr[58293]= -1836405100;
assign addr[58294]= -1659723983;
assign addr[58295]= -1449408469;
assign addr[58296]= -1209720613;
assign addr[58297]= -945517704;
assign addr[58298]= -662153826;
assign addr[58299]= -365371365;
assign addr[58300]= -61184634;
assign addr[58301]= 244242007;
assign addr[58302]= 544719071;
assign addr[58303]= 834157373;
assign addr[58304]= 1106691431;
assign addr[58305]= 1356798326;
assign addr[58306]= 1579409630;
assign addr[58307]= 1770014111;
assign addr[58308]= 1924749160;
assign addr[58309]= 2040479063;
assign addr[58310]= 2114858546;
assign addr[58311]= 2146380306;
assign addr[58312]= 2134405552;
assign addr[58313]= 2079176953;
assign addr[58314]= 1981813720;
assign addr[58315]= 1844288924;
assign addr[58316]= 1669389513;
assign addr[58317]= 1460659832;
assign addr[58318]= 1222329801;
assign addr[58319]= 959229189;
assign addr[58320]= 676689746;
assign addr[58321]= 380437148;
assign addr[58322]= 76474970;
assign addr[58323]= -229036977;
assign addr[58324]= -529907477;
assign addr[58325]= -820039373;
assign addr[58326]= -1093553126;
assign addr[58327]= -1344905966;
assign addr[58328]= -1569004214;
assign addr[58329]= -1761306505;
assign addr[58330]= -1917915825;
assign addr[58331]= -2035658475;
assign addr[58332]= -2112148396;
assign addr[58333]= -2145835515;
assign addr[58334]= -2136037160;
assign addr[58335]= -2082951896;
assign addr[58336]= -1987655498;
assign addr[58337]= -1852079154;
assign addr[58338]= -1678970324;
assign addr[58339]= -1471837070;
assign addr[58340]= -1234876957;
assign addr[58341]= -972891995;
assign addr[58342]= -691191324;
assign addr[58343]= -395483624;
assign addr[58344]= -91761426;
assign addr[58345]= 213820322;
assign addr[58346]= 515068990;
assign addr[58347]= 805879757;
assign addr[58348]= 1080359326;
assign addr[58349]= 1332945355;
assign addr[58350]= 1558519173;
assign addr[58351]= 1752509516;
assign addr[58352]= 1910985158;
assign addr[58353]= 2030734582;
assign addr[58354]= 2109331059;
assign addr[58355]= 2145181827;
assign addr[58356]= 2137560369;
assign addr[58357]= 2086621133;
assign addr[58358]= 1993396407;
assign addr[58359]= 1859775393;
assign addr[58360]= 1688465931;
assign addr[58361]= 1482939614;
assign addr[58362]= 1247361445;
assign addr[58363]= 986505429;
assign addr[58364]= 705657826;
assign addr[58365]= 410510029;
assign addr[58366]= 107043224;
assign addr[58367]= -198592817;
assign addr[58368]= -500204365;
assign addr[58369]= -791679244;
assign addr[58370]= -1067110699;
assign addr[58371]= -1320917099;
assign addr[58372]= -1547955041;
assign addr[58373]= -1743623590;
assign addr[58374]= -1903957513;
assign addr[58375]= -2025707632;
assign addr[58376]= -2106406677;
assign addr[58377]= -2144419275;
assign addr[58378]= -2138975100;
assign addr[58379]= -2090184478;
assign addr[58380]= -1999036154;
assign addr[58381]= -1867377253;
assign addr[58382]= -1697875851;
assign addr[58383]= -1493966902;
assign addr[58384]= -1259782632;
assign addr[58385]= -1000068799;
assign addr[58386]= -720088517;
assign addr[58387]= -425515602;
assign addr[58388]= -122319591;
assign addr[58389]= 183355234;
assign addr[58390]= 485314355;
assign addr[58391]= 777438554;
assign addr[58392]= 1053807919;
assign addr[58393]= 1308821808;
assign addr[58394]= 1537312353;
assign addr[58395]= 1734649179;
assign addr[58396]= 1896833245;
assign addr[58397]= 2020577882;
assign addr[58398]= 2103375398;
assign addr[58399]= 2143547897;
assign addr[58400]= 2140281282;
assign addr[58401]= 2093641749;
assign addr[58402]= 2004574453;
assign addr[58403]= 1874884346;
assign addr[58404]= 1707199606;
assign addr[58405]= 1504918373;
assign addr[58406]= 1272139887;
assign addr[58407]= 1013581418;
assign addr[58408]= 734482665;
assign addr[58409]= 440499581;
assign addr[58410]= 137589750;
assign addr[58411]= -168108346;
assign addr[58412]= -470399716;
assign addr[58413]= -763158411;
assign addr[58414]= -1040451659;
assign addr[58415]= -1296660098;
assign addr[58416]= -1526591649;
assign addr[58417]= -1725586737;
assign addr[58418]= -1889612716;
assign addr[58419]= -2015345591;
assign addr[58420]= -2100237377;
assign addr[58421]= -2142567738;
assign addr[58422]= -2141478848;
assign addr[58423]= -2096992772;
assign addr[58424]= -2010011024;
assign addr[58425]= -1882296293;
assign addr[58426]= -1716436725;
assign addr[58427]= -1515793473;
assign addr[58428]= -1284432584;
assign addr[58429]= -1027042599;
assign addr[58430]= -748839539;
assign addr[58431]= -455461206;
assign addr[58432]= -152852926;
assign addr[58433]= 152852926;
assign addr[58434]= 455461206;
assign addr[58435]= 748839539;
assign addr[58436]= 1027042599;
assign addr[58437]= 1284432584;
assign addr[58438]= 1515793473;
assign addr[58439]= 1716436725;
assign addr[58440]= 1882296293;
assign addr[58441]= 2010011024;
assign addr[58442]= 2096992772;
assign addr[58443]= 2141478848;
assign addr[58444]= 2142567738;
assign addr[58445]= 2100237377;
assign addr[58446]= 2015345591;
assign addr[58447]= 1889612716;
assign addr[58448]= 1725586737;
assign addr[58449]= 1526591649;
assign addr[58450]= 1296660098;
assign addr[58451]= 1040451659;
assign addr[58452]= 763158411;
assign addr[58453]= 470399716;
assign addr[58454]= 168108346;
assign addr[58455]= -137589750;
assign addr[58456]= -440499581;
assign addr[58457]= -734482665;
assign addr[58458]= -1013581418;
assign addr[58459]= -1272139887;
assign addr[58460]= -1504918373;
assign addr[58461]= -1707199606;
assign addr[58462]= -1874884346;
assign addr[58463]= -2004574453;
assign addr[58464]= -2093641749;
assign addr[58465]= -2140281282;
assign addr[58466]= -2143547897;
assign addr[58467]= -2103375398;
assign addr[58468]= -2020577882;
assign addr[58469]= -1896833245;
assign addr[58470]= -1734649179;
assign addr[58471]= -1537312353;
assign addr[58472]= -1308821808;
assign addr[58473]= -1053807919;
assign addr[58474]= -777438554;
assign addr[58475]= -485314355;
assign addr[58476]= -183355234;
assign addr[58477]= 122319591;
assign addr[58478]= 425515602;
assign addr[58479]= 720088517;
assign addr[58480]= 1000068799;
assign addr[58481]= 1259782632;
assign addr[58482]= 1493966902;
assign addr[58483]= 1697875851;
assign addr[58484]= 1867377253;
assign addr[58485]= 1999036154;
assign addr[58486]= 2090184478;
assign addr[58487]= 2138975100;
assign addr[58488]= 2144419275;
assign addr[58489]= 2106406677;
assign addr[58490]= 2025707632;
assign addr[58491]= 1903957513;
assign addr[58492]= 1743623590;
assign addr[58493]= 1547955041;
assign addr[58494]= 1320917099;
assign addr[58495]= 1067110699;
assign addr[58496]= 791679244;
assign addr[58497]= 500204365;
assign addr[58498]= 198592817;
assign addr[58499]= -107043224;
assign addr[58500]= -410510029;
assign addr[58501]= -705657826;
assign addr[58502]= -986505429;
assign addr[58503]= -1247361445;
assign addr[58504]= -1482939614;
assign addr[58505]= -1688465931;
assign addr[58506]= -1859775393;
assign addr[58507]= -1993396407;
assign addr[58508]= -2086621133;
assign addr[58509]= -2137560369;
assign addr[58510]= -2145181827;
assign addr[58511]= -2109331059;
assign addr[58512]= -2030734582;
assign addr[58513]= -1910985158;
assign addr[58514]= -1752509516;
assign addr[58515]= -1558519173;
assign addr[58516]= -1332945355;
assign addr[58517]= -1080359326;
assign addr[58518]= -805879757;
assign addr[58519]= -515068990;
assign addr[58520]= -213820322;
assign addr[58521]= 91761426;
assign addr[58522]= 395483624;
assign addr[58523]= 691191324;
assign addr[58524]= 972891995;
assign addr[58525]= 1234876957;
assign addr[58526]= 1471837070;
assign addr[58527]= 1678970324;
assign addr[58528]= 1852079154;
assign addr[58529]= 1987655498;
assign addr[58530]= 2082951896;
assign addr[58531]= 2136037160;
assign addr[58532]= 2145835515;
assign addr[58533]= 2112148396;
assign addr[58534]= 2035658475;
assign addr[58535]= 1917915825;
assign addr[58536]= 1761306505;
assign addr[58537]= 1569004214;
assign addr[58538]= 1344905966;
assign addr[58539]= 1093553126;
assign addr[58540]= 820039373;
assign addr[58541]= 529907477;
assign addr[58542]= 229036977;
assign addr[58543]= -76474970;
assign addr[58544]= -380437148;
assign addr[58545]= -676689746;
assign addr[58546]= -959229189;
assign addr[58547]= -1222329801;
assign addr[58548]= -1460659832;
assign addr[58549]= -1669389513;
assign addr[58550]= -1844288924;
assign addr[58551]= -1981813720;
assign addr[58552]= -2079176953;
assign addr[58553]= -2134405552;
assign addr[58554]= -2146380306;
assign addr[58555]= -2114858546;
assign addr[58556]= -2040479063;
assign addr[58557]= -1924749160;
assign addr[58558]= -1770014111;
assign addr[58559]= -1579409630;
assign addr[58560]= -1356798326;
assign addr[58561]= -1106691431;
assign addr[58562]= -834157373;
assign addr[58563]= -544719071;
assign addr[58564]= -244242007;
assign addr[58565]= 61184634;
assign addr[58566]= 365371365;
assign addr[58567]= 662153826;
assign addr[58568]= 945517704;
assign addr[58569]= 1209720613;
assign addr[58570]= 1449408469;
assign addr[58571]= 1659723983;
assign addr[58572]= 1836405100;
assign addr[58573]= 1975871368;
assign addr[58574]= 2075296495;
assign addr[58575]= 2132665626;
assign addr[58576]= 2146816171;
assign addr[58577]= 2117461370;
assign addr[58578]= 2045196100;
assign addr[58579]= 1931484818;
assign addr[58580]= 1778631892;
assign addr[58581]= 1589734894;
assign addr[58582]= 1368621831;
assign addr[58583]= 1119773573;
assign addr[58584]= 848233042;
assign addr[58585]= 559503022;
assign addr[58586]= 259434643;
assign addr[58587]= -45891193;
assign addr[58588]= -350287041;
assign addr[58589]= -647584304;
assign addr[58590]= -931758235;
assign addr[58591]= -1197050035;
assign addr[58592]= -1438083551;
assign addr[58593]= -1649974225;
assign addr[58594]= -1828428082;
assign addr[58595]= -1969828744;
assign addr[58596]= -2071310720;
assign addr[58597]= -2130817471;
assign addr[58598]= -2147143090;
assign addr[58599]= -2119956737;
assign addr[58600]= -2049809346;
assign addr[58601]= -1938122457;
assign addr[58602]= -1787159411;
assign addr[58603]= -1599979481;
assign addr[58604]= -1380375881;
assign addr[58605]= -1132798888;
assign addr[58606]= -862265664;
assign addr[58607]= -574258580;
assign addr[58608]= -274614114;
assign addr[58609]= 30595422;
assign addr[58610]= 335184940;
assign addr[58611]= 632981917;
assign addr[58612]= 917951481;
assign addr[58613]= 1184318708;
assign addr[58614]= 1426685652;
assign addr[58615]= 1640140734;
assign addr[58616]= 1820358275;
assign addr[58617]= 1963686155;
assign addr[58618]= 2067219829;
assign addr[58619]= 2128861181;
assign addr[58620]= 2147361045;
assign addr[58621]= 2122344521;
assign addr[58622]= 2054318569;
assign addr[58623]= 1944661739;
assign addr[58624]= 1795596234;
assign addr[58625]= 1610142873;
assign addr[58626]= 1392059879;
assign addr[58627]= 1145766716;
assign addr[58628]= 876254528;
assign addr[58629]= 588984994;
assign addr[58630]= 289779648;
assign addr[58631]= -15298099;
assign addr[58632]= -320065829;
assign addr[58633]= -618347408;
assign addr[58634]= -904098143;
assign addr[58635]= -1171527280;
assign addr[58636]= -1415215352;
assign addr[58637]= -1630224009;
assign addr[58638]= -1812196087;
assign addr[58639]= -1957443913;
assign addr[58640]= -2063024031;
assign addr[58641]= -2126796855;
assign addr[58642]= -2147470025;
assign addr[58643]= -2124624598;
assign addr[58644]= -2058723538;
assign addr[58645]= -1951102334;
assign addr[58646]= -1803941934;
assign addr[58647]= -1620224553;
assign addr[58648]= -1403673233;
assign addr[58649]= -1158676398;
assign addr[58650]= -890198924;
assign addr[58651]= -603681519;
assign addr[58652]= -304930476;
assign addr[58653]= 0;
assign addr[58654]= 304930476;
assign addr[58655]= 603681519;
assign addr[58656]= 890198924;
assign addr[58657]= 1158676398;
assign addr[58658]= 1403673233;
assign addr[58659]= 1620224553;
assign addr[58660]= 1803941934;
assign addr[58661]= 1951102334;
assign addr[58662]= 2058723538;
assign addr[58663]= 2124624598;
assign addr[58664]= 2147470025;
assign addr[58665]= 2126796855;
assign addr[58666]= 2063024031;
assign addr[58667]= 1957443913;
assign addr[58668]= 1812196087;
assign addr[58669]= 1630224009;
assign addr[58670]= 1415215352;
assign addr[58671]= 1171527280;
assign addr[58672]= 904098143;
assign addr[58673]= 618347408;
assign addr[58674]= 320065829;
assign addr[58675]= 15298099;
assign addr[58676]= -289779648;
assign addr[58677]= -588984994;
assign addr[58678]= -876254528;
assign addr[58679]= -1145766716;
assign addr[58680]= -1392059879;
assign addr[58681]= -1610142873;
assign addr[58682]= -1795596234;
assign addr[58683]= -1944661739;
assign addr[58684]= -2054318569;
assign addr[58685]= -2122344521;
assign addr[58686]= -2147361045;
assign addr[58687]= -2128861181;
assign addr[58688]= -2067219829;
assign addr[58689]= -1963686155;
assign addr[58690]= -1820358275;
assign addr[58691]= -1640140734;
assign addr[58692]= -1426685652;
assign addr[58693]= -1184318708;
assign addr[58694]= -917951481;
assign addr[58695]= -632981917;
assign addr[58696]= -335184940;
assign addr[58697]= -30595422;
assign addr[58698]= 274614114;
assign addr[58699]= 574258580;
assign addr[58700]= 862265664;
assign addr[58701]= 1132798888;
assign addr[58702]= 1380375881;
assign addr[58703]= 1599979481;
assign addr[58704]= 1787159411;
assign addr[58705]= 1938122457;
assign addr[58706]= 2049809346;
assign addr[58707]= 2119956737;
assign addr[58708]= 2147143090;
assign addr[58709]= 2130817471;
assign addr[58710]= 2071310720;
assign addr[58711]= 1969828744;
assign addr[58712]= 1828428082;
assign addr[58713]= 1649974225;
assign addr[58714]= 1438083551;
assign addr[58715]= 1197050035;
assign addr[58716]= 931758235;
assign addr[58717]= 647584304;
assign addr[58718]= 350287041;
assign addr[58719]= 45891193;
assign addr[58720]= -259434643;
assign addr[58721]= -559503022;
assign addr[58722]= -848233042;
assign addr[58723]= -1119773573;
assign addr[58724]= -1368621831;
assign addr[58725]= -1589734894;
assign addr[58726]= -1778631892;
assign addr[58727]= -1931484818;
assign addr[58728]= -2045196100;
assign addr[58729]= -2117461370;
assign addr[58730]= -2146816171;
assign addr[58731]= -2132665626;
assign addr[58732]= -2075296495;
assign addr[58733]= -1975871368;
assign addr[58734]= -1836405100;
assign addr[58735]= -1659723983;
assign addr[58736]= -1449408469;
assign addr[58737]= -1209720613;
assign addr[58738]= -945517704;
assign addr[58739]= -662153826;
assign addr[58740]= -365371365;
assign addr[58741]= -61184634;
assign addr[58742]= 244242007;
assign addr[58743]= 544719071;
assign addr[58744]= 834157373;
assign addr[58745]= 1106691431;
assign addr[58746]= 1356798326;
assign addr[58747]= 1579409630;
assign addr[58748]= 1770014111;
assign addr[58749]= 1924749160;
assign addr[58750]= 2040479063;
assign addr[58751]= 2114858546;
assign addr[58752]= 2146380306;
assign addr[58753]= 2134405552;
assign addr[58754]= 2079176953;
assign addr[58755]= 1981813720;
assign addr[58756]= 1844288924;
assign addr[58757]= 1669389513;
assign addr[58758]= 1460659832;
assign addr[58759]= 1222329801;
assign addr[58760]= 959229189;
assign addr[58761]= 676689746;
assign addr[58762]= 380437148;
assign addr[58763]= 76474970;
assign addr[58764]= -229036977;
assign addr[58765]= -529907477;
assign addr[58766]= -820039373;
assign addr[58767]= -1093553126;
assign addr[58768]= -1344905966;
assign addr[58769]= -1569004214;
assign addr[58770]= -1761306505;
assign addr[58771]= -1917915825;
assign addr[58772]= -2035658475;
assign addr[58773]= -2112148396;
assign addr[58774]= -2145835515;
assign addr[58775]= -2136037160;
assign addr[58776]= -2082951896;
assign addr[58777]= -1987655498;
assign addr[58778]= -1852079154;
assign addr[58779]= -1678970324;
assign addr[58780]= -1471837070;
assign addr[58781]= -1234876957;
assign addr[58782]= -972891995;
assign addr[58783]= -691191324;
assign addr[58784]= -395483624;
assign addr[58785]= -91761426;
assign addr[58786]= 213820322;
assign addr[58787]= 515068990;
assign addr[58788]= 805879757;
assign addr[58789]= 1080359326;
assign addr[58790]= 1332945355;
assign addr[58791]= 1558519173;
assign addr[58792]= 1752509516;
assign addr[58793]= 1910985158;
assign addr[58794]= 2030734582;
assign addr[58795]= 2109331059;
assign addr[58796]= 2145181827;
assign addr[58797]= 2137560369;
assign addr[58798]= 2086621133;
assign addr[58799]= 1993396407;
assign addr[58800]= 1859775393;
assign addr[58801]= 1688465931;
assign addr[58802]= 1482939614;
assign addr[58803]= 1247361445;
assign addr[58804]= 986505429;
assign addr[58805]= 705657826;
assign addr[58806]= 410510029;
assign addr[58807]= 107043224;
assign addr[58808]= -198592817;
assign addr[58809]= -500204365;
assign addr[58810]= -791679244;
assign addr[58811]= -1067110699;
assign addr[58812]= -1320917099;
assign addr[58813]= -1547955041;
assign addr[58814]= -1743623590;
assign addr[58815]= -1903957513;
assign addr[58816]= -2025707632;
assign addr[58817]= -2106406677;
assign addr[58818]= -2144419275;
assign addr[58819]= -2138975100;
assign addr[58820]= -2090184478;
assign addr[58821]= -1999036154;
assign addr[58822]= -1867377253;
assign addr[58823]= -1697875851;
assign addr[58824]= -1493966902;
assign addr[58825]= -1259782632;
assign addr[58826]= -1000068799;
assign addr[58827]= -720088517;
assign addr[58828]= -425515602;
assign addr[58829]= -122319591;
assign addr[58830]= 183355234;
assign addr[58831]= 485314355;
assign addr[58832]= 777438554;
assign addr[58833]= 1053807919;
assign addr[58834]= 1308821808;
assign addr[58835]= 1537312353;
assign addr[58836]= 1734649179;
assign addr[58837]= 1896833245;
assign addr[58838]= 2020577882;
assign addr[58839]= 2103375398;
assign addr[58840]= 2143547897;
assign addr[58841]= 2140281282;
assign addr[58842]= 2093641749;
assign addr[58843]= 2004574453;
assign addr[58844]= 1874884346;
assign addr[58845]= 1707199606;
assign addr[58846]= 1504918373;
assign addr[58847]= 1272139887;
assign addr[58848]= 1013581418;
assign addr[58849]= 734482665;
assign addr[58850]= 440499581;
assign addr[58851]= 137589750;
assign addr[58852]= -168108346;
assign addr[58853]= -470399716;
assign addr[58854]= -763158411;
assign addr[58855]= -1040451659;
assign addr[58856]= -1296660098;
assign addr[58857]= -1526591649;
assign addr[58858]= -1725586737;
assign addr[58859]= -1889612716;
assign addr[58860]= -2015345591;
assign addr[58861]= -2100237377;
assign addr[58862]= -2142567738;
assign addr[58863]= -2141478848;
assign addr[58864]= -2096992772;
assign addr[58865]= -2010011024;
assign addr[58866]= -1882296293;
assign addr[58867]= -1716436725;
assign addr[58868]= -1515793473;
assign addr[58869]= -1284432584;
assign addr[58870]= -1027042599;
assign addr[58871]= -748839539;
assign addr[58872]= -455461206;
assign addr[58873]= -152852926;
assign addr[58874]= 152852926;
assign addr[58875]= 455461206;
assign addr[58876]= 748839539;
assign addr[58877]= 1027042599;
assign addr[58878]= 1284432584;
assign addr[58879]= 1515793473;
assign addr[58880]= 1716436725;
assign addr[58881]= 1882296293;
assign addr[58882]= 2010011024;
assign addr[58883]= 2096992772;
assign addr[58884]= 2141478848;
assign addr[58885]= 2142567738;
assign addr[58886]= 2100237377;
assign addr[58887]= 2015345591;
assign addr[58888]= 1889612716;
assign addr[58889]= 1725586737;
assign addr[58890]= 1526591649;
assign addr[58891]= 1296660098;
assign addr[58892]= 1040451659;
assign addr[58893]= 763158411;
assign addr[58894]= 470399716;
assign addr[58895]= 168108346;
assign addr[58896]= -137589750;
assign addr[58897]= -440499581;
assign addr[58898]= -734482665;
assign addr[58899]= -1013581418;
assign addr[58900]= -1272139887;
assign addr[58901]= -1504918373;
assign addr[58902]= -1707199606;
assign addr[58903]= -1874884346;
assign addr[58904]= -2004574453;
assign addr[58905]= -2093641749;
assign addr[58906]= -2140281282;
assign addr[58907]= -2143547897;
assign addr[58908]= -2103375398;
assign addr[58909]= -2020577882;
assign addr[58910]= -1896833245;
assign addr[58911]= -1734649179;
assign addr[58912]= -1537312353;
assign addr[58913]= -1308821808;
assign addr[58914]= -1053807919;
assign addr[58915]= -777438554;
assign addr[58916]= -485314355;
assign addr[58917]= -183355234;
assign addr[58918]= 122319591;
assign addr[58919]= 425515602;
assign addr[58920]= 720088517;
assign addr[58921]= 1000068799;
assign addr[58922]= 1259782632;
assign addr[58923]= 1493966902;
assign addr[58924]= 1697875851;
assign addr[58925]= 1867377253;
assign addr[58926]= 1999036154;
assign addr[58927]= 2090184478;
assign addr[58928]= 2138975100;
assign addr[58929]= 2144419275;
assign addr[58930]= 2106406677;
assign addr[58931]= 2025707632;
assign addr[58932]= 1903957513;
assign addr[58933]= 1743623590;
assign addr[58934]= 1547955041;
assign addr[58935]= 1320917099;
assign addr[58936]= 1067110699;
assign addr[58937]= 791679244;
assign addr[58938]= 500204365;
assign addr[58939]= 198592817;
assign addr[58940]= -107043224;
assign addr[58941]= -410510029;
assign addr[58942]= -705657826;
assign addr[58943]= -986505429;
assign addr[58944]= -1247361445;
assign addr[58945]= -1482939614;
assign addr[58946]= -1688465931;
assign addr[58947]= -1859775393;
assign addr[58948]= -1993396407;
assign addr[58949]= -2086621133;
assign addr[58950]= -2137560369;
assign addr[58951]= -2145181827;
assign addr[58952]= -2109331059;
assign addr[58953]= -2030734582;
assign addr[58954]= -1910985158;
assign addr[58955]= -1752509516;
assign addr[58956]= -1558519173;
assign addr[58957]= -1332945355;
assign addr[58958]= -1080359326;
assign addr[58959]= -805879757;
assign addr[58960]= -515068990;
assign addr[58961]= -213820322;
assign addr[58962]= 91761426;
assign addr[58963]= 395483624;
assign addr[58964]= 691191324;
assign addr[58965]= 972891995;
assign addr[58966]= 1234876957;
assign addr[58967]= 1471837070;
assign addr[58968]= 1678970324;
assign addr[58969]= 1852079154;
assign addr[58970]= 1987655498;
assign addr[58971]= 2082951896;
assign addr[58972]= 2136037160;
assign addr[58973]= 2145835515;
assign addr[58974]= 2112148396;
assign addr[58975]= 2035658475;
assign addr[58976]= 1917915825;
assign addr[58977]= 1761306505;
assign addr[58978]= 1569004214;
assign addr[58979]= 1344905966;
assign addr[58980]= 1093553126;
assign addr[58981]= 820039373;
assign addr[58982]= 529907477;
assign addr[58983]= 229036977;
assign addr[58984]= -76474970;
assign addr[58985]= -380437148;
assign addr[58986]= -676689746;
assign addr[58987]= -959229189;
assign addr[58988]= -1222329801;
assign addr[58989]= -1460659832;
assign addr[58990]= -1669389513;
assign addr[58991]= -1844288924;
assign addr[58992]= -1981813720;
assign addr[58993]= -2079176953;
assign addr[58994]= -2134405552;
assign addr[58995]= -2146380306;
assign addr[58996]= -2114858546;
assign addr[58997]= -2040479063;
assign addr[58998]= -1924749160;
assign addr[58999]= -1770014111;
assign addr[59000]= -1579409630;
assign addr[59001]= -1356798326;
assign addr[59002]= -1106691431;
assign addr[59003]= -834157373;
assign addr[59004]= -544719071;
assign addr[59005]= -244242007;
assign addr[59006]= 61184634;
assign addr[59007]= 365371365;
assign addr[59008]= 662153826;
assign addr[59009]= 945517704;
assign addr[59010]= 1209720613;
assign addr[59011]= 1449408469;
assign addr[59012]= 1659723983;
assign addr[59013]= 1836405100;
assign addr[59014]= 1975871368;
assign addr[59015]= 2075296495;
assign addr[59016]= 2132665626;
assign addr[59017]= 2146816171;
assign addr[59018]= 2117461370;
assign addr[59019]= 2045196100;
assign addr[59020]= 1931484818;
assign addr[59021]= 1778631892;
assign addr[59022]= 1589734894;
assign addr[59023]= 1368621831;
assign addr[59024]= 1119773573;
assign addr[59025]= 848233042;
assign addr[59026]= 559503022;
assign addr[59027]= 259434643;
assign addr[59028]= -45891193;
assign addr[59029]= -350287041;
assign addr[59030]= -647584304;
assign addr[59031]= -931758235;
assign addr[59032]= -1197050035;
assign addr[59033]= -1438083551;
assign addr[59034]= -1649974225;
assign addr[59035]= -1828428082;
assign addr[59036]= -1969828744;
assign addr[59037]= -2071310720;
assign addr[59038]= -2130817471;
assign addr[59039]= -2147143090;
assign addr[59040]= -2119956737;
assign addr[59041]= -2049809346;
assign addr[59042]= -1938122457;
assign addr[59043]= -1787159411;
assign addr[59044]= -1599979481;
assign addr[59045]= -1380375881;
assign addr[59046]= -1132798888;
assign addr[59047]= -862265664;
assign addr[59048]= -574258580;
assign addr[59049]= -274614114;
assign addr[59050]= 30595422;
assign addr[59051]= 335184940;
assign addr[59052]= 632981917;
assign addr[59053]= 917951481;
assign addr[59054]= 1184318708;
assign addr[59055]= 1426685652;
assign addr[59056]= 1640140734;
assign addr[59057]= 1820358275;
assign addr[59058]= 1963686155;
assign addr[59059]= 2067219829;
assign addr[59060]= 2128861181;
assign addr[59061]= 2147361045;
assign addr[59062]= 2122344521;
assign addr[59063]= 2054318569;
assign addr[59064]= 1944661739;
assign addr[59065]= 1795596234;
assign addr[59066]= 1610142873;
assign addr[59067]= 1392059879;
assign addr[59068]= 1145766716;
assign addr[59069]= 876254528;
assign addr[59070]= 588984994;
assign addr[59071]= 289779648;
assign addr[59072]= -15298099;
assign addr[59073]= -320065829;
assign addr[59074]= -618347408;
assign addr[59075]= -904098143;
assign addr[59076]= -1171527280;
assign addr[59077]= -1415215352;
assign addr[59078]= -1630224009;
assign addr[59079]= -1812196087;
assign addr[59080]= -1957443913;
assign addr[59081]= -2063024031;
assign addr[59082]= -2126796855;
assign addr[59083]= -2147470025;
assign addr[59084]= -2124624598;
assign addr[59085]= -2058723538;
assign addr[59086]= -1951102334;
assign addr[59087]= -1803941934;
assign addr[59088]= -1620224553;
assign addr[59089]= -1403673233;
assign addr[59090]= -1158676398;
assign addr[59091]= -890198924;
assign addr[59092]= -603681519;
assign addr[59093]= -304930476;
assign addr[59094]= 0;
assign addr[59095]= 304930476;
assign addr[59096]= 603681519;
assign addr[59097]= 890198924;
assign addr[59098]= 1158676398;
assign addr[59099]= 1403673233;
assign addr[59100]= 1620224553;
assign addr[59101]= 1803941934;
assign addr[59102]= 1951102334;
assign addr[59103]= 2058723538;
assign addr[59104]= 2124624598;
assign addr[59105]= 2147470025;
assign addr[59106]= 2126796855;
assign addr[59107]= 2063024031;
assign addr[59108]= 1957443913;
assign addr[59109]= 1812196087;
assign addr[59110]= 1630224009;
assign addr[59111]= 1415215352;
assign addr[59112]= 1171527280;
assign addr[59113]= 904098143;
assign addr[59114]= 618347408;
assign addr[59115]= 320065829;
assign addr[59116]= 15298099;
assign addr[59117]= -289779648;
assign addr[59118]= -588984994;
assign addr[59119]= -876254528;
assign addr[59120]= -1145766716;
assign addr[59121]= -1392059879;
assign addr[59122]= -1610142873;
assign addr[59123]= -1795596234;
assign addr[59124]= -1944661739;
assign addr[59125]= -2054318569;
assign addr[59126]= -2122344521;
assign addr[59127]= -2147361045;
assign addr[59128]= -2128861181;
assign addr[59129]= -2067219829;
assign addr[59130]= -1963686155;
assign addr[59131]= -1820358275;
assign addr[59132]= -1640140734;
assign addr[59133]= -1426685652;
assign addr[59134]= -1184318708;
assign addr[59135]= -917951481;
assign addr[59136]= -632981917;
assign addr[59137]= -335184940;
assign addr[59138]= -30595422;
assign addr[59139]= 274614114;
assign addr[59140]= 574258580;
assign addr[59141]= 862265664;
assign addr[59142]= 1132798888;
assign addr[59143]= 1380375881;
assign addr[59144]= 1599979481;
assign addr[59145]= 1787159411;
assign addr[59146]= 1938122457;
assign addr[59147]= 2049809346;
assign addr[59148]= 2119956737;
assign addr[59149]= 2147143090;
assign addr[59150]= 2130817471;
assign addr[59151]= 2071310720;
assign addr[59152]= 1969828744;
assign addr[59153]= 1828428082;
assign addr[59154]= 1649974225;
assign addr[59155]= 1438083551;
assign addr[59156]= 1197050035;
assign addr[59157]= 931758235;
assign addr[59158]= 647584304;
assign addr[59159]= 350287041;
assign addr[59160]= 45891193;
assign addr[59161]= -259434643;
assign addr[59162]= -559503022;
assign addr[59163]= -848233042;
assign addr[59164]= -1119773573;
assign addr[59165]= -1368621831;
assign addr[59166]= -1589734894;
assign addr[59167]= -1778631892;
assign addr[59168]= -1931484818;
assign addr[59169]= -2045196100;
assign addr[59170]= -2117461370;
assign addr[59171]= -2146816171;
assign addr[59172]= -2132665626;
assign addr[59173]= -2075296495;
assign addr[59174]= -1975871368;
assign addr[59175]= -1836405100;
assign addr[59176]= -1659723983;
assign addr[59177]= -1449408469;
assign addr[59178]= -1209720613;
assign addr[59179]= -945517704;
assign addr[59180]= -662153826;
assign addr[59181]= -365371365;
assign addr[59182]= -61184634;
assign addr[59183]= 244242007;
assign addr[59184]= 544719071;
assign addr[59185]= 834157373;
assign addr[59186]= 1106691431;
assign addr[59187]= 1356798326;
assign addr[59188]= 1579409630;
assign addr[59189]= 1770014111;
assign addr[59190]= 1924749160;
assign addr[59191]= 2040479063;
assign addr[59192]= 2114858546;
assign addr[59193]= 2146380306;
assign addr[59194]= 2134405552;
assign addr[59195]= 2079176953;
assign addr[59196]= 1981813720;
assign addr[59197]= 1844288924;
assign addr[59198]= 1669389513;
assign addr[59199]= 1460659832;
assign addr[59200]= 1222329801;
assign addr[59201]= 959229189;
assign addr[59202]= 676689746;
assign addr[59203]= 380437148;
assign addr[59204]= 76474970;
assign addr[59205]= -229036977;
assign addr[59206]= -529907477;
assign addr[59207]= -820039373;
assign addr[59208]= -1093553126;
assign addr[59209]= -1344905966;
assign addr[59210]= -1569004214;
assign addr[59211]= -1761306505;
assign addr[59212]= -1917915825;
assign addr[59213]= -2035658475;
assign addr[59214]= -2112148396;
assign addr[59215]= -2145835515;
assign addr[59216]= -2136037160;
assign addr[59217]= -2082951896;
assign addr[59218]= -1987655498;
assign addr[59219]= -1852079154;
assign addr[59220]= -1678970324;
assign addr[59221]= -1471837070;
assign addr[59222]= -1234876957;
assign addr[59223]= -972891995;
assign addr[59224]= -691191324;
assign addr[59225]= -395483624;
assign addr[59226]= -91761426;
assign addr[59227]= 213820322;
assign addr[59228]= 515068990;
assign addr[59229]= 805879757;
assign addr[59230]= 1080359326;
assign addr[59231]= 1332945355;
assign addr[59232]= 1558519173;
assign addr[59233]= 1752509516;
assign addr[59234]= 1910985158;
assign addr[59235]= 2030734582;
assign addr[59236]= 2109331059;
assign addr[59237]= 2145181827;
assign addr[59238]= 2137560369;
assign addr[59239]= 2086621133;
assign addr[59240]= 1993396407;
assign addr[59241]= 1859775393;
assign addr[59242]= 1688465931;
assign addr[59243]= 1482939614;
assign addr[59244]= 1247361445;
assign addr[59245]= 986505429;
assign addr[59246]= 705657826;
assign addr[59247]= 410510029;
assign addr[59248]= 107043224;
assign addr[59249]= -198592817;
assign addr[59250]= -500204365;
assign addr[59251]= -791679244;
assign addr[59252]= -1067110699;
assign addr[59253]= -1320917099;
assign addr[59254]= -1547955041;
assign addr[59255]= -1743623590;
assign addr[59256]= -1903957513;
assign addr[59257]= -2025707632;
assign addr[59258]= -2106406677;
assign addr[59259]= -2144419275;
assign addr[59260]= -2138975100;
assign addr[59261]= -2090184478;
assign addr[59262]= -1999036154;
assign addr[59263]= -1867377253;
assign addr[59264]= -1697875851;
assign addr[59265]= -1493966902;
assign addr[59266]= -1259782632;
assign addr[59267]= -1000068799;
assign addr[59268]= -720088517;
assign addr[59269]= -425515602;
assign addr[59270]= -122319591;
assign addr[59271]= 183355234;
assign addr[59272]= 485314355;
assign addr[59273]= 777438554;
assign addr[59274]= 1053807919;
assign addr[59275]= 1308821808;
assign addr[59276]= 1537312353;
assign addr[59277]= 1734649179;
assign addr[59278]= 1896833245;
assign addr[59279]= 2020577882;
assign addr[59280]= 2103375398;
assign addr[59281]= 2143547897;
assign addr[59282]= 2140281282;
assign addr[59283]= 2093641749;
assign addr[59284]= 2004574453;
assign addr[59285]= 1874884346;
assign addr[59286]= 1707199606;
assign addr[59287]= 1504918373;
assign addr[59288]= 1272139887;
assign addr[59289]= 1013581418;
assign addr[59290]= 734482665;
assign addr[59291]= 440499581;
assign addr[59292]= 137589750;
assign addr[59293]= -168108346;
assign addr[59294]= -470399716;
assign addr[59295]= -763158411;
assign addr[59296]= -1040451659;
assign addr[59297]= -1296660098;
assign addr[59298]= -1526591649;
assign addr[59299]= -1725586737;
assign addr[59300]= -1889612716;
assign addr[59301]= -2015345591;
assign addr[59302]= -2100237377;
assign addr[59303]= -2142567738;
assign addr[59304]= -2141478848;
assign addr[59305]= -2096992772;
assign addr[59306]= -2010011024;
assign addr[59307]= -1882296293;
assign addr[59308]= -1716436725;
assign addr[59309]= -1515793473;
assign addr[59310]= -1284432584;
assign addr[59311]= -1027042599;
assign addr[59312]= -748839539;
assign addr[59313]= -455461206;
assign addr[59314]= -152852926;
assign addr[59315]= 152852926;
assign addr[59316]= 455461206;
assign addr[59317]= 748839539;
assign addr[59318]= 1027042599;
assign addr[59319]= 1284432584;
assign addr[59320]= 1515793473;
assign addr[59321]= 1716436725;
assign addr[59322]= 1882296293;
assign addr[59323]= 2010011024;
assign addr[59324]= 2096992772;
assign addr[59325]= 2141478848;
assign addr[59326]= 2142567738;
assign addr[59327]= 2100237377;
assign addr[59328]= 2015345591;
assign addr[59329]= 1889612716;
assign addr[59330]= 1725586737;
assign addr[59331]= 1526591649;
assign addr[59332]= 1296660098;
assign addr[59333]= 1040451659;
assign addr[59334]= 763158411;
assign addr[59335]= 470399716;
assign addr[59336]= 168108346;
assign addr[59337]= -137589750;
assign addr[59338]= -440499581;
assign addr[59339]= -734482665;
assign addr[59340]= -1013581418;
assign addr[59341]= -1272139887;
assign addr[59342]= -1504918373;
assign addr[59343]= -1707199606;
assign addr[59344]= -1874884346;
assign addr[59345]= -2004574453;
assign addr[59346]= -2093641749;
assign addr[59347]= -2140281282;
assign addr[59348]= -2143547897;
assign addr[59349]= -2103375398;
assign addr[59350]= -2020577882;
assign addr[59351]= -1896833245;
assign addr[59352]= -1734649179;
assign addr[59353]= -1537312353;
assign addr[59354]= -1308821808;
assign addr[59355]= -1053807919;
assign addr[59356]= -777438554;
assign addr[59357]= -485314355;
assign addr[59358]= -183355234;
assign addr[59359]= 122319591;
assign addr[59360]= 425515602;
assign addr[59361]= 720088517;
assign addr[59362]= 1000068799;
assign addr[59363]= 1259782632;
assign addr[59364]= 1493966902;
assign addr[59365]= 1697875851;
assign addr[59366]= 1867377253;
assign addr[59367]= 1999036154;
assign addr[59368]= 2090184478;
assign addr[59369]= 2138975100;
assign addr[59370]= 2144419275;
assign addr[59371]= 2106406677;
assign addr[59372]= 2025707632;
assign addr[59373]= 1903957513;
assign addr[59374]= 1743623590;
assign addr[59375]= 1547955041;
assign addr[59376]= 1320917099;
assign addr[59377]= 1067110699;
assign addr[59378]= 791679244;
assign addr[59379]= 500204365;
assign addr[59380]= 198592817;
assign addr[59381]= -107043224;
assign addr[59382]= -410510029;
assign addr[59383]= -705657826;
assign addr[59384]= -986505429;
assign addr[59385]= -1247361445;
assign addr[59386]= -1482939614;
assign addr[59387]= -1688465931;
assign addr[59388]= -1859775393;
assign addr[59389]= -1993396407;
assign addr[59390]= -2086621133;
assign addr[59391]= -2137560369;
assign addr[59392]= -2145181827;
assign addr[59393]= -2109331059;
assign addr[59394]= -2030734582;
assign addr[59395]= -1910985158;
assign addr[59396]= -1752509516;
assign addr[59397]= -1558519173;
assign addr[59398]= -1332945355;
assign addr[59399]= -1080359326;
assign addr[59400]= -805879757;
assign addr[59401]= -515068990;
assign addr[59402]= -213820322;
assign addr[59403]= 91761426;
assign addr[59404]= 395483624;
assign addr[59405]= 691191324;
assign addr[59406]= 972891995;
assign addr[59407]= 1234876957;
assign addr[59408]= 1471837070;
assign addr[59409]= 1678970324;
assign addr[59410]= 1852079154;
assign addr[59411]= 1987655498;
assign addr[59412]= 2082951896;
assign addr[59413]= 2136037160;
assign addr[59414]= 2145835515;
assign addr[59415]= 2112148396;
assign addr[59416]= 2035658475;
assign addr[59417]= 1917915825;
assign addr[59418]= 1761306505;
assign addr[59419]= 1569004214;
assign addr[59420]= 1344905966;
assign addr[59421]= 1093553126;
assign addr[59422]= 820039373;
assign addr[59423]= 529907477;
assign addr[59424]= 229036977;
assign addr[59425]= -76474970;
assign addr[59426]= -380437148;
assign addr[59427]= -676689746;
assign addr[59428]= -959229189;
assign addr[59429]= -1222329801;
assign addr[59430]= -1460659832;
assign addr[59431]= -1669389513;
assign addr[59432]= -1844288924;
assign addr[59433]= -1981813720;
assign addr[59434]= -2079176953;
assign addr[59435]= -2134405552;
assign addr[59436]= -2146380306;
assign addr[59437]= -2114858546;
assign addr[59438]= -2040479063;
assign addr[59439]= -1924749160;
assign addr[59440]= -1770014111;
assign addr[59441]= -1579409630;
assign addr[59442]= -1356798326;
assign addr[59443]= -1106691431;
assign addr[59444]= -834157373;
assign addr[59445]= -544719071;
assign addr[59446]= -244242007;
assign addr[59447]= 61184634;
assign addr[59448]= 365371365;
assign addr[59449]= 662153826;
assign addr[59450]= 945517704;
assign addr[59451]= 1209720613;
assign addr[59452]= 1449408469;
assign addr[59453]= 1659723983;
assign addr[59454]= 1836405100;
assign addr[59455]= 1975871368;
assign addr[59456]= 2075296495;
assign addr[59457]= 2132665626;
assign addr[59458]= 2146816171;
assign addr[59459]= 2117461370;
assign addr[59460]= 2045196100;
assign addr[59461]= 1931484818;
assign addr[59462]= 1778631892;
assign addr[59463]= 1589734894;
assign addr[59464]= 1368621831;
assign addr[59465]= 1119773573;
assign addr[59466]= 848233042;
assign addr[59467]= 559503022;
assign addr[59468]= 259434643;
assign addr[59469]= -45891193;
assign addr[59470]= -350287041;
assign addr[59471]= -647584304;
assign addr[59472]= -931758235;
assign addr[59473]= -1197050035;
assign addr[59474]= -1438083551;
assign addr[59475]= -1649974225;
assign addr[59476]= -1828428082;
assign addr[59477]= -1969828744;
assign addr[59478]= -2071310720;
assign addr[59479]= -2130817471;
assign addr[59480]= -2147143090;
assign addr[59481]= -2119956737;
assign addr[59482]= -2049809346;
assign addr[59483]= -1938122457;
assign addr[59484]= -1787159411;
assign addr[59485]= -1599979481;
assign addr[59486]= -1380375881;
assign addr[59487]= -1132798888;
assign addr[59488]= -862265664;
assign addr[59489]= -574258580;
assign addr[59490]= -274614114;
assign addr[59491]= 30595422;
assign addr[59492]= 335184940;
assign addr[59493]= 632981917;
assign addr[59494]= 917951481;
assign addr[59495]= 1184318708;
assign addr[59496]= 1426685652;
assign addr[59497]= 1640140734;
assign addr[59498]= 1820358275;
assign addr[59499]= 1963686155;
assign addr[59500]= 2067219829;
assign addr[59501]= 2128861181;
assign addr[59502]= 2147361045;
assign addr[59503]= 2122344521;
assign addr[59504]= 2054318569;
assign addr[59505]= 1944661739;
assign addr[59506]= 1795596234;
assign addr[59507]= 1610142873;
assign addr[59508]= 1392059879;
assign addr[59509]= 1145766716;
assign addr[59510]= 876254528;
assign addr[59511]= 588984994;
assign addr[59512]= 289779648;
assign addr[59513]= -15298099;
assign addr[59514]= -320065829;
assign addr[59515]= -618347408;
assign addr[59516]= -904098143;
assign addr[59517]= -1171527280;
assign addr[59518]= -1415215352;
assign addr[59519]= -1630224009;
assign addr[59520]= -1812196087;
assign addr[59521]= -1957443913;
assign addr[59522]= -2063024031;
assign addr[59523]= -2126796855;
assign addr[59524]= -2147470025;
assign addr[59525]= -2124624598;
assign addr[59526]= -2058723538;
assign addr[59527]= -1951102334;
assign addr[59528]= -1803941934;
assign addr[59529]= -1620224553;
assign addr[59530]= -1403673233;
assign addr[59531]= -1158676398;
assign addr[59532]= -890198924;
assign addr[59533]= -603681519;
assign addr[59534]= -304930476;
assign addr[59535]= 0;
assign addr[59536]= 304930476;
assign addr[59537]= 603681519;
assign addr[59538]= 890198924;
assign addr[59539]= 1158676398;
assign addr[59540]= 1403673233;
assign addr[59541]= 1620224553;
assign addr[59542]= 1803941934;
assign addr[59543]= 1951102334;
assign addr[59544]= 2058723538;
assign addr[59545]= 2124624598;
assign addr[59546]= 2147470025;
assign addr[59547]= 2126796855;
assign addr[59548]= 2063024031;
assign addr[59549]= 1957443913;
assign addr[59550]= 1812196087;
assign addr[59551]= 1630224009;
assign addr[59552]= 1415215352;
assign addr[59553]= 1171527280;
assign addr[59554]= 904098143;
assign addr[59555]= 618347408;
assign addr[59556]= 320065829;
assign addr[59557]= 15298099;
assign addr[59558]= -289779648;
assign addr[59559]= -588984994;
assign addr[59560]= -876254528;
assign addr[59561]= -1145766716;
assign addr[59562]= -1392059879;
assign addr[59563]= -1610142873;
assign addr[59564]= -1795596234;
assign addr[59565]= -1944661739;
assign addr[59566]= -2054318569;
assign addr[59567]= -2122344521;
assign addr[59568]= -2147361045;
assign addr[59569]= -2128861181;
assign addr[59570]= -2067219829;
assign addr[59571]= -1963686155;
assign addr[59572]= -1820358275;
assign addr[59573]= -1640140734;
assign addr[59574]= -1426685652;
assign addr[59575]= -1184318708;
assign addr[59576]= -917951481;
assign addr[59577]= -632981917;
assign addr[59578]= -335184940;
assign addr[59579]= -30595422;
assign addr[59580]= 274614114;
assign addr[59581]= 574258580;
assign addr[59582]= 862265664;
assign addr[59583]= 1132798888;
assign addr[59584]= 1380375881;
assign addr[59585]= 1599979481;
assign addr[59586]= 1787159411;
assign addr[59587]= 1938122457;
assign addr[59588]= 2049809346;
assign addr[59589]= 2119956737;
assign addr[59590]= 2147143090;
assign addr[59591]= 2130817471;
assign addr[59592]= 2071310720;
assign addr[59593]= 1969828744;
assign addr[59594]= 1828428082;
assign addr[59595]= 1649974225;
assign addr[59596]= 1438083551;
assign addr[59597]= 1197050035;
assign addr[59598]= 931758235;
assign addr[59599]= 647584304;
assign addr[59600]= 350287041;
assign addr[59601]= 45891193;
assign addr[59602]= -259434643;
assign addr[59603]= -559503022;
assign addr[59604]= -848233042;
assign addr[59605]= -1119773573;
assign addr[59606]= -1368621831;
assign addr[59607]= -1589734894;
assign addr[59608]= -1778631892;
assign addr[59609]= -1931484818;
assign addr[59610]= -2045196100;
assign addr[59611]= -2117461370;
assign addr[59612]= -2146816171;
assign addr[59613]= -2132665626;
assign addr[59614]= -2075296495;
assign addr[59615]= -1975871368;
assign addr[59616]= -1836405100;
assign addr[59617]= -1659723983;
assign addr[59618]= -1449408469;
assign addr[59619]= -1209720613;
assign addr[59620]= -945517704;
assign addr[59621]= -662153826;
assign addr[59622]= -365371365;
assign addr[59623]= -61184634;
assign addr[59624]= 244242007;
assign addr[59625]= 544719071;
assign addr[59626]= 834157373;
assign addr[59627]= 1106691431;
assign addr[59628]= 1356798326;
assign addr[59629]= 1579409630;
assign addr[59630]= 1770014111;
assign addr[59631]= 1924749160;
assign addr[59632]= 2040479063;
assign addr[59633]= 2114858546;
assign addr[59634]= 2146380306;
assign addr[59635]= 2134405552;
assign addr[59636]= 2079176953;
assign addr[59637]= 1981813720;
assign addr[59638]= 1844288924;
assign addr[59639]= 1669389513;
assign addr[59640]= 1460659832;
assign addr[59641]= 1222329801;
assign addr[59642]= 959229189;
assign addr[59643]= 676689746;
assign addr[59644]= 380437148;
assign addr[59645]= 76474970;
assign addr[59646]= -229036977;
assign addr[59647]= -529907477;
assign addr[59648]= -820039373;
assign addr[59649]= -1093553126;
assign addr[59650]= -1344905966;
assign addr[59651]= -1569004214;
assign addr[59652]= -1761306505;
assign addr[59653]= -1917915825;
assign addr[59654]= -2035658475;
assign addr[59655]= -2112148396;
assign addr[59656]= -2145835515;
assign addr[59657]= -2136037160;
assign addr[59658]= -2082951896;
assign addr[59659]= -1987655498;
assign addr[59660]= -1852079154;
assign addr[59661]= -1678970324;
assign addr[59662]= -1471837070;
assign addr[59663]= -1234876957;
assign addr[59664]= -972891995;
assign addr[59665]= -691191324;
assign addr[59666]= -395483624;
assign addr[59667]= -91761426;
assign addr[59668]= 213820322;
assign addr[59669]= 515068990;
assign addr[59670]= 805879757;
assign addr[59671]= 1080359326;
assign addr[59672]= 1332945355;
assign addr[59673]= 1558519173;
assign addr[59674]= 1752509516;
assign addr[59675]= 1910985158;
assign addr[59676]= 2030734582;
assign addr[59677]= 2109331059;
assign addr[59678]= 2145181827;
assign addr[59679]= 2137560369;
assign addr[59680]= 2086621133;
assign addr[59681]= 1993396407;
assign addr[59682]= 1859775393;
assign addr[59683]= 1688465931;
assign addr[59684]= 1482939614;
assign addr[59685]= 1247361445;
assign addr[59686]= 986505429;
assign addr[59687]= 705657826;
assign addr[59688]= 410510029;
assign addr[59689]= 107043224;
assign addr[59690]= -198592817;
assign addr[59691]= -500204365;
assign addr[59692]= -791679244;
assign addr[59693]= -1067110699;
assign addr[59694]= -1320917099;
assign addr[59695]= -1547955041;
assign addr[59696]= -1743623590;
assign addr[59697]= -1903957513;
assign addr[59698]= -2025707632;
assign addr[59699]= -2106406677;
assign addr[59700]= -2144419275;
assign addr[59701]= -2138975100;
assign addr[59702]= -2090184478;
assign addr[59703]= -1999036154;
assign addr[59704]= -1867377253;
assign addr[59705]= -1697875851;
assign addr[59706]= -1493966902;
assign addr[59707]= -1259782632;
assign addr[59708]= -1000068799;
assign addr[59709]= -720088517;
assign addr[59710]= -425515602;
assign addr[59711]= -122319591;
assign addr[59712]= 183355234;
assign addr[59713]= 485314355;
assign addr[59714]= 777438554;
assign addr[59715]= 1053807919;
assign addr[59716]= 1308821808;
assign addr[59717]= 1537312353;
assign addr[59718]= 1734649179;
assign addr[59719]= 1896833245;
assign addr[59720]= 2020577882;
assign addr[59721]= 2103375398;
assign addr[59722]= 2143547897;
assign addr[59723]= 2140281282;
assign addr[59724]= 2093641749;
assign addr[59725]= 2004574453;
assign addr[59726]= 1874884346;
assign addr[59727]= 1707199606;
assign addr[59728]= 1504918373;
assign addr[59729]= 1272139887;
assign addr[59730]= 1013581418;
assign addr[59731]= 734482665;
assign addr[59732]= 440499581;
assign addr[59733]= 137589750;
assign addr[59734]= -168108346;
assign addr[59735]= -470399716;
assign addr[59736]= -763158411;
assign addr[59737]= -1040451659;
assign addr[59738]= -1296660098;
assign addr[59739]= -1526591649;
assign addr[59740]= -1725586737;
assign addr[59741]= -1889612716;
assign addr[59742]= -2015345591;
assign addr[59743]= -2100237377;
assign addr[59744]= -2142567738;
assign addr[59745]= -2141478848;
assign addr[59746]= -2096992772;
assign addr[59747]= -2010011024;
assign addr[59748]= -1882296293;
assign addr[59749]= -1716436725;
assign addr[59750]= -1515793473;
assign addr[59751]= -1284432584;
assign addr[59752]= -1027042599;
assign addr[59753]= -748839539;
assign addr[59754]= -455461206;
assign addr[59755]= -152852926;
assign addr[59756]= 152852926;
assign addr[59757]= 455461206;
assign addr[59758]= 748839539;
assign addr[59759]= 1027042599;
assign addr[59760]= 1284432584;
assign addr[59761]= 1515793473;
assign addr[59762]= 1716436725;
assign addr[59763]= 1882296293;
assign addr[59764]= 2010011024;
assign addr[59765]= 2096992772;
assign addr[59766]= 2141478848;
assign addr[59767]= 2142567738;
assign addr[59768]= 2100237377;
assign addr[59769]= 2015345591;
assign addr[59770]= 1889612716;
assign addr[59771]= 1725586737;
assign addr[59772]= 1526591649;
assign addr[59773]= 1296660098;
assign addr[59774]= 1040451659;
assign addr[59775]= 763158411;
assign addr[59776]= 470399716;
assign addr[59777]= 168108346;
assign addr[59778]= -137589750;
assign addr[59779]= -440499581;
assign addr[59780]= -734482665;
assign addr[59781]= -1013581418;
assign addr[59782]= -1272139887;
assign addr[59783]= -1504918373;
assign addr[59784]= -1707199606;
assign addr[59785]= -1874884346;
assign addr[59786]= -2004574453;
assign addr[59787]= -2093641749;
assign addr[59788]= -2140281282;
assign addr[59789]= -2143547897;
assign addr[59790]= -2103375398;
assign addr[59791]= -2020577882;
assign addr[59792]= -1896833245;
assign addr[59793]= -1734649179;
assign addr[59794]= -1537312353;
assign addr[59795]= -1308821808;
assign addr[59796]= -1053807919;
assign addr[59797]= -777438554;
assign addr[59798]= -485314355;
assign addr[59799]= -183355234;
assign addr[59800]= 122319591;
assign addr[59801]= 425515602;
assign addr[59802]= 720088517;
assign addr[59803]= 1000068799;
assign addr[59804]= 1259782632;
assign addr[59805]= 1493966902;
assign addr[59806]= 1697875851;
assign addr[59807]= 1867377253;
assign addr[59808]= 1999036154;
assign addr[59809]= 2090184478;
assign addr[59810]= 2138975100;
assign addr[59811]= 2144419275;
assign addr[59812]= 2106406677;
assign addr[59813]= 2025707632;
assign addr[59814]= 1903957513;
assign addr[59815]= 1743623590;
assign addr[59816]= 1547955041;
assign addr[59817]= 1320917099;
assign addr[59818]= 1067110699;
assign addr[59819]= 791679244;
assign addr[59820]= 500204365;
assign addr[59821]= 198592817;
assign addr[59822]= -107043224;
assign addr[59823]= -410510029;
assign addr[59824]= -705657826;
assign addr[59825]= -986505429;
assign addr[59826]= -1247361445;
assign addr[59827]= -1482939614;
assign addr[59828]= -1688465931;
assign addr[59829]= -1859775393;
assign addr[59830]= -1993396407;
assign addr[59831]= -2086621133;
assign addr[59832]= -2137560369;
assign addr[59833]= -2145181827;
assign addr[59834]= -2109331059;
assign addr[59835]= -2030734582;
assign addr[59836]= -1910985158;
assign addr[59837]= -1752509516;
assign addr[59838]= -1558519173;
assign addr[59839]= -1332945355;
assign addr[59840]= -1080359326;
assign addr[59841]= -805879757;
assign addr[59842]= -515068990;
assign addr[59843]= -213820322;
assign addr[59844]= 91761426;
assign addr[59845]= 395483624;
assign addr[59846]= 691191324;
assign addr[59847]= 972891995;
assign addr[59848]= 1234876957;
assign addr[59849]= 1471837070;
assign addr[59850]= 1678970324;
assign addr[59851]= 1852079154;
assign addr[59852]= 1987655498;
assign addr[59853]= 2082951896;
assign addr[59854]= 2136037160;
assign addr[59855]= 2145835515;
assign addr[59856]= 2112148396;
assign addr[59857]= 2035658475;
assign addr[59858]= 1917915825;
assign addr[59859]= 1761306505;
assign addr[59860]= 1569004214;
assign addr[59861]= 1344905966;
assign addr[59862]= 1093553126;
assign addr[59863]= 820039373;
assign addr[59864]= 529907477;
assign addr[59865]= 229036977;
assign addr[59866]= -76474970;
assign addr[59867]= -380437148;
assign addr[59868]= -676689746;
assign addr[59869]= -959229189;
assign addr[59870]= -1222329801;
assign addr[59871]= -1460659832;
assign addr[59872]= -1669389513;
assign addr[59873]= -1844288924;
assign addr[59874]= -1981813720;
assign addr[59875]= -2079176953;
assign addr[59876]= -2134405552;
assign addr[59877]= -2146380306;
assign addr[59878]= -2114858546;
assign addr[59879]= -2040479063;
assign addr[59880]= -1924749160;
assign addr[59881]= -1770014111;
assign addr[59882]= -1579409630;
assign addr[59883]= -1356798326;
assign addr[59884]= -1106691431;
assign addr[59885]= -834157373;
assign addr[59886]= -544719071;
assign addr[59887]= -244242007;
assign addr[59888]= 61184634;
assign addr[59889]= 365371365;
assign addr[59890]= 662153826;
assign addr[59891]= 945517704;
assign addr[59892]= 1209720613;
assign addr[59893]= 1449408469;
assign addr[59894]= 1659723983;
assign addr[59895]= 1836405100;
assign addr[59896]= 1975871368;
assign addr[59897]= 2075296495;
assign addr[59898]= 2132665626;
assign addr[59899]= 2146816171;
assign addr[59900]= 2117461370;
assign addr[59901]= 2045196100;
assign addr[59902]= 1931484818;
assign addr[59903]= 1778631892;
assign addr[59904]= 1589734894;
assign addr[59905]= 1368621831;
assign addr[59906]= 1119773573;
assign addr[59907]= 848233042;
assign addr[59908]= 559503022;
assign addr[59909]= 259434643;
assign addr[59910]= -45891193;
assign addr[59911]= -350287041;
assign addr[59912]= -647584304;
assign addr[59913]= -931758235;
assign addr[59914]= -1197050035;
assign addr[59915]= -1438083551;
assign addr[59916]= -1649974225;
assign addr[59917]= -1828428082;
assign addr[59918]= -1969828744;
assign addr[59919]= -2071310720;
assign addr[59920]= -2130817471;
assign addr[59921]= -2147143090;
assign addr[59922]= -2119956737;
assign addr[59923]= -2049809346;
assign addr[59924]= -1938122457;
assign addr[59925]= -1787159411;
assign addr[59926]= -1599979481;
assign addr[59927]= -1380375881;
assign addr[59928]= -1132798888;
assign addr[59929]= -862265664;
assign addr[59930]= -574258580;
assign addr[59931]= -274614114;
assign addr[59932]= 30595422;
assign addr[59933]= 335184940;
assign addr[59934]= 632981917;
assign addr[59935]= 917951481;
assign addr[59936]= 1184318708;
assign addr[59937]= 1426685652;
assign addr[59938]= 1640140734;
assign addr[59939]= 1820358275;
assign addr[59940]= 1963686155;
assign addr[59941]= 2067219829;
assign addr[59942]= 2128861181;
assign addr[59943]= 2147361045;
assign addr[59944]= 2122344521;
assign addr[59945]= 2054318569;
assign addr[59946]= 1944661739;
assign addr[59947]= 1795596234;
assign addr[59948]= 1610142873;
assign addr[59949]= 1392059879;
assign addr[59950]= 1145766716;
assign addr[59951]= 876254528;
assign addr[59952]= 588984994;
assign addr[59953]= 289779648;
assign addr[59954]= -15298099;
assign addr[59955]= -320065829;
assign addr[59956]= -618347408;
assign addr[59957]= -904098143;
assign addr[59958]= -1171527280;
assign addr[59959]= -1415215352;
assign addr[59960]= -1630224009;
assign addr[59961]= -1812196087;
assign addr[59962]= -1957443913;
assign addr[59963]= -2063024031;
assign addr[59964]= -2126796855;
assign addr[59965]= -2147470025;
assign addr[59966]= -2124624598;
assign addr[59967]= -2058723538;
assign addr[59968]= -1951102334;
assign addr[59969]= -1803941934;
assign addr[59970]= -1620224553;
assign addr[59971]= -1403673233;
assign addr[59972]= -1158676398;
assign addr[59973]= -890198924;
assign addr[59974]= -603681519;
assign addr[59975]= -304930476;
assign addr[59976]= 0;
assign addr[59977]= 304930476;
assign addr[59978]= 603681519;
assign addr[59979]= 890198924;
assign addr[59980]= 1158676398;
assign addr[59981]= 1403673233;
assign addr[59982]= 1620224553;
assign addr[59983]= 1803941934;
assign addr[59984]= 1951102334;
assign addr[59985]= 2058723538;
assign addr[59986]= 2124624598;
assign addr[59987]= 2147470025;
assign addr[59988]= 2126796855;
assign addr[59989]= 2063024031;
assign addr[59990]= 1957443913;
assign addr[59991]= 1812196087;
assign addr[59992]= 1630224009;
assign addr[59993]= 1415215352;
assign addr[59994]= 1171527280;
assign addr[59995]= 904098143;
assign addr[59996]= 618347408;
assign addr[59997]= 320065829;
assign addr[59998]= 15298099;
assign addr[59999]= -289779648;
assign addr[60000]= -588984994;
assign addr[60001]= -876254528;
assign addr[60002]= -1145766716;
assign addr[60003]= -1392059879;
assign addr[60004]= -1610142873;
assign addr[60005]= -1795596234;
assign addr[60006]= -1944661739;
assign addr[60007]= -2054318569;
assign addr[60008]= -2122344521;
assign addr[60009]= -2147361045;
assign addr[60010]= -2128861181;
assign addr[60011]= -2067219829;
assign addr[60012]= -1963686155;
assign addr[60013]= -1820358275;
assign addr[60014]= -1640140734;
assign addr[60015]= -1426685652;
assign addr[60016]= -1184318708;
assign addr[60017]= -917951481;
assign addr[60018]= -632981917;
assign addr[60019]= -335184940;
assign addr[60020]= -30595422;
assign addr[60021]= 274614114;
assign addr[60022]= 574258580;
assign addr[60023]= 862265664;
assign addr[60024]= 1132798888;
assign addr[60025]= 1380375881;
assign addr[60026]= 1599979481;
assign addr[60027]= 1787159411;
assign addr[60028]= 1938122457;
assign addr[60029]= 2049809346;
assign addr[60030]= 2119956737;
assign addr[60031]= 2147143090;
assign addr[60032]= 2130817471;
assign addr[60033]= 2071310720;
assign addr[60034]= 1969828744;
assign addr[60035]= 1828428082;
assign addr[60036]= 1649974225;
assign addr[60037]= 1438083551;
assign addr[60038]= 1197050035;
assign addr[60039]= 931758235;
assign addr[60040]= 647584304;
assign addr[60041]= 350287041;
assign addr[60042]= 45891193;
assign addr[60043]= -259434643;
assign addr[60044]= -559503022;
assign addr[60045]= -848233042;
assign addr[60046]= -1119773573;
assign addr[60047]= -1368621831;
assign addr[60048]= -1589734894;
assign addr[60049]= -1778631892;
assign addr[60050]= -1931484818;
assign addr[60051]= -2045196100;
assign addr[60052]= -2117461370;
assign addr[60053]= -2146816171;
assign addr[60054]= -2132665626;
assign addr[60055]= -2075296495;
assign addr[60056]= -1975871368;
assign addr[60057]= -1836405100;
assign addr[60058]= -1659723983;
assign addr[60059]= -1449408469;
assign addr[60060]= -1209720613;
assign addr[60061]= -945517704;
assign addr[60062]= -662153826;
assign addr[60063]= -365371365;
assign addr[60064]= -61184634;
assign addr[60065]= 244242007;
assign addr[60066]= 544719071;
assign addr[60067]= 834157373;
assign addr[60068]= 1106691431;
assign addr[60069]= 1356798326;
assign addr[60070]= 1579409630;
assign addr[60071]= 1770014111;
assign addr[60072]= 1924749160;
assign addr[60073]= 2040479063;
assign addr[60074]= 2114858546;
assign addr[60075]= 2146380306;
assign addr[60076]= 2134405552;
assign addr[60077]= 2079176953;
assign addr[60078]= 1981813720;
assign addr[60079]= 1844288924;
assign addr[60080]= 1669389513;
assign addr[60081]= 1460659832;
assign addr[60082]= 1222329801;
assign addr[60083]= 959229189;
assign addr[60084]= 676689746;
assign addr[60085]= 380437148;
assign addr[60086]= 76474970;
assign addr[60087]= -229036977;
assign addr[60088]= -529907477;
assign addr[60089]= -820039373;
assign addr[60090]= -1093553126;
assign addr[60091]= -1344905966;
assign addr[60092]= -1569004214;
assign addr[60093]= -1761306505;
assign addr[60094]= -1917915825;
assign addr[60095]= -2035658475;
assign addr[60096]= -2112148396;
assign addr[60097]= -2145835515;
assign addr[60098]= -2136037160;
assign addr[60099]= -2082951896;
assign addr[60100]= -1987655498;
assign addr[60101]= -1852079154;
assign addr[60102]= -1678970324;
assign addr[60103]= -1471837070;
assign addr[60104]= -1234876957;
assign addr[60105]= -972891995;
assign addr[60106]= -691191324;
assign addr[60107]= -395483624;
assign addr[60108]= -91761426;
assign addr[60109]= 213820322;
assign addr[60110]= 515068990;
assign addr[60111]= 805879757;
assign addr[60112]= 1080359326;
assign addr[60113]= 1332945355;
assign addr[60114]= 1558519173;
assign addr[60115]= 1752509516;
assign addr[60116]= 1910985158;
assign addr[60117]= 2030734582;
assign addr[60118]= 2109331059;
assign addr[60119]= 2145181827;
assign addr[60120]= 2137560369;
assign addr[60121]= 2086621133;
assign addr[60122]= 1993396407;
assign addr[60123]= 1859775393;
assign addr[60124]= 1688465931;
assign addr[60125]= 1482939614;
assign addr[60126]= 1247361445;
assign addr[60127]= 986505429;
assign addr[60128]= 705657826;
assign addr[60129]= 410510029;
assign addr[60130]= 107043224;
assign addr[60131]= -198592817;
assign addr[60132]= -500204365;
assign addr[60133]= -791679244;
assign addr[60134]= -1067110699;
assign addr[60135]= -1320917099;
assign addr[60136]= -1547955041;
assign addr[60137]= -1743623590;
assign addr[60138]= -1903957513;
assign addr[60139]= -2025707632;
assign addr[60140]= -2106406677;
assign addr[60141]= -2144419275;
assign addr[60142]= -2138975100;
assign addr[60143]= -2090184478;
assign addr[60144]= -1999036154;
assign addr[60145]= -1867377253;
assign addr[60146]= -1697875851;
assign addr[60147]= -1493966902;
assign addr[60148]= -1259782632;
assign addr[60149]= -1000068799;
assign addr[60150]= -720088517;
assign addr[60151]= -425515602;
assign addr[60152]= -122319591;
assign addr[60153]= 183355234;
assign addr[60154]= 485314355;
assign addr[60155]= 777438554;
assign addr[60156]= 1053807919;
assign addr[60157]= 1308821808;
assign addr[60158]= 1537312353;
assign addr[60159]= 1734649179;
assign addr[60160]= 1896833245;
assign addr[60161]= 2020577882;
assign addr[60162]= 2103375398;
assign addr[60163]= 2143547897;
assign addr[60164]= 2140281282;
assign addr[60165]= 2093641749;
assign addr[60166]= 2004574453;
assign addr[60167]= 1874884346;
assign addr[60168]= 1707199606;
assign addr[60169]= 1504918373;
assign addr[60170]= 1272139887;
assign addr[60171]= 1013581418;
assign addr[60172]= 734482665;
assign addr[60173]= 440499581;
assign addr[60174]= 137589750;
assign addr[60175]= -168108346;
assign addr[60176]= -470399716;
assign addr[60177]= -763158411;
assign addr[60178]= -1040451659;
assign addr[60179]= -1296660098;
assign addr[60180]= -1526591649;
assign addr[60181]= -1725586737;
assign addr[60182]= -1889612716;
assign addr[60183]= -2015345591;
assign addr[60184]= -2100237377;
assign addr[60185]= -2142567738;
assign addr[60186]= -2141478848;
assign addr[60187]= -2096992772;
assign addr[60188]= -2010011024;
assign addr[60189]= -1882296293;
assign addr[60190]= -1716436725;
assign addr[60191]= -1515793473;
assign addr[60192]= -1284432584;
assign addr[60193]= -1027042599;
assign addr[60194]= -748839539;
assign addr[60195]= -455461206;
assign addr[60196]= -152852926;
assign addr[60197]= 152852926;
assign addr[60198]= 455461206;
assign addr[60199]= 748839539;
assign addr[60200]= 1027042599;
assign addr[60201]= 1284432584;
assign addr[60202]= 1515793473;
assign addr[60203]= 1716436725;
assign addr[60204]= 1882296293;
assign addr[60205]= 2010011024;
assign addr[60206]= 2096992772;
assign addr[60207]= 2141478848;
assign addr[60208]= 2142567738;
assign addr[60209]= 2100237377;
assign addr[60210]= 2015345591;
assign addr[60211]= 1889612716;
assign addr[60212]= 1725586737;
assign addr[60213]= 1526591649;
assign addr[60214]= 1296660098;
assign addr[60215]= 1040451659;
assign addr[60216]= 763158411;
assign addr[60217]= 470399716;
assign addr[60218]= 168108346;
assign addr[60219]= -137589750;
assign addr[60220]= -440499581;
assign addr[60221]= -734482665;
assign addr[60222]= -1013581418;
assign addr[60223]= -1272139887;
assign addr[60224]= -1504918373;
assign addr[60225]= -1707199606;
assign addr[60226]= -1874884346;
assign addr[60227]= -2004574453;
assign addr[60228]= -2093641749;
assign addr[60229]= -2140281282;
assign addr[60230]= -2143547897;
assign addr[60231]= -2103375398;
assign addr[60232]= -2020577882;
assign addr[60233]= -1896833245;
assign addr[60234]= -1734649179;
assign addr[60235]= -1537312353;
assign addr[60236]= -1308821808;
assign addr[60237]= -1053807919;
assign addr[60238]= -777438554;
assign addr[60239]= -485314355;
assign addr[60240]= -183355234;
assign addr[60241]= 122319591;
assign addr[60242]= 425515602;
assign addr[60243]= 720088517;
assign addr[60244]= 1000068799;
assign addr[60245]= 1259782632;
assign addr[60246]= 1493966902;
assign addr[60247]= 1697875851;
assign addr[60248]= 1867377253;
assign addr[60249]= 1999036154;
assign addr[60250]= 2090184478;
assign addr[60251]= 2138975100;
assign addr[60252]= 2144419275;
assign addr[60253]= 2106406677;
assign addr[60254]= 2025707632;
assign addr[60255]= 1903957513;
assign addr[60256]= 1743623590;
assign addr[60257]= 1547955041;
assign addr[60258]= 1320917099;
assign addr[60259]= 1067110699;
assign addr[60260]= 791679244;
assign addr[60261]= 500204365;
assign addr[60262]= 198592817;
assign addr[60263]= -107043224;
assign addr[60264]= -410510029;
assign addr[60265]= -705657826;
assign addr[60266]= -986505429;
assign addr[60267]= -1247361445;
assign addr[60268]= -1482939614;
assign addr[60269]= -1688465931;
assign addr[60270]= -1859775393;
assign addr[60271]= -1993396407;
assign addr[60272]= -2086621133;
assign addr[60273]= -2137560369;
assign addr[60274]= -2145181827;
assign addr[60275]= -2109331059;
assign addr[60276]= -2030734582;
assign addr[60277]= -1910985158;
assign addr[60278]= -1752509516;
assign addr[60279]= -1558519173;
assign addr[60280]= -1332945355;
assign addr[60281]= -1080359326;
assign addr[60282]= -805879757;
assign addr[60283]= -515068990;
assign addr[60284]= -213820322;
assign addr[60285]= 91761426;
assign addr[60286]= 395483624;
assign addr[60287]= 691191324;
assign addr[60288]= 972891995;
assign addr[60289]= 1234876957;
assign addr[60290]= 1471837070;
assign addr[60291]= 1678970324;
assign addr[60292]= 1852079154;
assign addr[60293]= 1987655498;
assign addr[60294]= 2082951896;
assign addr[60295]= 2136037160;
assign addr[60296]= 2145835515;
assign addr[60297]= 2112148396;
assign addr[60298]= 2035658475;
assign addr[60299]= 1917915825;
assign addr[60300]= 1761306505;
assign addr[60301]= 1569004214;
assign addr[60302]= 1344905966;
assign addr[60303]= 1093553126;
assign addr[60304]= 820039373;
assign addr[60305]= 529907477;
assign addr[60306]= 229036977;
assign addr[60307]= -76474970;
assign addr[60308]= -380437148;
assign addr[60309]= -676689746;
assign addr[60310]= -959229189;
assign addr[60311]= -1222329801;
assign addr[60312]= -1460659832;
assign addr[60313]= -1669389513;
assign addr[60314]= -1844288924;
assign addr[60315]= -1981813720;
assign addr[60316]= -2079176953;
assign addr[60317]= -2134405552;
assign addr[60318]= -2146380306;
assign addr[60319]= -2114858546;
assign addr[60320]= -2040479063;
assign addr[60321]= -1924749160;
assign addr[60322]= -1770014111;
assign addr[60323]= -1579409630;
assign addr[60324]= -1356798326;
assign addr[60325]= -1106691431;
assign addr[60326]= -834157373;
assign addr[60327]= -544719071;
assign addr[60328]= -244242007;
assign addr[60329]= 61184634;
assign addr[60330]= 365371365;
assign addr[60331]= 662153826;
assign addr[60332]= 945517704;
assign addr[60333]= 1209720613;
assign addr[60334]= 1449408469;
assign addr[60335]= 1659723983;
assign addr[60336]= 1836405100;
assign addr[60337]= 1975871368;
assign addr[60338]= 2075296495;
assign addr[60339]= 2132665626;
assign addr[60340]= 2146816171;
assign addr[60341]= 2117461370;
assign addr[60342]= 2045196100;
assign addr[60343]= 1931484818;
assign addr[60344]= 1778631892;
assign addr[60345]= 1589734894;
assign addr[60346]= 1368621831;
assign addr[60347]= 1119773573;
assign addr[60348]= 848233042;
assign addr[60349]= 559503022;
assign addr[60350]= 259434643;
assign addr[60351]= -45891193;
assign addr[60352]= -350287041;
assign addr[60353]= -647584304;
assign addr[60354]= -931758235;
assign addr[60355]= -1197050035;
assign addr[60356]= -1438083551;
assign addr[60357]= -1649974225;
assign addr[60358]= -1828428082;
assign addr[60359]= -1969828744;
assign addr[60360]= -2071310720;
assign addr[60361]= -2130817471;
assign addr[60362]= -2147143090;
assign addr[60363]= -2119956737;
assign addr[60364]= -2049809346;
assign addr[60365]= -1938122457;
assign addr[60366]= -1787159411;
assign addr[60367]= -1599979481;
assign addr[60368]= -1380375881;
assign addr[60369]= -1132798888;
assign addr[60370]= -862265664;
assign addr[60371]= -574258580;
assign addr[60372]= -274614114;
assign addr[60373]= 30595422;
assign addr[60374]= 335184940;
assign addr[60375]= 632981917;
assign addr[60376]= 917951481;
assign addr[60377]= 1184318708;
assign addr[60378]= 1426685652;
assign addr[60379]= 1640140734;
assign addr[60380]= 1820358275;
assign addr[60381]= 1963686155;
assign addr[60382]= 2067219829;
assign addr[60383]= 2128861181;
assign addr[60384]= 2147361045;
assign addr[60385]= 2122344521;
assign addr[60386]= 2054318569;
assign addr[60387]= 1944661739;
assign addr[60388]= 1795596234;
assign addr[60389]= 1610142873;
assign addr[60390]= 1392059879;
assign addr[60391]= 1145766716;
assign addr[60392]= 876254528;
assign addr[60393]= 588984994;
assign addr[60394]= 289779648;
assign addr[60395]= -15298099;
assign addr[60396]= -320065829;
assign addr[60397]= -618347408;
assign addr[60398]= -904098143;
assign addr[60399]= -1171527280;
assign addr[60400]= -1415215352;
assign addr[60401]= -1630224009;
assign addr[60402]= -1812196087;
assign addr[60403]= -1957443913;
assign addr[60404]= -2063024031;
assign addr[60405]= -2126796855;
assign addr[60406]= -2147470025;
assign addr[60407]= -2124624598;
assign addr[60408]= -2058723538;
assign addr[60409]= -1951102334;
assign addr[60410]= -1803941934;
assign addr[60411]= -1620224553;
assign addr[60412]= -1403673233;
assign addr[60413]= -1158676398;
assign addr[60414]= -890198924;
assign addr[60415]= -603681519;
assign addr[60416]= -304930476;
assign addr[60417]= 0;
assign addr[60418]= 304930476;
assign addr[60419]= 603681519;
assign addr[60420]= 890198924;
assign addr[60421]= 1158676398;
assign addr[60422]= 1403673233;
assign addr[60423]= 1620224553;
assign addr[60424]= 1803941934;
assign addr[60425]= 1951102334;
assign addr[60426]= 2058723538;
assign addr[60427]= 2124624598;
assign addr[60428]= 2147470025;
assign addr[60429]= 2126796855;
assign addr[60430]= 2063024031;
assign addr[60431]= 1957443913;
assign addr[60432]= 1812196087;
assign addr[60433]= 1630224009;
assign addr[60434]= 1415215352;
assign addr[60435]= 1171527280;
assign addr[60436]= 904098143;
assign addr[60437]= 618347408;
assign addr[60438]= 320065829;
assign addr[60439]= 15298099;
assign addr[60440]= -289779648;
assign addr[60441]= -588984994;
assign addr[60442]= -876254528;
assign addr[60443]= -1145766716;
assign addr[60444]= -1392059879;
assign addr[60445]= -1610142873;
assign addr[60446]= -1795596234;
assign addr[60447]= -1944661739;
assign addr[60448]= -2054318569;
assign addr[60449]= -2122344521;
assign addr[60450]= -2147361045;
assign addr[60451]= -2128861181;
assign addr[60452]= -2067219829;
assign addr[60453]= -1963686155;
assign addr[60454]= -1820358275;
assign addr[60455]= -1640140734;
assign addr[60456]= -1426685652;
assign addr[60457]= -1184318708;
assign addr[60458]= -917951481;
assign addr[60459]= -632981917;
assign addr[60460]= -335184940;
assign addr[60461]= -30595422;
assign addr[60462]= 274614114;
assign addr[60463]= 574258580;
assign addr[60464]= 862265664;
assign addr[60465]= 1132798888;
assign addr[60466]= 1380375881;
assign addr[60467]= 1599979481;
assign addr[60468]= 1787159411;
assign addr[60469]= 1938122457;
assign addr[60470]= 2049809346;
assign addr[60471]= 2119956737;
assign addr[60472]= 2147143090;
assign addr[60473]= 2130817471;
assign addr[60474]= 2071310720;
assign addr[60475]= 1969828744;
assign addr[60476]= 1828428082;
assign addr[60477]= 1649974225;
assign addr[60478]= 1438083551;
assign addr[60479]= 1197050035;
assign addr[60480]= 931758235;
assign addr[60481]= 647584304;
assign addr[60482]= 350287041;
assign addr[60483]= 45891193;
assign addr[60484]= -259434643;
assign addr[60485]= -559503022;
assign addr[60486]= -848233042;
assign addr[60487]= -1119773573;
assign addr[60488]= -1368621831;
assign addr[60489]= -1589734894;
assign addr[60490]= -1778631892;
assign addr[60491]= -1931484818;
assign addr[60492]= -2045196100;
assign addr[60493]= -2117461370;
assign addr[60494]= -2146816171;
assign addr[60495]= -2132665626;
assign addr[60496]= -2075296495;
assign addr[60497]= -1975871368;
assign addr[60498]= -1836405100;
assign addr[60499]= -1659723983;
assign addr[60500]= -1449408469;
assign addr[60501]= -1209720613;
assign addr[60502]= -945517704;
assign addr[60503]= -662153826;
assign addr[60504]= -365371365;
assign addr[60505]= -61184634;
assign addr[60506]= 244242007;
assign addr[60507]= 544719071;
assign addr[60508]= 834157373;
assign addr[60509]= 1106691431;
assign addr[60510]= 1356798326;
assign addr[60511]= 1579409630;
assign addr[60512]= 1770014111;
assign addr[60513]= 1924749160;
assign addr[60514]= 2040479063;
assign addr[60515]= 2114858546;
assign addr[60516]= 2146380306;
assign addr[60517]= 2134405552;
assign addr[60518]= 2079176953;
assign addr[60519]= 1981813720;
assign addr[60520]= 1844288924;
assign addr[60521]= 1669389513;
assign addr[60522]= 1460659832;
assign addr[60523]= 1222329801;
assign addr[60524]= 959229189;
assign addr[60525]= 676689746;
assign addr[60526]= 380437148;
assign addr[60527]= 76474970;
assign addr[60528]= -229036977;
assign addr[60529]= -529907477;
assign addr[60530]= -820039373;
assign addr[60531]= -1093553126;
assign addr[60532]= -1344905966;
assign addr[60533]= -1569004214;
assign addr[60534]= -1761306505;
assign addr[60535]= -1917915825;
assign addr[60536]= -2035658475;
assign addr[60537]= -2112148396;
assign addr[60538]= -2145835515;
assign addr[60539]= -2136037160;
assign addr[60540]= -2082951896;
assign addr[60541]= -1987655498;
assign addr[60542]= -1852079154;
assign addr[60543]= -1678970324;
assign addr[60544]= -1471837070;
assign addr[60545]= -1234876957;
assign addr[60546]= -972891995;
assign addr[60547]= -691191324;
assign addr[60548]= -395483624;
assign addr[60549]= -91761426;
assign addr[60550]= 213820322;
assign addr[60551]= 515068990;
assign addr[60552]= 805879757;
assign addr[60553]= 1080359326;
assign addr[60554]= 1332945355;
assign addr[60555]= 1558519173;
assign addr[60556]= 1752509516;
assign addr[60557]= 1910985158;
assign addr[60558]= 2030734582;
assign addr[60559]= 2109331059;
assign addr[60560]= 2145181827;
assign addr[60561]= 2137560369;
assign addr[60562]= 2086621133;
assign addr[60563]= 1993396407;
assign addr[60564]= 1859775393;
assign addr[60565]= 1688465931;
assign addr[60566]= 1482939614;
assign addr[60567]= 1247361445;
assign addr[60568]= 986505429;
assign addr[60569]= 705657826;
assign addr[60570]= 410510029;
assign addr[60571]= 107043224;
assign addr[60572]= -198592817;
assign addr[60573]= -500204365;
assign addr[60574]= -791679244;
assign addr[60575]= -1067110699;
assign addr[60576]= -1320917099;
assign addr[60577]= -1547955041;
assign addr[60578]= -1743623590;
assign addr[60579]= -1903957513;
assign addr[60580]= -2025707632;
assign addr[60581]= -2106406677;
assign addr[60582]= -2144419275;
assign addr[60583]= -2138975100;
assign addr[60584]= -2090184478;
assign addr[60585]= -1999036154;
assign addr[60586]= -1867377253;
assign addr[60587]= -1697875851;
assign addr[60588]= -1493966902;
assign addr[60589]= -1259782632;
assign addr[60590]= -1000068799;
assign addr[60591]= -720088517;
assign addr[60592]= -425515602;
assign addr[60593]= -122319591;
assign addr[60594]= 183355234;
assign addr[60595]= 485314355;
assign addr[60596]= 777438554;
assign addr[60597]= 1053807919;
assign addr[60598]= 1308821808;
assign addr[60599]= 1537312353;
assign addr[60600]= 1734649179;
assign addr[60601]= 1896833245;
assign addr[60602]= 2020577882;
assign addr[60603]= 2103375398;
assign addr[60604]= 2143547897;
assign addr[60605]= 2140281282;
assign addr[60606]= 2093641749;
assign addr[60607]= 2004574453;
assign addr[60608]= 1874884346;
assign addr[60609]= 1707199606;
assign addr[60610]= 1504918373;
assign addr[60611]= 1272139887;
assign addr[60612]= 1013581418;
assign addr[60613]= 734482665;
assign addr[60614]= 440499581;
assign addr[60615]= 137589750;
assign addr[60616]= -168108346;
assign addr[60617]= -470399716;
assign addr[60618]= -763158411;
assign addr[60619]= -1040451659;
assign addr[60620]= -1296660098;
assign addr[60621]= -1526591649;
assign addr[60622]= -1725586737;
assign addr[60623]= -1889612716;
assign addr[60624]= -2015345591;
assign addr[60625]= -2100237377;
assign addr[60626]= -2142567738;
assign addr[60627]= -2141478848;
assign addr[60628]= -2096992772;
assign addr[60629]= -2010011024;
assign addr[60630]= -1882296293;
assign addr[60631]= -1716436725;
assign addr[60632]= -1515793473;
assign addr[60633]= -1284432584;
assign addr[60634]= -1027042599;
assign addr[60635]= -748839539;
assign addr[60636]= -455461206;
assign addr[60637]= -152852926;
assign addr[60638]= 152852926;
assign addr[60639]= 455461206;
assign addr[60640]= 748839539;
assign addr[60641]= 1027042599;
assign addr[60642]= 1284432584;
assign addr[60643]= 1515793473;
assign addr[60644]= 1716436725;
assign addr[60645]= 1882296293;
assign addr[60646]= 2010011024;
assign addr[60647]= 2096992772;
assign addr[60648]= 2141478848;
assign addr[60649]= 2142567738;
assign addr[60650]= 2100237377;
assign addr[60651]= 2015345591;
assign addr[60652]= 1889612716;
assign addr[60653]= 1725586737;
assign addr[60654]= 1526591649;
assign addr[60655]= 1296660098;
assign addr[60656]= 1040451659;
assign addr[60657]= 763158411;
assign addr[60658]= 470399716;
assign addr[60659]= 168108346;
assign addr[60660]= -137589750;
assign addr[60661]= -440499581;
assign addr[60662]= -734482665;
assign addr[60663]= -1013581418;
assign addr[60664]= -1272139887;
assign addr[60665]= -1504918373;
assign addr[60666]= -1707199606;
assign addr[60667]= -1874884346;
assign addr[60668]= -2004574453;
assign addr[60669]= -2093641749;
assign addr[60670]= -2140281282;
assign addr[60671]= -2143547897;
assign addr[60672]= -2103375398;
assign addr[60673]= -2020577882;
assign addr[60674]= -1896833245;
assign addr[60675]= -1734649179;
assign addr[60676]= -1537312353;
assign addr[60677]= -1308821808;
assign addr[60678]= -1053807919;
assign addr[60679]= -777438554;
assign addr[60680]= -485314355;
assign addr[60681]= -183355234;
assign addr[60682]= 122319591;
assign addr[60683]= 425515602;
assign addr[60684]= 720088517;
assign addr[60685]= 1000068799;
assign addr[60686]= 1259782632;
assign addr[60687]= 1493966902;
assign addr[60688]= 1697875851;
assign addr[60689]= 1867377253;
assign addr[60690]= 1999036154;
assign addr[60691]= 2090184478;
assign addr[60692]= 2138975100;
assign addr[60693]= 2144419275;
assign addr[60694]= 2106406677;
assign addr[60695]= 2025707632;
assign addr[60696]= 1903957513;
assign addr[60697]= 1743623590;
assign addr[60698]= 1547955041;
assign addr[60699]= 1320917099;
assign addr[60700]= 1067110699;
assign addr[60701]= 791679244;
assign addr[60702]= 500204365;
assign addr[60703]= 198592817;
assign addr[60704]= -107043224;
assign addr[60705]= -410510029;
assign addr[60706]= -705657826;
assign addr[60707]= -986505429;
assign addr[60708]= -1247361445;
assign addr[60709]= -1482939614;
assign addr[60710]= -1688465931;
assign addr[60711]= -1859775393;
assign addr[60712]= -1993396407;
assign addr[60713]= -2086621133;
assign addr[60714]= -2137560369;
assign addr[60715]= -2145181827;
assign addr[60716]= -2109331059;
assign addr[60717]= -2030734582;
assign addr[60718]= -1910985158;
assign addr[60719]= -1752509516;
assign addr[60720]= -1558519173;
assign addr[60721]= -1332945355;
assign addr[60722]= -1080359326;
assign addr[60723]= -805879757;
assign addr[60724]= -515068990;
assign addr[60725]= -213820322;
assign addr[60726]= 91761426;
assign addr[60727]= 395483624;
assign addr[60728]= 691191324;
assign addr[60729]= 972891995;
assign addr[60730]= 1234876957;
assign addr[60731]= 1471837070;
assign addr[60732]= 1678970324;
assign addr[60733]= 1852079154;
assign addr[60734]= 1987655498;
assign addr[60735]= 2082951896;
assign addr[60736]= 2136037160;
assign addr[60737]= 2145835515;
assign addr[60738]= 2112148396;
assign addr[60739]= 2035658475;
assign addr[60740]= 1917915825;
assign addr[60741]= 1761306505;
assign addr[60742]= 1569004214;
assign addr[60743]= 1344905966;
assign addr[60744]= 1093553126;
assign addr[60745]= 820039373;
assign addr[60746]= 529907477;
assign addr[60747]= 229036977;
assign addr[60748]= -76474970;
assign addr[60749]= -380437148;
assign addr[60750]= -676689746;
assign addr[60751]= -959229189;
assign addr[60752]= -1222329801;
assign addr[60753]= -1460659832;
assign addr[60754]= -1669389513;
assign addr[60755]= -1844288924;
assign addr[60756]= -1981813720;
assign addr[60757]= -2079176953;
assign addr[60758]= -2134405552;
assign addr[60759]= -2146380306;
assign addr[60760]= -2114858546;
assign addr[60761]= -2040479063;
assign addr[60762]= -1924749160;
assign addr[60763]= -1770014111;
assign addr[60764]= -1579409630;
assign addr[60765]= -1356798326;
assign addr[60766]= -1106691431;
assign addr[60767]= -834157373;
assign addr[60768]= -544719071;
assign addr[60769]= -244242007;
assign addr[60770]= 61184634;
assign addr[60771]= 365371365;
assign addr[60772]= 662153826;
assign addr[60773]= 945517704;
assign addr[60774]= 1209720613;
assign addr[60775]= 1449408469;
assign addr[60776]= 1659723983;
assign addr[60777]= 1836405100;
assign addr[60778]= 1975871368;
assign addr[60779]= 2075296495;
assign addr[60780]= 2132665626;
assign addr[60781]= 2146816171;
assign addr[60782]= 2117461370;
assign addr[60783]= 2045196100;
assign addr[60784]= 1931484818;
assign addr[60785]= 1778631892;
assign addr[60786]= 1589734894;
assign addr[60787]= 1368621831;
assign addr[60788]= 1119773573;
assign addr[60789]= 848233042;
assign addr[60790]= 559503022;
assign addr[60791]= 259434643;
assign addr[60792]= -45891193;
assign addr[60793]= -350287041;
assign addr[60794]= -647584304;
assign addr[60795]= -931758235;
assign addr[60796]= -1197050035;
assign addr[60797]= -1438083551;
assign addr[60798]= -1649974225;
assign addr[60799]= -1828428082;
assign addr[60800]= -1969828744;
assign addr[60801]= -2071310720;
assign addr[60802]= -2130817471;
assign addr[60803]= -2147143090;
assign addr[60804]= -2119956737;
assign addr[60805]= -2049809346;
assign addr[60806]= -1938122457;
assign addr[60807]= -1787159411;
assign addr[60808]= -1599979481;
assign addr[60809]= -1380375881;
assign addr[60810]= -1132798888;
assign addr[60811]= -862265664;
assign addr[60812]= -574258580;
assign addr[60813]= -274614114;
assign addr[60814]= 30595422;
assign addr[60815]= 335184940;
assign addr[60816]= 632981917;
assign addr[60817]= 917951481;
assign addr[60818]= 1184318708;
assign addr[60819]= 1426685652;
assign addr[60820]= 1640140734;
assign addr[60821]= 1820358275;
assign addr[60822]= 1963686155;
assign addr[60823]= 2067219829;
assign addr[60824]= 2128861181;
assign addr[60825]= 2147361045;
assign addr[60826]= 2122344521;
assign addr[60827]= 2054318569;
assign addr[60828]= 1944661739;
assign addr[60829]= 1795596234;
assign addr[60830]= 1610142873;
assign addr[60831]= 1392059879;
assign addr[60832]= 1145766716;
assign addr[60833]= 876254528;
assign addr[60834]= 588984994;
assign addr[60835]= 289779648;
assign addr[60836]= -15298099;
assign addr[60837]= -320065829;
assign addr[60838]= -618347408;
assign addr[60839]= -904098143;
assign addr[60840]= -1171527280;
assign addr[60841]= -1415215352;
assign addr[60842]= -1630224009;
assign addr[60843]= -1812196087;
assign addr[60844]= -1957443913;
assign addr[60845]= -2063024031;
assign addr[60846]= -2126796855;
assign addr[60847]= -2147470025;
assign addr[60848]= -2124624598;
assign addr[60849]= -2058723538;
assign addr[60850]= -1951102334;
assign addr[60851]= -1803941934;
assign addr[60852]= -1620224553;
assign addr[60853]= -1403673233;
assign addr[60854]= -1158676398;
assign addr[60855]= -890198924;
assign addr[60856]= -603681519;
assign addr[60857]= -304930476;
assign addr[60858]= 0;
assign addr[60859]= 304930476;
assign addr[60860]= 603681519;
assign addr[60861]= 890198924;
assign addr[60862]= 1158676398;
assign addr[60863]= 1403673233;
assign addr[60864]= 1620224553;
assign addr[60865]= 1803941934;
assign addr[60866]= 1951102334;
assign addr[60867]= 2058723538;
assign addr[60868]= 2124624598;
assign addr[60869]= 2147470025;
assign addr[60870]= 2126796855;
assign addr[60871]= 2063024031;
assign addr[60872]= 1957443913;
assign addr[60873]= 1812196087;
assign addr[60874]= 1630224009;
assign addr[60875]= 1415215352;
assign addr[60876]= 1171527280;
assign addr[60877]= 904098143;
assign addr[60878]= 618347408;
assign addr[60879]= 320065829;
assign addr[60880]= 15298099;
assign addr[60881]= -289779648;
assign addr[60882]= -588984994;
assign addr[60883]= -876254528;
assign addr[60884]= -1145766716;
assign addr[60885]= -1392059879;
assign addr[60886]= -1610142873;
assign addr[60887]= -1795596234;
assign addr[60888]= -1944661739;
assign addr[60889]= -2054318569;
assign addr[60890]= -2122344521;
assign addr[60891]= -2147361045;
assign addr[60892]= -2128861181;
assign addr[60893]= -2067219829;
assign addr[60894]= -1963686155;
assign addr[60895]= -1820358275;
assign addr[60896]= -1640140734;
assign addr[60897]= -1426685652;
assign addr[60898]= -1184318708;
assign addr[60899]= -917951481;
assign addr[60900]= -632981917;
assign addr[60901]= -335184940;
assign addr[60902]= -30595422;
assign addr[60903]= 274614114;
assign addr[60904]= 574258580;
assign addr[60905]= 862265664;
assign addr[60906]= 1132798888;
assign addr[60907]= 1380375881;
assign addr[60908]= 1599979481;
assign addr[60909]= 1787159411;
assign addr[60910]= 1938122457;
assign addr[60911]= 2049809346;
assign addr[60912]= 2119956737;
assign addr[60913]= 2147143090;
assign addr[60914]= 2130817471;
assign addr[60915]= 2071310720;
assign addr[60916]= 1969828744;
assign addr[60917]= 1828428082;
assign addr[60918]= 1649974225;
assign addr[60919]= 1438083551;
assign addr[60920]= 1197050035;
assign addr[60921]= 931758235;
assign addr[60922]= 647584304;
assign addr[60923]= 350287041;
assign addr[60924]= 45891193;
assign addr[60925]= -259434643;
assign addr[60926]= -559503022;
assign addr[60927]= -848233042;
assign addr[60928]= -1119773573;
assign addr[60929]= -1368621831;
assign addr[60930]= -1589734894;
assign addr[60931]= -1778631892;
assign addr[60932]= -1931484818;
assign addr[60933]= -2045196100;
assign addr[60934]= -2117461370;
assign addr[60935]= -2146816171;
assign addr[60936]= -2132665626;
assign addr[60937]= -2075296495;
assign addr[60938]= -1975871368;
assign addr[60939]= -1836405100;
assign addr[60940]= -1659723983;
assign addr[60941]= -1449408469;
assign addr[60942]= -1209720613;
assign addr[60943]= -945517704;
assign addr[60944]= -662153826;
assign addr[60945]= -365371365;
assign addr[60946]= -61184634;
assign addr[60947]= 244242007;
assign addr[60948]= 544719071;
assign addr[60949]= 834157373;
assign addr[60950]= 1106691431;
assign addr[60951]= 1356798326;
assign addr[60952]= 1579409630;
assign addr[60953]= 1770014111;
assign addr[60954]= 1924749160;
assign addr[60955]= 2040479063;
assign addr[60956]= 2114858546;
assign addr[60957]= 2146380306;
assign addr[60958]= 2134405552;
assign addr[60959]= 2079176953;
assign addr[60960]= 1981813720;
assign addr[60961]= 1844288924;
assign addr[60962]= 1669389513;
assign addr[60963]= 1460659832;
assign addr[60964]= 1222329801;
assign addr[60965]= 959229189;
assign addr[60966]= 676689746;
assign addr[60967]= 380437148;
assign addr[60968]= 76474970;
assign addr[60969]= -229036977;
assign addr[60970]= -529907477;
assign addr[60971]= -820039373;
assign addr[60972]= -1093553126;
assign addr[60973]= -1344905966;
assign addr[60974]= -1569004214;
assign addr[60975]= -1761306505;
assign addr[60976]= -1917915825;
assign addr[60977]= -2035658475;
assign addr[60978]= -2112148396;
assign addr[60979]= -2145835515;
assign addr[60980]= -2136037160;
assign addr[60981]= -2082951896;
assign addr[60982]= -1987655498;
assign addr[60983]= -1852079154;
assign addr[60984]= -1678970324;
assign addr[60985]= -1471837070;
assign addr[60986]= -1234876957;
assign addr[60987]= -972891995;
assign addr[60988]= -691191324;
assign addr[60989]= -395483624;
assign addr[60990]= -91761426;
assign addr[60991]= 213820322;
assign addr[60992]= 515068990;
assign addr[60993]= 805879757;
assign addr[60994]= 1080359326;
assign addr[60995]= 1332945355;
assign addr[60996]= 1558519173;
assign addr[60997]= 1752509516;
assign addr[60998]= 1910985158;
assign addr[60999]= 2030734582;
assign addr[61000]= 2109331059;
assign addr[61001]= 2145181827;
assign addr[61002]= 2137560369;
assign addr[61003]= 2086621133;
assign addr[61004]= 1993396407;
assign addr[61005]= 1859775393;
assign addr[61006]= 1688465931;
assign addr[61007]= 1482939614;
assign addr[61008]= 1247361445;
assign addr[61009]= 986505429;
assign addr[61010]= 705657826;
assign addr[61011]= 410510029;
assign addr[61012]= 107043224;
assign addr[61013]= -198592817;
assign addr[61014]= -500204365;
assign addr[61015]= -791679244;
assign addr[61016]= -1067110699;
assign addr[61017]= -1320917099;
assign addr[61018]= -1547955041;
assign addr[61019]= -1743623590;
assign addr[61020]= -1903957513;
assign addr[61021]= -2025707632;
assign addr[61022]= -2106406677;
assign addr[61023]= -2144419275;
assign addr[61024]= -2138975100;
assign addr[61025]= -2090184478;
assign addr[61026]= -1999036154;
assign addr[61027]= -1867377253;
assign addr[61028]= -1697875851;
assign addr[61029]= -1493966902;
assign addr[61030]= -1259782632;
assign addr[61031]= -1000068799;
assign addr[61032]= -720088517;
assign addr[61033]= -425515602;
assign addr[61034]= -122319591;
assign addr[61035]= 183355234;
assign addr[61036]= 485314355;
assign addr[61037]= 777438554;
assign addr[61038]= 1053807919;
assign addr[61039]= 1308821808;
assign addr[61040]= 1537312353;
assign addr[61041]= 1734649179;
assign addr[61042]= 1896833245;
assign addr[61043]= 2020577882;
assign addr[61044]= 2103375398;
assign addr[61045]= 2143547897;
assign addr[61046]= 2140281282;
assign addr[61047]= 2093641749;
assign addr[61048]= 2004574453;
assign addr[61049]= 1874884346;
assign addr[61050]= 1707199606;
assign addr[61051]= 1504918373;
assign addr[61052]= 1272139887;
assign addr[61053]= 1013581418;
assign addr[61054]= 734482665;
assign addr[61055]= 440499581;
assign addr[61056]= 137589750;
assign addr[61057]= -168108346;
assign addr[61058]= -470399716;
assign addr[61059]= -763158411;
assign addr[61060]= -1040451659;
assign addr[61061]= -1296660098;
assign addr[61062]= -1526591649;
assign addr[61063]= -1725586737;
assign addr[61064]= -1889612716;
assign addr[61065]= -2015345591;
assign addr[61066]= -2100237377;
assign addr[61067]= -2142567738;
assign addr[61068]= -2141478848;
assign addr[61069]= -2096992772;
assign addr[61070]= -2010011024;
assign addr[61071]= -1882296293;
assign addr[61072]= -1716436725;
assign addr[61073]= -1515793473;
assign addr[61074]= -1284432584;
assign addr[61075]= -1027042599;
assign addr[61076]= -748839539;
assign addr[61077]= -455461206;
assign addr[61078]= -152852926;
assign addr[61079]= 152852926;
assign addr[61080]= 455461206;
assign addr[61081]= 748839539;
assign addr[61082]= 1027042599;
assign addr[61083]= 1284432584;
assign addr[61084]= 1515793473;
assign addr[61085]= 1716436725;
assign addr[61086]= 1882296293;
assign addr[61087]= 2010011024;
assign addr[61088]= 2096992772;
assign addr[61089]= 2141478848;
assign addr[61090]= 2142567738;
assign addr[61091]= 2100237377;
assign addr[61092]= 2015345591;
assign addr[61093]= 1889612716;
assign addr[61094]= 1725586737;
assign addr[61095]= 1526591649;
assign addr[61096]= 1296660098;
assign addr[61097]= 1040451659;
assign addr[61098]= 763158411;
assign addr[61099]= 470399716;
assign addr[61100]= 168108346;
assign addr[61101]= -137589750;
assign addr[61102]= -440499581;
assign addr[61103]= -734482665;
assign addr[61104]= -1013581418;
assign addr[61105]= -1272139887;
assign addr[61106]= -1504918373;
assign addr[61107]= -1707199606;
assign addr[61108]= -1874884346;
assign addr[61109]= -2004574453;
assign addr[61110]= -2093641749;
assign addr[61111]= -2140281282;
assign addr[61112]= -2143547897;
assign addr[61113]= -2103375398;
assign addr[61114]= -2020577882;
assign addr[61115]= -1896833245;
assign addr[61116]= -1734649179;
assign addr[61117]= -1537312353;
assign addr[61118]= -1308821808;
assign addr[61119]= -1053807919;
assign addr[61120]= -777438554;
assign addr[61121]= -485314355;
assign addr[61122]= -183355234;
assign addr[61123]= 122319591;
assign addr[61124]= 425515602;
assign addr[61125]= 720088517;
assign addr[61126]= 1000068799;
assign addr[61127]= 1259782632;
assign addr[61128]= 1493966902;
assign addr[61129]= 1697875851;
assign addr[61130]= 1867377253;
assign addr[61131]= 1999036154;
assign addr[61132]= 2090184478;
assign addr[61133]= 2138975100;
assign addr[61134]= 2144419275;
assign addr[61135]= 2106406677;
assign addr[61136]= 2025707632;
assign addr[61137]= 1903957513;
assign addr[61138]= 1743623590;
assign addr[61139]= 1547955041;
assign addr[61140]= 1320917099;
assign addr[61141]= 1067110699;
assign addr[61142]= 791679244;
assign addr[61143]= 500204365;
assign addr[61144]= 198592817;
assign addr[61145]= -107043224;
assign addr[61146]= -410510029;
assign addr[61147]= -705657826;
assign addr[61148]= -986505429;
assign addr[61149]= -1247361445;
assign addr[61150]= -1482939614;
assign addr[61151]= -1688465931;
assign addr[61152]= -1859775393;
assign addr[61153]= -1993396407;
assign addr[61154]= -2086621133;
assign addr[61155]= -2137560369;
assign addr[61156]= -2145181827;
assign addr[61157]= -2109331059;
assign addr[61158]= -2030734582;
assign addr[61159]= -1910985158;
assign addr[61160]= -1752509516;
assign addr[61161]= -1558519173;
assign addr[61162]= -1332945355;
assign addr[61163]= -1080359326;
assign addr[61164]= -805879757;
assign addr[61165]= -515068990;
assign addr[61166]= -213820322;
assign addr[61167]= 91761426;
assign addr[61168]= 395483624;
assign addr[61169]= 691191324;
assign addr[61170]= 972891995;
assign addr[61171]= 1234876957;
assign addr[61172]= 1471837070;
assign addr[61173]= 1678970324;
assign addr[61174]= 1852079154;
assign addr[61175]= 1987655498;
assign addr[61176]= 2082951896;
assign addr[61177]= 2136037160;
assign addr[61178]= 2145835515;
assign addr[61179]= 2112148396;
assign addr[61180]= 2035658475;
assign addr[61181]= 1917915825;
assign addr[61182]= 1761306505;
assign addr[61183]= 1569004214;
assign addr[61184]= 1344905966;
assign addr[61185]= 1093553126;
assign addr[61186]= 820039373;
assign addr[61187]= 529907477;
assign addr[61188]= 229036977;
assign addr[61189]= -76474970;
assign addr[61190]= -380437148;
assign addr[61191]= -676689746;
assign addr[61192]= -959229189;
assign addr[61193]= -1222329801;
assign addr[61194]= -1460659832;
assign addr[61195]= -1669389513;
assign addr[61196]= -1844288924;
assign addr[61197]= -1981813720;
assign addr[61198]= -2079176953;
assign addr[61199]= -2134405552;
assign addr[61200]= -2146380306;
assign addr[61201]= -2114858546;
assign addr[61202]= -2040479063;
assign addr[61203]= -1924749160;
assign addr[61204]= -1770014111;
assign addr[61205]= -1579409630;
assign addr[61206]= -1356798326;
assign addr[61207]= -1106691431;
assign addr[61208]= -834157373;
assign addr[61209]= -544719071;
assign addr[61210]= -244242007;
assign addr[61211]= 61184634;
assign addr[61212]= 365371365;
assign addr[61213]= 662153826;
assign addr[61214]= 945517704;
assign addr[61215]= 1209720613;
assign addr[61216]= 1449408469;
assign addr[61217]= 1659723983;
assign addr[61218]= 1836405100;
assign addr[61219]= 1975871368;
assign addr[61220]= 2075296495;
assign addr[61221]= 2132665626;
assign addr[61222]= 2146816171;
assign addr[61223]= 2117461370;
assign addr[61224]= 2045196100;
assign addr[61225]= 1931484818;
assign addr[61226]= 1778631892;
assign addr[61227]= 1589734894;
assign addr[61228]= 1368621831;
assign addr[61229]= 1119773573;
assign addr[61230]= 848233042;
assign addr[61231]= 559503022;
assign addr[61232]= 259434643;
assign addr[61233]= -45891193;
assign addr[61234]= -350287041;
assign addr[61235]= -647584304;
assign addr[61236]= -931758235;
assign addr[61237]= -1197050035;
assign addr[61238]= -1438083551;
assign addr[61239]= -1649974225;
assign addr[61240]= -1828428082;
assign addr[61241]= -1969828744;
assign addr[61242]= -2071310720;
assign addr[61243]= -2130817471;
assign addr[61244]= -2147143090;
assign addr[61245]= -2119956737;
assign addr[61246]= -2049809346;
assign addr[61247]= -1938122457;
assign addr[61248]= -1787159411;
assign addr[61249]= -1599979481;
assign addr[61250]= -1380375881;
assign addr[61251]= -1132798888;
assign addr[61252]= -862265664;
assign addr[61253]= -574258580;
assign addr[61254]= -274614114;
assign addr[61255]= 30595422;
assign addr[61256]= 335184940;
assign addr[61257]= 632981917;
assign addr[61258]= 917951481;
assign addr[61259]= 1184318708;
assign addr[61260]= 1426685652;
assign addr[61261]= 1640140734;
assign addr[61262]= 1820358275;
assign addr[61263]= 1963686155;
assign addr[61264]= 2067219829;
assign addr[61265]= 2128861181;
assign addr[61266]= 2147361045;
assign addr[61267]= 2122344521;
assign addr[61268]= 2054318569;
assign addr[61269]= 1944661739;
assign addr[61270]= 1795596234;
assign addr[61271]= 1610142873;
assign addr[61272]= 1392059879;
assign addr[61273]= 1145766716;
assign addr[61274]= 876254528;
assign addr[61275]= 588984994;
assign addr[61276]= 289779648;
assign addr[61277]= -15298099;
assign addr[61278]= -320065829;
assign addr[61279]= -618347408;
assign addr[61280]= -904098143;
assign addr[61281]= -1171527280;
assign addr[61282]= -1415215352;
assign addr[61283]= -1630224009;
assign addr[61284]= -1812196087;
assign addr[61285]= -1957443913;
assign addr[61286]= -2063024031;
assign addr[61287]= -2126796855;
assign addr[61288]= -2147470025;
assign addr[61289]= -2124624598;
assign addr[61290]= -2058723538;
assign addr[61291]= -1951102334;
assign addr[61292]= -1803941934;
assign addr[61293]= -1620224553;
assign addr[61294]= -1403673233;
assign addr[61295]= -1158676398;
assign addr[61296]= -890198924;
assign addr[61297]= -603681519;
assign addr[61298]= -304930476;
assign addr[61299]= 0;
assign addr[61300]= 304930476;
assign addr[61301]= 603681519;
assign addr[61302]= 890198924;
assign addr[61303]= 1158676398;
assign addr[61304]= 1403673233;
assign addr[61305]= 1620224553;
assign addr[61306]= 1803941934;
assign addr[61307]= 1951102334;
assign addr[61308]= 2058723538;
assign addr[61309]= 2124624598;
assign addr[61310]= 2147470025;
assign addr[61311]= 2126796855;
assign addr[61312]= 2063024031;
assign addr[61313]= 1957443913;
assign addr[61314]= 1812196087;
assign addr[61315]= 1630224009;
assign addr[61316]= 1415215352;
assign addr[61317]= 1171527280;
assign addr[61318]= 904098143;
assign addr[61319]= 618347408;
assign addr[61320]= 320065829;
assign addr[61321]= 15298099;
assign addr[61322]= -289779648;
assign addr[61323]= -588984994;
assign addr[61324]= -876254528;
assign addr[61325]= -1145766716;
assign addr[61326]= -1392059879;
assign addr[61327]= -1610142873;
assign addr[61328]= -1795596234;
assign addr[61329]= -1944661739;
assign addr[61330]= -2054318569;
assign addr[61331]= -2122344521;
assign addr[61332]= -2147361045;
assign addr[61333]= -2128861181;
assign addr[61334]= -2067219829;
assign addr[61335]= -1963686155;
assign addr[61336]= -1820358275;
assign addr[61337]= -1640140734;
assign addr[61338]= -1426685652;
assign addr[61339]= -1184318708;
assign addr[61340]= -917951481;
assign addr[61341]= -632981917;
assign addr[61342]= -335184940;
assign addr[61343]= -30595422;
assign addr[61344]= 274614114;
assign addr[61345]= 574258580;
assign addr[61346]= 862265664;
assign addr[61347]= 1132798888;
assign addr[61348]= 1380375881;
assign addr[61349]= 1599979481;
assign addr[61350]= 1787159411;
assign addr[61351]= 1938122457;
assign addr[61352]= 2049809346;
assign addr[61353]= 2119956737;
assign addr[61354]= 2147143090;
assign addr[61355]= 2130817471;
assign addr[61356]= 2071310720;
assign addr[61357]= 1969828744;
assign addr[61358]= 1828428082;
assign addr[61359]= 1649974225;
assign addr[61360]= 1438083551;
assign addr[61361]= 1197050035;
assign addr[61362]= 931758235;
assign addr[61363]= 647584304;
assign addr[61364]= 350287041;
assign addr[61365]= 45891193;
assign addr[61366]= -259434643;
assign addr[61367]= -559503022;
assign addr[61368]= -848233042;
assign addr[61369]= -1119773573;
assign addr[61370]= -1368621831;
assign addr[61371]= -1589734894;
assign addr[61372]= -1778631892;
assign addr[61373]= -1931484818;
assign addr[61374]= -2045196100;
assign addr[61375]= -2117461370;
assign addr[61376]= -2146816171;
assign addr[61377]= -2132665626;
assign addr[61378]= -2075296495;
assign addr[61379]= -1975871368;
assign addr[61380]= -1836405100;
assign addr[61381]= -1659723983;
assign addr[61382]= -1449408469;
assign addr[61383]= -1209720613;
assign addr[61384]= -945517704;
assign addr[61385]= -662153826;
assign addr[61386]= -365371365;
assign addr[61387]= -61184634;
assign addr[61388]= 244242007;
assign addr[61389]= 544719071;
assign addr[61390]= 834157373;
assign addr[61391]= 1106691431;
assign addr[61392]= 1356798326;
assign addr[61393]= 1579409630;
assign addr[61394]= 1770014111;
assign addr[61395]= 1924749160;
assign addr[61396]= 2040479063;
assign addr[61397]= 2114858546;
assign addr[61398]= 2146380306;
assign addr[61399]= 2134405552;
assign addr[61400]= 2079176953;
assign addr[61401]= 1981813720;
assign addr[61402]= 1844288924;
assign addr[61403]= 1669389513;
assign addr[61404]= 1460659832;
assign addr[61405]= 1222329801;
assign addr[61406]= 959229189;
assign addr[61407]= 676689746;
assign addr[61408]= 380437148;
assign addr[61409]= 76474970;
assign addr[61410]= -229036977;
assign addr[61411]= -529907477;
assign addr[61412]= -820039373;
assign addr[61413]= -1093553126;
assign addr[61414]= -1344905966;
assign addr[61415]= -1569004214;
assign addr[61416]= -1761306505;
assign addr[61417]= -1917915825;
assign addr[61418]= -2035658475;
assign addr[61419]= -2112148396;
assign addr[61420]= -2145835515;
assign addr[61421]= -2136037160;
assign addr[61422]= -2082951896;
assign addr[61423]= -1987655498;
assign addr[61424]= -1852079154;
assign addr[61425]= -1678970324;
assign addr[61426]= -1471837070;
assign addr[61427]= -1234876957;
assign addr[61428]= -972891995;
assign addr[61429]= -691191324;
assign addr[61430]= -395483624;
assign addr[61431]= -91761426;
assign addr[61432]= 213820322;
assign addr[61433]= 515068990;
assign addr[61434]= 805879757;
assign addr[61435]= 1080359326;
assign addr[61436]= 1332945355;
assign addr[61437]= 1558519173;
assign addr[61438]= 1752509516;
assign addr[61439]= 1910985158;
assign addr[61440]= 2030734582;
assign addr[61441]= 2109331059;
assign addr[61442]= 2145181827;
assign addr[61443]= 2137560369;
assign addr[61444]= 2086621133;
assign addr[61445]= 1993396407;
assign addr[61446]= 1859775393;
assign addr[61447]= 1688465931;
assign addr[61448]= 1482939614;
assign addr[61449]= 1247361445;
assign addr[61450]= 986505429;
assign addr[61451]= 705657826;
assign addr[61452]= 410510029;
assign addr[61453]= 107043224;
assign addr[61454]= -198592817;
assign addr[61455]= -500204365;
assign addr[61456]= -791679244;
assign addr[61457]= -1067110699;
assign addr[61458]= -1320917099;
assign addr[61459]= -1547955041;
assign addr[61460]= -1743623590;
assign addr[61461]= -1903957513;
assign addr[61462]= -2025707632;
assign addr[61463]= -2106406677;
assign addr[61464]= -2144419275;
assign addr[61465]= -2138975100;
assign addr[61466]= -2090184478;
assign addr[61467]= -1999036154;
assign addr[61468]= -1867377253;
assign addr[61469]= -1697875851;
assign addr[61470]= -1493966902;
assign addr[61471]= -1259782632;
assign addr[61472]= -1000068799;
assign addr[61473]= -720088517;
assign addr[61474]= -425515602;
assign addr[61475]= -122319591;
assign addr[61476]= 183355234;
assign addr[61477]= 485314355;
assign addr[61478]= 777438554;
assign addr[61479]= 1053807919;
assign addr[61480]= 1308821808;
assign addr[61481]= 1537312353;
assign addr[61482]= 1734649179;
assign addr[61483]= 1896833245;
assign addr[61484]= 2020577882;
assign addr[61485]= 2103375398;
assign addr[61486]= 2143547897;
assign addr[61487]= 2140281282;
assign addr[61488]= 2093641749;
assign addr[61489]= 2004574453;
assign addr[61490]= 1874884346;
assign addr[61491]= 1707199606;
assign addr[61492]= 1504918373;
assign addr[61493]= 1272139887;
assign addr[61494]= 1013581418;
assign addr[61495]= 734482665;
assign addr[61496]= 440499581;
assign addr[61497]= 137589750;
assign addr[61498]= -168108346;
assign addr[61499]= -470399716;
assign addr[61500]= -763158411;
assign addr[61501]= -1040451659;
assign addr[61502]= -1296660098;
assign addr[61503]= -1526591649;
assign addr[61504]= -1725586737;
assign addr[61505]= -1889612716;
assign addr[61506]= -2015345591;
assign addr[61507]= -2100237377;
assign addr[61508]= -2142567738;
assign addr[61509]= -2141478848;
assign addr[61510]= -2096992772;
assign addr[61511]= -2010011024;
assign addr[61512]= -1882296293;
assign addr[61513]= -1716436725;
assign addr[61514]= -1515793473;
assign addr[61515]= -1284432584;
assign addr[61516]= -1027042599;
assign addr[61517]= -748839539;
assign addr[61518]= -455461206;
assign addr[61519]= -152852926;
assign addr[61520]= 152852926;
assign addr[61521]= 455461206;
assign addr[61522]= 748839539;
assign addr[61523]= 1027042599;
assign addr[61524]= 1284432584;
assign addr[61525]= 1515793473;
assign addr[61526]= 1716436725;
assign addr[61527]= 1882296293;
assign addr[61528]= 2010011024;
assign addr[61529]= 2096992772;
assign addr[61530]= 2141478848;
assign addr[61531]= 2142567738;
assign addr[61532]= 2100237377;
assign addr[61533]= 2015345591;
assign addr[61534]= 1889612716;
assign addr[61535]= 1725586737;
assign addr[61536]= 1526591649;
assign addr[61537]= 1296660098;
assign addr[61538]= 1040451659;
assign addr[61539]= 763158411;
assign addr[61540]= 470399716;
assign addr[61541]= 168108346;
assign addr[61542]= -137589750;
assign addr[61543]= -440499581;
assign addr[61544]= -734482665;
assign addr[61545]= -1013581418;
assign addr[61546]= -1272139887;
assign addr[61547]= -1504918373;
assign addr[61548]= -1707199606;
assign addr[61549]= -1874884346;
assign addr[61550]= -2004574453;
assign addr[61551]= -2093641749;
assign addr[61552]= -2140281282;
assign addr[61553]= -2143547897;
assign addr[61554]= -2103375398;
assign addr[61555]= -2020577882;
assign addr[61556]= -1896833245;
assign addr[61557]= -1734649179;
assign addr[61558]= -1537312353;
assign addr[61559]= -1308821808;
assign addr[61560]= -1053807919;
assign addr[61561]= -777438554;
assign addr[61562]= -485314355;
assign addr[61563]= -183355234;
assign addr[61564]= 122319591;
assign addr[61565]= 425515602;
assign addr[61566]= 720088517;
assign addr[61567]= 1000068799;
assign addr[61568]= 1259782632;
assign addr[61569]= 1493966902;
assign addr[61570]= 1697875851;
assign addr[61571]= 1867377253;
assign addr[61572]= 1999036154;
assign addr[61573]= 2090184478;
assign addr[61574]= 2138975100;
assign addr[61575]= 2144419275;
assign addr[61576]= 2106406677;
assign addr[61577]= 2025707632;
assign addr[61578]= 1903957513;
assign addr[61579]= 1743623590;
assign addr[61580]= 1547955041;
assign addr[61581]= 1320917099;
assign addr[61582]= 1067110699;
assign addr[61583]= 791679244;
assign addr[61584]= 500204365;
assign addr[61585]= 198592817;
assign addr[61586]= -107043224;
assign addr[61587]= -410510029;
assign addr[61588]= -705657826;
assign addr[61589]= -986505429;
assign addr[61590]= -1247361445;
assign addr[61591]= -1482939614;
assign addr[61592]= -1688465931;
assign addr[61593]= -1859775393;
assign addr[61594]= -1993396407;
assign addr[61595]= -2086621133;
assign addr[61596]= -2137560369;
assign addr[61597]= -2145181827;
assign addr[61598]= -2109331059;
assign addr[61599]= -2030734582;
assign addr[61600]= -1910985158;
assign addr[61601]= -1752509516;
assign addr[61602]= -1558519173;
assign addr[61603]= -1332945355;
assign addr[61604]= -1080359326;
assign addr[61605]= -805879757;
assign addr[61606]= -515068990;
assign addr[61607]= -213820322;
assign addr[61608]= 91761426;
assign addr[61609]= 395483624;
assign addr[61610]= 691191324;
assign addr[61611]= 972891995;
assign addr[61612]= 1234876957;
assign addr[61613]= 1471837070;
assign addr[61614]= 1678970324;
assign addr[61615]= 1852079154;
assign addr[61616]= 1987655498;
assign addr[61617]= 2082951896;
assign addr[61618]= 2136037160;
assign addr[61619]= 2145835515;
assign addr[61620]= 2112148396;
assign addr[61621]= 2035658475;
assign addr[61622]= 1917915825;
assign addr[61623]= 1761306505;
assign addr[61624]= 1569004214;
assign addr[61625]= 1344905966;
assign addr[61626]= 1093553126;
assign addr[61627]= 820039373;
assign addr[61628]= 529907477;
assign addr[61629]= 229036977;
assign addr[61630]= -76474970;
assign addr[61631]= -380437148;
assign addr[61632]= -676689746;
assign addr[61633]= -959229189;
assign addr[61634]= -1222329801;
assign addr[61635]= -1460659832;
assign addr[61636]= -1669389513;
assign addr[61637]= -1844288924;
assign addr[61638]= -1981813720;
assign addr[61639]= -2079176953;
assign addr[61640]= -2134405552;
assign addr[61641]= -2146380306;
assign addr[61642]= -2114858546;
assign addr[61643]= -2040479063;
assign addr[61644]= -1924749160;
assign addr[61645]= -1770014111;
assign addr[61646]= -1579409630;
assign addr[61647]= -1356798326;
assign addr[61648]= -1106691431;
assign addr[61649]= -834157373;
assign addr[61650]= -544719071;
assign addr[61651]= -244242007;
assign addr[61652]= 61184634;
assign addr[61653]= 365371365;
assign addr[61654]= 662153826;
assign addr[61655]= 945517704;
assign addr[61656]= 1209720613;
assign addr[61657]= 1449408469;
assign addr[61658]= 1659723983;
assign addr[61659]= 1836405100;
assign addr[61660]= 1975871368;
assign addr[61661]= 2075296495;
assign addr[61662]= 2132665626;
assign addr[61663]= 2146816171;
assign addr[61664]= 2117461370;
assign addr[61665]= 2045196100;
assign addr[61666]= 1931484818;
assign addr[61667]= 1778631892;
assign addr[61668]= 1589734894;
assign addr[61669]= 1368621831;
assign addr[61670]= 1119773573;
assign addr[61671]= 848233042;
assign addr[61672]= 559503022;
assign addr[61673]= 259434643;
assign addr[61674]= -45891193;
assign addr[61675]= -350287041;
assign addr[61676]= -647584304;
assign addr[61677]= -931758235;
assign addr[61678]= -1197050035;
assign addr[61679]= -1438083551;
assign addr[61680]= -1649974225;
assign addr[61681]= -1828428082;
assign addr[61682]= -1969828744;
assign addr[61683]= -2071310720;
assign addr[61684]= -2130817471;
assign addr[61685]= -2147143090;
assign addr[61686]= -2119956737;
assign addr[61687]= -2049809346;
assign addr[61688]= -1938122457;
assign addr[61689]= -1787159411;
assign addr[61690]= -1599979481;
assign addr[61691]= -1380375881;
assign addr[61692]= -1132798888;
assign addr[61693]= -862265664;
assign addr[61694]= -574258580;
assign addr[61695]= -274614114;
assign addr[61696]= 30595422;
assign addr[61697]= 335184940;
assign addr[61698]= 632981917;
assign addr[61699]= 917951481;
assign addr[61700]= 1184318708;
assign addr[61701]= 1426685652;
assign addr[61702]= 1640140734;
assign addr[61703]= 1820358275;
assign addr[61704]= 1963686155;
assign addr[61705]= 2067219829;
assign addr[61706]= 2128861181;
assign addr[61707]= 2147361045;
assign addr[61708]= 2122344521;
assign addr[61709]= 2054318569;
assign addr[61710]= 1944661739;
assign addr[61711]= 1795596234;
assign addr[61712]= 1610142873;
assign addr[61713]= 1392059879;
assign addr[61714]= 1145766716;
assign addr[61715]= 876254528;
assign addr[61716]= 588984994;
assign addr[61717]= 289779648;
assign addr[61718]= -15298099;
assign addr[61719]= -320065829;
assign addr[61720]= -618347408;
assign addr[61721]= -904098143;
assign addr[61722]= -1171527280;
assign addr[61723]= -1415215352;
assign addr[61724]= -1630224009;
assign addr[61725]= -1812196087;
assign addr[61726]= -1957443913;
assign addr[61727]= -2063024031;
assign addr[61728]= -2126796855;
assign addr[61729]= -2147470025;
assign addr[61730]= -2124624598;
assign addr[61731]= -2058723538;
assign addr[61732]= -1951102334;
assign addr[61733]= -1803941934;
assign addr[61734]= -1620224553;
assign addr[61735]= -1403673233;
assign addr[61736]= -1158676398;
assign addr[61737]= -890198924;
assign addr[61738]= -603681519;
assign addr[61739]= -304930476;
assign addr[61740]= 0;
assign addr[61741]= 304930476;
assign addr[61742]= 603681519;
assign addr[61743]= 890198924;
assign addr[61744]= 1158676398;
assign addr[61745]= 1403673233;
assign addr[61746]= 1620224553;
assign addr[61747]= 1803941934;
assign addr[61748]= 1951102334;
assign addr[61749]= 2058723538;
assign addr[61750]= 2124624598;
assign addr[61751]= 2147470025;
assign addr[61752]= 2126796855;
assign addr[61753]= 2063024031;
assign addr[61754]= 1957443913;
assign addr[61755]= 1812196087;
assign addr[61756]= 1630224009;
assign addr[61757]= 1415215352;
assign addr[61758]= 1171527280;
assign addr[61759]= 904098143;
assign addr[61760]= 618347408;
assign addr[61761]= 320065829;
assign addr[61762]= 15298099;
assign addr[61763]= -289779648;
assign addr[61764]= -588984994;
assign addr[61765]= -876254528;
assign addr[61766]= -1145766716;
assign addr[61767]= -1392059879;
assign addr[61768]= -1610142873;
assign addr[61769]= -1795596234;
assign addr[61770]= -1944661739;
assign addr[61771]= -2054318569;
assign addr[61772]= -2122344521;
assign addr[61773]= -2147361045;
assign addr[61774]= -2128861181;
assign addr[61775]= -2067219829;
assign addr[61776]= -1963686155;
assign addr[61777]= -1820358275;
assign addr[61778]= -1640140734;
assign addr[61779]= -1426685652;
assign addr[61780]= -1184318708;
assign addr[61781]= -917951481;
assign addr[61782]= -632981917;
assign addr[61783]= -335184940;
assign addr[61784]= -30595422;
assign addr[61785]= 274614114;
assign addr[61786]= 574258580;
assign addr[61787]= 862265664;
assign addr[61788]= 1132798888;
assign addr[61789]= 1380375881;
assign addr[61790]= 1599979481;
assign addr[61791]= 1787159411;
assign addr[61792]= 1938122457;
assign addr[61793]= 2049809346;
assign addr[61794]= 2119956737;
assign addr[61795]= 2147143090;
assign addr[61796]= 2130817471;
assign addr[61797]= 2071310720;
assign addr[61798]= 1969828744;
assign addr[61799]= 1828428082;
assign addr[61800]= 1649974225;
assign addr[61801]= 1438083551;
assign addr[61802]= 1197050035;
assign addr[61803]= 931758235;
assign addr[61804]= 647584304;
assign addr[61805]= 350287041;
assign addr[61806]= 45891193;
assign addr[61807]= -259434643;
assign addr[61808]= -559503022;
assign addr[61809]= -848233042;
assign addr[61810]= -1119773573;
assign addr[61811]= -1368621831;
assign addr[61812]= -1589734894;
assign addr[61813]= -1778631892;
assign addr[61814]= -1931484818;
assign addr[61815]= -2045196100;
assign addr[61816]= -2117461370;
assign addr[61817]= -2146816171;
assign addr[61818]= -2132665626;
assign addr[61819]= -2075296495;
assign addr[61820]= -1975871368;
assign addr[61821]= -1836405100;
assign addr[61822]= -1659723983;
assign addr[61823]= -1449408469;
assign addr[61824]= -1209720613;
assign addr[61825]= -945517704;
assign addr[61826]= -662153826;
assign addr[61827]= -365371365;
assign addr[61828]= -61184634;
assign addr[61829]= 244242007;
assign addr[61830]= 544719071;
assign addr[61831]= 834157373;
assign addr[61832]= 1106691431;
assign addr[61833]= 1356798326;
assign addr[61834]= 1579409630;
assign addr[61835]= 1770014111;
assign addr[61836]= 1924749160;
assign addr[61837]= 2040479063;
assign addr[61838]= 2114858546;
assign addr[61839]= 2146380306;
assign addr[61840]= 2134405552;
assign addr[61841]= 2079176953;
assign addr[61842]= 1981813720;
assign addr[61843]= 1844288924;
assign addr[61844]= 1669389513;
assign addr[61845]= 1460659832;
assign addr[61846]= 1222329801;
assign addr[61847]= 959229189;
assign addr[61848]= 676689746;
assign addr[61849]= 380437148;
assign addr[61850]= 76474970;
assign addr[61851]= -229036977;
assign addr[61852]= -529907477;
assign addr[61853]= -820039373;
assign addr[61854]= -1093553126;
assign addr[61855]= -1344905966;
assign addr[61856]= -1569004214;
assign addr[61857]= -1761306505;
assign addr[61858]= -1917915825;
assign addr[61859]= -2035658475;
assign addr[61860]= -2112148396;
assign addr[61861]= -2145835515;
assign addr[61862]= -2136037160;
assign addr[61863]= -2082951896;
assign addr[61864]= -1987655498;
assign addr[61865]= -1852079154;
assign addr[61866]= -1678970324;
assign addr[61867]= -1471837070;
assign addr[61868]= -1234876957;
assign addr[61869]= -972891995;
assign addr[61870]= -691191324;
assign addr[61871]= -395483624;
assign addr[61872]= -91761426;
assign addr[61873]= 213820322;
assign addr[61874]= 515068990;
assign addr[61875]= 805879757;
assign addr[61876]= 1080359326;
assign addr[61877]= 1332945355;
assign addr[61878]= 1558519173;
assign addr[61879]= 1752509516;
assign addr[61880]= 1910985158;
assign addr[61881]= 2030734582;
assign addr[61882]= 2109331059;
assign addr[61883]= 2145181827;
assign addr[61884]= 2137560369;
assign addr[61885]= 2086621133;
assign addr[61886]= 1993396407;
assign addr[61887]= 1859775393;
assign addr[61888]= 1688465931;
assign addr[61889]= 1482939614;
assign addr[61890]= 1247361445;
assign addr[61891]= 986505429;
assign addr[61892]= 705657826;
assign addr[61893]= 410510029;
assign addr[61894]= 107043224;
assign addr[61895]= -198592817;
assign addr[61896]= -500204365;
assign addr[61897]= -791679244;
assign addr[61898]= -1067110699;
assign addr[61899]= -1320917099;
assign addr[61900]= -1547955041;
assign addr[61901]= -1743623590;
assign addr[61902]= -1903957513;
assign addr[61903]= -2025707632;
assign addr[61904]= -2106406677;
assign addr[61905]= -2144419275;
assign addr[61906]= -2138975100;
assign addr[61907]= -2090184478;
assign addr[61908]= -1999036154;
assign addr[61909]= -1867377253;
assign addr[61910]= -1697875851;
assign addr[61911]= -1493966902;
assign addr[61912]= -1259782632;
assign addr[61913]= -1000068799;
assign addr[61914]= -720088517;
assign addr[61915]= -425515602;
assign addr[61916]= -122319591;
assign addr[61917]= 183355234;
assign addr[61918]= 485314355;
assign addr[61919]= 777438554;
assign addr[61920]= 1053807919;
assign addr[61921]= 1308821808;
assign addr[61922]= 1537312353;
assign addr[61923]= 1734649179;
assign addr[61924]= 1896833245;
assign addr[61925]= 2020577882;
assign addr[61926]= 2103375398;
assign addr[61927]= 2143547897;
assign addr[61928]= 2140281282;
assign addr[61929]= 2093641749;
assign addr[61930]= 2004574453;
assign addr[61931]= 1874884346;
assign addr[61932]= 1707199606;
assign addr[61933]= 1504918373;
assign addr[61934]= 1272139887;
assign addr[61935]= 1013581418;
assign addr[61936]= 734482665;
assign addr[61937]= 440499581;
assign addr[61938]= 137589750;
assign addr[61939]= -168108346;
assign addr[61940]= -470399716;
assign addr[61941]= -763158411;
assign addr[61942]= -1040451659;
assign addr[61943]= -1296660098;
assign addr[61944]= -1526591649;
assign addr[61945]= -1725586737;
assign addr[61946]= -1889612716;
assign addr[61947]= -2015345591;
assign addr[61948]= -2100237377;
assign addr[61949]= -2142567738;
assign addr[61950]= -2141478848;
assign addr[61951]= -2096992772;
assign addr[61952]= -2010011024;
assign addr[61953]= -1882296293;
assign addr[61954]= -1716436725;
assign addr[61955]= -1515793473;
assign addr[61956]= -1284432584;
assign addr[61957]= -1027042599;
assign addr[61958]= -748839539;
assign addr[61959]= -455461206;
assign addr[61960]= -152852926;
assign addr[61961]= 152852926;
assign addr[61962]= 455461206;
assign addr[61963]= 748839539;
assign addr[61964]= 1027042599;
assign addr[61965]= 1284432584;
assign addr[61966]= 1515793473;
assign addr[61967]= 1716436725;
assign addr[61968]= 1882296293;
assign addr[61969]= 2010011024;
assign addr[61970]= 2096992772;
assign addr[61971]= 2141478848;
assign addr[61972]= 2142567738;
assign addr[61973]= 2100237377;
assign addr[61974]= 2015345591;
assign addr[61975]= 1889612716;
assign addr[61976]= 1725586737;
assign addr[61977]= 1526591649;
assign addr[61978]= 1296660098;
assign addr[61979]= 1040451659;
assign addr[61980]= 763158411;
assign addr[61981]= 470399716;
assign addr[61982]= 168108346;
assign addr[61983]= -137589750;
assign addr[61984]= -440499581;
assign addr[61985]= -734482665;
assign addr[61986]= -1013581418;
assign addr[61987]= -1272139887;
assign addr[61988]= -1504918373;
assign addr[61989]= -1707199606;
assign addr[61990]= -1874884346;
assign addr[61991]= -2004574453;
assign addr[61992]= -2093641749;
assign addr[61993]= -2140281282;
assign addr[61994]= -2143547897;
assign addr[61995]= -2103375398;
assign addr[61996]= -2020577882;
assign addr[61997]= -1896833245;
assign addr[61998]= -1734649179;
assign addr[61999]= -1537312353;
assign addr[62000]= -1308821808;
assign addr[62001]= -1053807919;
assign addr[62002]= -777438554;
assign addr[62003]= -485314355;
assign addr[62004]= -183355234;
assign addr[62005]= 122319591;
assign addr[62006]= 425515602;
assign addr[62007]= 720088517;
assign addr[62008]= 1000068799;
assign addr[62009]= 1259782632;
assign addr[62010]= 1493966902;
assign addr[62011]= 1697875851;
assign addr[62012]= 1867377253;
assign addr[62013]= 1999036154;
assign addr[62014]= 2090184478;
assign addr[62015]= 2138975100;
assign addr[62016]= 2144419275;
assign addr[62017]= 2106406677;
assign addr[62018]= 2025707632;
assign addr[62019]= 1903957513;
assign addr[62020]= 1743623590;
assign addr[62021]= 1547955041;
assign addr[62022]= 1320917099;
assign addr[62023]= 1067110699;
assign addr[62024]= 791679244;
assign addr[62025]= 500204365;
assign addr[62026]= 198592817;
assign addr[62027]= -107043224;
assign addr[62028]= -410510029;
assign addr[62029]= -705657826;
assign addr[62030]= -986505429;
assign addr[62031]= -1247361445;
assign addr[62032]= -1482939614;
assign addr[62033]= -1688465931;
assign addr[62034]= -1859775393;
assign addr[62035]= -1993396407;
assign addr[62036]= -2086621133;
assign addr[62037]= -2137560369;
assign addr[62038]= -2145181827;
assign addr[62039]= -2109331059;
assign addr[62040]= -2030734582;
assign addr[62041]= -1910985158;
assign addr[62042]= -1752509516;
assign addr[62043]= -1558519173;
assign addr[62044]= -1332945355;
assign addr[62045]= -1080359326;
assign addr[62046]= -805879757;
assign addr[62047]= -515068990;
assign addr[62048]= -213820322;
assign addr[62049]= 91761426;
assign addr[62050]= 395483624;
assign addr[62051]= 691191324;
assign addr[62052]= 972891995;
assign addr[62053]= 1234876957;
assign addr[62054]= 1471837070;
assign addr[62055]= 1678970324;
assign addr[62056]= 1852079154;
assign addr[62057]= 1987655498;
assign addr[62058]= 2082951896;
assign addr[62059]= 2136037160;
assign addr[62060]= 2145835515;
assign addr[62061]= 2112148396;
assign addr[62062]= 2035658475;
assign addr[62063]= 1917915825;
assign addr[62064]= 1761306505;
assign addr[62065]= 1569004214;
assign addr[62066]= 1344905966;
assign addr[62067]= 1093553126;
assign addr[62068]= 820039373;
assign addr[62069]= 529907477;
assign addr[62070]= 229036977;
assign addr[62071]= -76474970;
assign addr[62072]= -380437148;
assign addr[62073]= -676689746;
assign addr[62074]= -959229189;
assign addr[62075]= -1222329801;
assign addr[62076]= -1460659832;
assign addr[62077]= -1669389513;
assign addr[62078]= -1844288924;
assign addr[62079]= -1981813720;
assign addr[62080]= -2079176953;
assign addr[62081]= -2134405552;
assign addr[62082]= -2146380306;
assign addr[62083]= -2114858546;
assign addr[62084]= -2040479063;
assign addr[62085]= -1924749160;
assign addr[62086]= -1770014111;
assign addr[62087]= -1579409630;
assign addr[62088]= -1356798326;
assign addr[62089]= -1106691431;
assign addr[62090]= -834157373;
assign addr[62091]= -544719071;
assign addr[62092]= -244242007;
assign addr[62093]= 61184634;
assign addr[62094]= 365371365;
assign addr[62095]= 662153826;
assign addr[62096]= 945517704;
assign addr[62097]= 1209720613;
assign addr[62098]= 1449408469;
assign addr[62099]= 1659723983;
assign addr[62100]= 1836405100;
assign addr[62101]= 1975871368;
assign addr[62102]= 2075296495;
assign addr[62103]= 2132665626;
assign addr[62104]= 2146816171;
assign addr[62105]= 2117461370;
assign addr[62106]= 2045196100;
assign addr[62107]= 1931484818;
assign addr[62108]= 1778631892;
assign addr[62109]= 1589734894;
assign addr[62110]= 1368621831;
assign addr[62111]= 1119773573;
assign addr[62112]= 848233042;
assign addr[62113]= 559503022;
assign addr[62114]= 259434643;
assign addr[62115]= -45891193;
assign addr[62116]= -350287041;
assign addr[62117]= -647584304;
assign addr[62118]= -931758235;
assign addr[62119]= -1197050035;
assign addr[62120]= -1438083551;
assign addr[62121]= -1649974225;
assign addr[62122]= -1828428082;
assign addr[62123]= -1969828744;
assign addr[62124]= -2071310720;
assign addr[62125]= -2130817471;
assign addr[62126]= -2147143090;
assign addr[62127]= -2119956737;
assign addr[62128]= -2049809346;
assign addr[62129]= -1938122457;
assign addr[62130]= -1787159411;
assign addr[62131]= -1599979481;
assign addr[62132]= -1380375881;
assign addr[62133]= -1132798888;
assign addr[62134]= -862265664;
assign addr[62135]= -574258580;
assign addr[62136]= -274614114;
assign addr[62137]= 30595422;
assign addr[62138]= 335184940;
assign addr[62139]= 632981917;
assign addr[62140]= 917951481;
assign addr[62141]= 1184318708;
assign addr[62142]= 1426685652;
assign addr[62143]= 1640140734;
assign addr[62144]= 1820358275;
assign addr[62145]= 1963686155;
assign addr[62146]= 2067219829;
assign addr[62147]= 2128861181;
assign addr[62148]= 2147361045;
assign addr[62149]= 2122344521;
assign addr[62150]= 2054318569;
assign addr[62151]= 1944661739;
assign addr[62152]= 1795596234;
assign addr[62153]= 1610142873;
assign addr[62154]= 1392059879;
assign addr[62155]= 1145766716;
assign addr[62156]= 876254528;
assign addr[62157]= 588984994;
assign addr[62158]= 289779648;
assign addr[62159]= -15298099;
assign addr[62160]= -320065829;
assign addr[62161]= -618347408;
assign addr[62162]= -904098143;
assign addr[62163]= -1171527280;
assign addr[62164]= -1415215352;
assign addr[62165]= -1630224009;
assign addr[62166]= -1812196087;
assign addr[62167]= -1957443913;
assign addr[62168]= -2063024031;
assign addr[62169]= -2126796855;
assign addr[62170]= -2147470025;
assign addr[62171]= -2124624598;
assign addr[62172]= -2058723538;
assign addr[62173]= -1951102334;
assign addr[62174]= -1803941934;
assign addr[62175]= -1620224553;
assign addr[62176]= -1403673233;
assign addr[62177]= -1158676398;
assign addr[62178]= -890198924;
assign addr[62179]= -603681519;
assign addr[62180]= -304930476;
assign addr[62181]= 0;
assign addr[62182]= 304930476;
assign addr[62183]= 603681519;
assign addr[62184]= 890198924;
assign addr[62185]= 1158676398;
assign addr[62186]= 1403673233;
assign addr[62187]= 1620224553;
assign addr[62188]= 1803941934;
assign addr[62189]= 1951102334;
assign addr[62190]= 2058723538;
assign addr[62191]= 2124624598;
assign addr[62192]= 2147470025;
assign addr[62193]= 2126796855;
assign addr[62194]= 2063024031;
assign addr[62195]= 1957443913;
assign addr[62196]= 1812196087;
assign addr[62197]= 1630224009;
assign addr[62198]= 1415215352;
assign addr[62199]= 1171527280;
assign addr[62200]= 904098143;
assign addr[62201]= 618347408;
assign addr[62202]= 320065829;
assign addr[62203]= 15298099;
assign addr[62204]= -289779648;
assign addr[62205]= -588984994;
assign addr[62206]= -876254528;
assign addr[62207]= -1145766716;
assign addr[62208]= -1392059879;
assign addr[62209]= -1610142873;
assign addr[62210]= -1795596234;
assign addr[62211]= -1944661739;
assign addr[62212]= -2054318569;
assign addr[62213]= -2122344521;
assign addr[62214]= -2147361045;
assign addr[62215]= -2128861181;
assign addr[62216]= -2067219829;
assign addr[62217]= -1963686155;
assign addr[62218]= -1820358275;
assign addr[62219]= -1640140734;
assign addr[62220]= -1426685652;
assign addr[62221]= -1184318708;
assign addr[62222]= -917951481;
assign addr[62223]= -632981917;
assign addr[62224]= -335184940;
assign addr[62225]= -30595422;
assign addr[62226]= 274614114;
assign addr[62227]= 574258580;
assign addr[62228]= 862265664;
assign addr[62229]= 1132798888;
assign addr[62230]= 1380375881;
assign addr[62231]= 1599979481;
assign addr[62232]= 1787159411;
assign addr[62233]= 1938122457;
assign addr[62234]= 2049809346;
assign addr[62235]= 2119956737;
assign addr[62236]= 2147143090;
assign addr[62237]= 2130817471;
assign addr[62238]= 2071310720;
assign addr[62239]= 1969828744;
assign addr[62240]= 1828428082;
assign addr[62241]= 1649974225;
assign addr[62242]= 1438083551;
assign addr[62243]= 1197050035;
assign addr[62244]= 931758235;
assign addr[62245]= 647584304;
assign addr[62246]= 350287041;
assign addr[62247]= 45891193;
assign addr[62248]= -259434643;
assign addr[62249]= -559503022;
assign addr[62250]= -848233042;
assign addr[62251]= -1119773573;
assign addr[62252]= -1368621831;
assign addr[62253]= -1589734894;
assign addr[62254]= -1778631892;
assign addr[62255]= -1931484818;
assign addr[62256]= -2045196100;
assign addr[62257]= -2117461370;
assign addr[62258]= -2146816171;
assign addr[62259]= -2132665626;
assign addr[62260]= -2075296495;
assign addr[62261]= -1975871368;
assign addr[62262]= -1836405100;
assign addr[62263]= -1659723983;
assign addr[62264]= -1449408469;
assign addr[62265]= -1209720613;
assign addr[62266]= -945517704;
assign addr[62267]= -662153826;
assign addr[62268]= -365371365;
assign addr[62269]= -61184634;
assign addr[62270]= 244242007;
assign addr[62271]= 544719071;
assign addr[62272]= 834157373;
assign addr[62273]= 1106691431;
assign addr[62274]= 1356798326;
assign addr[62275]= 1579409630;
assign addr[62276]= 1770014111;
assign addr[62277]= 1924749160;
assign addr[62278]= 2040479063;
assign addr[62279]= 2114858546;
assign addr[62280]= 2146380306;
assign addr[62281]= 2134405552;
assign addr[62282]= 2079176953;
assign addr[62283]= 1981813720;
assign addr[62284]= 1844288924;
assign addr[62285]= 1669389513;
assign addr[62286]= 1460659832;
assign addr[62287]= 1222329801;
assign addr[62288]= 959229189;
assign addr[62289]= 676689746;
assign addr[62290]= 380437148;
assign addr[62291]= 76474970;
assign addr[62292]= -229036977;
assign addr[62293]= -529907477;
assign addr[62294]= -820039373;
assign addr[62295]= -1093553126;
assign addr[62296]= -1344905966;
assign addr[62297]= -1569004214;
assign addr[62298]= -1761306505;
assign addr[62299]= -1917915825;
assign addr[62300]= -2035658475;
assign addr[62301]= -2112148396;
assign addr[62302]= -2145835515;
assign addr[62303]= -2136037160;
assign addr[62304]= -2082951896;
assign addr[62305]= -1987655498;
assign addr[62306]= -1852079154;
assign addr[62307]= -1678970324;
assign addr[62308]= -1471837070;
assign addr[62309]= -1234876957;
assign addr[62310]= -972891995;
assign addr[62311]= -691191324;
assign addr[62312]= -395483624;
assign addr[62313]= -91761426;
assign addr[62314]= 213820322;
assign addr[62315]= 515068990;
assign addr[62316]= 805879757;
assign addr[62317]= 1080359326;
assign addr[62318]= 1332945355;
assign addr[62319]= 1558519173;
assign addr[62320]= 1752509516;
assign addr[62321]= 1910985158;
assign addr[62322]= 2030734582;
assign addr[62323]= 2109331059;
assign addr[62324]= 2145181827;
assign addr[62325]= 2137560369;
assign addr[62326]= 2086621133;
assign addr[62327]= 1993396407;
assign addr[62328]= 1859775393;
assign addr[62329]= 1688465931;
assign addr[62330]= 1482939614;
assign addr[62331]= 1247361445;
assign addr[62332]= 986505429;
assign addr[62333]= 705657826;
assign addr[62334]= 410510029;
assign addr[62335]= 107043224;
assign addr[62336]= -198592817;
assign addr[62337]= -500204365;
assign addr[62338]= -791679244;
assign addr[62339]= -1067110699;
assign addr[62340]= -1320917099;
assign addr[62341]= -1547955041;
assign addr[62342]= -1743623590;
assign addr[62343]= -1903957513;
assign addr[62344]= -2025707632;
assign addr[62345]= -2106406677;
assign addr[62346]= -2144419275;
assign addr[62347]= -2138975100;
assign addr[62348]= -2090184478;
assign addr[62349]= -1999036154;
assign addr[62350]= -1867377253;
assign addr[62351]= -1697875851;
assign addr[62352]= -1493966902;
assign addr[62353]= -1259782632;
assign addr[62354]= -1000068799;
assign addr[62355]= -720088517;
assign addr[62356]= -425515602;
assign addr[62357]= -122319591;
assign addr[62358]= 183355234;
assign addr[62359]= 485314355;
assign addr[62360]= 777438554;
assign addr[62361]= 1053807919;
assign addr[62362]= 1308821808;
assign addr[62363]= 1537312353;
assign addr[62364]= 1734649179;
assign addr[62365]= 1896833245;
assign addr[62366]= 2020577882;
assign addr[62367]= 2103375398;
assign addr[62368]= 2143547897;
assign addr[62369]= 2140281282;
assign addr[62370]= 2093641749;
assign addr[62371]= 2004574453;
assign addr[62372]= 1874884346;
assign addr[62373]= 1707199606;
assign addr[62374]= 1504918373;
assign addr[62375]= 1272139887;
assign addr[62376]= 1013581418;
assign addr[62377]= 734482665;
assign addr[62378]= 440499581;
assign addr[62379]= 137589750;
assign addr[62380]= -168108346;
assign addr[62381]= -470399716;
assign addr[62382]= -763158411;
assign addr[62383]= -1040451659;
assign addr[62384]= -1296660098;
assign addr[62385]= -1526591649;
assign addr[62386]= -1725586737;
assign addr[62387]= -1889612716;
assign addr[62388]= -2015345591;
assign addr[62389]= -2100237377;
assign addr[62390]= -2142567738;
assign addr[62391]= -2141478848;
assign addr[62392]= -2096992772;
assign addr[62393]= -2010011024;
assign addr[62394]= -1882296293;
assign addr[62395]= -1716436725;
assign addr[62396]= -1515793473;
assign addr[62397]= -1284432584;
assign addr[62398]= -1027042599;
assign addr[62399]= -748839539;
assign addr[62400]= -455461206;
assign addr[62401]= -152852926;
assign addr[62402]= 152852926;
assign addr[62403]= 455461206;
assign addr[62404]= 748839539;
assign addr[62405]= 1027042599;
assign addr[62406]= 1284432584;
assign addr[62407]= 1515793473;
assign addr[62408]= 1716436725;
assign addr[62409]= 1882296293;
assign addr[62410]= 2010011024;
assign addr[62411]= 2096992772;
assign addr[62412]= 2141478848;
assign addr[62413]= 2142567738;
assign addr[62414]= 2100237377;
assign addr[62415]= 2015345591;
assign addr[62416]= 1889612716;
assign addr[62417]= 1725586737;
assign addr[62418]= 1526591649;
assign addr[62419]= 1296660098;
assign addr[62420]= 1040451659;
assign addr[62421]= 763158411;
assign addr[62422]= 470399716;
assign addr[62423]= 168108346;
assign addr[62424]= -137589750;
assign addr[62425]= -440499581;
assign addr[62426]= -734482665;
assign addr[62427]= -1013581418;
assign addr[62428]= -1272139887;
assign addr[62429]= -1504918373;
assign addr[62430]= -1707199606;
assign addr[62431]= -1874884346;
assign addr[62432]= -2004574453;
assign addr[62433]= -2093641749;
assign addr[62434]= -2140281282;
assign addr[62435]= -2143547897;
assign addr[62436]= -2103375398;
assign addr[62437]= -2020577882;
assign addr[62438]= -1896833245;
assign addr[62439]= -1734649179;
assign addr[62440]= -1537312353;
assign addr[62441]= -1308821808;
assign addr[62442]= -1053807919;
assign addr[62443]= -777438554;
assign addr[62444]= -485314355;
assign addr[62445]= -183355234;
assign addr[62446]= 122319591;
assign addr[62447]= 425515602;
assign addr[62448]= 720088517;
assign addr[62449]= 1000068799;
assign addr[62450]= 1259782632;
assign addr[62451]= 1493966902;
assign addr[62452]= 1697875851;
assign addr[62453]= 1867377253;
assign addr[62454]= 1999036154;
assign addr[62455]= 2090184478;
assign addr[62456]= 2138975100;
assign addr[62457]= 2144419275;
assign addr[62458]= 2106406677;
assign addr[62459]= 2025707632;
assign addr[62460]= 1903957513;
assign addr[62461]= 1743623590;
assign addr[62462]= 1547955041;
assign addr[62463]= 1320917099;
assign addr[62464]= 1067110699;
assign addr[62465]= 791679244;
assign addr[62466]= 500204365;
assign addr[62467]= 198592817;
assign addr[62468]= -107043224;
assign addr[62469]= -410510029;
assign addr[62470]= -705657826;
assign addr[62471]= -986505429;
assign addr[62472]= -1247361445;
assign addr[62473]= -1482939614;
assign addr[62474]= -1688465931;
assign addr[62475]= -1859775393;
assign addr[62476]= -1993396407;
assign addr[62477]= -2086621133;
assign addr[62478]= -2137560369;
assign addr[62479]= -2145181827;
assign addr[62480]= -2109331059;
assign addr[62481]= -2030734582;
assign addr[62482]= -1910985158;
assign addr[62483]= -1752509516;
assign addr[62484]= -1558519173;
assign addr[62485]= -1332945355;
assign addr[62486]= -1080359326;
assign addr[62487]= -805879757;
assign addr[62488]= -515068990;
assign addr[62489]= -213820322;
assign addr[62490]= 91761426;
assign addr[62491]= 395483624;
assign addr[62492]= 691191324;
assign addr[62493]= 972891995;
assign addr[62494]= 1234876957;
assign addr[62495]= 1471837070;
assign addr[62496]= 1678970324;
assign addr[62497]= 1852079154;
assign addr[62498]= 1987655498;
assign addr[62499]= 2082951896;
assign addr[62500]= 2136037160;
assign addr[62501]= 2145835515;
assign addr[62502]= 2112148396;
assign addr[62503]= 2035658475;
assign addr[62504]= 1917915825;
assign addr[62505]= 1761306505;
assign addr[62506]= 1569004214;
assign addr[62507]= 1344905966;
assign addr[62508]= 1093553126;
assign addr[62509]= 820039373;
assign addr[62510]= 529907477;
assign addr[62511]= 229036977;
assign addr[62512]= -76474970;
assign addr[62513]= -380437148;
assign addr[62514]= -676689746;
assign addr[62515]= -959229189;
assign addr[62516]= -1222329801;
assign addr[62517]= -1460659832;
assign addr[62518]= -1669389513;
assign addr[62519]= -1844288924;
assign addr[62520]= -1981813720;
assign addr[62521]= -2079176953;
assign addr[62522]= -2134405552;
assign addr[62523]= -2146380306;
assign addr[62524]= -2114858546;
assign addr[62525]= -2040479063;
assign addr[62526]= -1924749160;
assign addr[62527]= -1770014111;
assign addr[62528]= -1579409630;
assign addr[62529]= -1356798326;
assign addr[62530]= -1106691431;
assign addr[62531]= -834157373;
assign addr[62532]= -544719071;
assign addr[62533]= -244242007;
assign addr[62534]= 61184634;
assign addr[62535]= 365371365;
assign addr[62536]= 662153826;
assign addr[62537]= 945517704;
assign addr[62538]= 1209720613;
assign addr[62539]= 1449408469;
assign addr[62540]= 1659723983;
assign addr[62541]= 1836405100;
assign addr[62542]= 1975871368;
assign addr[62543]= 2075296495;
assign addr[62544]= 2132665626;
assign addr[62545]= 2146816171;
assign addr[62546]= 2117461370;
assign addr[62547]= 2045196100;
assign addr[62548]= 1931484818;
assign addr[62549]= 1778631892;
assign addr[62550]= 1589734894;
assign addr[62551]= 1368621831;
assign addr[62552]= 1119773573;
assign addr[62553]= 848233042;
assign addr[62554]= 559503022;
assign addr[62555]= 259434643;
assign addr[62556]= -45891193;
assign addr[62557]= -350287041;
assign addr[62558]= -647584304;
assign addr[62559]= -931758235;
assign addr[62560]= -1197050035;
assign addr[62561]= -1438083551;
assign addr[62562]= -1649974225;
assign addr[62563]= -1828428082;
assign addr[62564]= -1969828744;
assign addr[62565]= -2071310720;
assign addr[62566]= -2130817471;
assign addr[62567]= -2147143090;
assign addr[62568]= -2119956737;
assign addr[62569]= -2049809346;
assign addr[62570]= -1938122457;
assign addr[62571]= -1787159411;
assign addr[62572]= -1599979481;
assign addr[62573]= -1380375881;
assign addr[62574]= -1132798888;
assign addr[62575]= -862265664;
assign addr[62576]= -574258580;
assign addr[62577]= -274614114;
assign addr[62578]= 30595422;
assign addr[62579]= 335184940;
assign addr[62580]= 632981917;
assign addr[62581]= 917951481;
assign addr[62582]= 1184318708;
assign addr[62583]= 1426685652;
assign addr[62584]= 1640140734;
assign addr[62585]= 1820358275;
assign addr[62586]= 1963686155;
assign addr[62587]= 2067219829;
assign addr[62588]= 2128861181;
assign addr[62589]= 2147361045;
assign addr[62590]= 2122344521;
assign addr[62591]= 2054318569;
assign addr[62592]= 1944661739;
assign addr[62593]= 1795596234;
assign addr[62594]= 1610142873;
assign addr[62595]= 1392059879;
assign addr[62596]= 1145766716;
assign addr[62597]= 876254528;
assign addr[62598]= 588984994;
assign addr[62599]= 289779648;
assign addr[62600]= -15298099;
assign addr[62601]= -320065829;
assign addr[62602]= -618347408;
assign addr[62603]= -904098143;
assign addr[62604]= -1171527280;
assign addr[62605]= -1415215352;
assign addr[62606]= -1630224009;
assign addr[62607]= -1812196087;
assign addr[62608]= -1957443913;
assign addr[62609]= -2063024031;
assign addr[62610]= -2126796855;
assign addr[62611]= -2147470025;
assign addr[62612]= -2124624598;
assign addr[62613]= -2058723538;
assign addr[62614]= -1951102334;
assign addr[62615]= -1803941934;
assign addr[62616]= -1620224553;
assign addr[62617]= -1403673233;
assign addr[62618]= -1158676398;
assign addr[62619]= -890198924;
assign addr[62620]= -603681519;
assign addr[62621]= -304930476;
assign addr[62622]= 0;
assign addr[62623]= 304930476;
assign addr[62624]= 603681519;
assign addr[62625]= 890198924;
assign addr[62626]= 1158676398;
assign addr[62627]= 1403673233;
assign addr[62628]= 1620224553;
assign addr[62629]= 1803941934;
assign addr[62630]= 1951102334;
assign addr[62631]= 2058723538;
assign addr[62632]= 2124624598;
assign addr[62633]= 2147470025;
assign addr[62634]= 2126796855;
assign addr[62635]= 2063024031;
assign addr[62636]= 1957443913;
assign addr[62637]= 1812196087;
assign addr[62638]= 1630224009;
assign addr[62639]= 1415215352;
assign addr[62640]= 1171527280;
assign addr[62641]= 904098143;
assign addr[62642]= 618347408;
assign addr[62643]= 320065829;
assign addr[62644]= 15298099;
assign addr[62645]= -289779648;
assign addr[62646]= -588984994;
assign addr[62647]= -876254528;
assign addr[62648]= -1145766716;
assign addr[62649]= -1392059879;
assign addr[62650]= -1610142873;
assign addr[62651]= -1795596234;
assign addr[62652]= -1944661739;
assign addr[62653]= -2054318569;
assign addr[62654]= -2122344521;
assign addr[62655]= -2147361045;
assign addr[62656]= -2128861181;
assign addr[62657]= -2067219829;
assign addr[62658]= -1963686155;
assign addr[62659]= -1820358275;
assign addr[62660]= -1640140734;
assign addr[62661]= -1426685652;
assign addr[62662]= -1184318708;
assign addr[62663]= -917951481;
assign addr[62664]= -632981917;
assign addr[62665]= -335184940;
assign addr[62666]= -30595422;
assign addr[62667]= 274614114;
assign addr[62668]= 574258580;
assign addr[62669]= 862265664;
assign addr[62670]= 1132798888;
assign addr[62671]= 1380375881;
assign addr[62672]= 1599979481;
assign addr[62673]= 1787159411;
assign addr[62674]= 1938122457;
assign addr[62675]= 2049809346;
assign addr[62676]= 2119956737;
assign addr[62677]= 2147143090;
assign addr[62678]= 2130817471;
assign addr[62679]= 2071310720;
assign addr[62680]= 1969828744;
assign addr[62681]= 1828428082;
assign addr[62682]= 1649974225;
assign addr[62683]= 1438083551;
assign addr[62684]= 1197050035;
assign addr[62685]= 931758235;
assign addr[62686]= 647584304;
assign addr[62687]= 350287041;
assign addr[62688]= 45891193;
assign addr[62689]= -259434643;
assign addr[62690]= -559503022;
assign addr[62691]= -848233042;
assign addr[62692]= -1119773573;
assign addr[62693]= -1368621831;
assign addr[62694]= -1589734894;
assign addr[62695]= -1778631892;
assign addr[62696]= -1931484818;
assign addr[62697]= -2045196100;
assign addr[62698]= -2117461370;
assign addr[62699]= -2146816171;
assign addr[62700]= -2132665626;
assign addr[62701]= -2075296495;
assign addr[62702]= -1975871368;
assign addr[62703]= -1836405100;
assign addr[62704]= -1659723983;
assign addr[62705]= -1449408469;
assign addr[62706]= -1209720613;
assign addr[62707]= -945517704;
assign addr[62708]= -662153826;
assign addr[62709]= -365371365;
assign addr[62710]= -61184634;
assign addr[62711]= 244242007;
assign addr[62712]= 544719071;
assign addr[62713]= 834157373;
assign addr[62714]= 1106691431;
assign addr[62715]= 1356798326;
assign addr[62716]= 1579409630;
assign addr[62717]= 1770014111;
assign addr[62718]= 1924749160;
assign addr[62719]= 2040479063;
assign addr[62720]= 2114858546;
assign addr[62721]= 2146380306;
assign addr[62722]= 2134405552;
assign addr[62723]= 2079176953;
assign addr[62724]= 1981813720;
assign addr[62725]= 1844288924;
assign addr[62726]= 1669389513;
assign addr[62727]= 1460659832;
assign addr[62728]= 1222329801;
assign addr[62729]= 959229189;
assign addr[62730]= 676689746;
assign addr[62731]= 380437148;
assign addr[62732]= 76474970;
assign addr[62733]= -229036977;
assign addr[62734]= -529907477;
assign addr[62735]= -820039373;
assign addr[62736]= -1093553126;
assign addr[62737]= -1344905966;
assign addr[62738]= -1569004214;
assign addr[62739]= -1761306505;
assign addr[62740]= -1917915825;
assign addr[62741]= -2035658475;
assign addr[62742]= -2112148396;
assign addr[62743]= -2145835515;
assign addr[62744]= -2136037160;
assign addr[62745]= -2082951896;
assign addr[62746]= -1987655498;
assign addr[62747]= -1852079154;
assign addr[62748]= -1678970324;
assign addr[62749]= -1471837070;
assign addr[62750]= -1234876957;
assign addr[62751]= -972891995;
assign addr[62752]= -691191324;
assign addr[62753]= -395483624;
assign addr[62754]= -91761426;
assign addr[62755]= 213820322;
assign addr[62756]= 515068990;
assign addr[62757]= 805879757;
assign addr[62758]= 1080359326;
assign addr[62759]= 1332945355;
assign addr[62760]= 1558519173;
assign addr[62761]= 1752509516;
assign addr[62762]= 1910985158;
assign addr[62763]= 2030734582;
assign addr[62764]= 2109331059;
assign addr[62765]= 2145181827;
assign addr[62766]= 2137560369;
assign addr[62767]= 2086621133;
assign addr[62768]= 1993396407;
assign addr[62769]= 1859775393;
assign addr[62770]= 1688465931;
assign addr[62771]= 1482939614;
assign addr[62772]= 1247361445;
assign addr[62773]= 986505429;
assign addr[62774]= 705657826;
assign addr[62775]= 410510029;
assign addr[62776]= 107043224;
assign addr[62777]= -198592817;
assign addr[62778]= -500204365;
assign addr[62779]= -791679244;
assign addr[62780]= -1067110699;
assign addr[62781]= -1320917099;
assign addr[62782]= -1547955041;
assign addr[62783]= -1743623590;
assign addr[62784]= -1903957513;
assign addr[62785]= -2025707632;
assign addr[62786]= -2106406677;
assign addr[62787]= -2144419275;
assign addr[62788]= -2138975100;
assign addr[62789]= -2090184478;
assign addr[62790]= -1999036154;
assign addr[62791]= -1867377253;
assign addr[62792]= -1697875851;
assign addr[62793]= -1493966902;
assign addr[62794]= -1259782632;
assign addr[62795]= -1000068799;
assign addr[62796]= -720088517;
assign addr[62797]= -425515602;
assign addr[62798]= -122319591;
assign addr[62799]= 183355234;
assign addr[62800]= 485314355;
assign addr[62801]= 777438554;
assign addr[62802]= 1053807919;
assign addr[62803]= 1308821808;
assign addr[62804]= 1537312353;
assign addr[62805]= 1734649179;
assign addr[62806]= 1896833245;
assign addr[62807]= 2020577882;
assign addr[62808]= 2103375398;
assign addr[62809]= 2143547897;
assign addr[62810]= 2140281282;
assign addr[62811]= 2093641749;
assign addr[62812]= 2004574453;
assign addr[62813]= 1874884346;
assign addr[62814]= 1707199606;
assign addr[62815]= 1504918373;
assign addr[62816]= 1272139887;
assign addr[62817]= 1013581418;
assign addr[62818]= 734482665;
assign addr[62819]= 440499581;
assign addr[62820]= 137589750;
assign addr[62821]= -168108346;
assign addr[62822]= -470399716;
assign addr[62823]= -763158411;
assign addr[62824]= -1040451659;
assign addr[62825]= -1296660098;
assign addr[62826]= -1526591649;
assign addr[62827]= -1725586737;
assign addr[62828]= -1889612716;
assign addr[62829]= -2015345591;
assign addr[62830]= -2100237377;
assign addr[62831]= -2142567738;
assign addr[62832]= -2141478848;
assign addr[62833]= -2096992772;
assign addr[62834]= -2010011024;
assign addr[62835]= -1882296293;
assign addr[62836]= -1716436725;
assign addr[62837]= -1515793473;
assign addr[62838]= -1284432584;
assign addr[62839]= -1027042599;
assign addr[62840]= -748839539;
assign addr[62841]= -455461206;
assign addr[62842]= -152852926;
assign addr[62843]= 152852926;
assign addr[62844]= 455461206;
assign addr[62845]= 748839539;
assign addr[62846]= 1027042599;
assign addr[62847]= 1284432584;
assign addr[62848]= 1515793473;
assign addr[62849]= 1716436725;
assign addr[62850]= 1882296293;
assign addr[62851]= 2010011024;
assign addr[62852]= 2096992772;
assign addr[62853]= 2141478848;
assign addr[62854]= 2142567738;
assign addr[62855]= 2100237377;
assign addr[62856]= 2015345591;
assign addr[62857]= 1889612716;
assign addr[62858]= 1725586737;
assign addr[62859]= 1526591649;
assign addr[62860]= 1296660098;
assign addr[62861]= 1040451659;
assign addr[62862]= 763158411;
assign addr[62863]= 470399716;
assign addr[62864]= 168108346;
assign addr[62865]= -137589750;
assign addr[62866]= -440499581;
assign addr[62867]= -734482665;
assign addr[62868]= -1013581418;
assign addr[62869]= -1272139887;
assign addr[62870]= -1504918373;
assign addr[62871]= -1707199606;
assign addr[62872]= -1874884346;
assign addr[62873]= -2004574453;
assign addr[62874]= -2093641749;
assign addr[62875]= -2140281282;
assign addr[62876]= -2143547897;
assign addr[62877]= -2103375398;
assign addr[62878]= -2020577882;
assign addr[62879]= -1896833245;
assign addr[62880]= -1734649179;
assign addr[62881]= -1537312353;
assign addr[62882]= -1308821808;
assign addr[62883]= -1053807919;
assign addr[62884]= -777438554;
assign addr[62885]= -485314355;
assign addr[62886]= -183355234;
assign addr[62887]= 122319591;
assign addr[62888]= 425515602;
assign addr[62889]= 720088517;
assign addr[62890]= 1000068799;
assign addr[62891]= 1259782632;
assign addr[62892]= 1493966902;
assign addr[62893]= 1697875851;
assign addr[62894]= 1867377253;
assign addr[62895]= 1999036154;
assign addr[62896]= 2090184478;
assign addr[62897]= 2138975100;
assign addr[62898]= 2144419275;
assign addr[62899]= 2106406677;
assign addr[62900]= 2025707632;
assign addr[62901]= 1903957513;
assign addr[62902]= 1743623590;
assign addr[62903]= 1547955041;
assign addr[62904]= 1320917099;
assign addr[62905]= 1067110699;
assign addr[62906]= 791679244;
assign addr[62907]= 500204365;
assign addr[62908]= 198592817;
assign addr[62909]= -107043224;
assign addr[62910]= -410510029;
assign addr[62911]= -705657826;
assign addr[62912]= -986505429;
assign addr[62913]= -1247361445;
assign addr[62914]= -1482939614;
assign addr[62915]= -1688465931;
assign addr[62916]= -1859775393;
assign addr[62917]= -1993396407;
assign addr[62918]= -2086621133;
assign addr[62919]= -2137560369;
assign addr[62920]= -2145181827;
assign addr[62921]= -2109331059;
assign addr[62922]= -2030734582;
assign addr[62923]= -1910985158;
assign addr[62924]= -1752509516;
assign addr[62925]= -1558519173;
assign addr[62926]= -1332945355;
assign addr[62927]= -1080359326;
assign addr[62928]= -805879757;
assign addr[62929]= -515068990;
assign addr[62930]= -213820322;
assign addr[62931]= 91761426;
assign addr[62932]= 395483624;
assign addr[62933]= 691191324;
assign addr[62934]= 972891995;
assign addr[62935]= 1234876957;
assign addr[62936]= 1471837070;
assign addr[62937]= 1678970324;
assign addr[62938]= 1852079154;
assign addr[62939]= 1987655498;
assign addr[62940]= 2082951896;
assign addr[62941]= 2136037160;
assign addr[62942]= 2145835515;
assign addr[62943]= 2112148396;
assign addr[62944]= 2035658475;
assign addr[62945]= 1917915825;
assign addr[62946]= 1761306505;
assign addr[62947]= 1569004214;
assign addr[62948]= 1344905966;
assign addr[62949]= 1093553126;
assign addr[62950]= 820039373;
assign addr[62951]= 529907477;
assign addr[62952]= 229036977;
assign addr[62953]= -76474970;
assign addr[62954]= -380437148;
assign addr[62955]= -676689746;
assign addr[62956]= -959229189;
assign addr[62957]= -1222329801;
assign addr[62958]= -1460659832;
assign addr[62959]= -1669389513;
assign addr[62960]= -1844288924;
assign addr[62961]= -1981813720;
assign addr[62962]= -2079176953;
assign addr[62963]= -2134405552;
assign addr[62964]= -2146380306;
assign addr[62965]= -2114858546;
assign addr[62966]= -2040479063;
assign addr[62967]= -1924749160;
assign addr[62968]= -1770014111;
assign addr[62969]= -1579409630;
assign addr[62970]= -1356798326;
assign addr[62971]= -1106691431;
assign addr[62972]= -834157373;
assign addr[62973]= -544719071;
assign addr[62974]= -244242007;
assign addr[62975]= 61184634;
assign addr[62976]= 365371365;
assign addr[62977]= 662153826;
assign addr[62978]= 945517704;
assign addr[62979]= 1209720613;
assign addr[62980]= 1449408469;
assign addr[62981]= 1659723983;
assign addr[62982]= 1836405100;
assign addr[62983]= 1975871368;
assign addr[62984]= 2075296495;
assign addr[62985]= 2132665626;
assign addr[62986]= 2146816171;
assign addr[62987]= 2117461370;
assign addr[62988]= 2045196100;
assign addr[62989]= 1931484818;
assign addr[62990]= 1778631892;
assign addr[62991]= 1589734894;
assign addr[62992]= 1368621831;
assign addr[62993]= 1119773573;
assign addr[62994]= 848233042;
assign addr[62995]= 559503022;
assign addr[62996]= 259434643;
assign addr[62997]= -45891193;
assign addr[62998]= -350287041;
assign addr[62999]= -647584304;
assign addr[63000]= -931758235;
assign addr[63001]= -1197050035;
assign addr[63002]= -1438083551;
assign addr[63003]= -1649974225;
assign addr[63004]= -1828428082;
assign addr[63005]= -1969828744;
assign addr[63006]= -2071310720;
assign addr[63007]= -2130817471;
assign addr[63008]= -2147143090;
assign addr[63009]= -2119956737;
assign addr[63010]= -2049809346;
assign addr[63011]= -1938122457;
assign addr[63012]= -1787159411;
assign addr[63013]= -1599979481;
assign addr[63014]= -1380375881;
assign addr[63015]= -1132798888;
assign addr[63016]= -862265664;
assign addr[63017]= -574258580;
assign addr[63018]= -274614114;
assign addr[63019]= 30595422;
assign addr[63020]= 335184940;
assign addr[63021]= 632981917;
assign addr[63022]= 917951481;
assign addr[63023]= 1184318708;
assign addr[63024]= 1426685652;
assign addr[63025]= 1640140734;
assign addr[63026]= 1820358275;
assign addr[63027]= 1963686155;
assign addr[63028]= 2067219829;
assign addr[63029]= 2128861181;
assign addr[63030]= 2147361045;
assign addr[63031]= 2122344521;
assign addr[63032]= 2054318569;
assign addr[63033]= 1944661739;
assign addr[63034]= 1795596234;
assign addr[63035]= 1610142873;
assign addr[63036]= 1392059879;
assign addr[63037]= 1145766716;
assign addr[63038]= 876254528;
assign addr[63039]= 588984994;
assign addr[63040]= 289779648;
assign addr[63041]= -15298099;
assign addr[63042]= -320065829;
assign addr[63043]= -618347408;
assign addr[63044]= -904098143;
assign addr[63045]= -1171527280;
assign addr[63046]= -1415215352;
assign addr[63047]= -1630224009;
assign addr[63048]= -1812196087;
assign addr[63049]= -1957443913;
assign addr[63050]= -2063024031;
assign addr[63051]= -2126796855;
assign addr[63052]= -2147470025;
assign addr[63053]= -2124624598;
assign addr[63054]= -2058723538;
assign addr[63055]= -1951102334;
assign addr[63056]= -1803941934;
assign addr[63057]= -1620224553;
assign addr[63058]= -1403673233;
assign addr[63059]= -1158676398;
assign addr[63060]= -890198924;
assign addr[63061]= -603681519;
assign addr[63062]= -304930476;
assign addr[63063]= 0;
assign addr[63064]= 304930476;
assign addr[63065]= 603681519;
assign addr[63066]= 890198924;
assign addr[63067]= 1158676398;
assign addr[63068]= 1403673233;
assign addr[63069]= 1620224553;
assign addr[63070]= 1803941934;
assign addr[63071]= 1951102334;
assign addr[63072]= 2058723538;
assign addr[63073]= 2124624598;
assign addr[63074]= 2147470025;
assign addr[63075]= 2126796855;
assign addr[63076]= 2063024031;
assign addr[63077]= 1957443913;
assign addr[63078]= 1812196087;
assign addr[63079]= 1630224009;
assign addr[63080]= 1415215352;
assign addr[63081]= 1171527280;
assign addr[63082]= 904098143;
assign addr[63083]= 618347408;
assign addr[63084]= 320065829;
assign addr[63085]= 15298099;
assign addr[63086]= -289779648;
assign addr[63087]= -588984994;
assign addr[63088]= -876254528;
assign addr[63089]= -1145766716;
assign addr[63090]= -1392059879;
assign addr[63091]= -1610142873;
assign addr[63092]= -1795596234;
assign addr[63093]= -1944661739;
assign addr[63094]= -2054318569;
assign addr[63095]= -2122344521;
assign addr[63096]= -2147361045;
assign addr[63097]= -2128861181;
assign addr[63098]= -2067219829;
assign addr[63099]= -1963686155;
assign addr[63100]= -1820358275;
assign addr[63101]= -1640140734;
assign addr[63102]= -1426685652;
assign addr[63103]= -1184318708;
assign addr[63104]= -917951481;
assign addr[63105]= -632981917;
assign addr[63106]= -335184940;
assign addr[63107]= -30595422;
assign addr[63108]= 274614114;
assign addr[63109]= 574258580;
assign addr[63110]= 862265664;
assign addr[63111]= 1132798888;
assign addr[63112]= 1380375881;
assign addr[63113]= 1599979481;
assign addr[63114]= 1787159411;
assign addr[63115]= 1938122457;
assign addr[63116]= 2049809346;
assign addr[63117]= 2119956737;
assign addr[63118]= 2147143090;
assign addr[63119]= 2130817471;
assign addr[63120]= 2071310720;
assign addr[63121]= 1969828744;
assign addr[63122]= 1828428082;
assign addr[63123]= 1649974225;
assign addr[63124]= 1438083551;
assign addr[63125]= 1197050035;
assign addr[63126]= 931758235;
assign addr[63127]= 647584304;
assign addr[63128]= 350287041;
assign addr[63129]= 45891193;
assign addr[63130]= -259434643;
assign addr[63131]= -559503022;
assign addr[63132]= -848233042;
assign addr[63133]= -1119773573;
assign addr[63134]= -1368621831;
assign addr[63135]= -1589734894;
assign addr[63136]= -1778631892;
assign addr[63137]= -1931484818;
assign addr[63138]= -2045196100;
assign addr[63139]= -2117461370;
assign addr[63140]= -2146816171;
assign addr[63141]= -2132665626;
assign addr[63142]= -2075296495;
assign addr[63143]= -1975871368;
assign addr[63144]= -1836405100;
assign addr[63145]= -1659723983;
assign addr[63146]= -1449408469;
assign addr[63147]= -1209720613;
assign addr[63148]= -945517704;
assign addr[63149]= -662153826;
assign addr[63150]= -365371365;
assign addr[63151]= -61184634;
assign addr[63152]= 244242007;
assign addr[63153]= 544719071;
assign addr[63154]= 834157373;
assign addr[63155]= 1106691431;
assign addr[63156]= 1356798326;
assign addr[63157]= 1579409630;
assign addr[63158]= 1770014111;
assign addr[63159]= 1924749160;
assign addr[63160]= 2040479063;
assign addr[63161]= 2114858546;
assign addr[63162]= 2146380306;
assign addr[63163]= 2134405552;
assign addr[63164]= 2079176953;
assign addr[63165]= 1981813720;
assign addr[63166]= 1844288924;
assign addr[63167]= 1669389513;
assign addr[63168]= 1460659832;
assign addr[63169]= 1222329801;
assign addr[63170]= 959229189;
assign addr[63171]= 676689746;
assign addr[63172]= 380437148;
assign addr[63173]= 76474970;
assign addr[63174]= -229036977;
assign addr[63175]= -529907477;
assign addr[63176]= -820039373;
assign addr[63177]= -1093553126;
assign addr[63178]= -1344905966;
assign addr[63179]= -1569004214;
assign addr[63180]= -1761306505;
assign addr[63181]= -1917915825;
assign addr[63182]= -2035658475;
assign addr[63183]= -2112148396;
assign addr[63184]= -2145835515;
assign addr[63185]= -2136037160;
assign addr[63186]= -2082951896;
assign addr[63187]= -1987655498;
assign addr[63188]= -1852079154;
assign addr[63189]= -1678970324;
assign addr[63190]= -1471837070;
assign addr[63191]= -1234876957;
assign addr[63192]= -972891995;
assign addr[63193]= -691191324;
assign addr[63194]= -395483624;
assign addr[63195]= -91761426;
assign addr[63196]= 213820322;
assign addr[63197]= 515068990;
assign addr[63198]= 805879757;
assign addr[63199]= 1080359326;
assign addr[63200]= 1332945355;
assign addr[63201]= 1558519173;
assign addr[63202]= 1752509516;
assign addr[63203]= 1910985158;
assign addr[63204]= 2030734582;
assign addr[63205]= 2109331059;
assign addr[63206]= 2145181827;
assign addr[63207]= 2137560369;
assign addr[63208]= 2086621133;
assign addr[63209]= 1993396407;
assign addr[63210]= 1859775393;
assign addr[63211]= 1688465931;
assign addr[63212]= 1482939614;
assign addr[63213]= 1247361445;
assign addr[63214]= 986505429;
assign addr[63215]= 705657826;
assign addr[63216]= 410510029;
assign addr[63217]= 107043224;
assign addr[63218]= -198592817;
assign addr[63219]= -500204365;
assign addr[63220]= -791679244;
assign addr[63221]= -1067110699;
assign addr[63222]= -1320917099;
assign addr[63223]= -1547955041;
assign addr[63224]= -1743623590;
assign addr[63225]= -1903957513;
assign addr[63226]= -2025707632;
assign addr[63227]= -2106406677;
assign addr[63228]= -2144419275;
assign addr[63229]= -2138975100;
assign addr[63230]= -2090184478;
assign addr[63231]= -1999036154;
assign addr[63232]= -1867377253;
assign addr[63233]= -1697875851;
assign addr[63234]= -1493966902;
assign addr[63235]= -1259782632;
assign addr[63236]= -1000068799;
assign addr[63237]= -720088517;
assign addr[63238]= -425515602;
assign addr[63239]= -122319591;
assign addr[63240]= 183355234;
assign addr[63241]= 485314355;
assign addr[63242]= 777438554;
assign addr[63243]= 1053807919;
assign addr[63244]= 1308821808;
assign addr[63245]= 1537312353;
assign addr[63246]= 1734649179;
assign addr[63247]= 1896833245;
assign addr[63248]= 2020577882;
assign addr[63249]= 2103375398;
assign addr[63250]= 2143547897;
assign addr[63251]= 2140281282;
assign addr[63252]= 2093641749;
assign addr[63253]= 2004574453;
assign addr[63254]= 1874884346;
assign addr[63255]= 1707199606;
assign addr[63256]= 1504918373;
assign addr[63257]= 1272139887;
assign addr[63258]= 1013581418;
assign addr[63259]= 734482665;
assign addr[63260]= 440499581;
assign addr[63261]= 137589750;
assign addr[63262]= -168108346;
assign addr[63263]= -470399716;
assign addr[63264]= -763158411;
assign addr[63265]= -1040451659;
assign addr[63266]= -1296660098;
assign addr[63267]= -1526591649;
assign addr[63268]= -1725586737;
assign addr[63269]= -1889612716;
assign addr[63270]= -2015345591;
assign addr[63271]= -2100237377;
assign addr[63272]= -2142567738;
assign addr[63273]= -2141478848;
assign addr[63274]= -2096992772;
assign addr[63275]= -2010011024;
assign addr[63276]= -1882296293;
assign addr[63277]= -1716436725;
assign addr[63278]= -1515793473;
assign addr[63279]= -1284432584;
assign addr[63280]= -1027042599;
assign addr[63281]= -748839539;
assign addr[63282]= -455461206;
assign addr[63283]= -152852926;
assign addr[63284]= 152852926;
assign addr[63285]= 455461206;
assign addr[63286]= 748839539;
assign addr[63287]= 1027042599;
assign addr[63288]= 1284432584;
assign addr[63289]= 1515793473;
assign addr[63290]= 1716436725;
assign addr[63291]= 1882296293;
assign addr[63292]= 2010011024;
assign addr[63293]= 2096992772;
assign addr[63294]= 2141478848;
assign addr[63295]= 2142567738;
assign addr[63296]= 2100237377;
assign addr[63297]= 2015345591;
assign addr[63298]= 1889612716;
assign addr[63299]= 1725586737;
assign addr[63300]= 1526591649;
assign addr[63301]= 1296660098;
assign addr[63302]= 1040451659;
assign addr[63303]= 763158411;
assign addr[63304]= 470399716;
assign addr[63305]= 168108346;
assign addr[63306]= -137589750;
assign addr[63307]= -440499581;
assign addr[63308]= -734482665;
assign addr[63309]= -1013581418;
assign addr[63310]= -1272139887;
assign addr[63311]= -1504918373;
assign addr[63312]= -1707199606;
assign addr[63313]= -1874884346;
assign addr[63314]= -2004574453;
assign addr[63315]= -2093641749;
assign addr[63316]= -2140281282;
assign addr[63317]= -2143547897;
assign addr[63318]= -2103375398;
assign addr[63319]= -2020577882;
assign addr[63320]= -1896833245;
assign addr[63321]= -1734649179;
assign addr[63322]= -1537312353;
assign addr[63323]= -1308821808;
assign addr[63324]= -1053807919;
assign addr[63325]= -777438554;
assign addr[63326]= -485314355;
assign addr[63327]= -183355234;
assign addr[63328]= 122319591;
assign addr[63329]= 425515602;
assign addr[63330]= 720088517;
assign addr[63331]= 1000068799;
assign addr[63332]= 1259782632;
assign addr[63333]= 1493966902;
assign addr[63334]= 1697875851;
assign addr[63335]= 1867377253;
assign addr[63336]= 1999036154;
assign addr[63337]= 2090184478;
assign addr[63338]= 2138975100;
assign addr[63339]= 2144419275;
assign addr[63340]= 2106406677;
assign addr[63341]= 2025707632;
assign addr[63342]= 1903957513;
assign addr[63343]= 1743623590;
assign addr[63344]= 1547955041;
assign addr[63345]= 1320917099;
assign addr[63346]= 1067110699;
assign addr[63347]= 791679244;
assign addr[63348]= 500204365;
assign addr[63349]= 198592817;
assign addr[63350]= -107043224;
assign addr[63351]= -410510029;
assign addr[63352]= -705657826;
assign addr[63353]= -986505429;
assign addr[63354]= -1247361445;
assign addr[63355]= -1482939614;
assign addr[63356]= -1688465931;
assign addr[63357]= -1859775393;
assign addr[63358]= -1993396407;
assign addr[63359]= -2086621133;
assign addr[63360]= -2137560369;
assign addr[63361]= -2145181827;
assign addr[63362]= -2109331059;
assign addr[63363]= -2030734582;
assign addr[63364]= -1910985158;
assign addr[63365]= -1752509516;
assign addr[63366]= -1558519173;
assign addr[63367]= -1332945355;
assign addr[63368]= -1080359326;
assign addr[63369]= -805879757;
assign addr[63370]= -515068990;
assign addr[63371]= -213820322;
assign addr[63372]= 91761426;
assign addr[63373]= 395483624;
assign addr[63374]= 691191324;
assign addr[63375]= 972891995;
assign addr[63376]= 1234876957;
assign addr[63377]= 1471837070;
assign addr[63378]= 1678970324;
assign addr[63379]= 1852079154;
assign addr[63380]= 1987655498;
assign addr[63381]= 2082951896;
assign addr[63382]= 2136037160;
assign addr[63383]= 2145835515;
assign addr[63384]= 2112148396;
assign addr[63385]= 2035658475;
assign addr[63386]= 1917915825;
assign addr[63387]= 1761306505;
assign addr[63388]= 1569004214;
assign addr[63389]= 1344905966;
assign addr[63390]= 1093553126;
assign addr[63391]= 820039373;
assign addr[63392]= 529907477;
assign addr[63393]= 229036977;
assign addr[63394]= -76474970;
assign addr[63395]= -380437148;
assign addr[63396]= -676689746;
assign addr[63397]= -959229189;
assign addr[63398]= -1222329801;
assign addr[63399]= -1460659832;
assign addr[63400]= -1669389513;
assign addr[63401]= -1844288924;
assign addr[63402]= -1981813720;
assign addr[63403]= -2079176953;
assign addr[63404]= -2134405552;
assign addr[63405]= -2146380306;
assign addr[63406]= -2114858546;
assign addr[63407]= -2040479063;
assign addr[63408]= -1924749160;
assign addr[63409]= -1770014111;
assign addr[63410]= -1579409630;
assign addr[63411]= -1356798326;
assign addr[63412]= -1106691431;
assign addr[63413]= -834157373;
assign addr[63414]= -544719071;
assign addr[63415]= -244242007;
assign addr[63416]= 61184634;
assign addr[63417]= 365371365;
assign addr[63418]= 662153826;
assign addr[63419]= 945517704;
assign addr[63420]= 1209720613;
assign addr[63421]= 1449408469;
assign addr[63422]= 1659723983;
assign addr[63423]= 1836405100;
assign addr[63424]= 1975871368;
assign addr[63425]= 2075296495;
assign addr[63426]= 2132665626;
assign addr[63427]= 2146816171;
assign addr[63428]= 2117461370;
assign addr[63429]= 2045196100;
assign addr[63430]= 1931484818;
assign addr[63431]= 1778631892;
assign addr[63432]= 1589734894;
assign addr[63433]= 1368621831;
assign addr[63434]= 1119773573;
assign addr[63435]= 848233042;
assign addr[63436]= 559503022;
assign addr[63437]= 259434643;
assign addr[63438]= -45891193;
assign addr[63439]= -350287041;
assign addr[63440]= -647584304;
assign addr[63441]= -931758235;
assign addr[63442]= -1197050035;
assign addr[63443]= -1438083551;
assign addr[63444]= -1649974225;
assign addr[63445]= -1828428082;
assign addr[63446]= -1969828744;
assign addr[63447]= -2071310720;
assign addr[63448]= -2130817471;
assign addr[63449]= -2147143090;
assign addr[63450]= -2119956737;
assign addr[63451]= -2049809346;
assign addr[63452]= -1938122457;
assign addr[63453]= -1787159411;
assign addr[63454]= -1599979481;
assign addr[63455]= -1380375881;
assign addr[63456]= -1132798888;
assign addr[63457]= -862265664;
assign addr[63458]= -574258580;
assign addr[63459]= -274614114;
assign addr[63460]= 30595422;
assign addr[63461]= 335184940;
assign addr[63462]= 632981917;
assign addr[63463]= 917951481;
assign addr[63464]= 1184318708;
assign addr[63465]= 1426685652;
assign addr[63466]= 1640140734;
assign addr[63467]= 1820358275;
assign addr[63468]= 1963686155;
assign addr[63469]= 2067219829;
assign addr[63470]= 2128861181;
assign addr[63471]= 2147361045;
assign addr[63472]= 2122344521;
assign addr[63473]= 2054318569;
assign addr[63474]= 1944661739;
assign addr[63475]= 1795596234;
assign addr[63476]= 1610142873;
assign addr[63477]= 1392059879;
assign addr[63478]= 1145766716;
assign addr[63479]= 876254528;
assign addr[63480]= 588984994;
assign addr[63481]= 289779648;
assign addr[63482]= -15298099;
assign addr[63483]= -320065829;
assign addr[63484]= -618347408;
assign addr[63485]= -904098143;
assign addr[63486]= -1171527280;
assign addr[63487]= -1415215352;
assign addr[63488]= -1630224009;
assign addr[63489]= -1812196087;
assign addr[63490]= -1957443913;
assign addr[63491]= -2063024031;
assign addr[63492]= -2126796855;
assign addr[63493]= -2147470025;
assign addr[63494]= -2124624598;
assign addr[63495]= -2058723538;
assign addr[63496]= -1951102334;
assign addr[63497]= -1803941934;
assign addr[63498]= -1620224553;
assign addr[63499]= -1403673233;
assign addr[63500]= -1158676398;
assign addr[63501]= -890198924;
assign addr[63502]= -603681519;
assign addr[63503]= -304930476;
assign addr[63504]= 0;
assign addr[63505]= 304930476;
assign addr[63506]= 603681519;
assign addr[63507]= 890198924;
assign addr[63508]= 1158676398;
assign addr[63509]= 1403673233;
assign addr[63510]= 1620224553;
assign addr[63511]= 1803941934;
assign addr[63512]= 1951102334;
assign addr[63513]= 2058723538;
assign addr[63514]= 2124624598;
assign addr[63515]= 2147470025;
assign addr[63516]= 2126796855;
assign addr[63517]= 2063024031;
assign addr[63518]= 1957443913;
assign addr[63519]= 1812196087;
assign addr[63520]= 1630224009;
assign addr[63521]= 1415215352;
assign addr[63522]= 1171527280;
assign addr[63523]= 904098143;
assign addr[63524]= 618347408;
assign addr[63525]= 320065829;
assign addr[63526]= 15298099;
assign addr[63527]= -289779648;
assign addr[63528]= -588984994;
assign addr[63529]= -876254528;
assign addr[63530]= -1145766716;
assign addr[63531]= -1392059879;
assign addr[63532]= -1610142873;
assign addr[63533]= -1795596234;
assign addr[63534]= -1944661739;
assign addr[63535]= -2054318569;
assign addr[63536]= -2122344521;
assign addr[63537]= -2147361045;
assign addr[63538]= -2128861181;
assign addr[63539]= -2067219829;
assign addr[63540]= -1963686155;
assign addr[63541]= -1820358275;
assign addr[63542]= -1640140734;
assign addr[63543]= -1426685652;
assign addr[63544]= -1184318708;
assign addr[63545]= -917951481;
assign addr[63546]= -632981917;
assign addr[63547]= -335184940;
assign addr[63548]= -30595422;
assign addr[63549]= 274614114;
assign addr[63550]= 574258580;
assign addr[63551]= 862265664;
assign addr[63552]= 1132798888;
assign addr[63553]= 1380375881;
assign addr[63554]= 1599979481;
assign addr[63555]= 1787159411;
assign addr[63556]= 1938122457;
assign addr[63557]= 2049809346;
assign addr[63558]= 2119956737;
assign addr[63559]= 2147143090;
assign addr[63560]= 2130817471;
assign addr[63561]= 2071310720;
assign addr[63562]= 1969828744;
assign addr[63563]= 1828428082;
assign addr[63564]= 1649974225;
assign addr[63565]= 1438083551;
assign addr[63566]= 1197050035;
assign addr[63567]= 931758235;
assign addr[63568]= 647584304;
assign addr[63569]= 350287041;
assign addr[63570]= 45891193;
assign addr[63571]= -259434643;
assign addr[63572]= -559503022;
assign addr[63573]= -848233042;
assign addr[63574]= -1119773573;
assign addr[63575]= -1368621831;
assign addr[63576]= -1589734894;
assign addr[63577]= -1778631892;
assign addr[63578]= -1931484818;
assign addr[63579]= -2045196100;
assign addr[63580]= -2117461370;
assign addr[63581]= -2146816171;
assign addr[63582]= -2132665626;
assign addr[63583]= -2075296495;
assign addr[63584]= -1975871368;
assign addr[63585]= -1836405100;
assign addr[63586]= -1659723983;
assign addr[63587]= -1449408469;
assign addr[63588]= -1209720613;
assign addr[63589]= -945517704;
assign addr[63590]= -662153826;
assign addr[63591]= -365371365;
assign addr[63592]= -61184634;
assign addr[63593]= 244242007;
assign addr[63594]= 544719071;
assign addr[63595]= 834157373;
assign addr[63596]= 1106691431;
assign addr[63597]= 1356798326;
assign addr[63598]= 1579409630;
assign addr[63599]= 1770014111;
assign addr[63600]= 1924749160;
assign addr[63601]= 2040479063;
assign addr[63602]= 2114858546;
assign addr[63603]= 2146380306;
assign addr[63604]= 2134405552;
assign addr[63605]= 2079176953;
assign addr[63606]= 1981813720;
assign addr[63607]= 1844288924;
assign addr[63608]= 1669389513;
assign addr[63609]= 1460659832;
assign addr[63610]= 1222329801;
assign addr[63611]= 959229189;
assign addr[63612]= 676689746;
assign addr[63613]= 380437148;
assign addr[63614]= 76474970;
assign addr[63615]= -229036977;
assign addr[63616]= -529907477;
assign addr[63617]= -820039373;
assign addr[63618]= -1093553126;
assign addr[63619]= -1344905966;
assign addr[63620]= -1569004214;
assign addr[63621]= -1761306505;
assign addr[63622]= -1917915825;
assign addr[63623]= -2035658475;
assign addr[63624]= -2112148396;
assign addr[63625]= -2145835515;
assign addr[63626]= -2136037160;
assign addr[63627]= -2082951896;
assign addr[63628]= -1987655498;
assign addr[63629]= -1852079154;
assign addr[63630]= -1678970324;
assign addr[63631]= -1471837070;
assign addr[63632]= -1234876957;
assign addr[63633]= -972891995;
assign addr[63634]= -691191324;
assign addr[63635]= -395483624;
assign addr[63636]= -91761426;
assign addr[63637]= 213820322;
assign addr[63638]= 515068990;
assign addr[63639]= 805879757;
assign addr[63640]= 1080359326;
assign addr[63641]= 1332945355;
assign addr[63642]= 1558519173;
assign addr[63643]= 1752509516;
assign addr[63644]= 1910985158;
assign addr[63645]= 2030734582;
assign addr[63646]= 2109331059;
assign addr[63647]= 2145181827;
assign addr[63648]= 2137560369;
assign addr[63649]= 2086621133;
assign addr[63650]= 1993396407;
assign addr[63651]= 1859775393;
assign addr[63652]= 1688465931;
assign addr[63653]= 1482939614;
assign addr[63654]= 1247361445;
assign addr[63655]= 986505429;
assign addr[63656]= 705657826;
assign addr[63657]= 410510029;
assign addr[63658]= 107043224;
assign addr[63659]= -198592817;
assign addr[63660]= -500204365;
assign addr[63661]= -791679244;
assign addr[63662]= -1067110699;
assign addr[63663]= -1320917099;
assign addr[63664]= -1547955041;
assign addr[63665]= -1743623590;
assign addr[63666]= -1903957513;
assign addr[63667]= -2025707632;
assign addr[63668]= -2106406677;
assign addr[63669]= -2144419275;
assign addr[63670]= -2138975100;
assign addr[63671]= -2090184478;
assign addr[63672]= -1999036154;
assign addr[63673]= -1867377253;
assign addr[63674]= -1697875851;
assign addr[63675]= -1493966902;
assign addr[63676]= -1259782632;
assign addr[63677]= -1000068799;
assign addr[63678]= -720088517;
assign addr[63679]= -425515602;
assign addr[63680]= -122319591;
assign addr[63681]= 183355234;
assign addr[63682]= 485314355;
assign addr[63683]= 777438554;
assign addr[63684]= 1053807919;
assign addr[63685]= 1308821808;
assign addr[63686]= 1537312353;
assign addr[63687]= 1734649179;
assign addr[63688]= 1896833245;
assign addr[63689]= 2020577882;
assign addr[63690]= 2103375398;
assign addr[63691]= 2143547897;
assign addr[63692]= 2140281282;
assign addr[63693]= 2093641749;
assign addr[63694]= 2004574453;
assign addr[63695]= 1874884346;
assign addr[63696]= 1707199606;
assign addr[63697]= 1504918373;
assign addr[63698]= 1272139887;
assign addr[63699]= 1013581418;
assign addr[63700]= 734482665;
assign addr[63701]= 440499581;
assign addr[63702]= 137589750;
assign addr[63703]= -168108346;
assign addr[63704]= -470399716;
assign addr[63705]= -763158411;
assign addr[63706]= -1040451659;
assign addr[63707]= -1296660098;
assign addr[63708]= -1526591649;
assign addr[63709]= -1725586737;
assign addr[63710]= -1889612716;
assign addr[63711]= -2015345591;
assign addr[63712]= -2100237377;
assign addr[63713]= -2142567738;
assign addr[63714]= -2141478848;
assign addr[63715]= -2096992772;
assign addr[63716]= -2010011024;
assign addr[63717]= -1882296293;
assign addr[63718]= -1716436725;
assign addr[63719]= -1515793473;
assign addr[63720]= -1284432584;
assign addr[63721]= -1027042599;
assign addr[63722]= -748839539;
assign addr[63723]= -455461206;
assign addr[63724]= -152852926;
assign addr[63725]= 152852926;
assign addr[63726]= 455461206;
assign addr[63727]= 748839539;
assign addr[63728]= 1027042599;
assign addr[63729]= 1284432584;
assign addr[63730]= 1515793473;
assign addr[63731]= 1716436725;
assign addr[63732]= 1882296293;
assign addr[63733]= 2010011024;
assign addr[63734]= 2096992772;
assign addr[63735]= 2141478848;
assign addr[63736]= 2142567738;
assign addr[63737]= 2100237377;
assign addr[63738]= 2015345591;
assign addr[63739]= 1889612716;
assign addr[63740]= 1725586737;
assign addr[63741]= 1526591649;
assign addr[63742]= 1296660098;
assign addr[63743]= 1040451659;
assign addr[63744]= 763158411;
assign addr[63745]= 470399716;
assign addr[63746]= 168108346;
assign addr[63747]= -137589750;
assign addr[63748]= -440499581;
assign addr[63749]= -734482665;
assign addr[63750]= -1013581418;
assign addr[63751]= -1272139887;
assign addr[63752]= -1504918373;
assign addr[63753]= -1707199606;
assign addr[63754]= -1874884346;
assign addr[63755]= -2004574453;
assign addr[63756]= -2093641749;
assign addr[63757]= -2140281282;
assign addr[63758]= -2143547897;
assign addr[63759]= -2103375398;
assign addr[63760]= -2020577882;
assign addr[63761]= -1896833245;
assign addr[63762]= -1734649179;
assign addr[63763]= -1537312353;
assign addr[63764]= -1308821808;
assign addr[63765]= -1053807919;
assign addr[63766]= -777438554;
assign addr[63767]= -485314355;
assign addr[63768]= -183355234;
assign addr[63769]= 122319591;
assign addr[63770]= 425515602;
assign addr[63771]= 720088517;
assign addr[63772]= 1000068799;
assign addr[63773]= 1259782632;
assign addr[63774]= 1493966902;
assign addr[63775]= 1697875851;
assign addr[63776]= 1867377253;
assign addr[63777]= 1999036154;
assign addr[63778]= 2090184478;
assign addr[63779]= 2138975100;
assign addr[63780]= 2144419275;
assign addr[63781]= 2106406677;
assign addr[63782]= 2025707632;
assign addr[63783]= 1903957513;
assign addr[63784]= 1743623590;
assign addr[63785]= 1547955041;
assign addr[63786]= 1320917099;
assign addr[63787]= 1067110699;
assign addr[63788]= 791679244;
assign addr[63789]= 500204365;
assign addr[63790]= 198592817;
assign addr[63791]= -107043224;
assign addr[63792]= -410510029;
assign addr[63793]= -705657826;
assign addr[63794]= -986505429;
assign addr[63795]= -1247361445;
assign addr[63796]= -1482939614;
assign addr[63797]= -1688465931;
assign addr[63798]= -1859775393;
assign addr[63799]= -1993396407;
assign addr[63800]= -2086621133;
assign addr[63801]= -2137560369;
assign addr[63802]= -2145181827;
assign addr[63803]= -2109331059;
assign addr[63804]= -2030734582;
assign addr[63805]= -1910985158;
assign addr[63806]= -1752509516;
assign addr[63807]= -1558519173;
assign addr[63808]= -1332945355;
assign addr[63809]= -1080359326;
assign addr[63810]= -805879757;
assign addr[63811]= -515068990;
assign addr[63812]= -213820322;
assign addr[63813]= 91761426;
assign addr[63814]= 395483624;
assign addr[63815]= 691191324;
assign addr[63816]= 972891995;
assign addr[63817]= 1234876957;
assign addr[63818]= 1471837070;
assign addr[63819]= 1678970324;
assign addr[63820]= 1852079154;
assign addr[63821]= 1987655498;
assign addr[63822]= 2082951896;
assign addr[63823]= 2136037160;
assign addr[63824]= 2145835515;
assign addr[63825]= 2112148396;
assign addr[63826]= 2035658475;
assign addr[63827]= 1917915825;
assign addr[63828]= 1761306505;
assign addr[63829]= 1569004214;
assign addr[63830]= 1344905966;
assign addr[63831]= 1093553126;
assign addr[63832]= 820039373;
assign addr[63833]= 529907477;
assign addr[63834]= 229036977;
assign addr[63835]= -76474970;
assign addr[63836]= -380437148;
assign addr[63837]= -676689746;
assign addr[63838]= -959229189;
assign addr[63839]= -1222329801;
assign addr[63840]= -1460659832;
assign addr[63841]= -1669389513;
assign addr[63842]= -1844288924;
assign addr[63843]= -1981813720;
assign addr[63844]= -2079176953;
assign addr[63845]= -2134405552;
assign addr[63846]= -2146380306;
assign addr[63847]= -2114858546;
assign addr[63848]= -2040479063;
assign addr[63849]= -1924749160;
assign addr[63850]= -1770014111;
assign addr[63851]= -1579409630;
assign addr[63852]= -1356798326;
assign addr[63853]= -1106691431;
assign addr[63854]= -834157373;
assign addr[63855]= -544719071;
assign addr[63856]= -244242007;
assign addr[63857]= 61184634;
assign addr[63858]= 365371365;
assign addr[63859]= 662153826;
assign addr[63860]= 945517704;
assign addr[63861]= 1209720613;
assign addr[63862]= 1449408469;
assign addr[63863]= 1659723983;
assign addr[63864]= 1836405100;
assign addr[63865]= 1975871368;
assign addr[63866]= 2075296495;
assign addr[63867]= 2132665626;
assign addr[63868]= 2146816171;
assign addr[63869]= 2117461370;
assign addr[63870]= 2045196100;
assign addr[63871]= 1931484818;
assign addr[63872]= 1778631892;
assign addr[63873]= 1589734894;
assign addr[63874]= 1368621831;
assign addr[63875]= 1119773573;
assign addr[63876]= 848233042;
assign addr[63877]= 559503022;
assign addr[63878]= 259434643;
assign addr[63879]= -45891193;
assign addr[63880]= -350287041;
assign addr[63881]= -647584304;
assign addr[63882]= -931758235;
assign addr[63883]= -1197050035;
assign addr[63884]= -1438083551;
assign addr[63885]= -1649974225;
assign addr[63886]= -1828428082;
assign addr[63887]= -1969828744;
assign addr[63888]= -2071310720;
assign addr[63889]= -2130817471;
assign addr[63890]= -2147143090;
assign addr[63891]= -2119956737;
assign addr[63892]= -2049809346;
assign addr[63893]= -1938122457;
assign addr[63894]= -1787159411;
assign addr[63895]= -1599979481;
assign addr[63896]= -1380375881;
assign addr[63897]= -1132798888;
assign addr[63898]= -862265664;
assign addr[63899]= -574258580;
assign addr[63900]= -274614114;
assign addr[63901]= 30595422;
assign addr[63902]= 335184940;
assign addr[63903]= 632981917;
assign addr[63904]= 917951481;
assign addr[63905]= 1184318708;
assign addr[63906]= 1426685652;
assign addr[63907]= 1640140734;
assign addr[63908]= 1820358275;
assign addr[63909]= 1963686155;
assign addr[63910]= 2067219829;
assign addr[63911]= 2128861181;
assign addr[63912]= 2147361045;
assign addr[63913]= 2122344521;
assign addr[63914]= 2054318569;
assign addr[63915]= 1944661739;
assign addr[63916]= 1795596234;
assign addr[63917]= 1610142873;
assign addr[63918]= 1392059879;
assign addr[63919]= 1145766716;
assign addr[63920]= 876254528;
assign addr[63921]= 588984994;
assign addr[63922]= 289779648;
assign addr[63923]= -15298099;
assign addr[63924]= -320065829;
assign addr[63925]= -618347408;
assign addr[63926]= -904098143;
assign addr[63927]= -1171527280;
assign addr[63928]= -1415215352;
assign addr[63929]= -1630224009;
assign addr[63930]= -1812196087;
assign addr[63931]= -1957443913;
assign addr[63932]= -2063024031;
assign addr[63933]= -2126796855;
assign addr[63934]= -2147470025;
assign addr[63935]= -2124624598;
assign addr[63936]= -2058723538;
assign addr[63937]= -1951102334;
assign addr[63938]= -1803941934;
assign addr[63939]= -1620224553;
assign addr[63940]= -1403673233;
assign addr[63941]= -1158676398;
assign addr[63942]= -890198924;
assign addr[63943]= -603681519;
assign addr[63944]= -304930476;
assign addr[63945]= 0;
assign addr[63946]= 304930476;
assign addr[63947]= 603681519;
assign addr[63948]= 890198924;
assign addr[63949]= 1158676398;
assign addr[63950]= 1403673233;
assign addr[63951]= 1620224553;
assign addr[63952]= 1803941934;
assign addr[63953]= 1951102334;
assign addr[63954]= 2058723538;
assign addr[63955]= 2124624598;
assign addr[63956]= 2147470025;
assign addr[63957]= 2126796855;
assign addr[63958]= 2063024031;
assign addr[63959]= 1957443913;
assign addr[63960]= 1812196087;
assign addr[63961]= 1630224009;
assign addr[63962]= 1415215352;
assign addr[63963]= 1171527280;
assign addr[63964]= 904098143;
assign addr[63965]= 618347408;
assign addr[63966]= 320065829;
assign addr[63967]= 15298099;
assign addr[63968]= -289779648;
assign addr[63969]= -588984994;
assign addr[63970]= -876254528;
assign addr[63971]= -1145766716;
assign addr[63972]= -1392059879;
assign addr[63973]= -1610142873;
assign addr[63974]= -1795596234;
assign addr[63975]= -1944661739;
assign addr[63976]= -2054318569;
assign addr[63977]= -2122344521;
assign addr[63978]= -2147361045;
assign addr[63979]= -2128861181;
assign addr[63980]= -2067219829;
assign addr[63981]= -1963686155;
assign addr[63982]= -1820358275;
assign addr[63983]= -1640140734;
assign addr[63984]= -1426685652;
assign addr[63985]= -1184318708;
assign addr[63986]= -917951481;
assign addr[63987]= -632981917;
assign addr[63988]= -335184940;
assign addr[63989]= -30595422;
assign addr[63990]= 274614114;
assign addr[63991]= 574258580;
assign addr[63992]= 862265664;
assign addr[63993]= 1132798888;
assign addr[63994]= 1380375881;
assign addr[63995]= 1599979481;
assign addr[63996]= 1787159411;
assign addr[63997]= 1938122457;
assign addr[63998]= 2049809346;
assign addr[63999]= 2119956737;
assign addr[64000]= 2147143090;
assign addr[64001]= 2130817471;
assign addr[64002]= 2071310720;
assign addr[64003]= 1969828744;
assign addr[64004]= 1828428082;
assign addr[64005]= 1649974225;
assign addr[64006]= 1438083551;
assign addr[64007]= 1197050035;
assign addr[64008]= 931758235;
assign addr[64009]= 647584304;
assign addr[64010]= 350287041;
assign addr[64011]= 45891193;
assign addr[64012]= -259434643;
assign addr[64013]= -559503022;
assign addr[64014]= -848233042;
assign addr[64015]= -1119773573;
assign addr[64016]= -1368621831;
assign addr[64017]= -1589734894;
assign addr[64018]= -1778631892;
assign addr[64019]= -1931484818;
assign addr[64020]= -2045196100;
assign addr[64021]= -2117461370;
assign addr[64022]= -2146816171;
assign addr[64023]= -2132665626;
assign addr[64024]= -2075296495;
assign addr[64025]= -1975871368;
assign addr[64026]= -1836405100;
assign addr[64027]= -1659723983;
assign addr[64028]= -1449408469;
assign addr[64029]= -1209720613;
assign addr[64030]= -945517704;
assign addr[64031]= -662153826;
assign addr[64032]= -365371365;
assign addr[64033]= -61184634;
assign addr[64034]= 244242007;
assign addr[64035]= 544719071;
assign addr[64036]= 834157373;
assign addr[64037]= 1106691431;
assign addr[64038]= 1356798326;
assign addr[64039]= 1579409630;
assign addr[64040]= 1770014111;
assign addr[64041]= 1924749160;
assign addr[64042]= 2040479063;
assign addr[64043]= 2114858546;
assign addr[64044]= 2146380306;
assign addr[64045]= 2134405552;
assign addr[64046]= 2079176953;
assign addr[64047]= 1981813720;
assign addr[64048]= 1844288924;
assign addr[64049]= 1669389513;
assign addr[64050]= 1460659832;
assign addr[64051]= 1222329801;
assign addr[64052]= 959229189;
assign addr[64053]= 676689746;
assign addr[64054]= 380437148;
assign addr[64055]= 76474970;
assign addr[64056]= -229036977;
assign addr[64057]= -529907477;
assign addr[64058]= -820039373;
assign addr[64059]= -1093553126;
assign addr[64060]= -1344905966;
assign addr[64061]= -1569004214;
assign addr[64062]= -1761306505;
assign addr[64063]= -1917915825;
assign addr[64064]= -2035658475;
assign addr[64065]= -2112148396;
assign addr[64066]= -2145835515;
assign addr[64067]= -2136037160;
assign addr[64068]= -2082951896;
assign addr[64069]= -1987655498;
assign addr[64070]= -1852079154;
assign addr[64071]= -1678970324;
assign addr[64072]= -1471837070;
assign addr[64073]= -1234876957;
assign addr[64074]= -972891995;
assign addr[64075]= -691191324;
assign addr[64076]= -395483624;
assign addr[64077]= -91761426;
assign addr[64078]= 213820322;
assign addr[64079]= 515068990;
assign addr[64080]= 805879757;
assign addr[64081]= 1080359326;
assign addr[64082]= 1332945355;
assign addr[64083]= 1558519173;
assign addr[64084]= 1752509516;
assign addr[64085]= 1910985158;
assign addr[64086]= 2030734582;
assign addr[64087]= 2109331059;
assign addr[64088]= 2145181827;
assign addr[64089]= 2137560369;
assign addr[64090]= 2086621133;
assign addr[64091]= 1993396407;
assign addr[64092]= 1859775393;
assign addr[64093]= 1688465931;
assign addr[64094]= 1482939614;
assign addr[64095]= 1247361445;
assign addr[64096]= 986505429;
assign addr[64097]= 705657826;
assign addr[64098]= 410510029;
assign addr[64099]= 107043224;
assign addr[64100]= -198592817;
assign addr[64101]= -500204365;
assign addr[64102]= -791679244;
assign addr[64103]= -1067110699;
assign addr[64104]= -1320917099;
assign addr[64105]= -1547955041;
assign addr[64106]= -1743623590;
assign addr[64107]= -1903957513;
assign addr[64108]= -2025707632;
assign addr[64109]= -2106406677;
assign addr[64110]= -2144419275;
assign addr[64111]= -2138975100;
assign addr[64112]= -2090184478;
assign addr[64113]= -1999036154;
assign addr[64114]= -1867377253;
assign addr[64115]= -1697875851;
assign addr[64116]= -1493966902;
assign addr[64117]= -1259782632;
assign addr[64118]= -1000068799;
assign addr[64119]= -720088517;
assign addr[64120]= -425515602;
assign addr[64121]= -122319591;
assign addr[64122]= 183355234;
assign addr[64123]= 485314355;
assign addr[64124]= 777438554;
assign addr[64125]= 1053807919;
assign addr[64126]= 1308821808;
assign addr[64127]= 1537312353;
assign addr[64128]= 1734649179;
assign addr[64129]= 1896833245;
assign addr[64130]= 2020577882;
assign addr[64131]= 2103375398;
assign addr[64132]= 2143547897;
assign addr[64133]= 2140281282;
assign addr[64134]= 2093641749;
assign addr[64135]= 2004574453;
assign addr[64136]= 1874884346;
assign addr[64137]= 1707199606;
assign addr[64138]= 1504918373;
assign addr[64139]= 1272139887;
assign addr[64140]= 1013581418;
assign addr[64141]= 734482665;
assign addr[64142]= 440499581;
assign addr[64143]= 137589750;
assign addr[64144]= -168108346;
assign addr[64145]= -470399716;
assign addr[64146]= -763158411;
assign addr[64147]= -1040451659;
assign addr[64148]= -1296660098;
assign addr[64149]= -1526591649;
assign addr[64150]= -1725586737;
assign addr[64151]= -1889612716;
assign addr[64152]= -2015345591;
assign addr[64153]= -2100237377;
assign addr[64154]= -2142567738;
assign addr[64155]= -2141478848;
assign addr[64156]= -2096992772;
assign addr[64157]= -2010011024;
assign addr[64158]= -1882296293;
assign addr[64159]= -1716436725;
assign addr[64160]= -1515793473;
assign addr[64161]= -1284432584;
assign addr[64162]= -1027042599;
assign addr[64163]= -748839539;
assign addr[64164]= -455461206;
assign addr[64165]= -152852926;
assign addr[64166]= 152852926;
assign addr[64167]= 455461206;
assign addr[64168]= 748839539;
assign addr[64169]= 1027042599;
assign addr[64170]= 1284432584;
assign addr[64171]= 1515793473;
assign addr[64172]= 1716436725;
assign addr[64173]= 1882296293;
assign addr[64174]= 2010011024;
assign addr[64175]= 2096992772;
assign addr[64176]= 2141478848;
assign addr[64177]= 2142567738;
assign addr[64178]= 2100237377;
assign addr[64179]= 2015345591;
assign addr[64180]= 1889612716;
assign addr[64181]= 1725586737;
assign addr[64182]= 1526591649;
assign addr[64183]= 1296660098;
assign addr[64184]= 1040451659;
assign addr[64185]= 763158411;
assign addr[64186]= 470399716;
assign addr[64187]= 168108346;
assign addr[64188]= -137589750;
assign addr[64189]= -440499581;
assign addr[64190]= -734482665;
assign addr[64191]= -1013581418;
assign addr[64192]= -1272139887;
assign addr[64193]= -1504918373;
assign addr[64194]= -1707199606;
assign addr[64195]= -1874884346;
assign addr[64196]= -2004574453;
assign addr[64197]= -2093641749;
assign addr[64198]= -2140281282;
assign addr[64199]= -2143547897;
assign addr[64200]= -2103375398;
assign addr[64201]= -2020577882;
assign addr[64202]= -1896833245;
assign addr[64203]= -1734649179;
assign addr[64204]= -1537312353;
assign addr[64205]= -1308821808;
assign addr[64206]= -1053807919;
assign addr[64207]= -777438554;
assign addr[64208]= -485314355;
assign addr[64209]= -183355234;
assign addr[64210]= 122319591;
assign addr[64211]= 425515602;
assign addr[64212]= 720088517;
assign addr[64213]= 1000068799;
assign addr[64214]= 1259782632;
assign addr[64215]= 1493966902;
assign addr[64216]= 1697875851;
assign addr[64217]= 1867377253;
assign addr[64218]= 1999036154;
assign addr[64219]= 2090184478;
assign addr[64220]= 2138975100;
assign addr[64221]= 2144419275;
assign addr[64222]= 2106406677;
assign addr[64223]= 2025707632;
assign addr[64224]= 1903957513;
assign addr[64225]= 1743623590;
assign addr[64226]= 1547955041;
assign addr[64227]= 1320917099;
assign addr[64228]= 1067110699;
assign addr[64229]= 791679244;
assign addr[64230]= 500204365;
assign addr[64231]= 198592817;
assign addr[64232]= -107043224;
assign addr[64233]= -410510029;
assign addr[64234]= -705657826;
assign addr[64235]= -986505429;
assign addr[64236]= -1247361445;
assign addr[64237]= -1482939614;
assign addr[64238]= -1688465931;
assign addr[64239]= -1859775393;
assign addr[64240]= -1993396407;
assign addr[64241]= -2086621133;
assign addr[64242]= -2137560369;
assign addr[64243]= -2145181827;
assign addr[64244]= -2109331059;
assign addr[64245]= -2030734582;
assign addr[64246]= -1910985158;
assign addr[64247]= -1752509516;
assign addr[64248]= -1558519173;
assign addr[64249]= -1332945355;
assign addr[64250]= -1080359326;
assign addr[64251]= -805879757;
assign addr[64252]= -515068990;
assign addr[64253]= -213820322;
assign addr[64254]= 91761426;
assign addr[64255]= 395483624;
assign addr[64256]= 691191324;
assign addr[64257]= 972891995;
assign addr[64258]= 1234876957;
assign addr[64259]= 1471837070;
assign addr[64260]= 1678970324;
assign addr[64261]= 1852079154;
assign addr[64262]= 1987655498;
assign addr[64263]= 2082951896;
assign addr[64264]= 2136037160;
assign addr[64265]= 2145835515;
assign addr[64266]= 2112148396;
assign addr[64267]= 2035658475;
assign addr[64268]= 1917915825;
assign addr[64269]= 1761306505;
assign addr[64270]= 1569004214;
assign addr[64271]= 1344905966;
assign addr[64272]= 1093553126;
assign addr[64273]= 820039373;
assign addr[64274]= 529907477;
assign addr[64275]= 229036977;
assign addr[64276]= -76474970;
assign addr[64277]= -380437148;
assign addr[64278]= -676689746;
assign addr[64279]= -959229189;
assign addr[64280]= -1222329801;
assign addr[64281]= -1460659832;
assign addr[64282]= -1669389513;
assign addr[64283]= -1844288924;
assign addr[64284]= -1981813720;
assign addr[64285]= -2079176953;
assign addr[64286]= -2134405552;
assign addr[64287]= -2146380306;
assign addr[64288]= -2114858546;
assign addr[64289]= -2040479063;
assign addr[64290]= -1924749160;
assign addr[64291]= -1770014111;
assign addr[64292]= -1579409630;
assign addr[64293]= -1356798326;
assign addr[64294]= -1106691431;
assign addr[64295]= -834157373;
assign addr[64296]= -544719071;
assign addr[64297]= -244242007;
assign addr[64298]= 61184634;
assign addr[64299]= 365371365;
assign addr[64300]= 662153826;
assign addr[64301]= 945517704;
assign addr[64302]= 1209720613;
assign addr[64303]= 1449408469;
assign addr[64304]= 1659723983;
assign addr[64305]= 1836405100;
assign addr[64306]= 1975871368;
assign addr[64307]= 2075296495;
assign addr[64308]= 2132665626;
assign addr[64309]= 2146816171;
assign addr[64310]= 2117461370;
assign addr[64311]= 2045196100;
assign addr[64312]= 1931484818;
assign addr[64313]= 1778631892;
assign addr[64314]= 1589734894;
assign addr[64315]= 1368621831;
assign addr[64316]= 1119773573;
assign addr[64317]= 848233042;
assign addr[64318]= 559503022;
assign addr[64319]= 259434643;
assign addr[64320]= -45891193;
assign addr[64321]= -350287041;
assign addr[64322]= -647584304;
assign addr[64323]= -931758235;
assign addr[64324]= -1197050035;
assign addr[64325]= -1438083551;
assign addr[64326]= -1649974225;
assign addr[64327]= -1828428082;
assign addr[64328]= -1969828744;
assign addr[64329]= -2071310720;
assign addr[64330]= -2130817471;
assign addr[64331]= -2147143090;
assign addr[64332]= -2119956737;
assign addr[64333]= -2049809346;
assign addr[64334]= -1938122457;
assign addr[64335]= -1787159411;
assign addr[64336]= -1599979481;
assign addr[64337]= -1380375881;
assign addr[64338]= -1132798888;
assign addr[64339]= -862265664;
assign addr[64340]= -574258580;
assign addr[64341]= -274614114;
assign addr[64342]= 30595422;
assign addr[64343]= 335184940;
assign addr[64344]= 632981917;
assign addr[64345]= 917951481;
assign addr[64346]= 1184318708;
assign addr[64347]= 1426685652;
assign addr[64348]= 1640140734;
assign addr[64349]= 1820358275;
assign addr[64350]= 1963686155;
assign addr[64351]= 2067219829;
assign addr[64352]= 2128861181;
assign addr[64353]= 2147361045;
assign addr[64354]= 2122344521;
assign addr[64355]= 2054318569;
assign addr[64356]= 1944661739;
assign addr[64357]= 1795596234;
assign addr[64358]= 1610142873;
assign addr[64359]= 1392059879;
assign addr[64360]= 1145766716;
assign addr[64361]= 876254528;
assign addr[64362]= 588984994;
assign addr[64363]= 289779648;
assign addr[64364]= -15298099;
assign addr[64365]= -320065829;
assign addr[64366]= -618347408;
assign addr[64367]= -904098143;
assign addr[64368]= -1171527280;
assign addr[64369]= -1415215352;
assign addr[64370]= -1630224009;
assign addr[64371]= -1812196087;
assign addr[64372]= -1957443913;
assign addr[64373]= -2063024031;
assign addr[64374]= -2126796855;
assign addr[64375]= -2147470025;
assign addr[64376]= -2124624598;
assign addr[64377]= -2058723538;
assign addr[64378]= -1951102334;
assign addr[64379]= -1803941934;
assign addr[64380]= -1620224553;
assign addr[64381]= -1403673233;
assign addr[64382]= -1158676398;
assign addr[64383]= -890198924;
assign addr[64384]= -603681519;
assign addr[64385]= -304930476;
assign addr[64386]= 0;
assign addr[64387]= 304930476;
assign addr[64388]= 603681519;
assign addr[64389]= 890198924;
assign addr[64390]= 1158676398;
assign addr[64391]= 1403673233;
assign addr[64392]= 1620224553;
assign addr[64393]= 1803941934;
assign addr[64394]= 1951102334;
assign addr[64395]= 2058723538;
assign addr[64396]= 2124624598;
assign addr[64397]= 2147470025;
assign addr[64398]= 2126796855;
assign addr[64399]= 2063024031;
assign addr[64400]= 1957443913;
assign addr[64401]= 1812196087;
assign addr[64402]= 1630224009;
assign addr[64403]= 1415215352;
assign addr[64404]= 1171527280;
assign addr[64405]= 904098143;
assign addr[64406]= 618347408;
assign addr[64407]= 320065829;
assign addr[64408]= 15298099;
assign addr[64409]= -289779648;
assign addr[64410]= -588984994;
assign addr[64411]= -876254528;
assign addr[64412]= -1145766716;
assign addr[64413]= -1392059879;
assign addr[64414]= -1610142873;
assign addr[64415]= -1795596234;
assign addr[64416]= -1944661739;
assign addr[64417]= -2054318569;
assign addr[64418]= -2122344521;
assign addr[64419]= -2147361045;
assign addr[64420]= -2128861181;
assign addr[64421]= -2067219829;
assign addr[64422]= -1963686155;
assign addr[64423]= -1820358275;
assign addr[64424]= -1640140734;
assign addr[64425]= -1426685652;
assign addr[64426]= -1184318708;
assign addr[64427]= -917951481;
assign addr[64428]= -632981917;
assign addr[64429]= -335184940;
assign addr[64430]= -30595422;
assign addr[64431]= 274614114;
assign addr[64432]= 574258580;
assign addr[64433]= 862265664;
assign addr[64434]= 1132798888;
assign addr[64435]= 1380375881;
assign addr[64436]= 1599979481;
assign addr[64437]= 1787159411;
assign addr[64438]= 1938122457;
assign addr[64439]= 2049809346;
assign addr[64440]= 2119956737;
assign addr[64441]= 2147143090;
assign addr[64442]= 2130817471;
assign addr[64443]= 2071310720;
assign addr[64444]= 1969828744;
assign addr[64445]= 1828428082;
assign addr[64446]= 1649974225;
assign addr[64447]= 1438083551;
assign addr[64448]= 1197050035;
assign addr[64449]= 931758235;
assign addr[64450]= 647584304;
assign addr[64451]= 350287041;
assign addr[64452]= 45891193;
assign addr[64453]= -259434643;
assign addr[64454]= -559503022;
assign addr[64455]= -848233042;
assign addr[64456]= -1119773573;
assign addr[64457]= -1368621831;
assign addr[64458]= -1589734894;
assign addr[64459]= -1778631892;
assign addr[64460]= -1931484818;
assign addr[64461]= -2045196100;
assign addr[64462]= -2117461370;
assign addr[64463]= -2146816171;
assign addr[64464]= -2132665626;
assign addr[64465]= -2075296495;
assign addr[64466]= -1975871368;
assign addr[64467]= -1836405100;
assign addr[64468]= -1659723983;
assign addr[64469]= -1449408469;
assign addr[64470]= -1209720613;
assign addr[64471]= -945517704;
assign addr[64472]= -662153826;
assign addr[64473]= -365371365;
assign addr[64474]= -61184634;
assign addr[64475]= 244242007;
assign addr[64476]= 544719071;
assign addr[64477]= 834157373;
assign addr[64478]= 1106691431;
assign addr[64479]= 1356798326;
assign addr[64480]= 1579409630;
assign addr[64481]= 1770014111;
assign addr[64482]= 1924749160;
assign addr[64483]= 2040479063;
assign addr[64484]= 2114858546;
assign addr[64485]= 2146380306;
assign addr[64486]= 2134405552;
assign addr[64487]= 2079176953;
assign addr[64488]= 1981813720;
assign addr[64489]= 1844288924;
assign addr[64490]= 1669389513;
assign addr[64491]= 1460659832;
assign addr[64492]= 1222329801;
assign addr[64493]= 959229189;
assign addr[64494]= 676689746;
assign addr[64495]= 380437148;
assign addr[64496]= 76474970;
assign addr[64497]= -229036977;
assign addr[64498]= -529907477;
assign addr[64499]= -820039373;
assign addr[64500]= -1093553126;
assign addr[64501]= -1344905966;
assign addr[64502]= -1569004214;
assign addr[64503]= -1761306505;
assign addr[64504]= -1917915825;
assign addr[64505]= -2035658475;
assign addr[64506]= -2112148396;
assign addr[64507]= -2145835515;
assign addr[64508]= -2136037160;
assign addr[64509]= -2082951896;
assign addr[64510]= -1987655498;
assign addr[64511]= -1852079154;
assign addr[64512]= -1678970324;
assign addr[64513]= -1471837070;
assign addr[64514]= -1234876957;
assign addr[64515]= -972891995;
assign addr[64516]= -691191324;
assign addr[64517]= -395483624;
assign addr[64518]= -91761426;
assign addr[64519]= 213820322;
assign addr[64520]= 515068990;
assign addr[64521]= 805879757;
assign addr[64522]= 1080359326;
assign addr[64523]= 1332945355;
assign addr[64524]= 1558519173;
assign addr[64525]= 1752509516;
assign addr[64526]= 1910985158;
assign addr[64527]= 2030734582;
assign addr[64528]= 2109331059;
assign addr[64529]= 2145181827;
assign addr[64530]= 2137560369;
assign addr[64531]= 2086621133;
assign addr[64532]= 1993396407;
assign addr[64533]= 1859775393;
assign addr[64534]= 1688465931;
assign addr[64535]= 1482939614;
assign addr[64536]= 1247361445;
assign addr[64537]= 986505429;
assign addr[64538]= 705657826;
assign addr[64539]= 410510029;
assign addr[64540]= 107043224;
assign addr[64541]= -198592817;
assign addr[64542]= -500204365;
assign addr[64543]= -791679244;
assign addr[64544]= -1067110699;
assign addr[64545]= -1320917099;
assign addr[64546]= -1547955041;
assign addr[64547]= -1743623590;
assign addr[64548]= -1903957513;
assign addr[64549]= -2025707632;
assign addr[64550]= -2106406677;
assign addr[64551]= -2144419275;
assign addr[64552]= -2138975100;
assign addr[64553]= -2090184478;
assign addr[64554]= -1999036154;
assign addr[64555]= -1867377253;
assign addr[64556]= -1697875851;
assign addr[64557]= -1493966902;
assign addr[64558]= -1259782632;
assign addr[64559]= -1000068799;
assign addr[64560]= -720088517;
assign addr[64561]= -425515602;
assign addr[64562]= -122319591;
assign addr[64563]= 183355234;
assign addr[64564]= 485314355;
assign addr[64565]= 777438554;
assign addr[64566]= 1053807919;
assign addr[64567]= 1308821808;
assign addr[64568]= 1537312353;
assign addr[64569]= 1734649179;
assign addr[64570]= 1896833245;
assign addr[64571]= 2020577882;
assign addr[64572]= 2103375398;
assign addr[64573]= 2143547897;
assign addr[64574]= 2140281282;
assign addr[64575]= 2093641749;
assign addr[64576]= 2004574453;
assign addr[64577]= 1874884346;
assign addr[64578]= 1707199606;
assign addr[64579]= 1504918373;
assign addr[64580]= 1272139887;
assign addr[64581]= 1013581418;
assign addr[64582]= 734482665;
assign addr[64583]= 440499581;
assign addr[64584]= 137589750;
assign addr[64585]= -168108346;
assign addr[64586]= -470399716;
assign addr[64587]= -763158411;
assign addr[64588]= -1040451659;
assign addr[64589]= -1296660098;
assign addr[64590]= -1526591649;
assign addr[64591]= -1725586737;
assign addr[64592]= -1889612716;
assign addr[64593]= -2015345591;
assign addr[64594]= -2100237377;
assign addr[64595]= -2142567738;
assign addr[64596]= -2141478848;
assign addr[64597]= -2096992772;
assign addr[64598]= -2010011024;
assign addr[64599]= -1882296293;
assign addr[64600]= -1716436725;
assign addr[64601]= -1515793473;
assign addr[64602]= -1284432584;
assign addr[64603]= -1027042599;
assign addr[64604]= -748839539;
assign addr[64605]= -455461206;
assign addr[64606]= -152852926;
assign addr[64607]= 152852926;
assign addr[64608]= 455461206;
assign addr[64609]= 748839539;
assign addr[64610]= 1027042599;
assign addr[64611]= 1284432584;
assign addr[64612]= 1515793473;
assign addr[64613]= 1716436725;
assign addr[64614]= 1882296293;
assign addr[64615]= 2010011024;
assign addr[64616]= 2096992772;
assign addr[64617]= 2141478848;
assign addr[64618]= 2142567738;
assign addr[64619]= 2100237377;
assign addr[64620]= 2015345591;
assign addr[64621]= 1889612716;
assign addr[64622]= 1725586737;
assign addr[64623]= 1526591649;
assign addr[64624]= 1296660098;
assign addr[64625]= 1040451659;
assign addr[64626]= 763158411;
assign addr[64627]= 470399716;
assign addr[64628]= 168108346;
assign addr[64629]= -137589750;
assign addr[64630]= -440499581;
assign addr[64631]= -734482665;
assign addr[64632]= -1013581418;
assign addr[64633]= -1272139887;
assign addr[64634]= -1504918373;
assign addr[64635]= -1707199606;
assign addr[64636]= -1874884346;
assign addr[64637]= -2004574453;
assign addr[64638]= -2093641749;
assign addr[64639]= -2140281282;
assign addr[64640]= -2143547897;
assign addr[64641]= -2103375398;
assign addr[64642]= -2020577882;
assign addr[64643]= -1896833245;
assign addr[64644]= -1734649179;
assign addr[64645]= -1537312353;
assign addr[64646]= -1308821808;
assign addr[64647]= -1053807919;
assign addr[64648]= -777438554;
assign addr[64649]= -485314355;
assign addr[64650]= -183355234;
assign addr[64651]= 122319591;
assign addr[64652]= 425515602;
assign addr[64653]= 720088517;
assign addr[64654]= 1000068799;
assign addr[64655]= 1259782632;
assign addr[64656]= 1493966902;
assign addr[64657]= 1697875851;
assign addr[64658]= 1867377253;
assign addr[64659]= 1999036154;
assign addr[64660]= 2090184478;
assign addr[64661]= 2138975100;
assign addr[64662]= 2144419275;
assign addr[64663]= 2106406677;
assign addr[64664]= 2025707632;
assign addr[64665]= 1903957513;
assign addr[64666]= 1743623590;
assign addr[64667]= 1547955041;
assign addr[64668]= 1320917099;
assign addr[64669]= 1067110699;
assign addr[64670]= 791679244;
assign addr[64671]= 500204365;
assign addr[64672]= 198592817;
assign addr[64673]= -107043224;
assign addr[64674]= -410510029;
assign addr[64675]= -705657826;
assign addr[64676]= -986505429;
assign addr[64677]= -1247361445;
assign addr[64678]= -1482939614;
assign addr[64679]= -1688465931;
assign addr[64680]= -1859775393;
assign addr[64681]= -1993396407;
assign addr[64682]= -2086621133;
assign addr[64683]= -2137560369;
assign addr[64684]= -2145181827;
assign addr[64685]= -2109331059;
assign addr[64686]= -2030734582;
assign addr[64687]= -1910985158;
assign addr[64688]= -1752509516;
assign addr[64689]= -1558519173;
assign addr[64690]= -1332945355;
assign addr[64691]= -1080359326;
assign addr[64692]= -805879757;
assign addr[64693]= -515068990;
assign addr[64694]= -213820322;
assign addr[64695]= 91761426;
assign addr[64696]= 395483624;
assign addr[64697]= 691191324;
assign addr[64698]= 972891995;
assign addr[64699]= 1234876957;
assign addr[64700]= 1471837070;
assign addr[64701]= 1678970324;
assign addr[64702]= 1852079154;
assign addr[64703]= 1987655498;
assign addr[64704]= 2082951896;
assign addr[64705]= 2136037160;
assign addr[64706]= 2145835515;
assign addr[64707]= 2112148396;
assign addr[64708]= 2035658475;
assign addr[64709]= 1917915825;
assign addr[64710]= 1761306505;
assign addr[64711]= 1569004214;
assign addr[64712]= 1344905966;
assign addr[64713]= 1093553126;
assign addr[64714]= 820039373;
assign addr[64715]= 529907477;
assign addr[64716]= 229036977;
assign addr[64717]= -76474970;
assign addr[64718]= -380437148;
assign addr[64719]= -676689746;
assign addr[64720]= -959229189;
assign addr[64721]= -1222329801;
assign addr[64722]= -1460659832;
assign addr[64723]= -1669389513;
assign addr[64724]= -1844288924;
assign addr[64725]= -1981813720;
assign addr[64726]= -2079176953;
assign addr[64727]= -2134405552;
assign addr[64728]= -2146380306;
assign addr[64729]= -2114858546;
assign addr[64730]= -2040479063;
assign addr[64731]= -1924749160;
assign addr[64732]= -1770014111;
assign addr[64733]= -1579409630;
assign addr[64734]= -1356798326;
assign addr[64735]= -1106691431;
assign addr[64736]= -834157373;
assign addr[64737]= -544719071;
assign addr[64738]= -244242007;
assign addr[64739]= 61184634;
assign addr[64740]= 365371365;
assign addr[64741]= 662153826;
assign addr[64742]= 945517704;
assign addr[64743]= 1209720613;
assign addr[64744]= 1449408469;
assign addr[64745]= 1659723983;
assign addr[64746]= 1836405100;
assign addr[64747]= 1975871368;
assign addr[64748]= 2075296495;
assign addr[64749]= 2132665626;
assign addr[64750]= 2146816171;
assign addr[64751]= 2117461370;
assign addr[64752]= 2045196100;
assign addr[64753]= 1931484818;
assign addr[64754]= 1778631892;
assign addr[64755]= 1589734894;
assign addr[64756]= 1368621831;
assign addr[64757]= 1119773573;
assign addr[64758]= 848233042;
assign addr[64759]= 559503022;
assign addr[64760]= 259434643;
assign addr[64761]= -45891193;
assign addr[64762]= -350287041;
assign addr[64763]= -647584304;
assign addr[64764]= -931758235;
assign addr[64765]= -1197050035;
assign addr[64766]= -1438083551;
assign addr[64767]= -1649974225;
assign addr[64768]= -1828428082;
assign addr[64769]= -1969828744;
assign addr[64770]= -2071310720;
assign addr[64771]= -2130817471;
assign addr[64772]= -2147143090;
assign addr[64773]= -2119956737;
assign addr[64774]= -2049809346;
assign addr[64775]= -1938122457;
assign addr[64776]= -1787159411;
assign addr[64777]= -1599979481;
assign addr[64778]= -1380375881;
assign addr[64779]= -1132798888;
assign addr[64780]= -862265664;
assign addr[64781]= -574258580;
assign addr[64782]= -274614114;
assign addr[64783]= 30595422;
assign addr[64784]= 335184940;
assign addr[64785]= 632981917;
assign addr[64786]= 917951481;
assign addr[64787]= 1184318708;
assign addr[64788]= 1426685652;
assign addr[64789]= 1640140734;
assign addr[64790]= 1820358275;
assign addr[64791]= 1963686155;
assign addr[64792]= 2067219829;
assign addr[64793]= 2128861181;
assign addr[64794]= 2147361045;
assign addr[64795]= 2122344521;
assign addr[64796]= 2054318569;
assign addr[64797]= 1944661739;
assign addr[64798]= 1795596234;
assign addr[64799]= 1610142873;
assign addr[64800]= 1392059879;
assign addr[64801]= 1145766716;
assign addr[64802]= 876254528;
assign addr[64803]= 588984994;
assign addr[64804]= 289779648;
assign addr[64805]= -15298099;
assign addr[64806]= -320065829;
assign addr[64807]= -618347408;
assign addr[64808]= -904098143;
assign addr[64809]= -1171527280;
assign addr[64810]= -1415215352;
assign addr[64811]= -1630224009;
assign addr[64812]= -1812196087;
assign addr[64813]= -1957443913;
assign addr[64814]= -2063024031;
assign addr[64815]= -2126796855;
assign addr[64816]= -2147470025;
assign addr[64817]= -2124624598;
assign addr[64818]= -2058723538;
assign addr[64819]= -1951102334;
assign addr[64820]= -1803941934;
assign addr[64821]= -1620224553;
assign addr[64822]= -1403673233;
assign addr[64823]= -1158676398;
assign addr[64824]= -890198924;
assign addr[64825]= -603681519;
assign addr[64826]= -304930476;
assign addr[64827]= 0;
assign addr[64828]= 304930476;
assign addr[64829]= 603681519;
assign addr[64830]= 890198924;
assign addr[64831]= 1158676398;
assign addr[64832]= 1403673233;
assign addr[64833]= 1620224553;
assign addr[64834]= 1803941934;
assign addr[64835]= 1951102334;
assign addr[64836]= 2058723538;
assign addr[64837]= 2124624598;
assign addr[64838]= 2147470025;
assign addr[64839]= 2126796855;
assign addr[64840]= 2063024031;
assign addr[64841]= 1957443913;
assign addr[64842]= 1812196087;
assign addr[64843]= 1630224009;
assign addr[64844]= 1415215352;
assign addr[64845]= 1171527280;
assign addr[64846]= 904098143;
assign addr[64847]= 618347408;
assign addr[64848]= 320065829;
assign addr[64849]= 15298099;
assign addr[64850]= -289779648;
assign addr[64851]= -588984994;
assign addr[64852]= -876254528;
assign addr[64853]= -1145766716;
assign addr[64854]= -1392059879;
assign addr[64855]= -1610142873;
assign addr[64856]= -1795596234;
assign addr[64857]= -1944661739;
assign addr[64858]= -2054318569;
assign addr[64859]= -2122344521;
assign addr[64860]= -2147361045;
assign addr[64861]= -2128861181;
assign addr[64862]= -2067219829;
assign addr[64863]= -1963686155;
assign addr[64864]= -1820358275;
assign addr[64865]= -1640140734;
assign addr[64866]= -1426685652;
assign addr[64867]= -1184318708;
assign addr[64868]= -917951481;
assign addr[64869]= -632981917;
assign addr[64870]= -335184940;
assign addr[64871]= -30595422;
assign addr[64872]= 274614114;
assign addr[64873]= 574258580;
assign addr[64874]= 862265664;
assign addr[64875]= 1132798888;
assign addr[64876]= 1380375881;
assign addr[64877]= 1599979481;
assign addr[64878]= 1787159411;
assign addr[64879]= 1938122457;
assign addr[64880]= 2049809346;
assign addr[64881]= 2119956737;
assign addr[64882]= 2147143090;
assign addr[64883]= 2130817471;
assign addr[64884]= 2071310720;
assign addr[64885]= 1969828744;
assign addr[64886]= 1828428082;
assign addr[64887]= 1649974225;
assign addr[64888]= 1438083551;
assign addr[64889]= 1197050035;
assign addr[64890]= 931758235;
assign addr[64891]= 647584304;
assign addr[64892]= 350287041;
assign addr[64893]= 45891193;
assign addr[64894]= -259434643;
assign addr[64895]= -559503022;
assign addr[64896]= -848233042;
assign addr[64897]= -1119773573;
assign addr[64898]= -1368621831;
assign addr[64899]= -1589734894;
assign addr[64900]= -1778631892;
assign addr[64901]= -1931484818;
assign addr[64902]= -2045196100;
assign addr[64903]= -2117461370;
assign addr[64904]= -2146816171;
assign addr[64905]= -2132665626;
assign addr[64906]= -2075296495;
assign addr[64907]= -1975871368;
assign addr[64908]= -1836405100;
assign addr[64909]= -1659723983;
assign addr[64910]= -1449408469;
assign addr[64911]= -1209720613;
assign addr[64912]= -945517704;
assign addr[64913]= -662153826;
assign addr[64914]= -365371365;
assign addr[64915]= -61184634;
assign addr[64916]= 244242007;
assign addr[64917]= 544719071;
assign addr[64918]= 834157373;
assign addr[64919]= 1106691431;
assign addr[64920]= 1356798326;
assign addr[64921]= 1579409630;
assign addr[64922]= 1770014111;
assign addr[64923]= 1924749160;
assign addr[64924]= 2040479063;
assign addr[64925]= 2114858546;
assign addr[64926]= 2146380306;
assign addr[64927]= 2134405552;
assign addr[64928]= 2079176953;
assign addr[64929]= 1981813720;
assign addr[64930]= 1844288924;
assign addr[64931]= 1669389513;
assign addr[64932]= 1460659832;
assign addr[64933]= 1222329801;
assign addr[64934]= 959229189;
assign addr[64935]= 676689746;
assign addr[64936]= 380437148;
assign addr[64937]= 76474970;
assign addr[64938]= -229036977;
assign addr[64939]= -529907477;
assign addr[64940]= -820039373;
assign addr[64941]= -1093553126;
assign addr[64942]= -1344905966;
assign addr[64943]= -1569004214;
assign addr[64944]= -1761306505;
assign addr[64945]= -1917915825;
assign addr[64946]= -2035658475;
assign addr[64947]= -2112148396;
assign addr[64948]= -2145835515;
assign addr[64949]= -2136037160;
assign addr[64950]= -2082951896;
assign addr[64951]= -1987655498;
assign addr[64952]= -1852079154;
assign addr[64953]= -1678970324;
assign addr[64954]= -1471837070;
assign addr[64955]= -1234876957;
assign addr[64956]= -972891995;
assign addr[64957]= -691191324;
assign addr[64958]= -395483624;
assign addr[64959]= -91761426;
assign addr[64960]= 213820322;
assign addr[64961]= 515068990;
assign addr[64962]= 805879757;
assign addr[64963]= 1080359326;
assign addr[64964]= 1332945355;
assign addr[64965]= 1558519173;
assign addr[64966]= 1752509516;
assign addr[64967]= 1910985158;
assign addr[64968]= 2030734582;
assign addr[64969]= 2109331059;
assign addr[64970]= 2145181827;
assign addr[64971]= 2137560369;
assign addr[64972]= 2086621133;
assign addr[64973]= 1993396407;
assign addr[64974]= 1859775393;
assign addr[64975]= 1688465931;
assign addr[64976]= 1482939614;
assign addr[64977]= 1247361445;
assign addr[64978]= 986505429;
assign addr[64979]= 705657826;
assign addr[64980]= 410510029;
assign addr[64981]= 107043224;
assign addr[64982]= -198592817;
assign addr[64983]= -500204365;
assign addr[64984]= -791679244;
assign addr[64985]= -1067110699;
assign addr[64986]= -1320917099;
assign addr[64987]= -1547955041;
assign addr[64988]= -1743623590;
assign addr[64989]= -1903957513;
assign addr[64990]= -2025707632;
assign addr[64991]= -2106406677;
assign addr[64992]= -2144419275;
assign addr[64993]= -2138975100;
assign addr[64994]= -2090184478;
assign addr[64995]= -1999036154;
assign addr[64996]= -1867377253;
assign addr[64997]= -1697875851;
assign addr[64998]= -1493966902;
assign addr[64999]= -1259782632;
assign addr[65000]= -1000068799;
assign addr[65001]= -720088517;
assign addr[65002]= -425515602;
assign addr[65003]= -122319591;
assign addr[65004]= 183355234;
assign addr[65005]= 485314355;
assign addr[65006]= 777438554;
assign addr[65007]= 1053807919;
assign addr[65008]= 1308821808;
assign addr[65009]= 1537312353;
assign addr[65010]= 1734649179;
assign addr[65011]= 1896833245;
assign addr[65012]= 2020577882;
assign addr[65013]= 2103375398;
assign addr[65014]= 2143547897;
assign addr[65015]= 2140281282;
assign addr[65016]= 2093641749;
assign addr[65017]= 2004574453;
assign addr[65018]= 1874884346;
assign addr[65019]= 1707199606;
assign addr[65020]= 1504918373;
assign addr[65021]= 1272139887;
assign addr[65022]= 1013581418;
assign addr[65023]= 734482665;
assign addr[65024]= 440499581;
assign addr[65025]= 137589750;
assign addr[65026]= -168108346;
assign addr[65027]= -470399716;
assign addr[65028]= -763158411;
assign addr[65029]= -1040451659;
assign addr[65030]= -1296660098;
assign addr[65031]= -1526591649;
assign addr[65032]= -1725586737;
assign addr[65033]= -1889612716;
assign addr[65034]= -2015345591;
assign addr[65035]= -2100237377;
assign addr[65036]= -2142567738;
assign addr[65037]= -2141478848;
assign addr[65038]= -2096992772;
assign addr[65039]= -2010011024;
assign addr[65040]= -1882296293;
assign addr[65041]= -1716436725;
assign addr[65042]= -1515793473;
assign addr[65043]= -1284432584;
assign addr[65044]= -1027042599;
assign addr[65045]= -748839539;
assign addr[65046]= -455461206;
assign addr[65047]= -152852926;
assign addr[65048]= 152852926;
assign addr[65049]= 455461206;
assign addr[65050]= 748839539;
assign addr[65051]= 1027042599;
assign addr[65052]= 1284432584;
assign addr[65053]= 1515793473;
assign addr[65054]= 1716436725;
assign addr[65055]= 1882296293;
assign addr[65056]= 2010011024;
assign addr[65057]= 2096992772;
assign addr[65058]= 2141478848;
assign addr[65059]= 2142567738;
assign addr[65060]= 2100237377;
assign addr[65061]= 2015345591;
assign addr[65062]= 1889612716;
assign addr[65063]= 1725586737;
assign addr[65064]= 1526591649;
assign addr[65065]= 1296660098;
assign addr[65066]= 1040451659;
assign addr[65067]= 763158411;
assign addr[65068]= 470399716;
assign addr[65069]= 168108346;
assign addr[65070]= -137589750;
assign addr[65071]= -440499581;
assign addr[65072]= -734482665;
assign addr[65073]= -1013581418;
assign addr[65074]= -1272139887;
assign addr[65075]= -1504918373;
assign addr[65076]= -1707199606;
assign addr[65077]= -1874884346;
assign addr[65078]= -2004574453;
assign addr[65079]= -2093641749;
assign addr[65080]= -2140281282;
assign addr[65081]= -2143547897;
assign addr[65082]= -2103375398;
assign addr[65083]= -2020577882;
assign addr[65084]= -1896833245;
assign addr[65085]= -1734649179;
assign addr[65086]= -1537312353;
assign addr[65087]= -1308821808;
assign addr[65088]= -1053807919;
assign addr[65089]= -777438554;
assign addr[65090]= -485314355;
assign addr[65091]= -183355234;
assign addr[65092]= 122319591;
assign addr[65093]= 425515602;
assign addr[65094]= 720088517;
assign addr[65095]= 1000068799;
assign addr[65096]= 1259782632;
assign addr[65097]= 1493966902;
assign addr[65098]= 1697875851;
assign addr[65099]= 1867377253;
assign addr[65100]= 1999036154;
assign addr[65101]= 2090184478;
assign addr[65102]= 2138975100;
assign addr[65103]= 2144419275;
assign addr[65104]= 2106406677;
assign addr[65105]= 2025707632;
assign addr[65106]= 1903957513;
assign addr[65107]= 1743623590;
assign addr[65108]= 1547955041;
assign addr[65109]= 1320917099;
assign addr[65110]= 1067110699;
assign addr[65111]= 791679244;
assign addr[65112]= 500204365;
assign addr[65113]= 198592817;
assign addr[65114]= -107043224;
assign addr[65115]= -410510029;
assign addr[65116]= -705657826;
assign addr[65117]= -986505429;
assign addr[65118]= -1247361445;
assign addr[65119]= -1482939614;
assign addr[65120]= -1688465931;
assign addr[65121]= -1859775393;
assign addr[65122]= -1993396407;
assign addr[65123]= -2086621133;
assign addr[65124]= -2137560369;
assign addr[65125]= -2145181827;
assign addr[65126]= -2109331059;
assign addr[65127]= -2030734582;
assign addr[65128]= -1910985158;
assign addr[65129]= -1752509516;
assign addr[65130]= -1558519173;
assign addr[65131]= -1332945355;
assign addr[65132]= -1080359326;
assign addr[65133]= -805879757;
assign addr[65134]= -515068990;
assign addr[65135]= -213820322;
assign addr[65136]= 91761426;
assign addr[65137]= 395483624;
assign addr[65138]= 691191324;
assign addr[65139]= 972891995;
assign addr[65140]= 1234876957;
assign addr[65141]= 1471837070;
assign addr[65142]= 1678970324;
assign addr[65143]= 1852079154;
assign addr[65144]= 1987655498;
assign addr[65145]= 2082951896;
assign addr[65146]= 2136037160;
assign addr[65147]= 2145835515;
assign addr[65148]= 2112148396;
assign addr[65149]= 2035658475;
assign addr[65150]= 1917915825;
assign addr[65151]= 1761306505;
assign addr[65152]= 1569004214;
assign addr[65153]= 1344905966;
assign addr[65154]= 1093553126;
assign addr[65155]= 820039373;
assign addr[65156]= 529907477;
assign addr[65157]= 229036977;
assign addr[65158]= -76474970;
assign addr[65159]= -380437148;
assign addr[65160]= -676689746;
assign addr[65161]= -959229189;
assign addr[65162]= -1222329801;
assign addr[65163]= -1460659832;
assign addr[65164]= -1669389513;
assign addr[65165]= -1844288924;
assign addr[65166]= -1981813720;
assign addr[65167]= -2079176953;
assign addr[65168]= -2134405552;
assign addr[65169]= -2146380306;
assign addr[65170]= -2114858546;
assign addr[65171]= -2040479063;
assign addr[65172]= -1924749160;
assign addr[65173]= -1770014111;
assign addr[65174]= -1579409630;
assign addr[65175]= -1356798326;
assign addr[65176]= -1106691431;
assign addr[65177]= -834157373;
assign addr[65178]= -544719071;
assign addr[65179]= -244242007;
assign addr[65180]= 61184634;
assign addr[65181]= 365371365;
assign addr[65182]= 662153826;
assign addr[65183]= 945517704;
assign addr[65184]= 1209720613;
assign addr[65185]= 1449408469;
assign addr[65186]= 1659723983;
assign addr[65187]= 1836405100;
assign addr[65188]= 1975871368;
assign addr[65189]= 2075296495;
assign addr[65190]= 2132665626;
assign addr[65191]= 2146816171;
assign addr[65192]= 2117461370;
assign addr[65193]= 2045196100;
assign addr[65194]= 1931484818;
assign addr[65195]= 1778631892;
assign addr[65196]= 1589734894;
assign addr[65197]= 1368621831;
assign addr[65198]= 1119773573;
assign addr[65199]= 848233042;
assign addr[65200]= 559503022;
assign addr[65201]= 259434643;
assign addr[65202]= -45891193;
assign addr[65203]= -350287041;
assign addr[65204]= -647584304;
assign addr[65205]= -931758235;
assign addr[65206]= -1197050035;
assign addr[65207]= -1438083551;
assign addr[65208]= -1649974225;
assign addr[65209]= -1828428082;
assign addr[65210]= -1969828744;
assign addr[65211]= -2071310720;
assign addr[65212]= -2130817471;
assign addr[65213]= -2147143090;
assign addr[65214]= -2119956737;
assign addr[65215]= -2049809346;
assign addr[65216]= -1938122457;
assign addr[65217]= -1787159411;
assign addr[65218]= -1599979481;
assign addr[65219]= -1380375881;
assign addr[65220]= -1132798888;
assign addr[65221]= -862265664;
assign addr[65222]= -574258580;
assign addr[65223]= -274614114;
assign addr[65224]= 30595422;
assign addr[65225]= 335184940;
assign addr[65226]= 632981917;
assign addr[65227]= 917951481;
assign addr[65228]= 1184318708;
assign addr[65229]= 1426685652;
assign addr[65230]= 1640140734;
assign addr[65231]= 1820358275;
assign addr[65232]= 1963686155;
assign addr[65233]= 2067219829;
assign addr[65234]= 2128861181;
assign addr[65235]= 2147361045;
assign addr[65236]= 2122344521;
assign addr[65237]= 2054318569;
assign addr[65238]= 1944661739;
assign addr[65239]= 1795596234;
assign addr[65240]= 1610142873;
assign addr[65241]= 1392059879;
assign addr[65242]= 1145766716;
assign addr[65243]= 876254528;
assign addr[65244]= 588984994;
assign addr[65245]= 289779648;
assign addr[65246]= -15298099;
assign addr[65247]= -320065829;
assign addr[65248]= -618347408;
assign addr[65249]= -904098143;
assign addr[65250]= -1171527280;
assign addr[65251]= -1415215352;
assign addr[65252]= -1630224009;
assign addr[65253]= -1812196087;
assign addr[65254]= -1957443913;
assign addr[65255]= -2063024031;
assign addr[65256]= -2126796855;
assign addr[65257]= -2147470025;
assign addr[65258]= -2124624598;
assign addr[65259]= -2058723538;
assign addr[65260]= -1951102334;
assign addr[65261]= -1803941934;
assign addr[65262]= -1620224553;
assign addr[65263]= -1403673233;
assign addr[65264]= -1158676398;
assign addr[65265]= -890198924;
assign addr[65266]= -603681519;
assign addr[65267]= -304930476;
assign addr[65268]= 0;
assign addr[65269]= 304930476;
assign addr[65270]= 603681519;
assign addr[65271]= 890198924;
assign addr[65272]= 1158676398;
assign addr[65273]= 1403673233;
assign addr[65274]= 1620224553;
assign addr[65275]= 1803941934;
assign addr[65276]= 1951102334;
assign addr[65277]= 2058723538;
assign addr[65278]= 2124624598;
assign addr[65279]= 2147470025;
assign addr[65280]= 2126796855;
assign addr[65281]= 2063024031;
assign addr[65282]= 1957443913;
assign addr[65283]= 1812196087;
assign addr[65284]= 1630224009;
assign addr[65285]= 1415215352;
assign addr[65286]= 1171527280;
assign addr[65287]= 904098143;
assign addr[65288]= 618347408;
assign addr[65289]= 320065829;
assign addr[65290]= 15298099;
assign addr[65291]= -289779648;
assign addr[65292]= -588984994;
assign addr[65293]= -876254528;
assign addr[65294]= -1145766716;
assign addr[65295]= -1392059879;
assign addr[65296]= -1610142873;
assign addr[65297]= -1795596234;
assign addr[65298]= -1944661739;
assign addr[65299]= -2054318569;
assign addr[65300]= -2122344521;
assign addr[65301]= -2147361045;
assign addr[65302]= -2128861181;
assign addr[65303]= -2067219829;
assign addr[65304]= -1963686155;
assign addr[65305]= -1820358275;
assign addr[65306]= -1640140734;
assign addr[65307]= -1426685652;
assign addr[65308]= -1184318708;
assign addr[65309]= -917951481;
assign addr[65310]= -632981917;
assign addr[65311]= -335184940;
assign addr[65312]= -30595422;
assign addr[65313]= 274614114;
assign addr[65314]= 574258580;
assign addr[65315]= 862265664;
assign addr[65316]= 1132798888;
assign addr[65317]= 1380375881;
assign addr[65318]= 1599979481;
assign addr[65319]= 1787159411;
assign addr[65320]= 1938122457;
assign addr[65321]= 2049809346;
assign addr[65322]= 2119956737;
assign addr[65323]= 2147143090;
assign addr[65324]= 2130817471;
assign addr[65325]= 2071310720;
assign addr[65326]= 1969828744;
assign addr[65327]= 1828428082;
assign addr[65328]= 1649974225;
assign addr[65329]= 1438083551;
assign addr[65330]= 1197050035;
assign addr[65331]= 931758235;
assign addr[65332]= 647584304;
assign addr[65333]= 350287041;
assign addr[65334]= 45891193;
assign addr[65335]= -259434643;
assign addr[65336]= -559503022;
assign addr[65337]= -848233042;
assign addr[65338]= -1119773573;
assign addr[65339]= -1368621831;
assign addr[65340]= -1589734894;
assign addr[65341]= -1778631892;
assign addr[65342]= -1931484818;
assign addr[65343]= -2045196100;
assign addr[65344]= -2117461370;
assign addr[65345]= -2146816171;
assign addr[65346]= -2132665626;
assign addr[65347]= -2075296495;
assign addr[65348]= -1975871368;
assign addr[65349]= -1836405100;
assign addr[65350]= -1659723983;
assign addr[65351]= -1449408469;
assign addr[65352]= -1209720613;
assign addr[65353]= -945517704;
assign addr[65354]= -662153826;
assign addr[65355]= -365371365;
assign addr[65356]= -61184634;
assign addr[65357]= 244242007;
assign addr[65358]= 544719071;
assign addr[65359]= 834157373;
assign addr[65360]= 1106691431;
assign addr[65361]= 1356798326;
assign addr[65362]= 1579409630;
assign addr[65363]= 1770014111;
assign addr[65364]= 1924749160;
assign addr[65365]= 2040479063;
assign addr[65366]= 2114858546;
assign addr[65367]= 2146380306;
assign addr[65368]= 2134405552;
assign addr[65369]= 2079176953;
assign addr[65370]= 1981813720;
assign addr[65371]= 1844288924;
assign addr[65372]= 1669389513;
assign addr[65373]= 1460659832;
assign addr[65374]= 1222329801;
assign addr[65375]= 959229189;
assign addr[65376]= 676689746;
assign addr[65377]= 380437148;
assign addr[65378]= 76474970;
assign addr[65379]= -229036977;
assign addr[65380]= -529907477;
assign addr[65381]= -820039373;
assign addr[65382]= -1093553126;
assign addr[65383]= -1344905966;
assign addr[65384]= -1569004214;
assign addr[65385]= -1761306505;
assign addr[65386]= -1917915825;
assign addr[65387]= -2035658475;
assign addr[65388]= -2112148396;
assign addr[65389]= -2145835515;
assign addr[65390]= -2136037160;
assign addr[65391]= -2082951896;
assign addr[65392]= -1987655498;
assign addr[65393]= -1852079154;
assign addr[65394]= -1678970324;
assign addr[65395]= -1471837070;
assign addr[65396]= -1234876957;
assign addr[65397]= -972891995;
assign addr[65398]= -691191324;
assign addr[65399]= -395483624;
assign addr[65400]= -91761426;
assign addr[65401]= 213820322;
assign addr[65402]= 515068990;
assign addr[65403]= 805879757;
assign addr[65404]= 1080359326;
assign addr[65405]= 1332945355;
assign addr[65406]= 1558519173;
assign addr[65407]= 1752509516;
assign addr[65408]= 1910985158;
assign addr[65409]= 2030734582;
assign addr[65410]= 2109331059;
assign addr[65411]= 2145181827;
assign addr[65412]= 2137560369;
assign addr[65413]= 2086621133;
assign addr[65414]= 1993396407;
assign addr[65415]= 1859775393;
assign addr[65416]= 1688465931;
assign addr[65417]= 1482939614;
assign addr[65418]= 1247361445;
assign addr[65419]= 986505429;
assign addr[65420]= 705657826;
assign addr[65421]= 410510029;
assign addr[65422]= 107043224;
assign addr[65423]= -198592817;
assign addr[65424]= -500204365;
assign addr[65425]= -791679244;
assign addr[65426]= -1067110699;
assign addr[65427]= -1320917099;
assign addr[65428]= -1547955041;
assign addr[65429]= -1743623590;
assign addr[65430]= -1903957513;
assign addr[65431]= -2025707632;
assign addr[65432]= -2106406677;
assign addr[65433]= -2144419275;
assign addr[65434]= -2138975100;
assign addr[65435]= -2090184478;
assign addr[65436]= -1999036154;
assign addr[65437]= -1867377253;
assign addr[65438]= -1697875851;
assign addr[65439]= -1493966902;
assign addr[65440]= -1259782632;
assign addr[65441]= -1000068799;
assign addr[65442]= -720088517;
assign addr[65443]= -425515602;
assign addr[65444]= -122319591;
assign addr[65445]= 183355234;
assign addr[65446]= 485314355;
assign addr[65447]= 777438554;
assign addr[65448]= 1053807919;
assign addr[65449]= 1308821808;
assign addr[65450]= 1537312353;
assign addr[65451]= 1734649179;
assign addr[65452]= 1896833245;
assign addr[65453]= 2020577882;
assign addr[65454]= 2103375398;
assign addr[65455]= 2143547897;
assign addr[65456]= 2140281282;
assign addr[65457]= 2093641749;
assign addr[65458]= 2004574453;
assign addr[65459]= 1874884346;
assign addr[65460]= 1707199606;
assign addr[65461]= 1504918373;
assign addr[65462]= 1272139887;
assign addr[65463]= 1013581418;
assign addr[65464]= 734482665;
assign addr[65465]= 440499581;
assign addr[65466]= 137589750;
assign addr[65467]= -168108346;
assign addr[65468]= -470399716;
assign addr[65469]= -763158411;
assign addr[65470]= -1040451659;
assign addr[65471]= -1296660098;
assign addr[65472]= -1526591649;
assign addr[65473]= -1725586737;
assign addr[65474]= -1889612716;
assign addr[65475]= -2015345591;
assign addr[65476]= -2100237377;
assign addr[65477]= -2142567738;
assign addr[65478]= -2141478848;
assign addr[65479]= -2096992772;
assign addr[65480]= -2010011024;
assign addr[65481]= -1882296293;
assign addr[65482]= -1716436725;
assign addr[65483]= -1515793473;
assign addr[65484]= -1284432584;
assign addr[65485]= -1027042599;
assign addr[65486]= -748839539;
assign addr[65487]= -455461206;
assign addr[65488]= -152852926;
assign addr[65489]= 152852926;
assign addr[65490]= 455461206;
assign addr[65491]= 748839539;
assign addr[65492]= 1027042599;
assign addr[65493]= 1284432584;
assign addr[65494]= 1515793473;
assign addr[65495]= 1716436725;
assign addr[65496]= 1882296293;
assign addr[65497]= 2010011024;
assign addr[65498]= 2096992772;
assign addr[65499]= 2141478848;
assign addr[65500]= 2142567738;
assign addr[65501]= 2100237377;
assign addr[65502]= 2015345591;
assign addr[65503]= 1889612716;
assign addr[65504]= 1725586737;
assign addr[65505]= 1526591649;
assign addr[65506]= 1296660098;
assign addr[65507]= 1040451659;
assign addr[65508]= 763158411;
assign addr[65509]= 470399716;
assign addr[65510]= 168108346;
assign addr[65511]= -137589750;
assign addr[65512]= -440499581;
assign addr[65513]= -734482665;
assign addr[65514]= -1013581418;
assign addr[65515]= -1272139887;
assign addr[65516]= -1504918373;
assign addr[65517]= -1707199606;
assign addr[65518]= -1874884346;
assign addr[65519]= -2004574453;
assign addr[65520]= -2093641749;
assign addr[65521]= -2140281282;
assign addr[65522]= -2143547897;
assign addr[65523]= -2103375398;
assign addr[65524]= -2020577882;
assign addr[65525]= -1896833245;
assign addr[65526]= -1734649179;
assign addr[65527]= -1537312353;
assign addr[65528]= -1308821808;
assign addr[65529]= -1053807919;
assign addr[65530]= -777438554;
assign addr[65531]= -485314355;
assign addr[65532]= -183355234;
assign addr[65533]= 122319591;
assign addr[65534]= 425515602;
assign addr[65535]= 720088517;
endmodule