module rompcm88(
	input clk,//45m
	input reset_n,
	output signed [31:0]addrout
);

wire signed [31:0]addr[0:65535];
reg [8:0]k;
wire lrck;
always @(posedge clk or negedge reset_n)begin
	if(reset_n ==0) 
	k = 0;
	
	else
	k <= k+1;

end
assign lrck = k[8];
reg [15:0]i;
always @(posedge lrck or negedge reset_n)begin
	if(reset_n ==0)begin
		i <= 0;
	//	addrout <= 32'd0;
		end
	
	else begin
		i <= i+1;
	//	addrout <= addr[i];
		end
end

assign addrout = addr[i];
assign addr[0]= 0;
assign addr[1]= 152852926;
assign addr[2]= 304930476;
assign addr[3]= 455461206;
assign addr[4]= 603681519;
assign addr[5]= 748839539;
assign addr[6]= 890198924;
assign addr[7]= 1027042599;
assign addr[8]= 1158676398;
assign addr[9]= 1284432584;
assign addr[10]= 1403673233;
assign addr[11]= 1515793473;
assign addr[12]= 1620224553;
assign addr[13]= 1716436725;
assign addr[14]= 1803941934;
assign addr[15]= 1882296293;
assign addr[16]= 1951102334;
assign addr[17]= 2010011024;
assign addr[18]= 2058723538;
assign addr[19]= 2096992772;
assign addr[20]= 2124624598;
assign addr[21]= 2141478848;
assign addr[22]= 2147470025;
assign addr[23]= 2142567738;
assign addr[24]= 2126796855;
assign addr[25]= 2100237377;
assign addr[26]= 2063024031;
assign addr[27]= 2015345591;
assign addr[28]= 1957443913;
assign addr[29]= 1889612716;
assign addr[30]= 1812196087;
assign addr[31]= 1725586737;
assign addr[32]= 1630224009;
assign addr[33]= 1526591649;
assign addr[34]= 1415215352;
assign addr[35]= 1296660098;
assign addr[36]= 1171527280;
assign addr[37]= 1040451659;
assign addr[38]= 904098143;
assign addr[39]= 763158411;
assign addr[40]= 618347408;
assign addr[41]= 470399716;
assign addr[42]= 320065829;
assign addr[43]= 168108346;
assign addr[44]= 15298099;
assign addr[45]= -137589750;
assign addr[46]= -289779648;
assign addr[47]= -440499581;
assign addr[48]= -588984994;
assign addr[49]= -734482665;
assign addr[50]= -876254528;
assign addr[51]= -1013581418;
assign addr[52]= -1145766716;
assign addr[53]= -1272139887;
assign addr[54]= -1392059879;
assign addr[55]= -1504918373;
assign addr[56]= -1610142873;
assign addr[57]= -1707199606;
assign addr[58]= -1795596234;
assign addr[59]= -1874884346;
assign addr[60]= -1944661739;
assign addr[61]= -2004574453;
assign addr[62]= -2054318569;
assign addr[63]= -2093641749;
assign addr[64]= -2122344521;
assign addr[65]= -2140281282;
assign addr[66]= -2147361045;
assign addr[67]= -2143547897;
assign addr[68]= -2128861181;
assign addr[69]= -2103375398;
assign addr[70]= -2067219829;
assign addr[71]= -2020577882;
assign addr[72]= -1963686155;
assign addr[73]= -1896833245;
assign addr[74]= -1820358275;
assign addr[75]= -1734649179;
assign addr[76]= -1640140734;
assign addr[77]= -1537312353;
assign addr[78]= -1426685652;
assign addr[79]= -1308821808;
assign addr[80]= -1184318708;
assign addr[81]= -1053807919;
assign addr[82]= -917951481;
assign addr[83]= -777438554;
assign addr[84]= -632981917;
assign addr[85]= -485314355;
assign addr[86]= -335184940;
assign addr[87]= -183355234;
assign addr[88]= -30595422;
assign addr[89]= 122319591;
assign addr[90]= 274614114;
assign addr[91]= 425515602;
assign addr[92]= 574258580;
assign addr[93]= 720088517;
assign addr[94]= 862265664;
assign addr[95]= 1000068799;
assign addr[96]= 1132798888;
assign addr[97]= 1259782632;
assign addr[98]= 1380375881;
assign addr[99]= 1493966902;
assign addr[100]= 1599979481;
assign addr[101]= 1697875851;
assign addr[102]= 1787159411;
assign addr[103]= 1867377253;
assign addr[104]= 1938122457;
assign addr[105]= 1999036154;
assign addr[106]= 2049809346;
assign addr[107]= 2090184478;
assign addr[108]= 2119956737;
assign addr[109]= 2138975100;
assign addr[110]= 2147143090;
assign addr[111]= 2144419275;
assign addr[112]= 2130817471;
assign addr[113]= 2106406677;
assign addr[114]= 2071310720;
assign addr[115]= 2025707632;
assign addr[116]= 1969828744;
assign addr[117]= 1903957513;
assign addr[118]= 1828428082;
assign addr[119]= 1743623590;
assign addr[120]= 1649974225;
assign addr[121]= 1547955041;
assign addr[122]= 1438083551;
assign addr[123]= 1320917099;
assign addr[124]= 1197050035;
assign addr[125]= 1067110699;
assign addr[126]= 931758235;
assign addr[127]= 791679244;
assign addr[128]= 647584304;
assign addr[129]= 500204365;
assign addr[130]= 350287041;
assign addr[131]= 198592817;
assign addr[132]= 45891193;
assign addr[133]= -107043224;
assign addr[134]= -259434643;
assign addr[135]= -410510029;
assign addr[136]= -559503022;
assign addr[137]= -705657826;
assign addr[138]= -848233042;
assign addr[139]= -986505429;
assign addr[140]= -1119773573;
assign addr[141]= -1247361445;
assign addr[142]= -1368621831;
assign addr[143]= -1482939614;
assign addr[144]= -1589734894;
assign addr[145]= -1688465931;
assign addr[146]= -1778631892;
assign addr[147]= -1859775393;
assign addr[148]= -1931484818;
assign addr[149]= -1993396407;
assign addr[150]= -2045196100;
assign addr[151]= -2086621133;
assign addr[152]= -2117461370;
assign addr[153]= -2137560369;
assign addr[154]= -2146816171;
assign addr[155]= -2145181827;
assign addr[156]= -2132665626;
assign addr[157]= -2109331059;
assign addr[158]= -2075296495;
assign addr[159]= -2030734582;
assign addr[160]= -1975871368;
assign addr[161]= -1910985158;
assign addr[162]= -1836405100;
assign addr[163]= -1752509516;
assign addr[164]= -1659723983;
assign addr[165]= -1558519173;
assign addr[166]= -1449408469;
assign addr[167]= -1332945355;
assign addr[168]= -1209720613;
assign addr[169]= -1080359326;
assign addr[170]= -945517704;
assign addr[171]= -805879757;
assign addr[172]= -662153826;
assign addr[173]= -515068990;
assign addr[174]= -365371365;
assign addr[175]= -213820322;
assign addr[176]= -61184634;
assign addr[177]= 91761426;
assign addr[178]= 244242007;
assign addr[179]= 395483624;
assign addr[180]= 544719071;
assign addr[181]= 691191324;
assign addr[182]= 834157373;
assign addr[183]= 972891995;
assign addr[184]= 1106691431;
assign addr[185]= 1234876957;
assign addr[186]= 1356798326;
assign addr[187]= 1471837070;
assign addr[188]= 1579409630;
assign addr[189]= 1678970324;
assign addr[190]= 1770014111;
assign addr[191]= 1852079154;
assign addr[192]= 1924749160;
assign addr[193]= 1987655498;
assign addr[194]= 2040479063;
assign addr[195]= 2082951896;
assign addr[196]= 2114858546;
assign addr[197]= 2136037160;
assign addr[198]= 2146380306;
assign addr[199]= 2145835515;
assign addr[200]= 2134405552;
assign addr[201]= 2112148396;
assign addr[202]= 2079176953;
assign addr[203]= 2035658475;
assign addr[204]= 1981813720;
assign addr[205]= 1917915825;
assign addr[206]= 1844288924;
assign addr[207]= 1761306505;
assign addr[208]= 1669389513;
assign addr[209]= 1569004214;
assign addr[210]= 1460659832;
assign addr[211]= 1344905966;
assign addr[212]= 1222329801;
assign addr[213]= 1093553126;
assign addr[214]= 959229189;
assign addr[215]= 820039373;
assign addr[216]= 676689746;
assign addr[217]= 529907477;
assign addr[218]= 380437148;
assign addr[219]= 229036977;
assign addr[220]= 76474970;
assign addr[221]= -76474970;
assign addr[222]= -229036977;
assign addr[223]= -380437148;
assign addr[224]= -529907477;
assign addr[225]= -676689746;
assign addr[226]= -820039373;
assign addr[227]= -959229189;
assign addr[228]= -1093553126;
assign addr[229]= -1222329801;
assign addr[230]= -1344905966;
assign addr[231]= -1460659832;
assign addr[232]= -1569004214;
assign addr[233]= -1669389513;
assign addr[234]= -1761306505;
assign addr[235]= -1844288924;
assign addr[236]= -1917915825;
assign addr[237]= -1981813720;
assign addr[238]= -2035658475;
assign addr[239]= -2079176953;
assign addr[240]= -2112148396;
assign addr[241]= -2134405552;
assign addr[242]= -2145835515;
assign addr[243]= -2146380306;
assign addr[244]= -2136037160;
assign addr[245]= -2114858546;
assign addr[246]= -2082951896;
assign addr[247]= -2040479063;
assign addr[248]= -1987655498;
assign addr[249]= -1924749160;
assign addr[250]= -1852079154;
assign addr[251]= -1770014111;
assign addr[252]= -1678970324;
assign addr[253]= -1579409630;
assign addr[254]= -1471837070;
assign addr[255]= -1356798326;
assign addr[256]= -1234876957;
assign addr[257]= -1106691431;
assign addr[258]= -972891995;
assign addr[259]= -834157373;
assign addr[260]= -691191324;
assign addr[261]= -544719071;
assign addr[262]= -395483624;
assign addr[263]= -244242007;
assign addr[264]= -91761426;
assign addr[265]= 61184634;
assign addr[266]= 213820322;
assign addr[267]= 365371365;
assign addr[268]= 515068990;
assign addr[269]= 662153826;
assign addr[270]= 805879757;
assign addr[271]= 945517704;
assign addr[272]= 1080359326;
assign addr[273]= 1209720613;
assign addr[274]= 1332945355;
assign addr[275]= 1449408469;
assign addr[276]= 1558519173;
assign addr[277]= 1659723983;
assign addr[278]= 1752509516;
assign addr[279]= 1836405100;
assign addr[280]= 1910985158;
assign addr[281]= 1975871368;
assign addr[282]= 2030734582;
assign addr[283]= 2075296495;
assign addr[284]= 2109331059;
assign addr[285]= 2132665626;
assign addr[286]= 2145181827;
assign addr[287]= 2146816171;
assign addr[288]= 2137560369;
assign addr[289]= 2117461370;
assign addr[290]= 2086621133;
assign addr[291]= 2045196100;
assign addr[292]= 1993396407;
assign addr[293]= 1931484818;
assign addr[294]= 1859775393;
assign addr[295]= 1778631892;
assign addr[296]= 1688465931;
assign addr[297]= 1589734894;
assign addr[298]= 1482939614;
assign addr[299]= 1368621831;
assign addr[300]= 1247361445;
assign addr[301]= 1119773573;
assign addr[302]= 986505429;
assign addr[303]= 848233042;
assign addr[304]= 705657826;
assign addr[305]= 559503022;
assign addr[306]= 410510029;
assign addr[307]= 259434643;
assign addr[308]= 107043224;
assign addr[309]= -45891193;
assign addr[310]= -198592817;
assign addr[311]= -350287041;
assign addr[312]= -500204365;
assign addr[313]= -647584304;
assign addr[314]= -791679244;
assign addr[315]= -931758235;
assign addr[316]= -1067110699;
assign addr[317]= -1197050035;
assign addr[318]= -1320917099;
assign addr[319]= -1438083551;
assign addr[320]= -1547955041;
assign addr[321]= -1649974225;
assign addr[322]= -1743623590;
assign addr[323]= -1828428082;
assign addr[324]= -1903957513;
assign addr[325]= -1969828744;
assign addr[326]= -2025707632;
assign addr[327]= -2071310720;
assign addr[328]= -2106406677;
assign addr[329]= -2130817471;
assign addr[330]= -2144419275;
assign addr[331]= -2147143090;
assign addr[332]= -2138975100;
assign addr[333]= -2119956737;
assign addr[334]= -2090184478;
assign addr[335]= -2049809346;
assign addr[336]= -1999036154;
assign addr[337]= -1938122457;
assign addr[338]= -1867377253;
assign addr[339]= -1787159411;
assign addr[340]= -1697875851;
assign addr[341]= -1599979481;
assign addr[342]= -1493966902;
assign addr[343]= -1380375881;
assign addr[344]= -1259782632;
assign addr[345]= -1132798888;
assign addr[346]= -1000068799;
assign addr[347]= -862265664;
assign addr[348]= -720088517;
assign addr[349]= -574258580;
assign addr[350]= -425515602;
assign addr[351]= -274614114;
assign addr[352]= -122319591;
assign addr[353]= 30595422;
assign addr[354]= 183355234;
assign addr[355]= 335184940;
assign addr[356]= 485314355;
assign addr[357]= 632981917;
assign addr[358]= 777438554;
assign addr[359]= 917951481;
assign addr[360]= 1053807919;
assign addr[361]= 1184318708;
assign addr[362]= 1308821808;
assign addr[363]= 1426685652;
assign addr[364]= 1537312353;
assign addr[365]= 1640140734;
assign addr[366]= 1734649179;
assign addr[367]= 1820358275;
assign addr[368]= 1896833245;
assign addr[369]= 1963686155;
assign addr[370]= 2020577882;
assign addr[371]= 2067219829;
assign addr[372]= 2103375398;
assign addr[373]= 2128861181;
assign addr[374]= 2143547897;
assign addr[375]= 2147361045;
assign addr[376]= 2140281282;
assign addr[377]= 2122344521;
assign addr[378]= 2093641749;
assign addr[379]= 2054318569;
assign addr[380]= 2004574453;
assign addr[381]= 1944661739;
assign addr[382]= 1874884346;
assign addr[383]= 1795596234;
assign addr[384]= 1707199606;
assign addr[385]= 1610142873;
assign addr[386]= 1504918373;
assign addr[387]= 1392059879;
assign addr[388]= 1272139887;
assign addr[389]= 1145766716;
assign addr[390]= 1013581418;
assign addr[391]= 876254528;
assign addr[392]= 734482665;
assign addr[393]= 588984994;
assign addr[394]= 440499581;
assign addr[395]= 289779648;
assign addr[396]= 137589750;
assign addr[397]= -15298099;
assign addr[398]= -168108346;
assign addr[399]= -320065829;
assign addr[400]= -470399716;
assign addr[401]= -618347408;
assign addr[402]= -763158411;
assign addr[403]= -904098143;
assign addr[404]= -1040451659;
assign addr[405]= -1171527280;
assign addr[406]= -1296660098;
assign addr[407]= -1415215352;
assign addr[408]= -1526591649;
assign addr[409]= -1630224009;
assign addr[410]= -1725586737;
assign addr[411]= -1812196087;
assign addr[412]= -1889612716;
assign addr[413]= -1957443913;
assign addr[414]= -2015345591;
assign addr[415]= -2063024031;
assign addr[416]= -2100237377;
assign addr[417]= -2126796855;
assign addr[418]= -2142567738;
assign addr[419]= -2147470025;
assign addr[420]= -2141478848;
assign addr[421]= -2124624598;
assign addr[422]= -2096992772;
assign addr[423]= -2058723538;
assign addr[424]= -2010011024;
assign addr[425]= -1951102334;
assign addr[426]= -1882296293;
assign addr[427]= -1803941934;
assign addr[428]= -1716436725;
assign addr[429]= -1620224553;
assign addr[430]= -1515793473;
assign addr[431]= -1403673233;
assign addr[432]= -1284432584;
assign addr[433]= -1158676398;
assign addr[434]= -1027042599;
assign addr[435]= -890198924;
assign addr[436]= -748839539;
assign addr[437]= -603681519;
assign addr[438]= -455461206;
assign addr[439]= -304930476;
assign addr[440]= -152852926;
assign addr[441]= 0;
assign addr[442]= 152852926;
assign addr[443]= 304930476;
assign addr[444]= 455461206;
assign addr[445]= 603681519;
assign addr[446]= 748839539;
assign addr[447]= 890198924;
assign addr[448]= 1027042599;
assign addr[449]= 1158676398;
assign addr[450]= 1284432584;
assign addr[451]= 1403673233;
assign addr[452]= 1515793473;
assign addr[453]= 1620224553;
assign addr[454]= 1716436725;
assign addr[455]= 1803941934;
assign addr[456]= 1882296293;
assign addr[457]= 1951102334;
assign addr[458]= 2010011024;
assign addr[459]= 2058723538;
assign addr[460]= 2096992772;
assign addr[461]= 2124624598;
assign addr[462]= 2141478848;
assign addr[463]= 2147470025;
assign addr[464]= 2142567738;
assign addr[465]= 2126796855;
assign addr[466]= 2100237377;
assign addr[467]= 2063024031;
assign addr[468]= 2015345591;
assign addr[469]= 1957443913;
assign addr[470]= 1889612716;
assign addr[471]= 1812196087;
assign addr[472]= 1725586737;
assign addr[473]= 1630224009;
assign addr[474]= 1526591649;
assign addr[475]= 1415215352;
assign addr[476]= 1296660098;
assign addr[477]= 1171527280;
assign addr[478]= 1040451659;
assign addr[479]= 904098143;
assign addr[480]= 763158411;
assign addr[481]= 618347408;
assign addr[482]= 470399716;
assign addr[483]= 320065829;
assign addr[484]= 168108346;
assign addr[485]= 15298099;
assign addr[486]= -137589750;
assign addr[487]= -289779648;
assign addr[488]= -440499581;
assign addr[489]= -588984994;
assign addr[490]= -734482665;
assign addr[491]= -876254528;
assign addr[492]= -1013581418;
assign addr[493]= -1145766716;
assign addr[494]= -1272139887;
assign addr[495]= -1392059879;
assign addr[496]= -1504918373;
assign addr[497]= -1610142873;
assign addr[498]= -1707199606;
assign addr[499]= -1795596234;
assign addr[500]= -1874884346;
assign addr[501]= -1944661739;
assign addr[502]= -2004574453;
assign addr[503]= -2054318569;
assign addr[504]= -2093641749;
assign addr[505]= -2122344521;
assign addr[506]= -2140281282;
assign addr[507]= -2147361045;
assign addr[508]= -2143547897;
assign addr[509]= -2128861181;
assign addr[510]= -2103375398;
assign addr[511]= -2067219829;
assign addr[512]= -2020577882;
assign addr[513]= -1963686155;
assign addr[514]= -1896833245;
assign addr[515]= -1820358275;
assign addr[516]= -1734649179;
assign addr[517]= -1640140734;
assign addr[518]= -1537312353;
assign addr[519]= -1426685652;
assign addr[520]= -1308821808;
assign addr[521]= -1184318708;
assign addr[522]= -1053807919;
assign addr[523]= -917951481;
assign addr[524]= -777438554;
assign addr[525]= -632981917;
assign addr[526]= -485314355;
assign addr[527]= -335184940;
assign addr[528]= -183355234;
assign addr[529]= -30595422;
assign addr[530]= 122319591;
assign addr[531]= 274614114;
assign addr[532]= 425515602;
assign addr[533]= 574258580;
assign addr[534]= 720088517;
assign addr[535]= 862265664;
assign addr[536]= 1000068799;
assign addr[537]= 1132798888;
assign addr[538]= 1259782632;
assign addr[539]= 1380375881;
assign addr[540]= 1493966902;
assign addr[541]= 1599979481;
assign addr[542]= 1697875851;
assign addr[543]= 1787159411;
assign addr[544]= 1867377253;
assign addr[545]= 1938122457;
assign addr[546]= 1999036154;
assign addr[547]= 2049809346;
assign addr[548]= 2090184478;
assign addr[549]= 2119956737;
assign addr[550]= 2138975100;
assign addr[551]= 2147143090;
assign addr[552]= 2144419275;
assign addr[553]= 2130817471;
assign addr[554]= 2106406677;
assign addr[555]= 2071310720;
assign addr[556]= 2025707632;
assign addr[557]= 1969828744;
assign addr[558]= 1903957513;
assign addr[559]= 1828428082;
assign addr[560]= 1743623590;
assign addr[561]= 1649974225;
assign addr[562]= 1547955041;
assign addr[563]= 1438083551;
assign addr[564]= 1320917099;
assign addr[565]= 1197050035;
assign addr[566]= 1067110699;
assign addr[567]= 931758235;
assign addr[568]= 791679244;
assign addr[569]= 647584304;
assign addr[570]= 500204365;
assign addr[571]= 350287041;
assign addr[572]= 198592817;
assign addr[573]= 45891193;
assign addr[574]= -107043224;
assign addr[575]= -259434643;
assign addr[576]= -410510029;
assign addr[577]= -559503022;
assign addr[578]= -705657826;
assign addr[579]= -848233042;
assign addr[580]= -986505429;
assign addr[581]= -1119773573;
assign addr[582]= -1247361445;
assign addr[583]= -1368621831;
assign addr[584]= -1482939614;
assign addr[585]= -1589734894;
assign addr[586]= -1688465931;
assign addr[587]= -1778631892;
assign addr[588]= -1859775393;
assign addr[589]= -1931484818;
assign addr[590]= -1993396407;
assign addr[591]= -2045196100;
assign addr[592]= -2086621133;
assign addr[593]= -2117461370;
assign addr[594]= -2137560369;
assign addr[595]= -2146816171;
assign addr[596]= -2145181827;
assign addr[597]= -2132665626;
assign addr[598]= -2109331059;
assign addr[599]= -2075296495;
assign addr[600]= -2030734582;
assign addr[601]= -1975871368;
assign addr[602]= -1910985158;
assign addr[603]= -1836405100;
assign addr[604]= -1752509516;
assign addr[605]= -1659723983;
assign addr[606]= -1558519173;
assign addr[607]= -1449408469;
assign addr[608]= -1332945355;
assign addr[609]= -1209720613;
assign addr[610]= -1080359326;
assign addr[611]= -945517704;
assign addr[612]= -805879757;
assign addr[613]= -662153826;
assign addr[614]= -515068990;
assign addr[615]= -365371365;
assign addr[616]= -213820322;
assign addr[617]= -61184634;
assign addr[618]= 91761426;
assign addr[619]= 244242007;
assign addr[620]= 395483624;
assign addr[621]= 544719071;
assign addr[622]= 691191324;
assign addr[623]= 834157373;
assign addr[624]= 972891995;
assign addr[625]= 1106691431;
assign addr[626]= 1234876957;
assign addr[627]= 1356798326;
assign addr[628]= 1471837070;
assign addr[629]= 1579409630;
assign addr[630]= 1678970324;
assign addr[631]= 1770014111;
assign addr[632]= 1852079154;
assign addr[633]= 1924749160;
assign addr[634]= 1987655498;
assign addr[635]= 2040479063;
assign addr[636]= 2082951896;
assign addr[637]= 2114858546;
assign addr[638]= 2136037160;
assign addr[639]= 2146380306;
assign addr[640]= 2145835515;
assign addr[641]= 2134405552;
assign addr[642]= 2112148396;
assign addr[643]= 2079176953;
assign addr[644]= 2035658475;
assign addr[645]= 1981813720;
assign addr[646]= 1917915825;
assign addr[647]= 1844288924;
assign addr[648]= 1761306505;
assign addr[649]= 1669389513;
assign addr[650]= 1569004214;
assign addr[651]= 1460659832;
assign addr[652]= 1344905966;
assign addr[653]= 1222329801;
assign addr[654]= 1093553126;
assign addr[655]= 959229189;
assign addr[656]= 820039373;
assign addr[657]= 676689746;
assign addr[658]= 529907477;
assign addr[659]= 380437148;
assign addr[660]= 229036977;
assign addr[661]= 76474970;
assign addr[662]= -76474970;
assign addr[663]= -229036977;
assign addr[664]= -380437148;
assign addr[665]= -529907477;
assign addr[666]= -676689746;
assign addr[667]= -820039373;
assign addr[668]= -959229189;
assign addr[669]= -1093553126;
assign addr[670]= -1222329801;
assign addr[671]= -1344905966;
assign addr[672]= -1460659832;
assign addr[673]= -1569004214;
assign addr[674]= -1669389513;
assign addr[675]= -1761306505;
assign addr[676]= -1844288924;
assign addr[677]= -1917915825;
assign addr[678]= -1981813720;
assign addr[679]= -2035658475;
assign addr[680]= -2079176953;
assign addr[681]= -2112148396;
assign addr[682]= -2134405552;
assign addr[683]= -2145835515;
assign addr[684]= -2146380306;
assign addr[685]= -2136037160;
assign addr[686]= -2114858546;
assign addr[687]= -2082951896;
assign addr[688]= -2040479063;
assign addr[689]= -1987655498;
assign addr[690]= -1924749160;
assign addr[691]= -1852079154;
assign addr[692]= -1770014111;
assign addr[693]= -1678970324;
assign addr[694]= -1579409630;
assign addr[695]= -1471837070;
assign addr[696]= -1356798326;
assign addr[697]= -1234876957;
assign addr[698]= -1106691431;
assign addr[699]= -972891995;
assign addr[700]= -834157373;
assign addr[701]= -691191324;
assign addr[702]= -544719071;
assign addr[703]= -395483624;
assign addr[704]= -244242007;
assign addr[705]= -91761426;
assign addr[706]= 61184634;
assign addr[707]= 213820322;
assign addr[708]= 365371365;
assign addr[709]= 515068990;
assign addr[710]= 662153826;
assign addr[711]= 805879757;
assign addr[712]= 945517704;
assign addr[713]= 1080359326;
assign addr[714]= 1209720613;
assign addr[715]= 1332945355;
assign addr[716]= 1449408469;
assign addr[717]= 1558519173;
assign addr[718]= 1659723983;
assign addr[719]= 1752509516;
assign addr[720]= 1836405100;
assign addr[721]= 1910985158;
assign addr[722]= 1975871368;
assign addr[723]= 2030734582;
assign addr[724]= 2075296495;
assign addr[725]= 2109331059;
assign addr[726]= 2132665626;
assign addr[727]= 2145181827;
assign addr[728]= 2146816171;
assign addr[729]= 2137560369;
assign addr[730]= 2117461370;
assign addr[731]= 2086621133;
assign addr[732]= 2045196100;
assign addr[733]= 1993396407;
assign addr[734]= 1931484818;
assign addr[735]= 1859775393;
assign addr[736]= 1778631892;
assign addr[737]= 1688465931;
assign addr[738]= 1589734894;
assign addr[739]= 1482939614;
assign addr[740]= 1368621831;
assign addr[741]= 1247361445;
assign addr[742]= 1119773573;
assign addr[743]= 986505429;
assign addr[744]= 848233042;
assign addr[745]= 705657826;
assign addr[746]= 559503022;
assign addr[747]= 410510029;
assign addr[748]= 259434643;
assign addr[749]= 107043224;
assign addr[750]= -45891193;
assign addr[751]= -198592817;
assign addr[752]= -350287041;
assign addr[753]= -500204365;
assign addr[754]= -647584304;
assign addr[755]= -791679244;
assign addr[756]= -931758235;
assign addr[757]= -1067110699;
assign addr[758]= -1197050035;
assign addr[759]= -1320917099;
assign addr[760]= -1438083551;
assign addr[761]= -1547955041;
assign addr[762]= -1649974225;
assign addr[763]= -1743623590;
assign addr[764]= -1828428082;
assign addr[765]= -1903957513;
assign addr[766]= -1969828744;
assign addr[767]= -2025707632;
assign addr[768]= -2071310720;
assign addr[769]= -2106406677;
assign addr[770]= -2130817471;
assign addr[771]= -2144419275;
assign addr[772]= -2147143090;
assign addr[773]= -2138975100;
assign addr[774]= -2119956737;
assign addr[775]= -2090184478;
assign addr[776]= -2049809346;
assign addr[777]= -1999036154;
assign addr[778]= -1938122457;
assign addr[779]= -1867377253;
assign addr[780]= -1787159411;
assign addr[781]= -1697875851;
assign addr[782]= -1599979481;
assign addr[783]= -1493966902;
assign addr[784]= -1380375881;
assign addr[785]= -1259782632;
assign addr[786]= -1132798888;
assign addr[787]= -1000068799;
assign addr[788]= -862265664;
assign addr[789]= -720088517;
assign addr[790]= -574258580;
assign addr[791]= -425515602;
assign addr[792]= -274614114;
assign addr[793]= -122319591;
assign addr[794]= 30595422;
assign addr[795]= 183355234;
assign addr[796]= 335184940;
assign addr[797]= 485314355;
assign addr[798]= 632981917;
assign addr[799]= 777438554;
assign addr[800]= 917951481;
assign addr[801]= 1053807919;
assign addr[802]= 1184318708;
assign addr[803]= 1308821808;
assign addr[804]= 1426685652;
assign addr[805]= 1537312353;
assign addr[806]= 1640140734;
assign addr[807]= 1734649179;
assign addr[808]= 1820358275;
assign addr[809]= 1896833245;
assign addr[810]= 1963686155;
assign addr[811]= 2020577882;
assign addr[812]= 2067219829;
assign addr[813]= 2103375398;
assign addr[814]= 2128861181;
assign addr[815]= 2143547897;
assign addr[816]= 2147361045;
assign addr[817]= 2140281282;
assign addr[818]= 2122344521;
assign addr[819]= 2093641749;
assign addr[820]= 2054318569;
assign addr[821]= 2004574453;
assign addr[822]= 1944661739;
assign addr[823]= 1874884346;
assign addr[824]= 1795596234;
assign addr[825]= 1707199606;
assign addr[826]= 1610142873;
assign addr[827]= 1504918373;
assign addr[828]= 1392059879;
assign addr[829]= 1272139887;
assign addr[830]= 1145766716;
assign addr[831]= 1013581418;
assign addr[832]= 876254528;
assign addr[833]= 734482665;
assign addr[834]= 588984994;
assign addr[835]= 440499581;
assign addr[836]= 289779648;
assign addr[837]= 137589750;
assign addr[838]= -15298099;
assign addr[839]= -168108346;
assign addr[840]= -320065829;
assign addr[841]= -470399716;
assign addr[842]= -618347408;
assign addr[843]= -763158411;
assign addr[844]= -904098143;
assign addr[845]= -1040451659;
assign addr[846]= -1171527280;
assign addr[847]= -1296660098;
assign addr[848]= -1415215352;
assign addr[849]= -1526591649;
assign addr[850]= -1630224009;
assign addr[851]= -1725586737;
assign addr[852]= -1812196087;
assign addr[853]= -1889612716;
assign addr[854]= -1957443913;
assign addr[855]= -2015345591;
assign addr[856]= -2063024031;
assign addr[857]= -2100237377;
assign addr[858]= -2126796855;
assign addr[859]= -2142567738;
assign addr[860]= -2147470025;
assign addr[861]= -2141478848;
assign addr[862]= -2124624598;
assign addr[863]= -2096992772;
assign addr[864]= -2058723538;
assign addr[865]= -2010011024;
assign addr[866]= -1951102334;
assign addr[867]= -1882296293;
assign addr[868]= -1803941934;
assign addr[869]= -1716436725;
assign addr[870]= -1620224553;
assign addr[871]= -1515793473;
assign addr[872]= -1403673233;
assign addr[873]= -1284432584;
assign addr[874]= -1158676398;
assign addr[875]= -1027042599;
assign addr[876]= -890198924;
assign addr[877]= -748839539;
assign addr[878]= -603681519;
assign addr[879]= -455461206;
assign addr[880]= -304930476;
assign addr[881]= -152852926;
assign addr[882]= 0;
assign addr[883]= 152852926;
assign addr[884]= 304930476;
assign addr[885]= 455461206;
assign addr[886]= 603681519;
assign addr[887]= 748839539;
assign addr[888]= 890198924;
assign addr[889]= 1027042599;
assign addr[890]= 1158676398;
assign addr[891]= 1284432584;
assign addr[892]= 1403673233;
assign addr[893]= 1515793473;
assign addr[894]= 1620224553;
assign addr[895]= 1716436725;
assign addr[896]= 1803941934;
assign addr[897]= 1882296293;
assign addr[898]= 1951102334;
assign addr[899]= 2010011024;
assign addr[900]= 2058723538;
assign addr[901]= 2096992772;
assign addr[902]= 2124624598;
assign addr[903]= 2141478848;
assign addr[904]= 2147470025;
assign addr[905]= 2142567738;
assign addr[906]= 2126796855;
assign addr[907]= 2100237377;
assign addr[908]= 2063024031;
assign addr[909]= 2015345591;
assign addr[910]= 1957443913;
assign addr[911]= 1889612716;
assign addr[912]= 1812196087;
assign addr[913]= 1725586737;
assign addr[914]= 1630224009;
assign addr[915]= 1526591649;
assign addr[916]= 1415215352;
assign addr[917]= 1296660098;
assign addr[918]= 1171527280;
assign addr[919]= 1040451659;
assign addr[920]= 904098143;
assign addr[921]= 763158411;
assign addr[922]= 618347408;
assign addr[923]= 470399716;
assign addr[924]= 320065829;
assign addr[925]= 168108346;
assign addr[926]= 15298099;
assign addr[927]= -137589750;
assign addr[928]= -289779648;
assign addr[929]= -440499581;
assign addr[930]= -588984994;
assign addr[931]= -734482665;
assign addr[932]= -876254528;
assign addr[933]= -1013581418;
assign addr[934]= -1145766716;
assign addr[935]= -1272139887;
assign addr[936]= -1392059879;
assign addr[937]= -1504918373;
assign addr[938]= -1610142873;
assign addr[939]= -1707199606;
assign addr[940]= -1795596234;
assign addr[941]= -1874884346;
assign addr[942]= -1944661739;
assign addr[943]= -2004574453;
assign addr[944]= -2054318569;
assign addr[945]= -2093641749;
assign addr[946]= -2122344521;
assign addr[947]= -2140281282;
assign addr[948]= -2147361045;
assign addr[949]= -2143547897;
assign addr[950]= -2128861181;
assign addr[951]= -2103375398;
assign addr[952]= -2067219829;
assign addr[953]= -2020577882;
assign addr[954]= -1963686155;
assign addr[955]= -1896833245;
assign addr[956]= -1820358275;
assign addr[957]= -1734649179;
assign addr[958]= -1640140734;
assign addr[959]= -1537312353;
assign addr[960]= -1426685652;
assign addr[961]= -1308821808;
assign addr[962]= -1184318708;
assign addr[963]= -1053807919;
assign addr[964]= -917951481;
assign addr[965]= -777438554;
assign addr[966]= -632981917;
assign addr[967]= -485314355;
assign addr[968]= -335184940;
assign addr[969]= -183355234;
assign addr[970]= -30595422;
assign addr[971]= 122319591;
assign addr[972]= 274614114;
assign addr[973]= 425515602;
assign addr[974]= 574258580;
assign addr[975]= 720088517;
assign addr[976]= 862265664;
assign addr[977]= 1000068799;
assign addr[978]= 1132798888;
assign addr[979]= 1259782632;
assign addr[980]= 1380375881;
assign addr[981]= 1493966902;
assign addr[982]= 1599979481;
assign addr[983]= 1697875851;
assign addr[984]= 1787159411;
assign addr[985]= 1867377253;
assign addr[986]= 1938122457;
assign addr[987]= 1999036154;
assign addr[988]= 2049809346;
assign addr[989]= 2090184478;
assign addr[990]= 2119956737;
assign addr[991]= 2138975100;
assign addr[992]= 2147143090;
assign addr[993]= 2144419275;
assign addr[994]= 2130817471;
assign addr[995]= 2106406677;
assign addr[996]= 2071310720;
assign addr[997]= 2025707632;
assign addr[998]= 1969828744;
assign addr[999]= 1903957513;
assign addr[1000]= 1828428082;
assign addr[1001]= 1743623590;
assign addr[1002]= 1649974225;
assign addr[1003]= 1547955041;
assign addr[1004]= 1438083551;
assign addr[1005]= 1320917099;
assign addr[1006]= 1197050035;
assign addr[1007]= 1067110699;
assign addr[1008]= 931758235;
assign addr[1009]= 791679244;
assign addr[1010]= 647584304;
assign addr[1011]= 500204365;
assign addr[1012]= 350287041;
assign addr[1013]= 198592817;
assign addr[1014]= 45891193;
assign addr[1015]= -107043224;
assign addr[1016]= -259434643;
assign addr[1017]= -410510029;
assign addr[1018]= -559503022;
assign addr[1019]= -705657826;
assign addr[1020]= -848233042;
assign addr[1021]= -986505429;
assign addr[1022]= -1119773573;
assign addr[1023]= -1247361445;
assign addr[1024]= -1368621831;
assign addr[1025]= -1482939614;
assign addr[1026]= -1589734894;
assign addr[1027]= -1688465931;
assign addr[1028]= -1778631892;
assign addr[1029]= -1859775393;
assign addr[1030]= -1931484818;
assign addr[1031]= -1993396407;
assign addr[1032]= -2045196100;
assign addr[1033]= -2086621133;
assign addr[1034]= -2117461370;
assign addr[1035]= -2137560369;
assign addr[1036]= -2146816171;
assign addr[1037]= -2145181827;
assign addr[1038]= -2132665626;
assign addr[1039]= -2109331059;
assign addr[1040]= -2075296495;
assign addr[1041]= -2030734582;
assign addr[1042]= -1975871368;
assign addr[1043]= -1910985158;
assign addr[1044]= -1836405100;
assign addr[1045]= -1752509516;
assign addr[1046]= -1659723983;
assign addr[1047]= -1558519173;
assign addr[1048]= -1449408469;
assign addr[1049]= -1332945355;
assign addr[1050]= -1209720613;
assign addr[1051]= -1080359326;
assign addr[1052]= -945517704;
assign addr[1053]= -805879757;
assign addr[1054]= -662153826;
assign addr[1055]= -515068990;
assign addr[1056]= -365371365;
assign addr[1057]= -213820322;
assign addr[1058]= -61184634;
assign addr[1059]= 91761426;
assign addr[1060]= 244242007;
assign addr[1061]= 395483624;
assign addr[1062]= 544719071;
assign addr[1063]= 691191324;
assign addr[1064]= 834157373;
assign addr[1065]= 972891995;
assign addr[1066]= 1106691431;
assign addr[1067]= 1234876957;
assign addr[1068]= 1356798326;
assign addr[1069]= 1471837070;
assign addr[1070]= 1579409630;
assign addr[1071]= 1678970324;
assign addr[1072]= 1770014111;
assign addr[1073]= 1852079154;
assign addr[1074]= 1924749160;
assign addr[1075]= 1987655498;
assign addr[1076]= 2040479063;
assign addr[1077]= 2082951896;
assign addr[1078]= 2114858546;
assign addr[1079]= 2136037160;
assign addr[1080]= 2146380306;
assign addr[1081]= 2145835515;
assign addr[1082]= 2134405552;
assign addr[1083]= 2112148396;
assign addr[1084]= 2079176953;
assign addr[1085]= 2035658475;
assign addr[1086]= 1981813720;
assign addr[1087]= 1917915825;
assign addr[1088]= 1844288924;
assign addr[1089]= 1761306505;
assign addr[1090]= 1669389513;
assign addr[1091]= 1569004214;
assign addr[1092]= 1460659832;
assign addr[1093]= 1344905966;
assign addr[1094]= 1222329801;
assign addr[1095]= 1093553126;
assign addr[1096]= 959229189;
assign addr[1097]= 820039373;
assign addr[1098]= 676689746;
assign addr[1099]= 529907477;
assign addr[1100]= 380437148;
assign addr[1101]= 229036977;
assign addr[1102]= 76474970;
assign addr[1103]= -76474970;
assign addr[1104]= -229036977;
assign addr[1105]= -380437148;
assign addr[1106]= -529907477;
assign addr[1107]= -676689746;
assign addr[1108]= -820039373;
assign addr[1109]= -959229189;
assign addr[1110]= -1093553126;
assign addr[1111]= -1222329801;
assign addr[1112]= -1344905966;
assign addr[1113]= -1460659832;
assign addr[1114]= -1569004214;
assign addr[1115]= -1669389513;
assign addr[1116]= -1761306505;
assign addr[1117]= -1844288924;
assign addr[1118]= -1917915825;
assign addr[1119]= -1981813720;
assign addr[1120]= -2035658475;
assign addr[1121]= -2079176953;
assign addr[1122]= -2112148396;
assign addr[1123]= -2134405552;
assign addr[1124]= -2145835515;
assign addr[1125]= -2146380306;
assign addr[1126]= -2136037160;
assign addr[1127]= -2114858546;
assign addr[1128]= -2082951896;
assign addr[1129]= -2040479063;
assign addr[1130]= -1987655498;
assign addr[1131]= -1924749160;
assign addr[1132]= -1852079154;
assign addr[1133]= -1770014111;
assign addr[1134]= -1678970324;
assign addr[1135]= -1579409630;
assign addr[1136]= -1471837070;
assign addr[1137]= -1356798326;
assign addr[1138]= -1234876957;
assign addr[1139]= -1106691431;
assign addr[1140]= -972891995;
assign addr[1141]= -834157373;
assign addr[1142]= -691191324;
assign addr[1143]= -544719071;
assign addr[1144]= -395483624;
assign addr[1145]= -244242007;
assign addr[1146]= -91761426;
assign addr[1147]= 61184634;
assign addr[1148]= 213820322;
assign addr[1149]= 365371365;
assign addr[1150]= 515068990;
assign addr[1151]= 662153826;
assign addr[1152]= 805879757;
assign addr[1153]= 945517704;
assign addr[1154]= 1080359326;
assign addr[1155]= 1209720613;
assign addr[1156]= 1332945355;
assign addr[1157]= 1449408469;
assign addr[1158]= 1558519173;
assign addr[1159]= 1659723983;
assign addr[1160]= 1752509516;
assign addr[1161]= 1836405100;
assign addr[1162]= 1910985158;
assign addr[1163]= 1975871368;
assign addr[1164]= 2030734582;
assign addr[1165]= 2075296495;
assign addr[1166]= 2109331059;
assign addr[1167]= 2132665626;
assign addr[1168]= 2145181827;
assign addr[1169]= 2146816171;
assign addr[1170]= 2137560369;
assign addr[1171]= 2117461370;
assign addr[1172]= 2086621133;
assign addr[1173]= 2045196100;
assign addr[1174]= 1993396407;
assign addr[1175]= 1931484818;
assign addr[1176]= 1859775393;
assign addr[1177]= 1778631892;
assign addr[1178]= 1688465931;
assign addr[1179]= 1589734894;
assign addr[1180]= 1482939614;
assign addr[1181]= 1368621831;
assign addr[1182]= 1247361445;
assign addr[1183]= 1119773573;
assign addr[1184]= 986505429;
assign addr[1185]= 848233042;
assign addr[1186]= 705657826;
assign addr[1187]= 559503022;
assign addr[1188]= 410510029;
assign addr[1189]= 259434643;
assign addr[1190]= 107043224;
assign addr[1191]= -45891193;
assign addr[1192]= -198592817;
assign addr[1193]= -350287041;
assign addr[1194]= -500204365;
assign addr[1195]= -647584304;
assign addr[1196]= -791679244;
assign addr[1197]= -931758235;
assign addr[1198]= -1067110699;
assign addr[1199]= -1197050035;
assign addr[1200]= -1320917099;
assign addr[1201]= -1438083551;
assign addr[1202]= -1547955041;
assign addr[1203]= -1649974225;
assign addr[1204]= -1743623590;
assign addr[1205]= -1828428082;
assign addr[1206]= -1903957513;
assign addr[1207]= -1969828744;
assign addr[1208]= -2025707632;
assign addr[1209]= -2071310720;
assign addr[1210]= -2106406677;
assign addr[1211]= -2130817471;
assign addr[1212]= -2144419275;
assign addr[1213]= -2147143090;
assign addr[1214]= -2138975100;
assign addr[1215]= -2119956737;
assign addr[1216]= -2090184478;
assign addr[1217]= -2049809346;
assign addr[1218]= -1999036154;
assign addr[1219]= -1938122457;
assign addr[1220]= -1867377253;
assign addr[1221]= -1787159411;
assign addr[1222]= -1697875851;
assign addr[1223]= -1599979481;
assign addr[1224]= -1493966902;
assign addr[1225]= -1380375881;
assign addr[1226]= -1259782632;
assign addr[1227]= -1132798888;
assign addr[1228]= -1000068799;
assign addr[1229]= -862265664;
assign addr[1230]= -720088517;
assign addr[1231]= -574258580;
assign addr[1232]= -425515602;
assign addr[1233]= -274614114;
assign addr[1234]= -122319591;
assign addr[1235]= 30595422;
assign addr[1236]= 183355234;
assign addr[1237]= 335184940;
assign addr[1238]= 485314355;
assign addr[1239]= 632981917;
assign addr[1240]= 777438554;
assign addr[1241]= 917951481;
assign addr[1242]= 1053807919;
assign addr[1243]= 1184318708;
assign addr[1244]= 1308821808;
assign addr[1245]= 1426685652;
assign addr[1246]= 1537312353;
assign addr[1247]= 1640140734;
assign addr[1248]= 1734649179;
assign addr[1249]= 1820358275;
assign addr[1250]= 1896833245;
assign addr[1251]= 1963686155;
assign addr[1252]= 2020577882;
assign addr[1253]= 2067219829;
assign addr[1254]= 2103375398;
assign addr[1255]= 2128861181;
assign addr[1256]= 2143547897;
assign addr[1257]= 2147361045;
assign addr[1258]= 2140281282;
assign addr[1259]= 2122344521;
assign addr[1260]= 2093641749;
assign addr[1261]= 2054318569;
assign addr[1262]= 2004574453;
assign addr[1263]= 1944661739;
assign addr[1264]= 1874884346;
assign addr[1265]= 1795596234;
assign addr[1266]= 1707199606;
assign addr[1267]= 1610142873;
assign addr[1268]= 1504918373;
assign addr[1269]= 1392059879;
assign addr[1270]= 1272139887;
assign addr[1271]= 1145766716;
assign addr[1272]= 1013581418;
assign addr[1273]= 876254528;
assign addr[1274]= 734482665;
assign addr[1275]= 588984994;
assign addr[1276]= 440499581;
assign addr[1277]= 289779648;
assign addr[1278]= 137589750;
assign addr[1279]= -15298099;
assign addr[1280]= -168108346;
assign addr[1281]= -320065829;
assign addr[1282]= -470399716;
assign addr[1283]= -618347408;
assign addr[1284]= -763158411;
assign addr[1285]= -904098143;
assign addr[1286]= -1040451659;
assign addr[1287]= -1171527280;
assign addr[1288]= -1296660098;
assign addr[1289]= -1415215352;
assign addr[1290]= -1526591649;
assign addr[1291]= -1630224009;
assign addr[1292]= -1725586737;
assign addr[1293]= -1812196087;
assign addr[1294]= -1889612716;
assign addr[1295]= -1957443913;
assign addr[1296]= -2015345591;
assign addr[1297]= -2063024031;
assign addr[1298]= -2100237377;
assign addr[1299]= -2126796855;
assign addr[1300]= -2142567738;
assign addr[1301]= -2147470025;
assign addr[1302]= -2141478848;
assign addr[1303]= -2124624598;
assign addr[1304]= -2096992772;
assign addr[1305]= -2058723538;
assign addr[1306]= -2010011024;
assign addr[1307]= -1951102334;
assign addr[1308]= -1882296293;
assign addr[1309]= -1803941934;
assign addr[1310]= -1716436725;
assign addr[1311]= -1620224553;
assign addr[1312]= -1515793473;
assign addr[1313]= -1403673233;
assign addr[1314]= -1284432584;
assign addr[1315]= -1158676398;
assign addr[1316]= -1027042599;
assign addr[1317]= -890198924;
assign addr[1318]= -748839539;
assign addr[1319]= -603681519;
assign addr[1320]= -455461206;
assign addr[1321]= -304930476;
assign addr[1322]= -152852926;
assign addr[1323]= 0;
assign addr[1324]= 152852926;
assign addr[1325]= 304930476;
assign addr[1326]= 455461206;
assign addr[1327]= 603681519;
assign addr[1328]= 748839539;
assign addr[1329]= 890198924;
assign addr[1330]= 1027042599;
assign addr[1331]= 1158676398;
assign addr[1332]= 1284432584;
assign addr[1333]= 1403673233;
assign addr[1334]= 1515793473;
assign addr[1335]= 1620224553;
assign addr[1336]= 1716436725;
assign addr[1337]= 1803941934;
assign addr[1338]= 1882296293;
assign addr[1339]= 1951102334;
assign addr[1340]= 2010011024;
assign addr[1341]= 2058723538;
assign addr[1342]= 2096992772;
assign addr[1343]= 2124624598;
assign addr[1344]= 2141478848;
assign addr[1345]= 2147470025;
assign addr[1346]= 2142567738;
assign addr[1347]= 2126796855;
assign addr[1348]= 2100237377;
assign addr[1349]= 2063024031;
assign addr[1350]= 2015345591;
assign addr[1351]= 1957443913;
assign addr[1352]= 1889612716;
assign addr[1353]= 1812196087;
assign addr[1354]= 1725586737;
assign addr[1355]= 1630224009;
assign addr[1356]= 1526591649;
assign addr[1357]= 1415215352;
assign addr[1358]= 1296660098;
assign addr[1359]= 1171527280;
assign addr[1360]= 1040451659;
assign addr[1361]= 904098143;
assign addr[1362]= 763158411;
assign addr[1363]= 618347408;
assign addr[1364]= 470399716;
assign addr[1365]= 320065829;
assign addr[1366]= 168108346;
assign addr[1367]= 15298099;
assign addr[1368]= -137589750;
assign addr[1369]= -289779648;
assign addr[1370]= -440499581;
assign addr[1371]= -588984994;
assign addr[1372]= -734482665;
assign addr[1373]= -876254528;
assign addr[1374]= -1013581418;
assign addr[1375]= -1145766716;
assign addr[1376]= -1272139887;
assign addr[1377]= -1392059879;
assign addr[1378]= -1504918373;
assign addr[1379]= -1610142873;
assign addr[1380]= -1707199606;
assign addr[1381]= -1795596234;
assign addr[1382]= -1874884346;
assign addr[1383]= -1944661739;
assign addr[1384]= -2004574453;
assign addr[1385]= -2054318569;
assign addr[1386]= -2093641749;
assign addr[1387]= -2122344521;
assign addr[1388]= -2140281282;
assign addr[1389]= -2147361045;
assign addr[1390]= -2143547897;
assign addr[1391]= -2128861181;
assign addr[1392]= -2103375398;
assign addr[1393]= -2067219829;
assign addr[1394]= -2020577882;
assign addr[1395]= -1963686155;
assign addr[1396]= -1896833245;
assign addr[1397]= -1820358275;
assign addr[1398]= -1734649179;
assign addr[1399]= -1640140734;
assign addr[1400]= -1537312353;
assign addr[1401]= -1426685652;
assign addr[1402]= -1308821808;
assign addr[1403]= -1184318708;
assign addr[1404]= -1053807919;
assign addr[1405]= -917951481;
assign addr[1406]= -777438554;
assign addr[1407]= -632981917;
assign addr[1408]= -485314355;
assign addr[1409]= -335184940;
assign addr[1410]= -183355234;
assign addr[1411]= -30595422;
assign addr[1412]= 122319591;
assign addr[1413]= 274614114;
assign addr[1414]= 425515602;
assign addr[1415]= 574258580;
assign addr[1416]= 720088517;
assign addr[1417]= 862265664;
assign addr[1418]= 1000068799;
assign addr[1419]= 1132798888;
assign addr[1420]= 1259782632;
assign addr[1421]= 1380375881;
assign addr[1422]= 1493966902;
assign addr[1423]= 1599979481;
assign addr[1424]= 1697875851;
assign addr[1425]= 1787159411;
assign addr[1426]= 1867377253;
assign addr[1427]= 1938122457;
assign addr[1428]= 1999036154;
assign addr[1429]= 2049809346;
assign addr[1430]= 2090184478;
assign addr[1431]= 2119956737;
assign addr[1432]= 2138975100;
assign addr[1433]= 2147143090;
assign addr[1434]= 2144419275;
assign addr[1435]= 2130817471;
assign addr[1436]= 2106406677;
assign addr[1437]= 2071310720;
assign addr[1438]= 2025707632;
assign addr[1439]= 1969828744;
assign addr[1440]= 1903957513;
assign addr[1441]= 1828428082;
assign addr[1442]= 1743623590;
assign addr[1443]= 1649974225;
assign addr[1444]= 1547955041;
assign addr[1445]= 1438083551;
assign addr[1446]= 1320917099;
assign addr[1447]= 1197050035;
assign addr[1448]= 1067110699;
assign addr[1449]= 931758235;
assign addr[1450]= 791679244;
assign addr[1451]= 647584304;
assign addr[1452]= 500204365;
assign addr[1453]= 350287041;
assign addr[1454]= 198592817;
assign addr[1455]= 45891193;
assign addr[1456]= -107043224;
assign addr[1457]= -259434643;
assign addr[1458]= -410510029;
assign addr[1459]= -559503022;
assign addr[1460]= -705657826;
assign addr[1461]= -848233042;
assign addr[1462]= -986505429;
assign addr[1463]= -1119773573;
assign addr[1464]= -1247361445;
assign addr[1465]= -1368621831;
assign addr[1466]= -1482939614;
assign addr[1467]= -1589734894;
assign addr[1468]= -1688465931;
assign addr[1469]= -1778631892;
assign addr[1470]= -1859775393;
assign addr[1471]= -1931484818;
assign addr[1472]= -1993396407;
assign addr[1473]= -2045196100;
assign addr[1474]= -2086621133;
assign addr[1475]= -2117461370;
assign addr[1476]= -2137560369;
assign addr[1477]= -2146816171;
assign addr[1478]= -2145181827;
assign addr[1479]= -2132665626;
assign addr[1480]= -2109331059;
assign addr[1481]= -2075296495;
assign addr[1482]= -2030734582;
assign addr[1483]= -1975871368;
assign addr[1484]= -1910985158;
assign addr[1485]= -1836405100;
assign addr[1486]= -1752509516;
assign addr[1487]= -1659723983;
assign addr[1488]= -1558519173;
assign addr[1489]= -1449408469;
assign addr[1490]= -1332945355;
assign addr[1491]= -1209720613;
assign addr[1492]= -1080359326;
assign addr[1493]= -945517704;
assign addr[1494]= -805879757;
assign addr[1495]= -662153826;
assign addr[1496]= -515068990;
assign addr[1497]= -365371365;
assign addr[1498]= -213820322;
assign addr[1499]= -61184634;
assign addr[1500]= 91761426;
assign addr[1501]= 244242007;
assign addr[1502]= 395483624;
assign addr[1503]= 544719071;
assign addr[1504]= 691191324;
assign addr[1505]= 834157373;
assign addr[1506]= 972891995;
assign addr[1507]= 1106691431;
assign addr[1508]= 1234876957;
assign addr[1509]= 1356798326;
assign addr[1510]= 1471837070;
assign addr[1511]= 1579409630;
assign addr[1512]= 1678970324;
assign addr[1513]= 1770014111;
assign addr[1514]= 1852079154;
assign addr[1515]= 1924749160;
assign addr[1516]= 1987655498;
assign addr[1517]= 2040479063;
assign addr[1518]= 2082951896;
assign addr[1519]= 2114858546;
assign addr[1520]= 2136037160;
assign addr[1521]= 2146380306;
assign addr[1522]= 2145835515;
assign addr[1523]= 2134405552;
assign addr[1524]= 2112148396;
assign addr[1525]= 2079176953;
assign addr[1526]= 2035658475;
assign addr[1527]= 1981813720;
assign addr[1528]= 1917915825;
assign addr[1529]= 1844288924;
assign addr[1530]= 1761306505;
assign addr[1531]= 1669389513;
assign addr[1532]= 1569004214;
assign addr[1533]= 1460659832;
assign addr[1534]= 1344905966;
assign addr[1535]= 1222329801;
assign addr[1536]= 1093553126;
assign addr[1537]= 959229189;
assign addr[1538]= 820039373;
assign addr[1539]= 676689746;
assign addr[1540]= 529907477;
assign addr[1541]= 380437148;
assign addr[1542]= 229036977;
assign addr[1543]= 76474970;
assign addr[1544]= -76474970;
assign addr[1545]= -229036977;
assign addr[1546]= -380437148;
assign addr[1547]= -529907477;
assign addr[1548]= -676689746;
assign addr[1549]= -820039373;
assign addr[1550]= -959229189;
assign addr[1551]= -1093553126;
assign addr[1552]= -1222329801;
assign addr[1553]= -1344905966;
assign addr[1554]= -1460659832;
assign addr[1555]= -1569004214;
assign addr[1556]= -1669389513;
assign addr[1557]= -1761306505;
assign addr[1558]= -1844288924;
assign addr[1559]= -1917915825;
assign addr[1560]= -1981813720;
assign addr[1561]= -2035658475;
assign addr[1562]= -2079176953;
assign addr[1563]= -2112148396;
assign addr[1564]= -2134405552;
assign addr[1565]= -2145835515;
assign addr[1566]= -2146380306;
assign addr[1567]= -2136037160;
assign addr[1568]= -2114858546;
assign addr[1569]= -2082951896;
assign addr[1570]= -2040479063;
assign addr[1571]= -1987655498;
assign addr[1572]= -1924749160;
assign addr[1573]= -1852079154;
assign addr[1574]= -1770014111;
assign addr[1575]= -1678970324;
assign addr[1576]= -1579409630;
assign addr[1577]= -1471837070;
assign addr[1578]= -1356798326;
assign addr[1579]= -1234876957;
assign addr[1580]= -1106691431;
assign addr[1581]= -972891995;
assign addr[1582]= -834157373;
assign addr[1583]= -691191324;
assign addr[1584]= -544719071;
assign addr[1585]= -395483624;
assign addr[1586]= -244242007;
assign addr[1587]= -91761426;
assign addr[1588]= 61184634;
assign addr[1589]= 213820322;
assign addr[1590]= 365371365;
assign addr[1591]= 515068990;
assign addr[1592]= 662153826;
assign addr[1593]= 805879757;
assign addr[1594]= 945517704;
assign addr[1595]= 1080359326;
assign addr[1596]= 1209720613;
assign addr[1597]= 1332945355;
assign addr[1598]= 1449408469;
assign addr[1599]= 1558519173;
assign addr[1600]= 1659723983;
assign addr[1601]= 1752509516;
assign addr[1602]= 1836405100;
assign addr[1603]= 1910985158;
assign addr[1604]= 1975871368;
assign addr[1605]= 2030734582;
assign addr[1606]= 2075296495;
assign addr[1607]= 2109331059;
assign addr[1608]= 2132665626;
assign addr[1609]= 2145181827;
assign addr[1610]= 2146816171;
assign addr[1611]= 2137560369;
assign addr[1612]= 2117461370;
assign addr[1613]= 2086621133;
assign addr[1614]= 2045196100;
assign addr[1615]= 1993396407;
assign addr[1616]= 1931484818;
assign addr[1617]= 1859775393;
assign addr[1618]= 1778631892;
assign addr[1619]= 1688465931;
assign addr[1620]= 1589734894;
assign addr[1621]= 1482939614;
assign addr[1622]= 1368621831;
assign addr[1623]= 1247361445;
assign addr[1624]= 1119773573;
assign addr[1625]= 986505429;
assign addr[1626]= 848233042;
assign addr[1627]= 705657826;
assign addr[1628]= 559503022;
assign addr[1629]= 410510029;
assign addr[1630]= 259434643;
assign addr[1631]= 107043224;
assign addr[1632]= -45891193;
assign addr[1633]= -198592817;
assign addr[1634]= -350287041;
assign addr[1635]= -500204365;
assign addr[1636]= -647584304;
assign addr[1637]= -791679244;
assign addr[1638]= -931758235;
assign addr[1639]= -1067110699;
assign addr[1640]= -1197050035;
assign addr[1641]= -1320917099;
assign addr[1642]= -1438083551;
assign addr[1643]= -1547955041;
assign addr[1644]= -1649974225;
assign addr[1645]= -1743623590;
assign addr[1646]= -1828428082;
assign addr[1647]= -1903957513;
assign addr[1648]= -1969828744;
assign addr[1649]= -2025707632;
assign addr[1650]= -2071310720;
assign addr[1651]= -2106406677;
assign addr[1652]= -2130817471;
assign addr[1653]= -2144419275;
assign addr[1654]= -2147143090;
assign addr[1655]= -2138975100;
assign addr[1656]= -2119956737;
assign addr[1657]= -2090184478;
assign addr[1658]= -2049809346;
assign addr[1659]= -1999036154;
assign addr[1660]= -1938122457;
assign addr[1661]= -1867377253;
assign addr[1662]= -1787159411;
assign addr[1663]= -1697875851;
assign addr[1664]= -1599979481;
assign addr[1665]= -1493966902;
assign addr[1666]= -1380375881;
assign addr[1667]= -1259782632;
assign addr[1668]= -1132798888;
assign addr[1669]= -1000068799;
assign addr[1670]= -862265664;
assign addr[1671]= -720088517;
assign addr[1672]= -574258580;
assign addr[1673]= -425515602;
assign addr[1674]= -274614114;
assign addr[1675]= -122319591;
assign addr[1676]= 30595422;
assign addr[1677]= 183355234;
assign addr[1678]= 335184940;
assign addr[1679]= 485314355;
assign addr[1680]= 632981917;
assign addr[1681]= 777438554;
assign addr[1682]= 917951481;
assign addr[1683]= 1053807919;
assign addr[1684]= 1184318708;
assign addr[1685]= 1308821808;
assign addr[1686]= 1426685652;
assign addr[1687]= 1537312353;
assign addr[1688]= 1640140734;
assign addr[1689]= 1734649179;
assign addr[1690]= 1820358275;
assign addr[1691]= 1896833245;
assign addr[1692]= 1963686155;
assign addr[1693]= 2020577882;
assign addr[1694]= 2067219829;
assign addr[1695]= 2103375398;
assign addr[1696]= 2128861181;
assign addr[1697]= 2143547897;
assign addr[1698]= 2147361045;
assign addr[1699]= 2140281282;
assign addr[1700]= 2122344521;
assign addr[1701]= 2093641749;
assign addr[1702]= 2054318569;
assign addr[1703]= 2004574453;
assign addr[1704]= 1944661739;
assign addr[1705]= 1874884346;
assign addr[1706]= 1795596234;
assign addr[1707]= 1707199606;
assign addr[1708]= 1610142873;
assign addr[1709]= 1504918373;
assign addr[1710]= 1392059879;
assign addr[1711]= 1272139887;
assign addr[1712]= 1145766716;
assign addr[1713]= 1013581418;
assign addr[1714]= 876254528;
assign addr[1715]= 734482665;
assign addr[1716]= 588984994;
assign addr[1717]= 440499581;
assign addr[1718]= 289779648;
assign addr[1719]= 137589750;
assign addr[1720]= -15298099;
assign addr[1721]= -168108346;
assign addr[1722]= -320065829;
assign addr[1723]= -470399716;
assign addr[1724]= -618347408;
assign addr[1725]= -763158411;
assign addr[1726]= -904098143;
assign addr[1727]= -1040451659;
assign addr[1728]= -1171527280;
assign addr[1729]= -1296660098;
assign addr[1730]= -1415215352;
assign addr[1731]= -1526591649;
assign addr[1732]= -1630224009;
assign addr[1733]= -1725586737;
assign addr[1734]= -1812196087;
assign addr[1735]= -1889612716;
assign addr[1736]= -1957443913;
assign addr[1737]= -2015345591;
assign addr[1738]= -2063024031;
assign addr[1739]= -2100237377;
assign addr[1740]= -2126796855;
assign addr[1741]= -2142567738;
assign addr[1742]= -2147470025;
assign addr[1743]= -2141478848;
assign addr[1744]= -2124624598;
assign addr[1745]= -2096992772;
assign addr[1746]= -2058723538;
assign addr[1747]= -2010011024;
assign addr[1748]= -1951102334;
assign addr[1749]= -1882296293;
assign addr[1750]= -1803941934;
assign addr[1751]= -1716436725;
assign addr[1752]= -1620224553;
assign addr[1753]= -1515793473;
assign addr[1754]= -1403673233;
assign addr[1755]= -1284432584;
assign addr[1756]= -1158676398;
assign addr[1757]= -1027042599;
assign addr[1758]= -890198924;
assign addr[1759]= -748839539;
assign addr[1760]= -603681519;
assign addr[1761]= -455461206;
assign addr[1762]= -304930476;
assign addr[1763]= -152852926;
assign addr[1764]= 0;
assign addr[1765]= 152852926;
assign addr[1766]= 304930476;
assign addr[1767]= 455461206;
assign addr[1768]= 603681519;
assign addr[1769]= 748839539;
assign addr[1770]= 890198924;
assign addr[1771]= 1027042599;
assign addr[1772]= 1158676398;
assign addr[1773]= 1284432584;
assign addr[1774]= 1403673233;
assign addr[1775]= 1515793473;
assign addr[1776]= 1620224553;
assign addr[1777]= 1716436725;
assign addr[1778]= 1803941934;
assign addr[1779]= 1882296293;
assign addr[1780]= 1951102334;
assign addr[1781]= 2010011024;
assign addr[1782]= 2058723538;
assign addr[1783]= 2096992772;
assign addr[1784]= 2124624598;
assign addr[1785]= 2141478848;
assign addr[1786]= 2147470025;
assign addr[1787]= 2142567738;
assign addr[1788]= 2126796855;
assign addr[1789]= 2100237377;
assign addr[1790]= 2063024031;
assign addr[1791]= 2015345591;
assign addr[1792]= 1957443913;
assign addr[1793]= 1889612716;
assign addr[1794]= 1812196087;
assign addr[1795]= 1725586737;
assign addr[1796]= 1630224009;
assign addr[1797]= 1526591649;
assign addr[1798]= 1415215352;
assign addr[1799]= 1296660098;
assign addr[1800]= 1171527280;
assign addr[1801]= 1040451659;
assign addr[1802]= 904098143;
assign addr[1803]= 763158411;
assign addr[1804]= 618347408;
assign addr[1805]= 470399716;
assign addr[1806]= 320065829;
assign addr[1807]= 168108346;
assign addr[1808]= 15298099;
assign addr[1809]= -137589750;
assign addr[1810]= -289779648;
assign addr[1811]= -440499581;
assign addr[1812]= -588984994;
assign addr[1813]= -734482665;
assign addr[1814]= -876254528;
assign addr[1815]= -1013581418;
assign addr[1816]= -1145766716;
assign addr[1817]= -1272139887;
assign addr[1818]= -1392059879;
assign addr[1819]= -1504918373;
assign addr[1820]= -1610142873;
assign addr[1821]= -1707199606;
assign addr[1822]= -1795596234;
assign addr[1823]= -1874884346;
assign addr[1824]= -1944661739;
assign addr[1825]= -2004574453;
assign addr[1826]= -2054318569;
assign addr[1827]= -2093641749;
assign addr[1828]= -2122344521;
assign addr[1829]= -2140281282;
assign addr[1830]= -2147361045;
assign addr[1831]= -2143547897;
assign addr[1832]= -2128861181;
assign addr[1833]= -2103375398;
assign addr[1834]= -2067219829;
assign addr[1835]= -2020577882;
assign addr[1836]= -1963686155;
assign addr[1837]= -1896833245;
assign addr[1838]= -1820358275;
assign addr[1839]= -1734649179;
assign addr[1840]= -1640140734;
assign addr[1841]= -1537312353;
assign addr[1842]= -1426685652;
assign addr[1843]= -1308821808;
assign addr[1844]= -1184318708;
assign addr[1845]= -1053807919;
assign addr[1846]= -917951481;
assign addr[1847]= -777438554;
assign addr[1848]= -632981917;
assign addr[1849]= -485314355;
assign addr[1850]= -335184940;
assign addr[1851]= -183355234;
assign addr[1852]= -30595422;
assign addr[1853]= 122319591;
assign addr[1854]= 274614114;
assign addr[1855]= 425515602;
assign addr[1856]= 574258580;
assign addr[1857]= 720088517;
assign addr[1858]= 862265664;
assign addr[1859]= 1000068799;
assign addr[1860]= 1132798888;
assign addr[1861]= 1259782632;
assign addr[1862]= 1380375881;
assign addr[1863]= 1493966902;
assign addr[1864]= 1599979481;
assign addr[1865]= 1697875851;
assign addr[1866]= 1787159411;
assign addr[1867]= 1867377253;
assign addr[1868]= 1938122457;
assign addr[1869]= 1999036154;
assign addr[1870]= 2049809346;
assign addr[1871]= 2090184478;
assign addr[1872]= 2119956737;
assign addr[1873]= 2138975100;
assign addr[1874]= 2147143090;
assign addr[1875]= 2144419275;
assign addr[1876]= 2130817471;
assign addr[1877]= 2106406677;
assign addr[1878]= 2071310720;
assign addr[1879]= 2025707632;
assign addr[1880]= 1969828744;
assign addr[1881]= 1903957513;
assign addr[1882]= 1828428082;
assign addr[1883]= 1743623590;
assign addr[1884]= 1649974225;
assign addr[1885]= 1547955041;
assign addr[1886]= 1438083551;
assign addr[1887]= 1320917099;
assign addr[1888]= 1197050035;
assign addr[1889]= 1067110699;
assign addr[1890]= 931758235;
assign addr[1891]= 791679244;
assign addr[1892]= 647584304;
assign addr[1893]= 500204365;
assign addr[1894]= 350287041;
assign addr[1895]= 198592817;
assign addr[1896]= 45891193;
assign addr[1897]= -107043224;
assign addr[1898]= -259434643;
assign addr[1899]= -410510029;
assign addr[1900]= -559503022;
assign addr[1901]= -705657826;
assign addr[1902]= -848233042;
assign addr[1903]= -986505429;
assign addr[1904]= -1119773573;
assign addr[1905]= -1247361445;
assign addr[1906]= -1368621831;
assign addr[1907]= -1482939614;
assign addr[1908]= -1589734894;
assign addr[1909]= -1688465931;
assign addr[1910]= -1778631892;
assign addr[1911]= -1859775393;
assign addr[1912]= -1931484818;
assign addr[1913]= -1993396407;
assign addr[1914]= -2045196100;
assign addr[1915]= -2086621133;
assign addr[1916]= -2117461370;
assign addr[1917]= -2137560369;
assign addr[1918]= -2146816171;
assign addr[1919]= -2145181827;
assign addr[1920]= -2132665626;
assign addr[1921]= -2109331059;
assign addr[1922]= -2075296495;
assign addr[1923]= -2030734582;
assign addr[1924]= -1975871368;
assign addr[1925]= -1910985158;
assign addr[1926]= -1836405100;
assign addr[1927]= -1752509516;
assign addr[1928]= -1659723983;
assign addr[1929]= -1558519173;
assign addr[1930]= -1449408469;
assign addr[1931]= -1332945355;
assign addr[1932]= -1209720613;
assign addr[1933]= -1080359326;
assign addr[1934]= -945517704;
assign addr[1935]= -805879757;
assign addr[1936]= -662153826;
assign addr[1937]= -515068990;
assign addr[1938]= -365371365;
assign addr[1939]= -213820322;
assign addr[1940]= -61184634;
assign addr[1941]= 91761426;
assign addr[1942]= 244242007;
assign addr[1943]= 395483624;
assign addr[1944]= 544719071;
assign addr[1945]= 691191324;
assign addr[1946]= 834157373;
assign addr[1947]= 972891995;
assign addr[1948]= 1106691431;
assign addr[1949]= 1234876957;
assign addr[1950]= 1356798326;
assign addr[1951]= 1471837070;
assign addr[1952]= 1579409630;
assign addr[1953]= 1678970324;
assign addr[1954]= 1770014111;
assign addr[1955]= 1852079154;
assign addr[1956]= 1924749160;
assign addr[1957]= 1987655498;
assign addr[1958]= 2040479063;
assign addr[1959]= 2082951896;
assign addr[1960]= 2114858546;
assign addr[1961]= 2136037160;
assign addr[1962]= 2146380306;
assign addr[1963]= 2145835515;
assign addr[1964]= 2134405552;
assign addr[1965]= 2112148396;
assign addr[1966]= 2079176953;
assign addr[1967]= 2035658475;
assign addr[1968]= 1981813720;
assign addr[1969]= 1917915825;
assign addr[1970]= 1844288924;
assign addr[1971]= 1761306505;
assign addr[1972]= 1669389513;
assign addr[1973]= 1569004214;
assign addr[1974]= 1460659832;
assign addr[1975]= 1344905966;
assign addr[1976]= 1222329801;
assign addr[1977]= 1093553126;
assign addr[1978]= 959229189;
assign addr[1979]= 820039373;
assign addr[1980]= 676689746;
assign addr[1981]= 529907477;
assign addr[1982]= 380437148;
assign addr[1983]= 229036977;
assign addr[1984]= 76474970;
assign addr[1985]= -76474970;
assign addr[1986]= -229036977;
assign addr[1987]= -380437148;
assign addr[1988]= -529907477;
assign addr[1989]= -676689746;
assign addr[1990]= -820039373;
assign addr[1991]= -959229189;
assign addr[1992]= -1093553126;
assign addr[1993]= -1222329801;
assign addr[1994]= -1344905966;
assign addr[1995]= -1460659832;
assign addr[1996]= -1569004214;
assign addr[1997]= -1669389513;
assign addr[1998]= -1761306505;
assign addr[1999]= -1844288924;
assign addr[2000]= -1917915825;
assign addr[2001]= -1981813720;
assign addr[2002]= -2035658475;
assign addr[2003]= -2079176953;
assign addr[2004]= -2112148396;
assign addr[2005]= -2134405552;
assign addr[2006]= -2145835515;
assign addr[2007]= -2146380306;
assign addr[2008]= -2136037160;
assign addr[2009]= -2114858546;
assign addr[2010]= -2082951896;
assign addr[2011]= -2040479063;
assign addr[2012]= -1987655498;
assign addr[2013]= -1924749160;
assign addr[2014]= -1852079154;
assign addr[2015]= -1770014111;
assign addr[2016]= -1678970324;
assign addr[2017]= -1579409630;
assign addr[2018]= -1471837070;
assign addr[2019]= -1356798326;
assign addr[2020]= -1234876957;
assign addr[2021]= -1106691431;
assign addr[2022]= -972891995;
assign addr[2023]= -834157373;
assign addr[2024]= -691191324;
assign addr[2025]= -544719071;
assign addr[2026]= -395483624;
assign addr[2027]= -244242007;
assign addr[2028]= -91761426;
assign addr[2029]= 61184634;
assign addr[2030]= 213820322;
assign addr[2031]= 365371365;
assign addr[2032]= 515068990;
assign addr[2033]= 662153826;
assign addr[2034]= 805879757;
assign addr[2035]= 945517704;
assign addr[2036]= 1080359326;
assign addr[2037]= 1209720613;
assign addr[2038]= 1332945355;
assign addr[2039]= 1449408469;
assign addr[2040]= 1558519173;
assign addr[2041]= 1659723983;
assign addr[2042]= 1752509516;
assign addr[2043]= 1836405100;
assign addr[2044]= 1910985158;
assign addr[2045]= 1975871368;
assign addr[2046]= 2030734582;
assign addr[2047]= 2075296495;
assign addr[2048]= 2109331059;
assign addr[2049]= 2132665626;
assign addr[2050]= 2145181827;
assign addr[2051]= 2146816171;
assign addr[2052]= 2137560369;
assign addr[2053]= 2117461370;
assign addr[2054]= 2086621133;
assign addr[2055]= 2045196100;
assign addr[2056]= 1993396407;
assign addr[2057]= 1931484818;
assign addr[2058]= 1859775393;
assign addr[2059]= 1778631892;
assign addr[2060]= 1688465931;
assign addr[2061]= 1589734894;
assign addr[2062]= 1482939614;
assign addr[2063]= 1368621831;
assign addr[2064]= 1247361445;
assign addr[2065]= 1119773573;
assign addr[2066]= 986505429;
assign addr[2067]= 848233042;
assign addr[2068]= 705657826;
assign addr[2069]= 559503022;
assign addr[2070]= 410510029;
assign addr[2071]= 259434643;
assign addr[2072]= 107043224;
assign addr[2073]= -45891193;
assign addr[2074]= -198592817;
assign addr[2075]= -350287041;
assign addr[2076]= -500204365;
assign addr[2077]= -647584304;
assign addr[2078]= -791679244;
assign addr[2079]= -931758235;
assign addr[2080]= -1067110699;
assign addr[2081]= -1197050035;
assign addr[2082]= -1320917099;
assign addr[2083]= -1438083551;
assign addr[2084]= -1547955041;
assign addr[2085]= -1649974225;
assign addr[2086]= -1743623590;
assign addr[2087]= -1828428082;
assign addr[2088]= -1903957513;
assign addr[2089]= -1969828744;
assign addr[2090]= -2025707632;
assign addr[2091]= -2071310720;
assign addr[2092]= -2106406677;
assign addr[2093]= -2130817471;
assign addr[2094]= -2144419275;
assign addr[2095]= -2147143090;
assign addr[2096]= -2138975100;
assign addr[2097]= -2119956737;
assign addr[2098]= -2090184478;
assign addr[2099]= -2049809346;
assign addr[2100]= -1999036154;
assign addr[2101]= -1938122457;
assign addr[2102]= -1867377253;
assign addr[2103]= -1787159411;
assign addr[2104]= -1697875851;
assign addr[2105]= -1599979481;
assign addr[2106]= -1493966902;
assign addr[2107]= -1380375881;
assign addr[2108]= -1259782632;
assign addr[2109]= -1132798888;
assign addr[2110]= -1000068799;
assign addr[2111]= -862265664;
assign addr[2112]= -720088517;
assign addr[2113]= -574258580;
assign addr[2114]= -425515602;
assign addr[2115]= -274614114;
assign addr[2116]= -122319591;
assign addr[2117]= 30595422;
assign addr[2118]= 183355234;
assign addr[2119]= 335184940;
assign addr[2120]= 485314355;
assign addr[2121]= 632981917;
assign addr[2122]= 777438554;
assign addr[2123]= 917951481;
assign addr[2124]= 1053807919;
assign addr[2125]= 1184318708;
assign addr[2126]= 1308821808;
assign addr[2127]= 1426685652;
assign addr[2128]= 1537312353;
assign addr[2129]= 1640140734;
assign addr[2130]= 1734649179;
assign addr[2131]= 1820358275;
assign addr[2132]= 1896833245;
assign addr[2133]= 1963686155;
assign addr[2134]= 2020577882;
assign addr[2135]= 2067219829;
assign addr[2136]= 2103375398;
assign addr[2137]= 2128861181;
assign addr[2138]= 2143547897;
assign addr[2139]= 2147361045;
assign addr[2140]= 2140281282;
assign addr[2141]= 2122344521;
assign addr[2142]= 2093641749;
assign addr[2143]= 2054318569;
assign addr[2144]= 2004574453;
assign addr[2145]= 1944661739;
assign addr[2146]= 1874884346;
assign addr[2147]= 1795596234;
assign addr[2148]= 1707199606;
assign addr[2149]= 1610142873;
assign addr[2150]= 1504918373;
assign addr[2151]= 1392059879;
assign addr[2152]= 1272139887;
assign addr[2153]= 1145766716;
assign addr[2154]= 1013581418;
assign addr[2155]= 876254528;
assign addr[2156]= 734482665;
assign addr[2157]= 588984994;
assign addr[2158]= 440499581;
assign addr[2159]= 289779648;
assign addr[2160]= 137589750;
assign addr[2161]= -15298099;
assign addr[2162]= -168108346;
assign addr[2163]= -320065829;
assign addr[2164]= -470399716;
assign addr[2165]= -618347408;
assign addr[2166]= -763158411;
assign addr[2167]= -904098143;
assign addr[2168]= -1040451659;
assign addr[2169]= -1171527280;
assign addr[2170]= -1296660098;
assign addr[2171]= -1415215352;
assign addr[2172]= -1526591649;
assign addr[2173]= -1630224009;
assign addr[2174]= -1725586737;
assign addr[2175]= -1812196087;
assign addr[2176]= -1889612716;
assign addr[2177]= -1957443913;
assign addr[2178]= -2015345591;
assign addr[2179]= -2063024031;
assign addr[2180]= -2100237377;
assign addr[2181]= -2126796855;
assign addr[2182]= -2142567738;
assign addr[2183]= -2147470025;
assign addr[2184]= -2141478848;
assign addr[2185]= -2124624598;
assign addr[2186]= -2096992772;
assign addr[2187]= -2058723538;
assign addr[2188]= -2010011024;
assign addr[2189]= -1951102334;
assign addr[2190]= -1882296293;
assign addr[2191]= -1803941934;
assign addr[2192]= -1716436725;
assign addr[2193]= -1620224553;
assign addr[2194]= -1515793473;
assign addr[2195]= -1403673233;
assign addr[2196]= -1284432584;
assign addr[2197]= -1158676398;
assign addr[2198]= -1027042599;
assign addr[2199]= -890198924;
assign addr[2200]= -748839539;
assign addr[2201]= -603681519;
assign addr[2202]= -455461206;
assign addr[2203]= -304930476;
assign addr[2204]= -152852926;
assign addr[2205]= 0;
assign addr[2206]= 152852926;
assign addr[2207]= 304930476;
assign addr[2208]= 455461206;
assign addr[2209]= 603681519;
assign addr[2210]= 748839539;
assign addr[2211]= 890198924;
assign addr[2212]= 1027042599;
assign addr[2213]= 1158676398;
assign addr[2214]= 1284432584;
assign addr[2215]= 1403673233;
assign addr[2216]= 1515793473;
assign addr[2217]= 1620224553;
assign addr[2218]= 1716436725;
assign addr[2219]= 1803941934;
assign addr[2220]= 1882296293;
assign addr[2221]= 1951102334;
assign addr[2222]= 2010011024;
assign addr[2223]= 2058723538;
assign addr[2224]= 2096992772;
assign addr[2225]= 2124624598;
assign addr[2226]= 2141478848;
assign addr[2227]= 2147470025;
assign addr[2228]= 2142567738;
assign addr[2229]= 2126796855;
assign addr[2230]= 2100237377;
assign addr[2231]= 2063024031;
assign addr[2232]= 2015345591;
assign addr[2233]= 1957443913;
assign addr[2234]= 1889612716;
assign addr[2235]= 1812196087;
assign addr[2236]= 1725586737;
assign addr[2237]= 1630224009;
assign addr[2238]= 1526591649;
assign addr[2239]= 1415215352;
assign addr[2240]= 1296660098;
assign addr[2241]= 1171527280;
assign addr[2242]= 1040451659;
assign addr[2243]= 904098143;
assign addr[2244]= 763158411;
assign addr[2245]= 618347408;
assign addr[2246]= 470399716;
assign addr[2247]= 320065829;
assign addr[2248]= 168108346;
assign addr[2249]= 15298099;
assign addr[2250]= -137589750;
assign addr[2251]= -289779648;
assign addr[2252]= -440499581;
assign addr[2253]= -588984994;
assign addr[2254]= -734482665;
assign addr[2255]= -876254528;
assign addr[2256]= -1013581418;
assign addr[2257]= -1145766716;
assign addr[2258]= -1272139887;
assign addr[2259]= -1392059879;
assign addr[2260]= -1504918373;
assign addr[2261]= -1610142873;
assign addr[2262]= -1707199606;
assign addr[2263]= -1795596234;
assign addr[2264]= -1874884346;
assign addr[2265]= -1944661739;
assign addr[2266]= -2004574453;
assign addr[2267]= -2054318569;
assign addr[2268]= -2093641749;
assign addr[2269]= -2122344521;
assign addr[2270]= -2140281282;
assign addr[2271]= -2147361045;
assign addr[2272]= -2143547897;
assign addr[2273]= -2128861181;
assign addr[2274]= -2103375398;
assign addr[2275]= -2067219829;
assign addr[2276]= -2020577882;
assign addr[2277]= -1963686155;
assign addr[2278]= -1896833245;
assign addr[2279]= -1820358275;
assign addr[2280]= -1734649179;
assign addr[2281]= -1640140734;
assign addr[2282]= -1537312353;
assign addr[2283]= -1426685652;
assign addr[2284]= -1308821808;
assign addr[2285]= -1184318708;
assign addr[2286]= -1053807919;
assign addr[2287]= -917951481;
assign addr[2288]= -777438554;
assign addr[2289]= -632981917;
assign addr[2290]= -485314355;
assign addr[2291]= -335184940;
assign addr[2292]= -183355234;
assign addr[2293]= -30595422;
assign addr[2294]= 122319591;
assign addr[2295]= 274614114;
assign addr[2296]= 425515602;
assign addr[2297]= 574258580;
assign addr[2298]= 720088517;
assign addr[2299]= 862265664;
assign addr[2300]= 1000068799;
assign addr[2301]= 1132798888;
assign addr[2302]= 1259782632;
assign addr[2303]= 1380375881;
assign addr[2304]= 1493966902;
assign addr[2305]= 1599979481;
assign addr[2306]= 1697875851;
assign addr[2307]= 1787159411;
assign addr[2308]= 1867377253;
assign addr[2309]= 1938122457;
assign addr[2310]= 1999036154;
assign addr[2311]= 2049809346;
assign addr[2312]= 2090184478;
assign addr[2313]= 2119956737;
assign addr[2314]= 2138975100;
assign addr[2315]= 2147143090;
assign addr[2316]= 2144419275;
assign addr[2317]= 2130817471;
assign addr[2318]= 2106406677;
assign addr[2319]= 2071310720;
assign addr[2320]= 2025707632;
assign addr[2321]= 1969828744;
assign addr[2322]= 1903957513;
assign addr[2323]= 1828428082;
assign addr[2324]= 1743623590;
assign addr[2325]= 1649974225;
assign addr[2326]= 1547955041;
assign addr[2327]= 1438083551;
assign addr[2328]= 1320917099;
assign addr[2329]= 1197050035;
assign addr[2330]= 1067110699;
assign addr[2331]= 931758235;
assign addr[2332]= 791679244;
assign addr[2333]= 647584304;
assign addr[2334]= 500204365;
assign addr[2335]= 350287041;
assign addr[2336]= 198592817;
assign addr[2337]= 45891193;
assign addr[2338]= -107043224;
assign addr[2339]= -259434643;
assign addr[2340]= -410510029;
assign addr[2341]= -559503022;
assign addr[2342]= -705657826;
assign addr[2343]= -848233042;
assign addr[2344]= -986505429;
assign addr[2345]= -1119773573;
assign addr[2346]= -1247361445;
assign addr[2347]= -1368621831;
assign addr[2348]= -1482939614;
assign addr[2349]= -1589734894;
assign addr[2350]= -1688465931;
assign addr[2351]= -1778631892;
assign addr[2352]= -1859775393;
assign addr[2353]= -1931484818;
assign addr[2354]= -1993396407;
assign addr[2355]= -2045196100;
assign addr[2356]= -2086621133;
assign addr[2357]= -2117461370;
assign addr[2358]= -2137560369;
assign addr[2359]= -2146816171;
assign addr[2360]= -2145181827;
assign addr[2361]= -2132665626;
assign addr[2362]= -2109331059;
assign addr[2363]= -2075296495;
assign addr[2364]= -2030734582;
assign addr[2365]= -1975871368;
assign addr[2366]= -1910985158;
assign addr[2367]= -1836405100;
assign addr[2368]= -1752509516;
assign addr[2369]= -1659723983;
assign addr[2370]= -1558519173;
assign addr[2371]= -1449408469;
assign addr[2372]= -1332945355;
assign addr[2373]= -1209720613;
assign addr[2374]= -1080359326;
assign addr[2375]= -945517704;
assign addr[2376]= -805879757;
assign addr[2377]= -662153826;
assign addr[2378]= -515068990;
assign addr[2379]= -365371365;
assign addr[2380]= -213820322;
assign addr[2381]= -61184634;
assign addr[2382]= 91761426;
assign addr[2383]= 244242007;
assign addr[2384]= 395483624;
assign addr[2385]= 544719071;
assign addr[2386]= 691191324;
assign addr[2387]= 834157373;
assign addr[2388]= 972891995;
assign addr[2389]= 1106691431;
assign addr[2390]= 1234876957;
assign addr[2391]= 1356798326;
assign addr[2392]= 1471837070;
assign addr[2393]= 1579409630;
assign addr[2394]= 1678970324;
assign addr[2395]= 1770014111;
assign addr[2396]= 1852079154;
assign addr[2397]= 1924749160;
assign addr[2398]= 1987655498;
assign addr[2399]= 2040479063;
assign addr[2400]= 2082951896;
assign addr[2401]= 2114858546;
assign addr[2402]= 2136037160;
assign addr[2403]= 2146380306;
assign addr[2404]= 2145835515;
assign addr[2405]= 2134405552;
assign addr[2406]= 2112148396;
assign addr[2407]= 2079176953;
assign addr[2408]= 2035658475;
assign addr[2409]= 1981813720;
assign addr[2410]= 1917915825;
assign addr[2411]= 1844288924;
assign addr[2412]= 1761306505;
assign addr[2413]= 1669389513;
assign addr[2414]= 1569004214;
assign addr[2415]= 1460659832;
assign addr[2416]= 1344905966;
assign addr[2417]= 1222329801;
assign addr[2418]= 1093553126;
assign addr[2419]= 959229189;
assign addr[2420]= 820039373;
assign addr[2421]= 676689746;
assign addr[2422]= 529907477;
assign addr[2423]= 380437148;
assign addr[2424]= 229036977;
assign addr[2425]= 76474970;
assign addr[2426]= -76474970;
assign addr[2427]= -229036977;
assign addr[2428]= -380437148;
assign addr[2429]= -529907477;
assign addr[2430]= -676689746;
assign addr[2431]= -820039373;
assign addr[2432]= -959229189;
assign addr[2433]= -1093553126;
assign addr[2434]= -1222329801;
assign addr[2435]= -1344905966;
assign addr[2436]= -1460659832;
assign addr[2437]= -1569004214;
assign addr[2438]= -1669389513;
assign addr[2439]= -1761306505;
assign addr[2440]= -1844288924;
assign addr[2441]= -1917915825;
assign addr[2442]= -1981813720;
assign addr[2443]= -2035658475;
assign addr[2444]= -2079176953;
assign addr[2445]= -2112148396;
assign addr[2446]= -2134405552;
assign addr[2447]= -2145835515;
assign addr[2448]= -2146380306;
assign addr[2449]= -2136037160;
assign addr[2450]= -2114858546;
assign addr[2451]= -2082951896;
assign addr[2452]= -2040479063;
assign addr[2453]= -1987655498;
assign addr[2454]= -1924749160;
assign addr[2455]= -1852079154;
assign addr[2456]= -1770014111;
assign addr[2457]= -1678970324;
assign addr[2458]= -1579409630;
assign addr[2459]= -1471837070;
assign addr[2460]= -1356798326;
assign addr[2461]= -1234876957;
assign addr[2462]= -1106691431;
assign addr[2463]= -972891995;
assign addr[2464]= -834157373;
assign addr[2465]= -691191324;
assign addr[2466]= -544719071;
assign addr[2467]= -395483624;
assign addr[2468]= -244242007;
assign addr[2469]= -91761426;
assign addr[2470]= 61184634;
assign addr[2471]= 213820322;
assign addr[2472]= 365371365;
assign addr[2473]= 515068990;
assign addr[2474]= 662153826;
assign addr[2475]= 805879757;
assign addr[2476]= 945517704;
assign addr[2477]= 1080359326;
assign addr[2478]= 1209720613;
assign addr[2479]= 1332945355;
assign addr[2480]= 1449408469;
assign addr[2481]= 1558519173;
assign addr[2482]= 1659723983;
assign addr[2483]= 1752509516;
assign addr[2484]= 1836405100;
assign addr[2485]= 1910985158;
assign addr[2486]= 1975871368;
assign addr[2487]= 2030734582;
assign addr[2488]= 2075296495;
assign addr[2489]= 2109331059;
assign addr[2490]= 2132665626;
assign addr[2491]= 2145181827;
assign addr[2492]= 2146816171;
assign addr[2493]= 2137560369;
assign addr[2494]= 2117461370;
assign addr[2495]= 2086621133;
assign addr[2496]= 2045196100;
assign addr[2497]= 1993396407;
assign addr[2498]= 1931484818;
assign addr[2499]= 1859775393;
assign addr[2500]= 1778631892;
assign addr[2501]= 1688465931;
assign addr[2502]= 1589734894;
assign addr[2503]= 1482939614;
assign addr[2504]= 1368621831;
assign addr[2505]= 1247361445;
assign addr[2506]= 1119773573;
assign addr[2507]= 986505429;
assign addr[2508]= 848233042;
assign addr[2509]= 705657826;
assign addr[2510]= 559503022;
assign addr[2511]= 410510029;
assign addr[2512]= 259434643;
assign addr[2513]= 107043224;
assign addr[2514]= -45891193;
assign addr[2515]= -198592817;
assign addr[2516]= -350287041;
assign addr[2517]= -500204365;
assign addr[2518]= -647584304;
assign addr[2519]= -791679244;
assign addr[2520]= -931758235;
assign addr[2521]= -1067110699;
assign addr[2522]= -1197050035;
assign addr[2523]= -1320917099;
assign addr[2524]= -1438083551;
assign addr[2525]= -1547955041;
assign addr[2526]= -1649974225;
assign addr[2527]= -1743623590;
assign addr[2528]= -1828428082;
assign addr[2529]= -1903957513;
assign addr[2530]= -1969828744;
assign addr[2531]= -2025707632;
assign addr[2532]= -2071310720;
assign addr[2533]= -2106406677;
assign addr[2534]= -2130817471;
assign addr[2535]= -2144419275;
assign addr[2536]= -2147143090;
assign addr[2537]= -2138975100;
assign addr[2538]= -2119956737;
assign addr[2539]= -2090184478;
assign addr[2540]= -2049809346;
assign addr[2541]= -1999036154;
assign addr[2542]= -1938122457;
assign addr[2543]= -1867377253;
assign addr[2544]= -1787159411;
assign addr[2545]= -1697875851;
assign addr[2546]= -1599979481;
assign addr[2547]= -1493966902;
assign addr[2548]= -1380375881;
assign addr[2549]= -1259782632;
assign addr[2550]= -1132798888;
assign addr[2551]= -1000068799;
assign addr[2552]= -862265664;
assign addr[2553]= -720088517;
assign addr[2554]= -574258580;
assign addr[2555]= -425515602;
assign addr[2556]= -274614114;
assign addr[2557]= -122319591;
assign addr[2558]= 30595422;
assign addr[2559]= 183355234;
assign addr[2560]= 335184940;
assign addr[2561]= 485314355;
assign addr[2562]= 632981917;
assign addr[2563]= 777438554;
assign addr[2564]= 917951481;
assign addr[2565]= 1053807919;
assign addr[2566]= 1184318708;
assign addr[2567]= 1308821808;
assign addr[2568]= 1426685652;
assign addr[2569]= 1537312353;
assign addr[2570]= 1640140734;
assign addr[2571]= 1734649179;
assign addr[2572]= 1820358275;
assign addr[2573]= 1896833245;
assign addr[2574]= 1963686155;
assign addr[2575]= 2020577882;
assign addr[2576]= 2067219829;
assign addr[2577]= 2103375398;
assign addr[2578]= 2128861181;
assign addr[2579]= 2143547897;
assign addr[2580]= 2147361045;
assign addr[2581]= 2140281282;
assign addr[2582]= 2122344521;
assign addr[2583]= 2093641749;
assign addr[2584]= 2054318569;
assign addr[2585]= 2004574453;
assign addr[2586]= 1944661739;
assign addr[2587]= 1874884346;
assign addr[2588]= 1795596234;
assign addr[2589]= 1707199606;
assign addr[2590]= 1610142873;
assign addr[2591]= 1504918373;
assign addr[2592]= 1392059879;
assign addr[2593]= 1272139887;
assign addr[2594]= 1145766716;
assign addr[2595]= 1013581418;
assign addr[2596]= 876254528;
assign addr[2597]= 734482665;
assign addr[2598]= 588984994;
assign addr[2599]= 440499581;
assign addr[2600]= 289779648;
assign addr[2601]= 137589750;
assign addr[2602]= -15298099;
assign addr[2603]= -168108346;
assign addr[2604]= -320065829;
assign addr[2605]= -470399716;
assign addr[2606]= -618347408;
assign addr[2607]= -763158411;
assign addr[2608]= -904098143;
assign addr[2609]= -1040451659;
assign addr[2610]= -1171527280;
assign addr[2611]= -1296660098;
assign addr[2612]= -1415215352;
assign addr[2613]= -1526591649;
assign addr[2614]= -1630224009;
assign addr[2615]= -1725586737;
assign addr[2616]= -1812196087;
assign addr[2617]= -1889612716;
assign addr[2618]= -1957443913;
assign addr[2619]= -2015345591;
assign addr[2620]= -2063024031;
assign addr[2621]= -2100237377;
assign addr[2622]= -2126796855;
assign addr[2623]= -2142567738;
assign addr[2624]= -2147470025;
assign addr[2625]= -2141478848;
assign addr[2626]= -2124624598;
assign addr[2627]= -2096992772;
assign addr[2628]= -2058723538;
assign addr[2629]= -2010011024;
assign addr[2630]= -1951102334;
assign addr[2631]= -1882296293;
assign addr[2632]= -1803941934;
assign addr[2633]= -1716436725;
assign addr[2634]= -1620224553;
assign addr[2635]= -1515793473;
assign addr[2636]= -1403673233;
assign addr[2637]= -1284432584;
assign addr[2638]= -1158676398;
assign addr[2639]= -1027042599;
assign addr[2640]= -890198924;
assign addr[2641]= -748839539;
assign addr[2642]= -603681519;
assign addr[2643]= -455461206;
assign addr[2644]= -304930476;
assign addr[2645]= -152852926;
assign addr[2646]= 0;
assign addr[2647]= 152852926;
assign addr[2648]= 304930476;
assign addr[2649]= 455461206;
assign addr[2650]= 603681519;
assign addr[2651]= 748839539;
assign addr[2652]= 890198924;
assign addr[2653]= 1027042599;
assign addr[2654]= 1158676398;
assign addr[2655]= 1284432584;
assign addr[2656]= 1403673233;
assign addr[2657]= 1515793473;
assign addr[2658]= 1620224553;
assign addr[2659]= 1716436725;
assign addr[2660]= 1803941934;
assign addr[2661]= 1882296293;
assign addr[2662]= 1951102334;
assign addr[2663]= 2010011024;
assign addr[2664]= 2058723538;
assign addr[2665]= 2096992772;
assign addr[2666]= 2124624598;
assign addr[2667]= 2141478848;
assign addr[2668]= 2147470025;
assign addr[2669]= 2142567738;
assign addr[2670]= 2126796855;
assign addr[2671]= 2100237377;
assign addr[2672]= 2063024031;
assign addr[2673]= 2015345591;
assign addr[2674]= 1957443913;
assign addr[2675]= 1889612716;
assign addr[2676]= 1812196087;
assign addr[2677]= 1725586737;
assign addr[2678]= 1630224009;
assign addr[2679]= 1526591649;
assign addr[2680]= 1415215352;
assign addr[2681]= 1296660098;
assign addr[2682]= 1171527280;
assign addr[2683]= 1040451659;
assign addr[2684]= 904098143;
assign addr[2685]= 763158411;
assign addr[2686]= 618347408;
assign addr[2687]= 470399716;
assign addr[2688]= 320065829;
assign addr[2689]= 168108346;
assign addr[2690]= 15298099;
assign addr[2691]= -137589750;
assign addr[2692]= -289779648;
assign addr[2693]= -440499581;
assign addr[2694]= -588984994;
assign addr[2695]= -734482665;
assign addr[2696]= -876254528;
assign addr[2697]= -1013581418;
assign addr[2698]= -1145766716;
assign addr[2699]= -1272139887;
assign addr[2700]= -1392059879;
assign addr[2701]= -1504918373;
assign addr[2702]= -1610142873;
assign addr[2703]= -1707199606;
assign addr[2704]= -1795596234;
assign addr[2705]= -1874884346;
assign addr[2706]= -1944661739;
assign addr[2707]= -2004574453;
assign addr[2708]= -2054318569;
assign addr[2709]= -2093641749;
assign addr[2710]= -2122344521;
assign addr[2711]= -2140281282;
assign addr[2712]= -2147361045;
assign addr[2713]= -2143547897;
assign addr[2714]= -2128861181;
assign addr[2715]= -2103375398;
assign addr[2716]= -2067219829;
assign addr[2717]= -2020577882;
assign addr[2718]= -1963686155;
assign addr[2719]= -1896833245;
assign addr[2720]= -1820358275;
assign addr[2721]= -1734649179;
assign addr[2722]= -1640140734;
assign addr[2723]= -1537312353;
assign addr[2724]= -1426685652;
assign addr[2725]= -1308821808;
assign addr[2726]= -1184318708;
assign addr[2727]= -1053807919;
assign addr[2728]= -917951481;
assign addr[2729]= -777438554;
assign addr[2730]= -632981917;
assign addr[2731]= -485314355;
assign addr[2732]= -335184940;
assign addr[2733]= -183355234;
assign addr[2734]= -30595422;
assign addr[2735]= 122319591;
assign addr[2736]= 274614114;
assign addr[2737]= 425515602;
assign addr[2738]= 574258580;
assign addr[2739]= 720088517;
assign addr[2740]= 862265664;
assign addr[2741]= 1000068799;
assign addr[2742]= 1132798888;
assign addr[2743]= 1259782632;
assign addr[2744]= 1380375881;
assign addr[2745]= 1493966902;
assign addr[2746]= 1599979481;
assign addr[2747]= 1697875851;
assign addr[2748]= 1787159411;
assign addr[2749]= 1867377253;
assign addr[2750]= 1938122457;
assign addr[2751]= 1999036154;
assign addr[2752]= 2049809346;
assign addr[2753]= 2090184478;
assign addr[2754]= 2119956737;
assign addr[2755]= 2138975100;
assign addr[2756]= 2147143090;
assign addr[2757]= 2144419275;
assign addr[2758]= 2130817471;
assign addr[2759]= 2106406677;
assign addr[2760]= 2071310720;
assign addr[2761]= 2025707632;
assign addr[2762]= 1969828744;
assign addr[2763]= 1903957513;
assign addr[2764]= 1828428082;
assign addr[2765]= 1743623590;
assign addr[2766]= 1649974225;
assign addr[2767]= 1547955041;
assign addr[2768]= 1438083551;
assign addr[2769]= 1320917099;
assign addr[2770]= 1197050035;
assign addr[2771]= 1067110699;
assign addr[2772]= 931758235;
assign addr[2773]= 791679244;
assign addr[2774]= 647584304;
assign addr[2775]= 500204365;
assign addr[2776]= 350287041;
assign addr[2777]= 198592817;
assign addr[2778]= 45891193;
assign addr[2779]= -107043224;
assign addr[2780]= -259434643;
assign addr[2781]= -410510029;
assign addr[2782]= -559503022;
assign addr[2783]= -705657826;
assign addr[2784]= -848233042;
assign addr[2785]= -986505429;
assign addr[2786]= -1119773573;
assign addr[2787]= -1247361445;
assign addr[2788]= -1368621831;
assign addr[2789]= -1482939614;
assign addr[2790]= -1589734894;
assign addr[2791]= -1688465931;
assign addr[2792]= -1778631892;
assign addr[2793]= -1859775393;
assign addr[2794]= -1931484818;
assign addr[2795]= -1993396407;
assign addr[2796]= -2045196100;
assign addr[2797]= -2086621133;
assign addr[2798]= -2117461370;
assign addr[2799]= -2137560369;
assign addr[2800]= -2146816171;
assign addr[2801]= -2145181827;
assign addr[2802]= -2132665626;
assign addr[2803]= -2109331059;
assign addr[2804]= -2075296495;
assign addr[2805]= -2030734582;
assign addr[2806]= -1975871368;
assign addr[2807]= -1910985158;
assign addr[2808]= -1836405100;
assign addr[2809]= -1752509516;
assign addr[2810]= -1659723983;
assign addr[2811]= -1558519173;
assign addr[2812]= -1449408469;
assign addr[2813]= -1332945355;
assign addr[2814]= -1209720613;
assign addr[2815]= -1080359326;
assign addr[2816]= -945517704;
assign addr[2817]= -805879757;
assign addr[2818]= -662153826;
assign addr[2819]= -515068990;
assign addr[2820]= -365371365;
assign addr[2821]= -213820322;
assign addr[2822]= -61184634;
assign addr[2823]= 91761426;
assign addr[2824]= 244242007;
assign addr[2825]= 395483624;
assign addr[2826]= 544719071;
assign addr[2827]= 691191324;
assign addr[2828]= 834157373;
assign addr[2829]= 972891995;
assign addr[2830]= 1106691431;
assign addr[2831]= 1234876957;
assign addr[2832]= 1356798326;
assign addr[2833]= 1471837070;
assign addr[2834]= 1579409630;
assign addr[2835]= 1678970324;
assign addr[2836]= 1770014111;
assign addr[2837]= 1852079154;
assign addr[2838]= 1924749160;
assign addr[2839]= 1987655498;
assign addr[2840]= 2040479063;
assign addr[2841]= 2082951896;
assign addr[2842]= 2114858546;
assign addr[2843]= 2136037160;
assign addr[2844]= 2146380306;
assign addr[2845]= 2145835515;
assign addr[2846]= 2134405552;
assign addr[2847]= 2112148396;
assign addr[2848]= 2079176953;
assign addr[2849]= 2035658475;
assign addr[2850]= 1981813720;
assign addr[2851]= 1917915825;
assign addr[2852]= 1844288924;
assign addr[2853]= 1761306505;
assign addr[2854]= 1669389513;
assign addr[2855]= 1569004214;
assign addr[2856]= 1460659832;
assign addr[2857]= 1344905966;
assign addr[2858]= 1222329801;
assign addr[2859]= 1093553126;
assign addr[2860]= 959229189;
assign addr[2861]= 820039373;
assign addr[2862]= 676689746;
assign addr[2863]= 529907477;
assign addr[2864]= 380437148;
assign addr[2865]= 229036977;
assign addr[2866]= 76474970;
assign addr[2867]= -76474970;
assign addr[2868]= -229036977;
assign addr[2869]= -380437148;
assign addr[2870]= -529907477;
assign addr[2871]= -676689746;
assign addr[2872]= -820039373;
assign addr[2873]= -959229189;
assign addr[2874]= -1093553126;
assign addr[2875]= -1222329801;
assign addr[2876]= -1344905966;
assign addr[2877]= -1460659832;
assign addr[2878]= -1569004214;
assign addr[2879]= -1669389513;
assign addr[2880]= -1761306505;
assign addr[2881]= -1844288924;
assign addr[2882]= -1917915825;
assign addr[2883]= -1981813720;
assign addr[2884]= -2035658475;
assign addr[2885]= -2079176953;
assign addr[2886]= -2112148396;
assign addr[2887]= -2134405552;
assign addr[2888]= -2145835515;
assign addr[2889]= -2146380306;
assign addr[2890]= -2136037160;
assign addr[2891]= -2114858546;
assign addr[2892]= -2082951896;
assign addr[2893]= -2040479063;
assign addr[2894]= -1987655498;
assign addr[2895]= -1924749160;
assign addr[2896]= -1852079154;
assign addr[2897]= -1770014111;
assign addr[2898]= -1678970324;
assign addr[2899]= -1579409630;
assign addr[2900]= -1471837070;
assign addr[2901]= -1356798326;
assign addr[2902]= -1234876957;
assign addr[2903]= -1106691431;
assign addr[2904]= -972891995;
assign addr[2905]= -834157373;
assign addr[2906]= -691191324;
assign addr[2907]= -544719071;
assign addr[2908]= -395483624;
assign addr[2909]= -244242007;
assign addr[2910]= -91761426;
assign addr[2911]= 61184634;
assign addr[2912]= 213820322;
assign addr[2913]= 365371365;
assign addr[2914]= 515068990;
assign addr[2915]= 662153826;
assign addr[2916]= 805879757;
assign addr[2917]= 945517704;
assign addr[2918]= 1080359326;
assign addr[2919]= 1209720613;
assign addr[2920]= 1332945355;
assign addr[2921]= 1449408469;
assign addr[2922]= 1558519173;
assign addr[2923]= 1659723983;
assign addr[2924]= 1752509516;
assign addr[2925]= 1836405100;
assign addr[2926]= 1910985158;
assign addr[2927]= 1975871368;
assign addr[2928]= 2030734582;
assign addr[2929]= 2075296495;
assign addr[2930]= 2109331059;
assign addr[2931]= 2132665626;
assign addr[2932]= 2145181827;
assign addr[2933]= 2146816171;
assign addr[2934]= 2137560369;
assign addr[2935]= 2117461370;
assign addr[2936]= 2086621133;
assign addr[2937]= 2045196100;
assign addr[2938]= 1993396407;
assign addr[2939]= 1931484818;
assign addr[2940]= 1859775393;
assign addr[2941]= 1778631892;
assign addr[2942]= 1688465931;
assign addr[2943]= 1589734894;
assign addr[2944]= 1482939614;
assign addr[2945]= 1368621831;
assign addr[2946]= 1247361445;
assign addr[2947]= 1119773573;
assign addr[2948]= 986505429;
assign addr[2949]= 848233042;
assign addr[2950]= 705657826;
assign addr[2951]= 559503022;
assign addr[2952]= 410510029;
assign addr[2953]= 259434643;
assign addr[2954]= 107043224;
assign addr[2955]= -45891193;
assign addr[2956]= -198592817;
assign addr[2957]= -350287041;
assign addr[2958]= -500204365;
assign addr[2959]= -647584304;
assign addr[2960]= -791679244;
assign addr[2961]= -931758235;
assign addr[2962]= -1067110699;
assign addr[2963]= -1197050035;
assign addr[2964]= -1320917099;
assign addr[2965]= -1438083551;
assign addr[2966]= -1547955041;
assign addr[2967]= -1649974225;
assign addr[2968]= -1743623590;
assign addr[2969]= -1828428082;
assign addr[2970]= -1903957513;
assign addr[2971]= -1969828744;
assign addr[2972]= -2025707632;
assign addr[2973]= -2071310720;
assign addr[2974]= -2106406677;
assign addr[2975]= -2130817471;
assign addr[2976]= -2144419275;
assign addr[2977]= -2147143090;
assign addr[2978]= -2138975100;
assign addr[2979]= -2119956737;
assign addr[2980]= -2090184478;
assign addr[2981]= -2049809346;
assign addr[2982]= -1999036154;
assign addr[2983]= -1938122457;
assign addr[2984]= -1867377253;
assign addr[2985]= -1787159411;
assign addr[2986]= -1697875851;
assign addr[2987]= -1599979481;
assign addr[2988]= -1493966902;
assign addr[2989]= -1380375881;
assign addr[2990]= -1259782632;
assign addr[2991]= -1132798888;
assign addr[2992]= -1000068799;
assign addr[2993]= -862265664;
assign addr[2994]= -720088517;
assign addr[2995]= -574258580;
assign addr[2996]= -425515602;
assign addr[2997]= -274614114;
assign addr[2998]= -122319591;
assign addr[2999]= 30595422;
assign addr[3000]= 183355234;
assign addr[3001]= 335184940;
assign addr[3002]= 485314355;
assign addr[3003]= 632981917;
assign addr[3004]= 777438554;
assign addr[3005]= 917951481;
assign addr[3006]= 1053807919;
assign addr[3007]= 1184318708;
assign addr[3008]= 1308821808;
assign addr[3009]= 1426685652;
assign addr[3010]= 1537312353;
assign addr[3011]= 1640140734;
assign addr[3012]= 1734649179;
assign addr[3013]= 1820358275;
assign addr[3014]= 1896833245;
assign addr[3015]= 1963686155;
assign addr[3016]= 2020577882;
assign addr[3017]= 2067219829;
assign addr[3018]= 2103375398;
assign addr[3019]= 2128861181;
assign addr[3020]= 2143547897;
assign addr[3021]= 2147361045;
assign addr[3022]= 2140281282;
assign addr[3023]= 2122344521;
assign addr[3024]= 2093641749;
assign addr[3025]= 2054318569;
assign addr[3026]= 2004574453;
assign addr[3027]= 1944661739;
assign addr[3028]= 1874884346;
assign addr[3029]= 1795596234;
assign addr[3030]= 1707199606;
assign addr[3031]= 1610142873;
assign addr[3032]= 1504918373;
assign addr[3033]= 1392059879;
assign addr[3034]= 1272139887;
assign addr[3035]= 1145766716;
assign addr[3036]= 1013581418;
assign addr[3037]= 876254528;
assign addr[3038]= 734482665;
assign addr[3039]= 588984994;
assign addr[3040]= 440499581;
assign addr[3041]= 289779648;
assign addr[3042]= 137589750;
assign addr[3043]= -15298099;
assign addr[3044]= -168108346;
assign addr[3045]= -320065829;
assign addr[3046]= -470399716;
assign addr[3047]= -618347408;
assign addr[3048]= -763158411;
assign addr[3049]= -904098143;
assign addr[3050]= -1040451659;
assign addr[3051]= -1171527280;
assign addr[3052]= -1296660098;
assign addr[3053]= -1415215352;
assign addr[3054]= -1526591649;
assign addr[3055]= -1630224009;
assign addr[3056]= -1725586737;
assign addr[3057]= -1812196087;
assign addr[3058]= -1889612716;
assign addr[3059]= -1957443913;
assign addr[3060]= -2015345591;
assign addr[3061]= -2063024031;
assign addr[3062]= -2100237377;
assign addr[3063]= -2126796855;
assign addr[3064]= -2142567738;
assign addr[3065]= -2147470025;
assign addr[3066]= -2141478848;
assign addr[3067]= -2124624598;
assign addr[3068]= -2096992772;
assign addr[3069]= -2058723538;
assign addr[3070]= -2010011024;
assign addr[3071]= -1951102334;
assign addr[3072]= -1882296293;
assign addr[3073]= -1803941934;
assign addr[3074]= -1716436725;
assign addr[3075]= -1620224553;
assign addr[3076]= -1515793473;
assign addr[3077]= -1403673233;
assign addr[3078]= -1284432584;
assign addr[3079]= -1158676398;
assign addr[3080]= -1027042599;
assign addr[3081]= -890198924;
assign addr[3082]= -748839539;
assign addr[3083]= -603681519;
assign addr[3084]= -455461206;
assign addr[3085]= -304930476;
assign addr[3086]= -152852926;
assign addr[3087]= 0;
assign addr[3088]= 152852926;
assign addr[3089]= 304930476;
assign addr[3090]= 455461206;
assign addr[3091]= 603681519;
assign addr[3092]= 748839539;
assign addr[3093]= 890198924;
assign addr[3094]= 1027042599;
assign addr[3095]= 1158676398;
assign addr[3096]= 1284432584;
assign addr[3097]= 1403673233;
assign addr[3098]= 1515793473;
assign addr[3099]= 1620224553;
assign addr[3100]= 1716436725;
assign addr[3101]= 1803941934;
assign addr[3102]= 1882296293;
assign addr[3103]= 1951102334;
assign addr[3104]= 2010011024;
assign addr[3105]= 2058723538;
assign addr[3106]= 2096992772;
assign addr[3107]= 2124624598;
assign addr[3108]= 2141478848;
assign addr[3109]= 2147470025;
assign addr[3110]= 2142567738;
assign addr[3111]= 2126796855;
assign addr[3112]= 2100237377;
assign addr[3113]= 2063024031;
assign addr[3114]= 2015345591;
assign addr[3115]= 1957443913;
assign addr[3116]= 1889612716;
assign addr[3117]= 1812196087;
assign addr[3118]= 1725586737;
assign addr[3119]= 1630224009;
assign addr[3120]= 1526591649;
assign addr[3121]= 1415215352;
assign addr[3122]= 1296660098;
assign addr[3123]= 1171527280;
assign addr[3124]= 1040451659;
assign addr[3125]= 904098143;
assign addr[3126]= 763158411;
assign addr[3127]= 618347408;
assign addr[3128]= 470399716;
assign addr[3129]= 320065829;
assign addr[3130]= 168108346;
assign addr[3131]= 15298099;
assign addr[3132]= -137589750;
assign addr[3133]= -289779648;
assign addr[3134]= -440499581;
assign addr[3135]= -588984994;
assign addr[3136]= -734482665;
assign addr[3137]= -876254528;
assign addr[3138]= -1013581418;
assign addr[3139]= -1145766716;
assign addr[3140]= -1272139887;
assign addr[3141]= -1392059879;
assign addr[3142]= -1504918373;
assign addr[3143]= -1610142873;
assign addr[3144]= -1707199606;
assign addr[3145]= -1795596234;
assign addr[3146]= -1874884346;
assign addr[3147]= -1944661739;
assign addr[3148]= -2004574453;
assign addr[3149]= -2054318569;
assign addr[3150]= -2093641749;
assign addr[3151]= -2122344521;
assign addr[3152]= -2140281282;
assign addr[3153]= -2147361045;
assign addr[3154]= -2143547897;
assign addr[3155]= -2128861181;
assign addr[3156]= -2103375398;
assign addr[3157]= -2067219829;
assign addr[3158]= -2020577882;
assign addr[3159]= -1963686155;
assign addr[3160]= -1896833245;
assign addr[3161]= -1820358275;
assign addr[3162]= -1734649179;
assign addr[3163]= -1640140734;
assign addr[3164]= -1537312353;
assign addr[3165]= -1426685652;
assign addr[3166]= -1308821808;
assign addr[3167]= -1184318708;
assign addr[3168]= -1053807919;
assign addr[3169]= -917951481;
assign addr[3170]= -777438554;
assign addr[3171]= -632981917;
assign addr[3172]= -485314355;
assign addr[3173]= -335184940;
assign addr[3174]= -183355234;
assign addr[3175]= -30595422;
assign addr[3176]= 122319591;
assign addr[3177]= 274614114;
assign addr[3178]= 425515602;
assign addr[3179]= 574258580;
assign addr[3180]= 720088517;
assign addr[3181]= 862265664;
assign addr[3182]= 1000068799;
assign addr[3183]= 1132798888;
assign addr[3184]= 1259782632;
assign addr[3185]= 1380375881;
assign addr[3186]= 1493966902;
assign addr[3187]= 1599979481;
assign addr[3188]= 1697875851;
assign addr[3189]= 1787159411;
assign addr[3190]= 1867377253;
assign addr[3191]= 1938122457;
assign addr[3192]= 1999036154;
assign addr[3193]= 2049809346;
assign addr[3194]= 2090184478;
assign addr[3195]= 2119956737;
assign addr[3196]= 2138975100;
assign addr[3197]= 2147143090;
assign addr[3198]= 2144419275;
assign addr[3199]= 2130817471;
assign addr[3200]= 2106406677;
assign addr[3201]= 2071310720;
assign addr[3202]= 2025707632;
assign addr[3203]= 1969828744;
assign addr[3204]= 1903957513;
assign addr[3205]= 1828428082;
assign addr[3206]= 1743623590;
assign addr[3207]= 1649974225;
assign addr[3208]= 1547955041;
assign addr[3209]= 1438083551;
assign addr[3210]= 1320917099;
assign addr[3211]= 1197050035;
assign addr[3212]= 1067110699;
assign addr[3213]= 931758235;
assign addr[3214]= 791679244;
assign addr[3215]= 647584304;
assign addr[3216]= 500204365;
assign addr[3217]= 350287041;
assign addr[3218]= 198592817;
assign addr[3219]= 45891193;
assign addr[3220]= -107043224;
assign addr[3221]= -259434643;
assign addr[3222]= -410510029;
assign addr[3223]= -559503022;
assign addr[3224]= -705657826;
assign addr[3225]= -848233042;
assign addr[3226]= -986505429;
assign addr[3227]= -1119773573;
assign addr[3228]= -1247361445;
assign addr[3229]= -1368621831;
assign addr[3230]= -1482939614;
assign addr[3231]= -1589734894;
assign addr[3232]= -1688465931;
assign addr[3233]= -1778631892;
assign addr[3234]= -1859775393;
assign addr[3235]= -1931484818;
assign addr[3236]= -1993396407;
assign addr[3237]= -2045196100;
assign addr[3238]= -2086621133;
assign addr[3239]= -2117461370;
assign addr[3240]= -2137560369;
assign addr[3241]= -2146816171;
assign addr[3242]= -2145181827;
assign addr[3243]= -2132665626;
assign addr[3244]= -2109331059;
assign addr[3245]= -2075296495;
assign addr[3246]= -2030734582;
assign addr[3247]= -1975871368;
assign addr[3248]= -1910985158;
assign addr[3249]= -1836405100;
assign addr[3250]= -1752509516;
assign addr[3251]= -1659723983;
assign addr[3252]= -1558519173;
assign addr[3253]= -1449408469;
assign addr[3254]= -1332945355;
assign addr[3255]= -1209720613;
assign addr[3256]= -1080359326;
assign addr[3257]= -945517704;
assign addr[3258]= -805879757;
assign addr[3259]= -662153826;
assign addr[3260]= -515068990;
assign addr[3261]= -365371365;
assign addr[3262]= -213820322;
assign addr[3263]= -61184634;
assign addr[3264]= 91761426;
assign addr[3265]= 244242007;
assign addr[3266]= 395483624;
assign addr[3267]= 544719071;
assign addr[3268]= 691191324;
assign addr[3269]= 834157373;
assign addr[3270]= 972891995;
assign addr[3271]= 1106691431;
assign addr[3272]= 1234876957;
assign addr[3273]= 1356798326;
assign addr[3274]= 1471837070;
assign addr[3275]= 1579409630;
assign addr[3276]= 1678970324;
assign addr[3277]= 1770014111;
assign addr[3278]= 1852079154;
assign addr[3279]= 1924749160;
assign addr[3280]= 1987655498;
assign addr[3281]= 2040479063;
assign addr[3282]= 2082951896;
assign addr[3283]= 2114858546;
assign addr[3284]= 2136037160;
assign addr[3285]= 2146380306;
assign addr[3286]= 2145835515;
assign addr[3287]= 2134405552;
assign addr[3288]= 2112148396;
assign addr[3289]= 2079176953;
assign addr[3290]= 2035658475;
assign addr[3291]= 1981813720;
assign addr[3292]= 1917915825;
assign addr[3293]= 1844288924;
assign addr[3294]= 1761306505;
assign addr[3295]= 1669389513;
assign addr[3296]= 1569004214;
assign addr[3297]= 1460659832;
assign addr[3298]= 1344905966;
assign addr[3299]= 1222329801;
assign addr[3300]= 1093553126;
assign addr[3301]= 959229189;
assign addr[3302]= 820039373;
assign addr[3303]= 676689746;
assign addr[3304]= 529907477;
assign addr[3305]= 380437148;
assign addr[3306]= 229036977;
assign addr[3307]= 76474970;
assign addr[3308]= -76474970;
assign addr[3309]= -229036977;
assign addr[3310]= -380437148;
assign addr[3311]= -529907477;
assign addr[3312]= -676689746;
assign addr[3313]= -820039373;
assign addr[3314]= -959229189;
assign addr[3315]= -1093553126;
assign addr[3316]= -1222329801;
assign addr[3317]= -1344905966;
assign addr[3318]= -1460659832;
assign addr[3319]= -1569004214;
assign addr[3320]= -1669389513;
assign addr[3321]= -1761306505;
assign addr[3322]= -1844288924;
assign addr[3323]= -1917915825;
assign addr[3324]= -1981813720;
assign addr[3325]= -2035658475;
assign addr[3326]= -2079176953;
assign addr[3327]= -2112148396;
assign addr[3328]= -2134405552;
assign addr[3329]= -2145835515;
assign addr[3330]= -2146380306;
assign addr[3331]= -2136037160;
assign addr[3332]= -2114858546;
assign addr[3333]= -2082951896;
assign addr[3334]= -2040479063;
assign addr[3335]= -1987655498;
assign addr[3336]= -1924749160;
assign addr[3337]= -1852079154;
assign addr[3338]= -1770014111;
assign addr[3339]= -1678970324;
assign addr[3340]= -1579409630;
assign addr[3341]= -1471837070;
assign addr[3342]= -1356798326;
assign addr[3343]= -1234876957;
assign addr[3344]= -1106691431;
assign addr[3345]= -972891995;
assign addr[3346]= -834157373;
assign addr[3347]= -691191324;
assign addr[3348]= -544719071;
assign addr[3349]= -395483624;
assign addr[3350]= -244242007;
assign addr[3351]= -91761426;
assign addr[3352]= 61184634;
assign addr[3353]= 213820322;
assign addr[3354]= 365371365;
assign addr[3355]= 515068990;
assign addr[3356]= 662153826;
assign addr[3357]= 805879757;
assign addr[3358]= 945517704;
assign addr[3359]= 1080359326;
assign addr[3360]= 1209720613;
assign addr[3361]= 1332945355;
assign addr[3362]= 1449408469;
assign addr[3363]= 1558519173;
assign addr[3364]= 1659723983;
assign addr[3365]= 1752509516;
assign addr[3366]= 1836405100;
assign addr[3367]= 1910985158;
assign addr[3368]= 1975871368;
assign addr[3369]= 2030734582;
assign addr[3370]= 2075296495;
assign addr[3371]= 2109331059;
assign addr[3372]= 2132665626;
assign addr[3373]= 2145181827;
assign addr[3374]= 2146816171;
assign addr[3375]= 2137560369;
assign addr[3376]= 2117461370;
assign addr[3377]= 2086621133;
assign addr[3378]= 2045196100;
assign addr[3379]= 1993396407;
assign addr[3380]= 1931484818;
assign addr[3381]= 1859775393;
assign addr[3382]= 1778631892;
assign addr[3383]= 1688465931;
assign addr[3384]= 1589734894;
assign addr[3385]= 1482939614;
assign addr[3386]= 1368621831;
assign addr[3387]= 1247361445;
assign addr[3388]= 1119773573;
assign addr[3389]= 986505429;
assign addr[3390]= 848233042;
assign addr[3391]= 705657826;
assign addr[3392]= 559503022;
assign addr[3393]= 410510029;
assign addr[3394]= 259434643;
assign addr[3395]= 107043224;
assign addr[3396]= -45891193;
assign addr[3397]= -198592817;
assign addr[3398]= -350287041;
assign addr[3399]= -500204365;
assign addr[3400]= -647584304;
assign addr[3401]= -791679244;
assign addr[3402]= -931758235;
assign addr[3403]= -1067110699;
assign addr[3404]= -1197050035;
assign addr[3405]= -1320917099;
assign addr[3406]= -1438083551;
assign addr[3407]= -1547955041;
assign addr[3408]= -1649974225;
assign addr[3409]= -1743623590;
assign addr[3410]= -1828428082;
assign addr[3411]= -1903957513;
assign addr[3412]= -1969828744;
assign addr[3413]= -2025707632;
assign addr[3414]= -2071310720;
assign addr[3415]= -2106406677;
assign addr[3416]= -2130817471;
assign addr[3417]= -2144419275;
assign addr[3418]= -2147143090;
assign addr[3419]= -2138975100;
assign addr[3420]= -2119956737;
assign addr[3421]= -2090184478;
assign addr[3422]= -2049809346;
assign addr[3423]= -1999036154;
assign addr[3424]= -1938122457;
assign addr[3425]= -1867377253;
assign addr[3426]= -1787159411;
assign addr[3427]= -1697875851;
assign addr[3428]= -1599979481;
assign addr[3429]= -1493966902;
assign addr[3430]= -1380375881;
assign addr[3431]= -1259782632;
assign addr[3432]= -1132798888;
assign addr[3433]= -1000068799;
assign addr[3434]= -862265664;
assign addr[3435]= -720088517;
assign addr[3436]= -574258580;
assign addr[3437]= -425515602;
assign addr[3438]= -274614114;
assign addr[3439]= -122319591;
assign addr[3440]= 30595422;
assign addr[3441]= 183355234;
assign addr[3442]= 335184940;
assign addr[3443]= 485314355;
assign addr[3444]= 632981917;
assign addr[3445]= 777438554;
assign addr[3446]= 917951481;
assign addr[3447]= 1053807919;
assign addr[3448]= 1184318708;
assign addr[3449]= 1308821808;
assign addr[3450]= 1426685652;
assign addr[3451]= 1537312353;
assign addr[3452]= 1640140734;
assign addr[3453]= 1734649179;
assign addr[3454]= 1820358275;
assign addr[3455]= 1896833245;
assign addr[3456]= 1963686155;
assign addr[3457]= 2020577882;
assign addr[3458]= 2067219829;
assign addr[3459]= 2103375398;
assign addr[3460]= 2128861181;
assign addr[3461]= 2143547897;
assign addr[3462]= 2147361045;
assign addr[3463]= 2140281282;
assign addr[3464]= 2122344521;
assign addr[3465]= 2093641749;
assign addr[3466]= 2054318569;
assign addr[3467]= 2004574453;
assign addr[3468]= 1944661739;
assign addr[3469]= 1874884346;
assign addr[3470]= 1795596234;
assign addr[3471]= 1707199606;
assign addr[3472]= 1610142873;
assign addr[3473]= 1504918373;
assign addr[3474]= 1392059879;
assign addr[3475]= 1272139887;
assign addr[3476]= 1145766716;
assign addr[3477]= 1013581418;
assign addr[3478]= 876254528;
assign addr[3479]= 734482665;
assign addr[3480]= 588984994;
assign addr[3481]= 440499581;
assign addr[3482]= 289779648;
assign addr[3483]= 137589750;
assign addr[3484]= -15298099;
assign addr[3485]= -168108346;
assign addr[3486]= -320065829;
assign addr[3487]= -470399716;
assign addr[3488]= -618347408;
assign addr[3489]= -763158411;
assign addr[3490]= -904098143;
assign addr[3491]= -1040451659;
assign addr[3492]= -1171527280;
assign addr[3493]= -1296660098;
assign addr[3494]= -1415215352;
assign addr[3495]= -1526591649;
assign addr[3496]= -1630224009;
assign addr[3497]= -1725586737;
assign addr[3498]= -1812196087;
assign addr[3499]= -1889612716;
assign addr[3500]= -1957443913;
assign addr[3501]= -2015345591;
assign addr[3502]= -2063024031;
assign addr[3503]= -2100237377;
assign addr[3504]= -2126796855;
assign addr[3505]= -2142567738;
assign addr[3506]= -2147470025;
assign addr[3507]= -2141478848;
assign addr[3508]= -2124624598;
assign addr[3509]= -2096992772;
assign addr[3510]= -2058723538;
assign addr[3511]= -2010011024;
assign addr[3512]= -1951102334;
assign addr[3513]= -1882296293;
assign addr[3514]= -1803941934;
assign addr[3515]= -1716436725;
assign addr[3516]= -1620224553;
assign addr[3517]= -1515793473;
assign addr[3518]= -1403673233;
assign addr[3519]= -1284432584;
assign addr[3520]= -1158676398;
assign addr[3521]= -1027042599;
assign addr[3522]= -890198924;
assign addr[3523]= -748839539;
assign addr[3524]= -603681519;
assign addr[3525]= -455461206;
assign addr[3526]= -304930476;
assign addr[3527]= -152852926;
assign addr[3528]= 0;
assign addr[3529]= 152852926;
assign addr[3530]= 304930476;
assign addr[3531]= 455461206;
assign addr[3532]= 603681519;
assign addr[3533]= 748839539;
assign addr[3534]= 890198924;
assign addr[3535]= 1027042599;
assign addr[3536]= 1158676398;
assign addr[3537]= 1284432584;
assign addr[3538]= 1403673233;
assign addr[3539]= 1515793473;
assign addr[3540]= 1620224553;
assign addr[3541]= 1716436725;
assign addr[3542]= 1803941934;
assign addr[3543]= 1882296293;
assign addr[3544]= 1951102334;
assign addr[3545]= 2010011024;
assign addr[3546]= 2058723538;
assign addr[3547]= 2096992772;
assign addr[3548]= 2124624598;
assign addr[3549]= 2141478848;
assign addr[3550]= 2147470025;
assign addr[3551]= 2142567738;
assign addr[3552]= 2126796855;
assign addr[3553]= 2100237377;
assign addr[3554]= 2063024031;
assign addr[3555]= 2015345591;
assign addr[3556]= 1957443913;
assign addr[3557]= 1889612716;
assign addr[3558]= 1812196087;
assign addr[3559]= 1725586737;
assign addr[3560]= 1630224009;
assign addr[3561]= 1526591649;
assign addr[3562]= 1415215352;
assign addr[3563]= 1296660098;
assign addr[3564]= 1171527280;
assign addr[3565]= 1040451659;
assign addr[3566]= 904098143;
assign addr[3567]= 763158411;
assign addr[3568]= 618347408;
assign addr[3569]= 470399716;
assign addr[3570]= 320065829;
assign addr[3571]= 168108346;
assign addr[3572]= 15298099;
assign addr[3573]= -137589750;
assign addr[3574]= -289779648;
assign addr[3575]= -440499581;
assign addr[3576]= -588984994;
assign addr[3577]= -734482665;
assign addr[3578]= -876254528;
assign addr[3579]= -1013581418;
assign addr[3580]= -1145766716;
assign addr[3581]= -1272139887;
assign addr[3582]= -1392059879;
assign addr[3583]= -1504918373;
assign addr[3584]= -1610142873;
assign addr[3585]= -1707199606;
assign addr[3586]= -1795596234;
assign addr[3587]= -1874884346;
assign addr[3588]= -1944661739;
assign addr[3589]= -2004574453;
assign addr[3590]= -2054318569;
assign addr[3591]= -2093641749;
assign addr[3592]= -2122344521;
assign addr[3593]= -2140281282;
assign addr[3594]= -2147361045;
assign addr[3595]= -2143547897;
assign addr[3596]= -2128861181;
assign addr[3597]= -2103375398;
assign addr[3598]= -2067219829;
assign addr[3599]= -2020577882;
assign addr[3600]= -1963686155;
assign addr[3601]= -1896833245;
assign addr[3602]= -1820358275;
assign addr[3603]= -1734649179;
assign addr[3604]= -1640140734;
assign addr[3605]= -1537312353;
assign addr[3606]= -1426685652;
assign addr[3607]= -1308821808;
assign addr[3608]= -1184318708;
assign addr[3609]= -1053807919;
assign addr[3610]= -917951481;
assign addr[3611]= -777438554;
assign addr[3612]= -632981917;
assign addr[3613]= -485314355;
assign addr[3614]= -335184940;
assign addr[3615]= -183355234;
assign addr[3616]= -30595422;
assign addr[3617]= 122319591;
assign addr[3618]= 274614114;
assign addr[3619]= 425515602;
assign addr[3620]= 574258580;
assign addr[3621]= 720088517;
assign addr[3622]= 862265664;
assign addr[3623]= 1000068799;
assign addr[3624]= 1132798888;
assign addr[3625]= 1259782632;
assign addr[3626]= 1380375881;
assign addr[3627]= 1493966902;
assign addr[3628]= 1599979481;
assign addr[3629]= 1697875851;
assign addr[3630]= 1787159411;
assign addr[3631]= 1867377253;
assign addr[3632]= 1938122457;
assign addr[3633]= 1999036154;
assign addr[3634]= 2049809346;
assign addr[3635]= 2090184478;
assign addr[3636]= 2119956737;
assign addr[3637]= 2138975100;
assign addr[3638]= 2147143090;
assign addr[3639]= 2144419275;
assign addr[3640]= 2130817471;
assign addr[3641]= 2106406677;
assign addr[3642]= 2071310720;
assign addr[3643]= 2025707632;
assign addr[3644]= 1969828744;
assign addr[3645]= 1903957513;
assign addr[3646]= 1828428082;
assign addr[3647]= 1743623590;
assign addr[3648]= 1649974225;
assign addr[3649]= 1547955041;
assign addr[3650]= 1438083551;
assign addr[3651]= 1320917099;
assign addr[3652]= 1197050035;
assign addr[3653]= 1067110699;
assign addr[3654]= 931758235;
assign addr[3655]= 791679244;
assign addr[3656]= 647584304;
assign addr[3657]= 500204365;
assign addr[3658]= 350287041;
assign addr[3659]= 198592817;
assign addr[3660]= 45891193;
assign addr[3661]= -107043224;
assign addr[3662]= -259434643;
assign addr[3663]= -410510029;
assign addr[3664]= -559503022;
assign addr[3665]= -705657826;
assign addr[3666]= -848233042;
assign addr[3667]= -986505429;
assign addr[3668]= -1119773573;
assign addr[3669]= -1247361445;
assign addr[3670]= -1368621831;
assign addr[3671]= -1482939614;
assign addr[3672]= -1589734894;
assign addr[3673]= -1688465931;
assign addr[3674]= -1778631892;
assign addr[3675]= -1859775393;
assign addr[3676]= -1931484818;
assign addr[3677]= -1993396407;
assign addr[3678]= -2045196100;
assign addr[3679]= -2086621133;
assign addr[3680]= -2117461370;
assign addr[3681]= -2137560369;
assign addr[3682]= -2146816171;
assign addr[3683]= -2145181827;
assign addr[3684]= -2132665626;
assign addr[3685]= -2109331059;
assign addr[3686]= -2075296495;
assign addr[3687]= -2030734582;
assign addr[3688]= -1975871368;
assign addr[3689]= -1910985158;
assign addr[3690]= -1836405100;
assign addr[3691]= -1752509516;
assign addr[3692]= -1659723983;
assign addr[3693]= -1558519173;
assign addr[3694]= -1449408469;
assign addr[3695]= -1332945355;
assign addr[3696]= -1209720613;
assign addr[3697]= -1080359326;
assign addr[3698]= -945517704;
assign addr[3699]= -805879757;
assign addr[3700]= -662153826;
assign addr[3701]= -515068990;
assign addr[3702]= -365371365;
assign addr[3703]= -213820322;
assign addr[3704]= -61184634;
assign addr[3705]= 91761426;
assign addr[3706]= 244242007;
assign addr[3707]= 395483624;
assign addr[3708]= 544719071;
assign addr[3709]= 691191324;
assign addr[3710]= 834157373;
assign addr[3711]= 972891995;
assign addr[3712]= 1106691431;
assign addr[3713]= 1234876957;
assign addr[3714]= 1356798326;
assign addr[3715]= 1471837070;
assign addr[3716]= 1579409630;
assign addr[3717]= 1678970324;
assign addr[3718]= 1770014111;
assign addr[3719]= 1852079154;
assign addr[3720]= 1924749160;
assign addr[3721]= 1987655498;
assign addr[3722]= 2040479063;
assign addr[3723]= 2082951896;
assign addr[3724]= 2114858546;
assign addr[3725]= 2136037160;
assign addr[3726]= 2146380306;
assign addr[3727]= 2145835515;
assign addr[3728]= 2134405552;
assign addr[3729]= 2112148396;
assign addr[3730]= 2079176953;
assign addr[3731]= 2035658475;
assign addr[3732]= 1981813720;
assign addr[3733]= 1917915825;
assign addr[3734]= 1844288924;
assign addr[3735]= 1761306505;
assign addr[3736]= 1669389513;
assign addr[3737]= 1569004214;
assign addr[3738]= 1460659832;
assign addr[3739]= 1344905966;
assign addr[3740]= 1222329801;
assign addr[3741]= 1093553126;
assign addr[3742]= 959229189;
assign addr[3743]= 820039373;
assign addr[3744]= 676689746;
assign addr[3745]= 529907477;
assign addr[3746]= 380437148;
assign addr[3747]= 229036977;
assign addr[3748]= 76474970;
assign addr[3749]= -76474970;
assign addr[3750]= -229036977;
assign addr[3751]= -380437148;
assign addr[3752]= -529907477;
assign addr[3753]= -676689746;
assign addr[3754]= -820039373;
assign addr[3755]= -959229189;
assign addr[3756]= -1093553126;
assign addr[3757]= -1222329801;
assign addr[3758]= -1344905966;
assign addr[3759]= -1460659832;
assign addr[3760]= -1569004214;
assign addr[3761]= -1669389513;
assign addr[3762]= -1761306505;
assign addr[3763]= -1844288924;
assign addr[3764]= -1917915825;
assign addr[3765]= -1981813720;
assign addr[3766]= -2035658475;
assign addr[3767]= -2079176953;
assign addr[3768]= -2112148396;
assign addr[3769]= -2134405552;
assign addr[3770]= -2145835515;
assign addr[3771]= -2146380306;
assign addr[3772]= -2136037160;
assign addr[3773]= -2114858546;
assign addr[3774]= -2082951896;
assign addr[3775]= -2040479063;
assign addr[3776]= -1987655498;
assign addr[3777]= -1924749160;
assign addr[3778]= -1852079154;
assign addr[3779]= -1770014111;
assign addr[3780]= -1678970324;
assign addr[3781]= -1579409630;
assign addr[3782]= -1471837070;
assign addr[3783]= -1356798326;
assign addr[3784]= -1234876957;
assign addr[3785]= -1106691431;
assign addr[3786]= -972891995;
assign addr[3787]= -834157373;
assign addr[3788]= -691191324;
assign addr[3789]= -544719071;
assign addr[3790]= -395483624;
assign addr[3791]= -244242007;
assign addr[3792]= -91761426;
assign addr[3793]= 61184634;
assign addr[3794]= 213820322;
assign addr[3795]= 365371365;
assign addr[3796]= 515068990;
assign addr[3797]= 662153826;
assign addr[3798]= 805879757;
assign addr[3799]= 945517704;
assign addr[3800]= 1080359326;
assign addr[3801]= 1209720613;
assign addr[3802]= 1332945355;
assign addr[3803]= 1449408469;
assign addr[3804]= 1558519173;
assign addr[3805]= 1659723983;
assign addr[3806]= 1752509516;
assign addr[3807]= 1836405100;
assign addr[3808]= 1910985158;
assign addr[3809]= 1975871368;
assign addr[3810]= 2030734582;
assign addr[3811]= 2075296495;
assign addr[3812]= 2109331059;
assign addr[3813]= 2132665626;
assign addr[3814]= 2145181827;
assign addr[3815]= 2146816171;
assign addr[3816]= 2137560369;
assign addr[3817]= 2117461370;
assign addr[3818]= 2086621133;
assign addr[3819]= 2045196100;
assign addr[3820]= 1993396407;
assign addr[3821]= 1931484818;
assign addr[3822]= 1859775393;
assign addr[3823]= 1778631892;
assign addr[3824]= 1688465931;
assign addr[3825]= 1589734894;
assign addr[3826]= 1482939614;
assign addr[3827]= 1368621831;
assign addr[3828]= 1247361445;
assign addr[3829]= 1119773573;
assign addr[3830]= 986505429;
assign addr[3831]= 848233042;
assign addr[3832]= 705657826;
assign addr[3833]= 559503022;
assign addr[3834]= 410510029;
assign addr[3835]= 259434643;
assign addr[3836]= 107043224;
assign addr[3837]= -45891193;
assign addr[3838]= -198592817;
assign addr[3839]= -350287041;
assign addr[3840]= -500204365;
assign addr[3841]= -647584304;
assign addr[3842]= -791679244;
assign addr[3843]= -931758235;
assign addr[3844]= -1067110699;
assign addr[3845]= -1197050035;
assign addr[3846]= -1320917099;
assign addr[3847]= -1438083551;
assign addr[3848]= -1547955041;
assign addr[3849]= -1649974225;
assign addr[3850]= -1743623590;
assign addr[3851]= -1828428082;
assign addr[3852]= -1903957513;
assign addr[3853]= -1969828744;
assign addr[3854]= -2025707632;
assign addr[3855]= -2071310720;
assign addr[3856]= -2106406677;
assign addr[3857]= -2130817471;
assign addr[3858]= -2144419275;
assign addr[3859]= -2147143090;
assign addr[3860]= -2138975100;
assign addr[3861]= -2119956737;
assign addr[3862]= -2090184478;
assign addr[3863]= -2049809346;
assign addr[3864]= -1999036154;
assign addr[3865]= -1938122457;
assign addr[3866]= -1867377253;
assign addr[3867]= -1787159411;
assign addr[3868]= -1697875851;
assign addr[3869]= -1599979481;
assign addr[3870]= -1493966902;
assign addr[3871]= -1380375881;
assign addr[3872]= -1259782632;
assign addr[3873]= -1132798888;
assign addr[3874]= -1000068799;
assign addr[3875]= -862265664;
assign addr[3876]= -720088517;
assign addr[3877]= -574258580;
assign addr[3878]= -425515602;
assign addr[3879]= -274614114;
assign addr[3880]= -122319591;
assign addr[3881]= 30595422;
assign addr[3882]= 183355234;
assign addr[3883]= 335184940;
assign addr[3884]= 485314355;
assign addr[3885]= 632981917;
assign addr[3886]= 777438554;
assign addr[3887]= 917951481;
assign addr[3888]= 1053807919;
assign addr[3889]= 1184318708;
assign addr[3890]= 1308821808;
assign addr[3891]= 1426685652;
assign addr[3892]= 1537312353;
assign addr[3893]= 1640140734;
assign addr[3894]= 1734649179;
assign addr[3895]= 1820358275;
assign addr[3896]= 1896833245;
assign addr[3897]= 1963686155;
assign addr[3898]= 2020577882;
assign addr[3899]= 2067219829;
assign addr[3900]= 2103375398;
assign addr[3901]= 2128861181;
assign addr[3902]= 2143547897;
assign addr[3903]= 2147361045;
assign addr[3904]= 2140281282;
assign addr[3905]= 2122344521;
assign addr[3906]= 2093641749;
assign addr[3907]= 2054318569;
assign addr[3908]= 2004574453;
assign addr[3909]= 1944661739;
assign addr[3910]= 1874884346;
assign addr[3911]= 1795596234;
assign addr[3912]= 1707199606;
assign addr[3913]= 1610142873;
assign addr[3914]= 1504918373;
assign addr[3915]= 1392059879;
assign addr[3916]= 1272139887;
assign addr[3917]= 1145766716;
assign addr[3918]= 1013581418;
assign addr[3919]= 876254528;
assign addr[3920]= 734482665;
assign addr[3921]= 588984994;
assign addr[3922]= 440499581;
assign addr[3923]= 289779648;
assign addr[3924]= 137589750;
assign addr[3925]= -15298099;
assign addr[3926]= -168108346;
assign addr[3927]= -320065829;
assign addr[3928]= -470399716;
assign addr[3929]= -618347408;
assign addr[3930]= -763158411;
assign addr[3931]= -904098143;
assign addr[3932]= -1040451659;
assign addr[3933]= -1171527280;
assign addr[3934]= -1296660098;
assign addr[3935]= -1415215352;
assign addr[3936]= -1526591649;
assign addr[3937]= -1630224009;
assign addr[3938]= -1725586737;
assign addr[3939]= -1812196087;
assign addr[3940]= -1889612716;
assign addr[3941]= -1957443913;
assign addr[3942]= -2015345591;
assign addr[3943]= -2063024031;
assign addr[3944]= -2100237377;
assign addr[3945]= -2126796855;
assign addr[3946]= -2142567738;
assign addr[3947]= -2147470025;
assign addr[3948]= -2141478848;
assign addr[3949]= -2124624598;
assign addr[3950]= -2096992772;
assign addr[3951]= -2058723538;
assign addr[3952]= -2010011024;
assign addr[3953]= -1951102334;
assign addr[3954]= -1882296293;
assign addr[3955]= -1803941934;
assign addr[3956]= -1716436725;
assign addr[3957]= -1620224553;
assign addr[3958]= -1515793473;
assign addr[3959]= -1403673233;
assign addr[3960]= -1284432584;
assign addr[3961]= -1158676398;
assign addr[3962]= -1027042599;
assign addr[3963]= -890198924;
assign addr[3964]= -748839539;
assign addr[3965]= -603681519;
assign addr[3966]= -455461206;
assign addr[3967]= -304930476;
assign addr[3968]= -152852926;
assign addr[3969]= 0;
assign addr[3970]= 152852926;
assign addr[3971]= 304930476;
assign addr[3972]= 455461206;
assign addr[3973]= 603681519;
assign addr[3974]= 748839539;
assign addr[3975]= 890198924;
assign addr[3976]= 1027042599;
assign addr[3977]= 1158676398;
assign addr[3978]= 1284432584;
assign addr[3979]= 1403673233;
assign addr[3980]= 1515793473;
assign addr[3981]= 1620224553;
assign addr[3982]= 1716436725;
assign addr[3983]= 1803941934;
assign addr[3984]= 1882296293;
assign addr[3985]= 1951102334;
assign addr[3986]= 2010011024;
assign addr[3987]= 2058723538;
assign addr[3988]= 2096992772;
assign addr[3989]= 2124624598;
assign addr[3990]= 2141478848;
assign addr[3991]= 2147470025;
assign addr[3992]= 2142567738;
assign addr[3993]= 2126796855;
assign addr[3994]= 2100237377;
assign addr[3995]= 2063024031;
assign addr[3996]= 2015345591;
assign addr[3997]= 1957443913;
assign addr[3998]= 1889612716;
assign addr[3999]= 1812196087;
assign addr[4000]= 1725586737;
assign addr[4001]= 1630224009;
assign addr[4002]= 1526591649;
assign addr[4003]= 1415215352;
assign addr[4004]= 1296660098;
assign addr[4005]= 1171527280;
assign addr[4006]= 1040451659;
assign addr[4007]= 904098143;
assign addr[4008]= 763158411;
assign addr[4009]= 618347408;
assign addr[4010]= 470399716;
assign addr[4011]= 320065829;
assign addr[4012]= 168108346;
assign addr[4013]= 15298099;
assign addr[4014]= -137589750;
assign addr[4015]= -289779648;
assign addr[4016]= -440499581;
assign addr[4017]= -588984994;
assign addr[4018]= -734482665;
assign addr[4019]= -876254528;
assign addr[4020]= -1013581418;
assign addr[4021]= -1145766716;
assign addr[4022]= -1272139887;
assign addr[4023]= -1392059879;
assign addr[4024]= -1504918373;
assign addr[4025]= -1610142873;
assign addr[4026]= -1707199606;
assign addr[4027]= -1795596234;
assign addr[4028]= -1874884346;
assign addr[4029]= -1944661739;
assign addr[4030]= -2004574453;
assign addr[4031]= -2054318569;
assign addr[4032]= -2093641749;
assign addr[4033]= -2122344521;
assign addr[4034]= -2140281282;
assign addr[4035]= -2147361045;
assign addr[4036]= -2143547897;
assign addr[4037]= -2128861181;
assign addr[4038]= -2103375398;
assign addr[4039]= -2067219829;
assign addr[4040]= -2020577882;
assign addr[4041]= -1963686155;
assign addr[4042]= -1896833245;
assign addr[4043]= -1820358275;
assign addr[4044]= -1734649179;
assign addr[4045]= -1640140734;
assign addr[4046]= -1537312353;
assign addr[4047]= -1426685652;
assign addr[4048]= -1308821808;
assign addr[4049]= -1184318708;
assign addr[4050]= -1053807919;
assign addr[4051]= -917951481;
assign addr[4052]= -777438554;
assign addr[4053]= -632981917;
assign addr[4054]= -485314355;
assign addr[4055]= -335184940;
assign addr[4056]= -183355234;
assign addr[4057]= -30595422;
assign addr[4058]= 122319591;
assign addr[4059]= 274614114;
assign addr[4060]= 425515602;
assign addr[4061]= 574258580;
assign addr[4062]= 720088517;
assign addr[4063]= 862265664;
assign addr[4064]= 1000068799;
assign addr[4065]= 1132798888;
assign addr[4066]= 1259782632;
assign addr[4067]= 1380375881;
assign addr[4068]= 1493966902;
assign addr[4069]= 1599979481;
assign addr[4070]= 1697875851;
assign addr[4071]= 1787159411;
assign addr[4072]= 1867377253;
assign addr[4073]= 1938122457;
assign addr[4074]= 1999036154;
assign addr[4075]= 2049809346;
assign addr[4076]= 2090184478;
assign addr[4077]= 2119956737;
assign addr[4078]= 2138975100;
assign addr[4079]= 2147143090;
assign addr[4080]= 2144419275;
assign addr[4081]= 2130817471;
assign addr[4082]= 2106406677;
assign addr[4083]= 2071310720;
assign addr[4084]= 2025707632;
assign addr[4085]= 1969828744;
assign addr[4086]= 1903957513;
assign addr[4087]= 1828428082;
assign addr[4088]= 1743623590;
assign addr[4089]= 1649974225;
assign addr[4090]= 1547955041;
assign addr[4091]= 1438083551;
assign addr[4092]= 1320917099;
assign addr[4093]= 1197050035;
assign addr[4094]= 1067110699;
assign addr[4095]= 931758235;
assign addr[4096]= 791679244;
assign addr[4097]= 647584304;
assign addr[4098]= 500204365;
assign addr[4099]= 350287041;
assign addr[4100]= 198592817;
assign addr[4101]= 45891193;
assign addr[4102]= -107043224;
assign addr[4103]= -259434643;
assign addr[4104]= -410510029;
assign addr[4105]= -559503022;
assign addr[4106]= -705657826;
assign addr[4107]= -848233042;
assign addr[4108]= -986505429;
assign addr[4109]= -1119773573;
assign addr[4110]= -1247361445;
assign addr[4111]= -1368621831;
assign addr[4112]= -1482939614;
assign addr[4113]= -1589734894;
assign addr[4114]= -1688465931;
assign addr[4115]= -1778631892;
assign addr[4116]= -1859775393;
assign addr[4117]= -1931484818;
assign addr[4118]= -1993396407;
assign addr[4119]= -2045196100;
assign addr[4120]= -2086621133;
assign addr[4121]= -2117461370;
assign addr[4122]= -2137560369;
assign addr[4123]= -2146816171;
assign addr[4124]= -2145181827;
assign addr[4125]= -2132665626;
assign addr[4126]= -2109331059;
assign addr[4127]= -2075296495;
assign addr[4128]= -2030734582;
assign addr[4129]= -1975871368;
assign addr[4130]= -1910985158;
assign addr[4131]= -1836405100;
assign addr[4132]= -1752509516;
assign addr[4133]= -1659723983;
assign addr[4134]= -1558519173;
assign addr[4135]= -1449408469;
assign addr[4136]= -1332945355;
assign addr[4137]= -1209720613;
assign addr[4138]= -1080359326;
assign addr[4139]= -945517704;
assign addr[4140]= -805879757;
assign addr[4141]= -662153826;
assign addr[4142]= -515068990;
assign addr[4143]= -365371365;
assign addr[4144]= -213820322;
assign addr[4145]= -61184634;
assign addr[4146]= 91761426;
assign addr[4147]= 244242007;
assign addr[4148]= 395483624;
assign addr[4149]= 544719071;
assign addr[4150]= 691191324;
assign addr[4151]= 834157373;
assign addr[4152]= 972891995;
assign addr[4153]= 1106691431;
assign addr[4154]= 1234876957;
assign addr[4155]= 1356798326;
assign addr[4156]= 1471837070;
assign addr[4157]= 1579409630;
assign addr[4158]= 1678970324;
assign addr[4159]= 1770014111;
assign addr[4160]= 1852079154;
assign addr[4161]= 1924749160;
assign addr[4162]= 1987655498;
assign addr[4163]= 2040479063;
assign addr[4164]= 2082951896;
assign addr[4165]= 2114858546;
assign addr[4166]= 2136037160;
assign addr[4167]= 2146380306;
assign addr[4168]= 2145835515;
assign addr[4169]= 2134405552;
assign addr[4170]= 2112148396;
assign addr[4171]= 2079176953;
assign addr[4172]= 2035658475;
assign addr[4173]= 1981813720;
assign addr[4174]= 1917915825;
assign addr[4175]= 1844288924;
assign addr[4176]= 1761306505;
assign addr[4177]= 1669389513;
assign addr[4178]= 1569004214;
assign addr[4179]= 1460659832;
assign addr[4180]= 1344905966;
assign addr[4181]= 1222329801;
assign addr[4182]= 1093553126;
assign addr[4183]= 959229189;
assign addr[4184]= 820039373;
assign addr[4185]= 676689746;
assign addr[4186]= 529907477;
assign addr[4187]= 380437148;
assign addr[4188]= 229036977;
assign addr[4189]= 76474970;
assign addr[4190]= -76474970;
assign addr[4191]= -229036977;
assign addr[4192]= -380437148;
assign addr[4193]= -529907477;
assign addr[4194]= -676689746;
assign addr[4195]= -820039373;
assign addr[4196]= -959229189;
assign addr[4197]= -1093553126;
assign addr[4198]= -1222329801;
assign addr[4199]= -1344905966;
assign addr[4200]= -1460659832;
assign addr[4201]= -1569004214;
assign addr[4202]= -1669389513;
assign addr[4203]= -1761306505;
assign addr[4204]= -1844288924;
assign addr[4205]= -1917915825;
assign addr[4206]= -1981813720;
assign addr[4207]= -2035658475;
assign addr[4208]= -2079176953;
assign addr[4209]= -2112148396;
assign addr[4210]= -2134405552;
assign addr[4211]= -2145835515;
assign addr[4212]= -2146380306;
assign addr[4213]= -2136037160;
assign addr[4214]= -2114858546;
assign addr[4215]= -2082951896;
assign addr[4216]= -2040479063;
assign addr[4217]= -1987655498;
assign addr[4218]= -1924749160;
assign addr[4219]= -1852079154;
assign addr[4220]= -1770014111;
assign addr[4221]= -1678970324;
assign addr[4222]= -1579409630;
assign addr[4223]= -1471837070;
assign addr[4224]= -1356798326;
assign addr[4225]= -1234876957;
assign addr[4226]= -1106691431;
assign addr[4227]= -972891995;
assign addr[4228]= -834157373;
assign addr[4229]= -691191324;
assign addr[4230]= -544719071;
assign addr[4231]= -395483624;
assign addr[4232]= -244242007;
assign addr[4233]= -91761426;
assign addr[4234]= 61184634;
assign addr[4235]= 213820322;
assign addr[4236]= 365371365;
assign addr[4237]= 515068990;
assign addr[4238]= 662153826;
assign addr[4239]= 805879757;
assign addr[4240]= 945517704;
assign addr[4241]= 1080359326;
assign addr[4242]= 1209720613;
assign addr[4243]= 1332945355;
assign addr[4244]= 1449408469;
assign addr[4245]= 1558519173;
assign addr[4246]= 1659723983;
assign addr[4247]= 1752509516;
assign addr[4248]= 1836405100;
assign addr[4249]= 1910985158;
assign addr[4250]= 1975871368;
assign addr[4251]= 2030734582;
assign addr[4252]= 2075296495;
assign addr[4253]= 2109331059;
assign addr[4254]= 2132665626;
assign addr[4255]= 2145181827;
assign addr[4256]= 2146816171;
assign addr[4257]= 2137560369;
assign addr[4258]= 2117461370;
assign addr[4259]= 2086621133;
assign addr[4260]= 2045196100;
assign addr[4261]= 1993396407;
assign addr[4262]= 1931484818;
assign addr[4263]= 1859775393;
assign addr[4264]= 1778631892;
assign addr[4265]= 1688465931;
assign addr[4266]= 1589734894;
assign addr[4267]= 1482939614;
assign addr[4268]= 1368621831;
assign addr[4269]= 1247361445;
assign addr[4270]= 1119773573;
assign addr[4271]= 986505429;
assign addr[4272]= 848233042;
assign addr[4273]= 705657826;
assign addr[4274]= 559503022;
assign addr[4275]= 410510029;
assign addr[4276]= 259434643;
assign addr[4277]= 107043224;
assign addr[4278]= -45891193;
assign addr[4279]= -198592817;
assign addr[4280]= -350287041;
assign addr[4281]= -500204365;
assign addr[4282]= -647584304;
assign addr[4283]= -791679244;
assign addr[4284]= -931758235;
assign addr[4285]= -1067110699;
assign addr[4286]= -1197050035;
assign addr[4287]= -1320917099;
assign addr[4288]= -1438083551;
assign addr[4289]= -1547955041;
assign addr[4290]= -1649974225;
assign addr[4291]= -1743623590;
assign addr[4292]= -1828428082;
assign addr[4293]= -1903957513;
assign addr[4294]= -1969828744;
assign addr[4295]= -2025707632;
assign addr[4296]= -2071310720;
assign addr[4297]= -2106406677;
assign addr[4298]= -2130817471;
assign addr[4299]= -2144419275;
assign addr[4300]= -2147143090;
assign addr[4301]= -2138975100;
assign addr[4302]= -2119956737;
assign addr[4303]= -2090184478;
assign addr[4304]= -2049809346;
assign addr[4305]= -1999036154;
assign addr[4306]= -1938122457;
assign addr[4307]= -1867377253;
assign addr[4308]= -1787159411;
assign addr[4309]= -1697875851;
assign addr[4310]= -1599979481;
assign addr[4311]= -1493966902;
assign addr[4312]= -1380375881;
assign addr[4313]= -1259782632;
assign addr[4314]= -1132798888;
assign addr[4315]= -1000068799;
assign addr[4316]= -862265664;
assign addr[4317]= -720088517;
assign addr[4318]= -574258580;
assign addr[4319]= -425515602;
assign addr[4320]= -274614114;
assign addr[4321]= -122319591;
assign addr[4322]= 30595422;
assign addr[4323]= 183355234;
assign addr[4324]= 335184940;
assign addr[4325]= 485314355;
assign addr[4326]= 632981917;
assign addr[4327]= 777438554;
assign addr[4328]= 917951481;
assign addr[4329]= 1053807919;
assign addr[4330]= 1184318708;
assign addr[4331]= 1308821808;
assign addr[4332]= 1426685652;
assign addr[4333]= 1537312353;
assign addr[4334]= 1640140734;
assign addr[4335]= 1734649179;
assign addr[4336]= 1820358275;
assign addr[4337]= 1896833245;
assign addr[4338]= 1963686155;
assign addr[4339]= 2020577882;
assign addr[4340]= 2067219829;
assign addr[4341]= 2103375398;
assign addr[4342]= 2128861181;
assign addr[4343]= 2143547897;
assign addr[4344]= 2147361045;
assign addr[4345]= 2140281282;
assign addr[4346]= 2122344521;
assign addr[4347]= 2093641749;
assign addr[4348]= 2054318569;
assign addr[4349]= 2004574453;
assign addr[4350]= 1944661739;
assign addr[4351]= 1874884346;
assign addr[4352]= 1795596234;
assign addr[4353]= 1707199606;
assign addr[4354]= 1610142873;
assign addr[4355]= 1504918373;
assign addr[4356]= 1392059879;
assign addr[4357]= 1272139887;
assign addr[4358]= 1145766716;
assign addr[4359]= 1013581418;
assign addr[4360]= 876254528;
assign addr[4361]= 734482665;
assign addr[4362]= 588984994;
assign addr[4363]= 440499581;
assign addr[4364]= 289779648;
assign addr[4365]= 137589750;
assign addr[4366]= -15298099;
assign addr[4367]= -168108346;
assign addr[4368]= -320065829;
assign addr[4369]= -470399716;
assign addr[4370]= -618347408;
assign addr[4371]= -763158411;
assign addr[4372]= -904098143;
assign addr[4373]= -1040451659;
assign addr[4374]= -1171527280;
assign addr[4375]= -1296660098;
assign addr[4376]= -1415215352;
assign addr[4377]= -1526591649;
assign addr[4378]= -1630224009;
assign addr[4379]= -1725586737;
assign addr[4380]= -1812196087;
assign addr[4381]= -1889612716;
assign addr[4382]= -1957443913;
assign addr[4383]= -2015345591;
assign addr[4384]= -2063024031;
assign addr[4385]= -2100237377;
assign addr[4386]= -2126796855;
assign addr[4387]= -2142567738;
assign addr[4388]= -2147470025;
assign addr[4389]= -2141478848;
assign addr[4390]= -2124624598;
assign addr[4391]= -2096992772;
assign addr[4392]= -2058723538;
assign addr[4393]= -2010011024;
assign addr[4394]= -1951102334;
assign addr[4395]= -1882296293;
assign addr[4396]= -1803941934;
assign addr[4397]= -1716436725;
assign addr[4398]= -1620224553;
assign addr[4399]= -1515793473;
assign addr[4400]= -1403673233;
assign addr[4401]= -1284432584;
assign addr[4402]= -1158676398;
assign addr[4403]= -1027042599;
assign addr[4404]= -890198924;
assign addr[4405]= -748839539;
assign addr[4406]= -603681519;
assign addr[4407]= -455461206;
assign addr[4408]= -304930476;
assign addr[4409]= -152852926;
assign addr[4410]= 0;
assign addr[4411]= 152852926;
assign addr[4412]= 304930476;
assign addr[4413]= 455461206;
assign addr[4414]= 603681519;
assign addr[4415]= 748839539;
assign addr[4416]= 890198924;
assign addr[4417]= 1027042599;
assign addr[4418]= 1158676398;
assign addr[4419]= 1284432584;
assign addr[4420]= 1403673233;
assign addr[4421]= 1515793473;
assign addr[4422]= 1620224553;
assign addr[4423]= 1716436725;
assign addr[4424]= 1803941934;
assign addr[4425]= 1882296293;
assign addr[4426]= 1951102334;
assign addr[4427]= 2010011024;
assign addr[4428]= 2058723538;
assign addr[4429]= 2096992772;
assign addr[4430]= 2124624598;
assign addr[4431]= 2141478848;
assign addr[4432]= 2147470025;
assign addr[4433]= 2142567738;
assign addr[4434]= 2126796855;
assign addr[4435]= 2100237377;
assign addr[4436]= 2063024031;
assign addr[4437]= 2015345591;
assign addr[4438]= 1957443913;
assign addr[4439]= 1889612716;
assign addr[4440]= 1812196087;
assign addr[4441]= 1725586737;
assign addr[4442]= 1630224009;
assign addr[4443]= 1526591649;
assign addr[4444]= 1415215352;
assign addr[4445]= 1296660098;
assign addr[4446]= 1171527280;
assign addr[4447]= 1040451659;
assign addr[4448]= 904098143;
assign addr[4449]= 763158411;
assign addr[4450]= 618347408;
assign addr[4451]= 470399716;
assign addr[4452]= 320065829;
assign addr[4453]= 168108346;
assign addr[4454]= 15298099;
assign addr[4455]= -137589750;
assign addr[4456]= -289779648;
assign addr[4457]= -440499581;
assign addr[4458]= -588984994;
assign addr[4459]= -734482665;
assign addr[4460]= -876254528;
assign addr[4461]= -1013581418;
assign addr[4462]= -1145766716;
assign addr[4463]= -1272139887;
assign addr[4464]= -1392059879;
assign addr[4465]= -1504918373;
assign addr[4466]= -1610142873;
assign addr[4467]= -1707199606;
assign addr[4468]= -1795596234;
assign addr[4469]= -1874884346;
assign addr[4470]= -1944661739;
assign addr[4471]= -2004574453;
assign addr[4472]= -2054318569;
assign addr[4473]= -2093641749;
assign addr[4474]= -2122344521;
assign addr[4475]= -2140281282;
assign addr[4476]= -2147361045;
assign addr[4477]= -2143547897;
assign addr[4478]= -2128861181;
assign addr[4479]= -2103375398;
assign addr[4480]= -2067219829;
assign addr[4481]= -2020577882;
assign addr[4482]= -1963686155;
assign addr[4483]= -1896833245;
assign addr[4484]= -1820358275;
assign addr[4485]= -1734649179;
assign addr[4486]= -1640140734;
assign addr[4487]= -1537312353;
assign addr[4488]= -1426685652;
assign addr[4489]= -1308821808;
assign addr[4490]= -1184318708;
assign addr[4491]= -1053807919;
assign addr[4492]= -917951481;
assign addr[4493]= -777438554;
assign addr[4494]= -632981917;
assign addr[4495]= -485314355;
assign addr[4496]= -335184940;
assign addr[4497]= -183355234;
assign addr[4498]= -30595422;
assign addr[4499]= 122319591;
assign addr[4500]= 274614114;
assign addr[4501]= 425515602;
assign addr[4502]= 574258580;
assign addr[4503]= 720088517;
assign addr[4504]= 862265664;
assign addr[4505]= 1000068799;
assign addr[4506]= 1132798888;
assign addr[4507]= 1259782632;
assign addr[4508]= 1380375881;
assign addr[4509]= 1493966902;
assign addr[4510]= 1599979481;
assign addr[4511]= 1697875851;
assign addr[4512]= 1787159411;
assign addr[4513]= 1867377253;
assign addr[4514]= 1938122457;
assign addr[4515]= 1999036154;
assign addr[4516]= 2049809346;
assign addr[4517]= 2090184478;
assign addr[4518]= 2119956737;
assign addr[4519]= 2138975100;
assign addr[4520]= 2147143090;
assign addr[4521]= 2144419275;
assign addr[4522]= 2130817471;
assign addr[4523]= 2106406677;
assign addr[4524]= 2071310720;
assign addr[4525]= 2025707632;
assign addr[4526]= 1969828744;
assign addr[4527]= 1903957513;
assign addr[4528]= 1828428082;
assign addr[4529]= 1743623590;
assign addr[4530]= 1649974225;
assign addr[4531]= 1547955041;
assign addr[4532]= 1438083551;
assign addr[4533]= 1320917099;
assign addr[4534]= 1197050035;
assign addr[4535]= 1067110699;
assign addr[4536]= 931758235;
assign addr[4537]= 791679244;
assign addr[4538]= 647584304;
assign addr[4539]= 500204365;
assign addr[4540]= 350287041;
assign addr[4541]= 198592817;
assign addr[4542]= 45891193;
assign addr[4543]= -107043224;
assign addr[4544]= -259434643;
assign addr[4545]= -410510029;
assign addr[4546]= -559503022;
assign addr[4547]= -705657826;
assign addr[4548]= -848233042;
assign addr[4549]= -986505429;
assign addr[4550]= -1119773573;
assign addr[4551]= -1247361445;
assign addr[4552]= -1368621831;
assign addr[4553]= -1482939614;
assign addr[4554]= -1589734894;
assign addr[4555]= -1688465931;
assign addr[4556]= -1778631892;
assign addr[4557]= -1859775393;
assign addr[4558]= -1931484818;
assign addr[4559]= -1993396407;
assign addr[4560]= -2045196100;
assign addr[4561]= -2086621133;
assign addr[4562]= -2117461370;
assign addr[4563]= -2137560369;
assign addr[4564]= -2146816171;
assign addr[4565]= -2145181827;
assign addr[4566]= -2132665626;
assign addr[4567]= -2109331059;
assign addr[4568]= -2075296495;
assign addr[4569]= -2030734582;
assign addr[4570]= -1975871368;
assign addr[4571]= -1910985158;
assign addr[4572]= -1836405100;
assign addr[4573]= -1752509516;
assign addr[4574]= -1659723983;
assign addr[4575]= -1558519173;
assign addr[4576]= -1449408469;
assign addr[4577]= -1332945355;
assign addr[4578]= -1209720613;
assign addr[4579]= -1080359326;
assign addr[4580]= -945517704;
assign addr[4581]= -805879757;
assign addr[4582]= -662153826;
assign addr[4583]= -515068990;
assign addr[4584]= -365371365;
assign addr[4585]= -213820322;
assign addr[4586]= -61184634;
assign addr[4587]= 91761426;
assign addr[4588]= 244242007;
assign addr[4589]= 395483624;
assign addr[4590]= 544719071;
assign addr[4591]= 691191324;
assign addr[4592]= 834157373;
assign addr[4593]= 972891995;
assign addr[4594]= 1106691431;
assign addr[4595]= 1234876957;
assign addr[4596]= 1356798326;
assign addr[4597]= 1471837070;
assign addr[4598]= 1579409630;
assign addr[4599]= 1678970324;
assign addr[4600]= 1770014111;
assign addr[4601]= 1852079154;
assign addr[4602]= 1924749160;
assign addr[4603]= 1987655498;
assign addr[4604]= 2040479063;
assign addr[4605]= 2082951896;
assign addr[4606]= 2114858546;
assign addr[4607]= 2136037160;
assign addr[4608]= 2146380306;
assign addr[4609]= 2145835515;
assign addr[4610]= 2134405552;
assign addr[4611]= 2112148396;
assign addr[4612]= 2079176953;
assign addr[4613]= 2035658475;
assign addr[4614]= 1981813720;
assign addr[4615]= 1917915825;
assign addr[4616]= 1844288924;
assign addr[4617]= 1761306505;
assign addr[4618]= 1669389513;
assign addr[4619]= 1569004214;
assign addr[4620]= 1460659832;
assign addr[4621]= 1344905966;
assign addr[4622]= 1222329801;
assign addr[4623]= 1093553126;
assign addr[4624]= 959229189;
assign addr[4625]= 820039373;
assign addr[4626]= 676689746;
assign addr[4627]= 529907477;
assign addr[4628]= 380437148;
assign addr[4629]= 229036977;
assign addr[4630]= 76474970;
assign addr[4631]= -76474970;
assign addr[4632]= -229036977;
assign addr[4633]= -380437148;
assign addr[4634]= -529907477;
assign addr[4635]= -676689746;
assign addr[4636]= -820039373;
assign addr[4637]= -959229189;
assign addr[4638]= -1093553126;
assign addr[4639]= -1222329801;
assign addr[4640]= -1344905966;
assign addr[4641]= -1460659832;
assign addr[4642]= -1569004214;
assign addr[4643]= -1669389513;
assign addr[4644]= -1761306505;
assign addr[4645]= -1844288924;
assign addr[4646]= -1917915825;
assign addr[4647]= -1981813720;
assign addr[4648]= -2035658475;
assign addr[4649]= -2079176953;
assign addr[4650]= -2112148396;
assign addr[4651]= -2134405552;
assign addr[4652]= -2145835515;
assign addr[4653]= -2146380306;
assign addr[4654]= -2136037160;
assign addr[4655]= -2114858546;
assign addr[4656]= -2082951896;
assign addr[4657]= -2040479063;
assign addr[4658]= -1987655498;
assign addr[4659]= -1924749160;
assign addr[4660]= -1852079154;
assign addr[4661]= -1770014111;
assign addr[4662]= -1678970324;
assign addr[4663]= -1579409630;
assign addr[4664]= -1471837070;
assign addr[4665]= -1356798326;
assign addr[4666]= -1234876957;
assign addr[4667]= -1106691431;
assign addr[4668]= -972891995;
assign addr[4669]= -834157373;
assign addr[4670]= -691191324;
assign addr[4671]= -544719071;
assign addr[4672]= -395483624;
assign addr[4673]= -244242007;
assign addr[4674]= -91761426;
assign addr[4675]= 61184634;
assign addr[4676]= 213820322;
assign addr[4677]= 365371365;
assign addr[4678]= 515068990;
assign addr[4679]= 662153826;
assign addr[4680]= 805879757;
assign addr[4681]= 945517704;
assign addr[4682]= 1080359326;
assign addr[4683]= 1209720613;
assign addr[4684]= 1332945355;
assign addr[4685]= 1449408469;
assign addr[4686]= 1558519173;
assign addr[4687]= 1659723983;
assign addr[4688]= 1752509516;
assign addr[4689]= 1836405100;
assign addr[4690]= 1910985158;
assign addr[4691]= 1975871368;
assign addr[4692]= 2030734582;
assign addr[4693]= 2075296495;
assign addr[4694]= 2109331059;
assign addr[4695]= 2132665626;
assign addr[4696]= 2145181827;
assign addr[4697]= 2146816171;
assign addr[4698]= 2137560369;
assign addr[4699]= 2117461370;
assign addr[4700]= 2086621133;
assign addr[4701]= 2045196100;
assign addr[4702]= 1993396407;
assign addr[4703]= 1931484818;
assign addr[4704]= 1859775393;
assign addr[4705]= 1778631892;
assign addr[4706]= 1688465931;
assign addr[4707]= 1589734894;
assign addr[4708]= 1482939614;
assign addr[4709]= 1368621831;
assign addr[4710]= 1247361445;
assign addr[4711]= 1119773573;
assign addr[4712]= 986505429;
assign addr[4713]= 848233042;
assign addr[4714]= 705657826;
assign addr[4715]= 559503022;
assign addr[4716]= 410510029;
assign addr[4717]= 259434643;
assign addr[4718]= 107043224;
assign addr[4719]= -45891193;
assign addr[4720]= -198592817;
assign addr[4721]= -350287041;
assign addr[4722]= -500204365;
assign addr[4723]= -647584304;
assign addr[4724]= -791679244;
assign addr[4725]= -931758235;
assign addr[4726]= -1067110699;
assign addr[4727]= -1197050035;
assign addr[4728]= -1320917099;
assign addr[4729]= -1438083551;
assign addr[4730]= -1547955041;
assign addr[4731]= -1649974225;
assign addr[4732]= -1743623590;
assign addr[4733]= -1828428082;
assign addr[4734]= -1903957513;
assign addr[4735]= -1969828744;
assign addr[4736]= -2025707632;
assign addr[4737]= -2071310720;
assign addr[4738]= -2106406677;
assign addr[4739]= -2130817471;
assign addr[4740]= -2144419275;
assign addr[4741]= -2147143090;
assign addr[4742]= -2138975100;
assign addr[4743]= -2119956737;
assign addr[4744]= -2090184478;
assign addr[4745]= -2049809346;
assign addr[4746]= -1999036154;
assign addr[4747]= -1938122457;
assign addr[4748]= -1867377253;
assign addr[4749]= -1787159411;
assign addr[4750]= -1697875851;
assign addr[4751]= -1599979481;
assign addr[4752]= -1493966902;
assign addr[4753]= -1380375881;
assign addr[4754]= -1259782632;
assign addr[4755]= -1132798888;
assign addr[4756]= -1000068799;
assign addr[4757]= -862265664;
assign addr[4758]= -720088517;
assign addr[4759]= -574258580;
assign addr[4760]= -425515602;
assign addr[4761]= -274614114;
assign addr[4762]= -122319591;
assign addr[4763]= 30595422;
assign addr[4764]= 183355234;
assign addr[4765]= 335184940;
assign addr[4766]= 485314355;
assign addr[4767]= 632981917;
assign addr[4768]= 777438554;
assign addr[4769]= 917951481;
assign addr[4770]= 1053807919;
assign addr[4771]= 1184318708;
assign addr[4772]= 1308821808;
assign addr[4773]= 1426685652;
assign addr[4774]= 1537312353;
assign addr[4775]= 1640140734;
assign addr[4776]= 1734649179;
assign addr[4777]= 1820358275;
assign addr[4778]= 1896833245;
assign addr[4779]= 1963686155;
assign addr[4780]= 2020577882;
assign addr[4781]= 2067219829;
assign addr[4782]= 2103375398;
assign addr[4783]= 2128861181;
assign addr[4784]= 2143547897;
assign addr[4785]= 2147361045;
assign addr[4786]= 2140281282;
assign addr[4787]= 2122344521;
assign addr[4788]= 2093641749;
assign addr[4789]= 2054318569;
assign addr[4790]= 2004574453;
assign addr[4791]= 1944661739;
assign addr[4792]= 1874884346;
assign addr[4793]= 1795596234;
assign addr[4794]= 1707199606;
assign addr[4795]= 1610142873;
assign addr[4796]= 1504918373;
assign addr[4797]= 1392059879;
assign addr[4798]= 1272139887;
assign addr[4799]= 1145766716;
assign addr[4800]= 1013581418;
assign addr[4801]= 876254528;
assign addr[4802]= 734482665;
assign addr[4803]= 588984994;
assign addr[4804]= 440499581;
assign addr[4805]= 289779648;
assign addr[4806]= 137589750;
assign addr[4807]= -15298099;
assign addr[4808]= -168108346;
assign addr[4809]= -320065829;
assign addr[4810]= -470399716;
assign addr[4811]= -618347408;
assign addr[4812]= -763158411;
assign addr[4813]= -904098143;
assign addr[4814]= -1040451659;
assign addr[4815]= -1171527280;
assign addr[4816]= -1296660098;
assign addr[4817]= -1415215352;
assign addr[4818]= -1526591649;
assign addr[4819]= -1630224009;
assign addr[4820]= -1725586737;
assign addr[4821]= -1812196087;
assign addr[4822]= -1889612716;
assign addr[4823]= -1957443913;
assign addr[4824]= -2015345591;
assign addr[4825]= -2063024031;
assign addr[4826]= -2100237377;
assign addr[4827]= -2126796855;
assign addr[4828]= -2142567738;
assign addr[4829]= -2147470025;
assign addr[4830]= -2141478848;
assign addr[4831]= -2124624598;
assign addr[4832]= -2096992772;
assign addr[4833]= -2058723538;
assign addr[4834]= -2010011024;
assign addr[4835]= -1951102334;
assign addr[4836]= -1882296293;
assign addr[4837]= -1803941934;
assign addr[4838]= -1716436725;
assign addr[4839]= -1620224553;
assign addr[4840]= -1515793473;
assign addr[4841]= -1403673233;
assign addr[4842]= -1284432584;
assign addr[4843]= -1158676398;
assign addr[4844]= -1027042599;
assign addr[4845]= -890198924;
assign addr[4846]= -748839539;
assign addr[4847]= -603681519;
assign addr[4848]= -455461206;
assign addr[4849]= -304930476;
assign addr[4850]= -152852926;
assign addr[4851]= 0;
assign addr[4852]= 152852926;
assign addr[4853]= 304930476;
assign addr[4854]= 455461206;
assign addr[4855]= 603681519;
assign addr[4856]= 748839539;
assign addr[4857]= 890198924;
assign addr[4858]= 1027042599;
assign addr[4859]= 1158676398;
assign addr[4860]= 1284432584;
assign addr[4861]= 1403673233;
assign addr[4862]= 1515793473;
assign addr[4863]= 1620224553;
assign addr[4864]= 1716436725;
assign addr[4865]= 1803941934;
assign addr[4866]= 1882296293;
assign addr[4867]= 1951102334;
assign addr[4868]= 2010011024;
assign addr[4869]= 2058723538;
assign addr[4870]= 2096992772;
assign addr[4871]= 2124624598;
assign addr[4872]= 2141478848;
assign addr[4873]= 2147470025;
assign addr[4874]= 2142567738;
assign addr[4875]= 2126796855;
assign addr[4876]= 2100237377;
assign addr[4877]= 2063024031;
assign addr[4878]= 2015345591;
assign addr[4879]= 1957443913;
assign addr[4880]= 1889612716;
assign addr[4881]= 1812196087;
assign addr[4882]= 1725586737;
assign addr[4883]= 1630224009;
assign addr[4884]= 1526591649;
assign addr[4885]= 1415215352;
assign addr[4886]= 1296660098;
assign addr[4887]= 1171527280;
assign addr[4888]= 1040451659;
assign addr[4889]= 904098143;
assign addr[4890]= 763158411;
assign addr[4891]= 618347408;
assign addr[4892]= 470399716;
assign addr[4893]= 320065829;
assign addr[4894]= 168108346;
assign addr[4895]= 15298099;
assign addr[4896]= -137589750;
assign addr[4897]= -289779648;
assign addr[4898]= -440499581;
assign addr[4899]= -588984994;
assign addr[4900]= -734482665;
assign addr[4901]= -876254528;
assign addr[4902]= -1013581418;
assign addr[4903]= -1145766716;
assign addr[4904]= -1272139887;
assign addr[4905]= -1392059879;
assign addr[4906]= -1504918373;
assign addr[4907]= -1610142873;
assign addr[4908]= -1707199606;
assign addr[4909]= -1795596234;
assign addr[4910]= -1874884346;
assign addr[4911]= -1944661739;
assign addr[4912]= -2004574453;
assign addr[4913]= -2054318569;
assign addr[4914]= -2093641749;
assign addr[4915]= -2122344521;
assign addr[4916]= -2140281282;
assign addr[4917]= -2147361045;
assign addr[4918]= -2143547897;
assign addr[4919]= -2128861181;
assign addr[4920]= -2103375398;
assign addr[4921]= -2067219829;
assign addr[4922]= -2020577882;
assign addr[4923]= -1963686155;
assign addr[4924]= -1896833245;
assign addr[4925]= -1820358275;
assign addr[4926]= -1734649179;
assign addr[4927]= -1640140734;
assign addr[4928]= -1537312353;
assign addr[4929]= -1426685652;
assign addr[4930]= -1308821808;
assign addr[4931]= -1184318708;
assign addr[4932]= -1053807919;
assign addr[4933]= -917951481;
assign addr[4934]= -777438554;
assign addr[4935]= -632981917;
assign addr[4936]= -485314355;
assign addr[4937]= -335184940;
assign addr[4938]= -183355234;
assign addr[4939]= -30595422;
assign addr[4940]= 122319591;
assign addr[4941]= 274614114;
assign addr[4942]= 425515602;
assign addr[4943]= 574258580;
assign addr[4944]= 720088517;
assign addr[4945]= 862265664;
assign addr[4946]= 1000068799;
assign addr[4947]= 1132798888;
assign addr[4948]= 1259782632;
assign addr[4949]= 1380375881;
assign addr[4950]= 1493966902;
assign addr[4951]= 1599979481;
assign addr[4952]= 1697875851;
assign addr[4953]= 1787159411;
assign addr[4954]= 1867377253;
assign addr[4955]= 1938122457;
assign addr[4956]= 1999036154;
assign addr[4957]= 2049809346;
assign addr[4958]= 2090184478;
assign addr[4959]= 2119956737;
assign addr[4960]= 2138975100;
assign addr[4961]= 2147143090;
assign addr[4962]= 2144419275;
assign addr[4963]= 2130817471;
assign addr[4964]= 2106406677;
assign addr[4965]= 2071310720;
assign addr[4966]= 2025707632;
assign addr[4967]= 1969828744;
assign addr[4968]= 1903957513;
assign addr[4969]= 1828428082;
assign addr[4970]= 1743623590;
assign addr[4971]= 1649974225;
assign addr[4972]= 1547955041;
assign addr[4973]= 1438083551;
assign addr[4974]= 1320917099;
assign addr[4975]= 1197050035;
assign addr[4976]= 1067110699;
assign addr[4977]= 931758235;
assign addr[4978]= 791679244;
assign addr[4979]= 647584304;
assign addr[4980]= 500204365;
assign addr[4981]= 350287041;
assign addr[4982]= 198592817;
assign addr[4983]= 45891193;
assign addr[4984]= -107043224;
assign addr[4985]= -259434643;
assign addr[4986]= -410510029;
assign addr[4987]= -559503022;
assign addr[4988]= -705657826;
assign addr[4989]= -848233042;
assign addr[4990]= -986505429;
assign addr[4991]= -1119773573;
assign addr[4992]= -1247361445;
assign addr[4993]= -1368621831;
assign addr[4994]= -1482939614;
assign addr[4995]= -1589734894;
assign addr[4996]= -1688465931;
assign addr[4997]= -1778631892;
assign addr[4998]= -1859775393;
assign addr[4999]= -1931484818;
assign addr[5000]= -1993396407;
assign addr[5001]= -2045196100;
assign addr[5002]= -2086621133;
assign addr[5003]= -2117461370;
assign addr[5004]= -2137560369;
assign addr[5005]= -2146816171;
assign addr[5006]= -2145181827;
assign addr[5007]= -2132665626;
assign addr[5008]= -2109331059;
assign addr[5009]= -2075296495;
assign addr[5010]= -2030734582;
assign addr[5011]= -1975871368;
assign addr[5012]= -1910985158;
assign addr[5013]= -1836405100;
assign addr[5014]= -1752509516;
assign addr[5015]= -1659723983;
assign addr[5016]= -1558519173;
assign addr[5017]= -1449408469;
assign addr[5018]= -1332945355;
assign addr[5019]= -1209720613;
assign addr[5020]= -1080359326;
assign addr[5021]= -945517704;
assign addr[5022]= -805879757;
assign addr[5023]= -662153826;
assign addr[5024]= -515068990;
assign addr[5025]= -365371365;
assign addr[5026]= -213820322;
assign addr[5027]= -61184634;
assign addr[5028]= 91761426;
assign addr[5029]= 244242007;
assign addr[5030]= 395483624;
assign addr[5031]= 544719071;
assign addr[5032]= 691191324;
assign addr[5033]= 834157373;
assign addr[5034]= 972891995;
assign addr[5035]= 1106691431;
assign addr[5036]= 1234876957;
assign addr[5037]= 1356798326;
assign addr[5038]= 1471837070;
assign addr[5039]= 1579409630;
assign addr[5040]= 1678970324;
assign addr[5041]= 1770014111;
assign addr[5042]= 1852079154;
assign addr[5043]= 1924749160;
assign addr[5044]= 1987655498;
assign addr[5045]= 2040479063;
assign addr[5046]= 2082951896;
assign addr[5047]= 2114858546;
assign addr[5048]= 2136037160;
assign addr[5049]= 2146380306;
assign addr[5050]= 2145835515;
assign addr[5051]= 2134405552;
assign addr[5052]= 2112148396;
assign addr[5053]= 2079176953;
assign addr[5054]= 2035658475;
assign addr[5055]= 1981813720;
assign addr[5056]= 1917915825;
assign addr[5057]= 1844288924;
assign addr[5058]= 1761306505;
assign addr[5059]= 1669389513;
assign addr[5060]= 1569004214;
assign addr[5061]= 1460659832;
assign addr[5062]= 1344905966;
assign addr[5063]= 1222329801;
assign addr[5064]= 1093553126;
assign addr[5065]= 959229189;
assign addr[5066]= 820039373;
assign addr[5067]= 676689746;
assign addr[5068]= 529907477;
assign addr[5069]= 380437148;
assign addr[5070]= 229036977;
assign addr[5071]= 76474970;
assign addr[5072]= -76474970;
assign addr[5073]= -229036977;
assign addr[5074]= -380437148;
assign addr[5075]= -529907477;
assign addr[5076]= -676689746;
assign addr[5077]= -820039373;
assign addr[5078]= -959229189;
assign addr[5079]= -1093553126;
assign addr[5080]= -1222329801;
assign addr[5081]= -1344905966;
assign addr[5082]= -1460659832;
assign addr[5083]= -1569004214;
assign addr[5084]= -1669389513;
assign addr[5085]= -1761306505;
assign addr[5086]= -1844288924;
assign addr[5087]= -1917915825;
assign addr[5088]= -1981813720;
assign addr[5089]= -2035658475;
assign addr[5090]= -2079176953;
assign addr[5091]= -2112148396;
assign addr[5092]= -2134405552;
assign addr[5093]= -2145835515;
assign addr[5094]= -2146380306;
assign addr[5095]= -2136037160;
assign addr[5096]= -2114858546;
assign addr[5097]= -2082951896;
assign addr[5098]= -2040479063;
assign addr[5099]= -1987655498;
assign addr[5100]= -1924749160;
assign addr[5101]= -1852079154;
assign addr[5102]= -1770014111;
assign addr[5103]= -1678970324;
assign addr[5104]= -1579409630;
assign addr[5105]= -1471837070;
assign addr[5106]= -1356798326;
assign addr[5107]= -1234876957;
assign addr[5108]= -1106691431;
assign addr[5109]= -972891995;
assign addr[5110]= -834157373;
assign addr[5111]= -691191324;
assign addr[5112]= -544719071;
assign addr[5113]= -395483624;
assign addr[5114]= -244242007;
assign addr[5115]= -91761426;
assign addr[5116]= 61184634;
assign addr[5117]= 213820322;
assign addr[5118]= 365371365;
assign addr[5119]= 515068990;
assign addr[5120]= 662153826;
assign addr[5121]= 805879757;
assign addr[5122]= 945517704;
assign addr[5123]= 1080359326;
assign addr[5124]= 1209720613;
assign addr[5125]= 1332945355;
assign addr[5126]= 1449408469;
assign addr[5127]= 1558519173;
assign addr[5128]= 1659723983;
assign addr[5129]= 1752509516;
assign addr[5130]= 1836405100;
assign addr[5131]= 1910985158;
assign addr[5132]= 1975871368;
assign addr[5133]= 2030734582;
assign addr[5134]= 2075296495;
assign addr[5135]= 2109331059;
assign addr[5136]= 2132665626;
assign addr[5137]= 2145181827;
assign addr[5138]= 2146816171;
assign addr[5139]= 2137560369;
assign addr[5140]= 2117461370;
assign addr[5141]= 2086621133;
assign addr[5142]= 2045196100;
assign addr[5143]= 1993396407;
assign addr[5144]= 1931484818;
assign addr[5145]= 1859775393;
assign addr[5146]= 1778631892;
assign addr[5147]= 1688465931;
assign addr[5148]= 1589734894;
assign addr[5149]= 1482939614;
assign addr[5150]= 1368621831;
assign addr[5151]= 1247361445;
assign addr[5152]= 1119773573;
assign addr[5153]= 986505429;
assign addr[5154]= 848233042;
assign addr[5155]= 705657826;
assign addr[5156]= 559503022;
assign addr[5157]= 410510029;
assign addr[5158]= 259434643;
assign addr[5159]= 107043224;
assign addr[5160]= -45891193;
assign addr[5161]= -198592817;
assign addr[5162]= -350287041;
assign addr[5163]= -500204365;
assign addr[5164]= -647584304;
assign addr[5165]= -791679244;
assign addr[5166]= -931758235;
assign addr[5167]= -1067110699;
assign addr[5168]= -1197050035;
assign addr[5169]= -1320917099;
assign addr[5170]= -1438083551;
assign addr[5171]= -1547955041;
assign addr[5172]= -1649974225;
assign addr[5173]= -1743623590;
assign addr[5174]= -1828428082;
assign addr[5175]= -1903957513;
assign addr[5176]= -1969828744;
assign addr[5177]= -2025707632;
assign addr[5178]= -2071310720;
assign addr[5179]= -2106406677;
assign addr[5180]= -2130817471;
assign addr[5181]= -2144419275;
assign addr[5182]= -2147143090;
assign addr[5183]= -2138975100;
assign addr[5184]= -2119956737;
assign addr[5185]= -2090184478;
assign addr[5186]= -2049809346;
assign addr[5187]= -1999036154;
assign addr[5188]= -1938122457;
assign addr[5189]= -1867377253;
assign addr[5190]= -1787159411;
assign addr[5191]= -1697875851;
assign addr[5192]= -1599979481;
assign addr[5193]= -1493966902;
assign addr[5194]= -1380375881;
assign addr[5195]= -1259782632;
assign addr[5196]= -1132798888;
assign addr[5197]= -1000068799;
assign addr[5198]= -862265664;
assign addr[5199]= -720088517;
assign addr[5200]= -574258580;
assign addr[5201]= -425515602;
assign addr[5202]= -274614114;
assign addr[5203]= -122319591;
assign addr[5204]= 30595422;
assign addr[5205]= 183355234;
assign addr[5206]= 335184940;
assign addr[5207]= 485314355;
assign addr[5208]= 632981917;
assign addr[5209]= 777438554;
assign addr[5210]= 917951481;
assign addr[5211]= 1053807919;
assign addr[5212]= 1184318708;
assign addr[5213]= 1308821808;
assign addr[5214]= 1426685652;
assign addr[5215]= 1537312353;
assign addr[5216]= 1640140734;
assign addr[5217]= 1734649179;
assign addr[5218]= 1820358275;
assign addr[5219]= 1896833245;
assign addr[5220]= 1963686155;
assign addr[5221]= 2020577882;
assign addr[5222]= 2067219829;
assign addr[5223]= 2103375398;
assign addr[5224]= 2128861181;
assign addr[5225]= 2143547897;
assign addr[5226]= 2147361045;
assign addr[5227]= 2140281282;
assign addr[5228]= 2122344521;
assign addr[5229]= 2093641749;
assign addr[5230]= 2054318569;
assign addr[5231]= 2004574453;
assign addr[5232]= 1944661739;
assign addr[5233]= 1874884346;
assign addr[5234]= 1795596234;
assign addr[5235]= 1707199606;
assign addr[5236]= 1610142873;
assign addr[5237]= 1504918373;
assign addr[5238]= 1392059879;
assign addr[5239]= 1272139887;
assign addr[5240]= 1145766716;
assign addr[5241]= 1013581418;
assign addr[5242]= 876254528;
assign addr[5243]= 734482665;
assign addr[5244]= 588984994;
assign addr[5245]= 440499581;
assign addr[5246]= 289779648;
assign addr[5247]= 137589750;
assign addr[5248]= -15298099;
assign addr[5249]= -168108346;
assign addr[5250]= -320065829;
assign addr[5251]= -470399716;
assign addr[5252]= -618347408;
assign addr[5253]= -763158411;
assign addr[5254]= -904098143;
assign addr[5255]= -1040451659;
assign addr[5256]= -1171527280;
assign addr[5257]= -1296660098;
assign addr[5258]= -1415215352;
assign addr[5259]= -1526591649;
assign addr[5260]= -1630224009;
assign addr[5261]= -1725586737;
assign addr[5262]= -1812196087;
assign addr[5263]= -1889612716;
assign addr[5264]= -1957443913;
assign addr[5265]= -2015345591;
assign addr[5266]= -2063024031;
assign addr[5267]= -2100237377;
assign addr[5268]= -2126796855;
assign addr[5269]= -2142567738;
assign addr[5270]= -2147470025;
assign addr[5271]= -2141478848;
assign addr[5272]= -2124624598;
assign addr[5273]= -2096992772;
assign addr[5274]= -2058723538;
assign addr[5275]= -2010011024;
assign addr[5276]= -1951102334;
assign addr[5277]= -1882296293;
assign addr[5278]= -1803941934;
assign addr[5279]= -1716436725;
assign addr[5280]= -1620224553;
assign addr[5281]= -1515793473;
assign addr[5282]= -1403673233;
assign addr[5283]= -1284432584;
assign addr[5284]= -1158676398;
assign addr[5285]= -1027042599;
assign addr[5286]= -890198924;
assign addr[5287]= -748839539;
assign addr[5288]= -603681519;
assign addr[5289]= -455461206;
assign addr[5290]= -304930476;
assign addr[5291]= -152852926;
assign addr[5292]= 0;
assign addr[5293]= 152852926;
assign addr[5294]= 304930476;
assign addr[5295]= 455461206;
assign addr[5296]= 603681519;
assign addr[5297]= 748839539;
assign addr[5298]= 890198924;
assign addr[5299]= 1027042599;
assign addr[5300]= 1158676398;
assign addr[5301]= 1284432584;
assign addr[5302]= 1403673233;
assign addr[5303]= 1515793473;
assign addr[5304]= 1620224553;
assign addr[5305]= 1716436725;
assign addr[5306]= 1803941934;
assign addr[5307]= 1882296293;
assign addr[5308]= 1951102334;
assign addr[5309]= 2010011024;
assign addr[5310]= 2058723538;
assign addr[5311]= 2096992772;
assign addr[5312]= 2124624598;
assign addr[5313]= 2141478848;
assign addr[5314]= 2147470025;
assign addr[5315]= 2142567738;
assign addr[5316]= 2126796855;
assign addr[5317]= 2100237377;
assign addr[5318]= 2063024031;
assign addr[5319]= 2015345591;
assign addr[5320]= 1957443913;
assign addr[5321]= 1889612716;
assign addr[5322]= 1812196087;
assign addr[5323]= 1725586737;
assign addr[5324]= 1630224009;
assign addr[5325]= 1526591649;
assign addr[5326]= 1415215352;
assign addr[5327]= 1296660098;
assign addr[5328]= 1171527280;
assign addr[5329]= 1040451659;
assign addr[5330]= 904098143;
assign addr[5331]= 763158411;
assign addr[5332]= 618347408;
assign addr[5333]= 470399716;
assign addr[5334]= 320065829;
assign addr[5335]= 168108346;
assign addr[5336]= 15298099;
assign addr[5337]= -137589750;
assign addr[5338]= -289779648;
assign addr[5339]= -440499581;
assign addr[5340]= -588984994;
assign addr[5341]= -734482665;
assign addr[5342]= -876254528;
assign addr[5343]= -1013581418;
assign addr[5344]= -1145766716;
assign addr[5345]= -1272139887;
assign addr[5346]= -1392059879;
assign addr[5347]= -1504918373;
assign addr[5348]= -1610142873;
assign addr[5349]= -1707199606;
assign addr[5350]= -1795596234;
assign addr[5351]= -1874884346;
assign addr[5352]= -1944661739;
assign addr[5353]= -2004574453;
assign addr[5354]= -2054318569;
assign addr[5355]= -2093641749;
assign addr[5356]= -2122344521;
assign addr[5357]= -2140281282;
assign addr[5358]= -2147361045;
assign addr[5359]= -2143547897;
assign addr[5360]= -2128861181;
assign addr[5361]= -2103375398;
assign addr[5362]= -2067219829;
assign addr[5363]= -2020577882;
assign addr[5364]= -1963686155;
assign addr[5365]= -1896833245;
assign addr[5366]= -1820358275;
assign addr[5367]= -1734649179;
assign addr[5368]= -1640140734;
assign addr[5369]= -1537312353;
assign addr[5370]= -1426685652;
assign addr[5371]= -1308821808;
assign addr[5372]= -1184318708;
assign addr[5373]= -1053807919;
assign addr[5374]= -917951481;
assign addr[5375]= -777438554;
assign addr[5376]= -632981917;
assign addr[5377]= -485314355;
assign addr[5378]= -335184940;
assign addr[5379]= -183355234;
assign addr[5380]= -30595422;
assign addr[5381]= 122319591;
assign addr[5382]= 274614114;
assign addr[5383]= 425515602;
assign addr[5384]= 574258580;
assign addr[5385]= 720088517;
assign addr[5386]= 862265664;
assign addr[5387]= 1000068799;
assign addr[5388]= 1132798888;
assign addr[5389]= 1259782632;
assign addr[5390]= 1380375881;
assign addr[5391]= 1493966902;
assign addr[5392]= 1599979481;
assign addr[5393]= 1697875851;
assign addr[5394]= 1787159411;
assign addr[5395]= 1867377253;
assign addr[5396]= 1938122457;
assign addr[5397]= 1999036154;
assign addr[5398]= 2049809346;
assign addr[5399]= 2090184478;
assign addr[5400]= 2119956737;
assign addr[5401]= 2138975100;
assign addr[5402]= 2147143090;
assign addr[5403]= 2144419275;
assign addr[5404]= 2130817471;
assign addr[5405]= 2106406677;
assign addr[5406]= 2071310720;
assign addr[5407]= 2025707632;
assign addr[5408]= 1969828744;
assign addr[5409]= 1903957513;
assign addr[5410]= 1828428082;
assign addr[5411]= 1743623590;
assign addr[5412]= 1649974225;
assign addr[5413]= 1547955041;
assign addr[5414]= 1438083551;
assign addr[5415]= 1320917099;
assign addr[5416]= 1197050035;
assign addr[5417]= 1067110699;
assign addr[5418]= 931758235;
assign addr[5419]= 791679244;
assign addr[5420]= 647584304;
assign addr[5421]= 500204365;
assign addr[5422]= 350287041;
assign addr[5423]= 198592817;
assign addr[5424]= 45891193;
assign addr[5425]= -107043224;
assign addr[5426]= -259434643;
assign addr[5427]= -410510029;
assign addr[5428]= -559503022;
assign addr[5429]= -705657826;
assign addr[5430]= -848233042;
assign addr[5431]= -986505429;
assign addr[5432]= -1119773573;
assign addr[5433]= -1247361445;
assign addr[5434]= -1368621831;
assign addr[5435]= -1482939614;
assign addr[5436]= -1589734894;
assign addr[5437]= -1688465931;
assign addr[5438]= -1778631892;
assign addr[5439]= -1859775393;
assign addr[5440]= -1931484818;
assign addr[5441]= -1993396407;
assign addr[5442]= -2045196100;
assign addr[5443]= -2086621133;
assign addr[5444]= -2117461370;
assign addr[5445]= -2137560369;
assign addr[5446]= -2146816171;
assign addr[5447]= -2145181827;
assign addr[5448]= -2132665626;
assign addr[5449]= -2109331059;
assign addr[5450]= -2075296495;
assign addr[5451]= -2030734582;
assign addr[5452]= -1975871368;
assign addr[5453]= -1910985158;
assign addr[5454]= -1836405100;
assign addr[5455]= -1752509516;
assign addr[5456]= -1659723983;
assign addr[5457]= -1558519173;
assign addr[5458]= -1449408469;
assign addr[5459]= -1332945355;
assign addr[5460]= -1209720613;
assign addr[5461]= -1080359326;
assign addr[5462]= -945517704;
assign addr[5463]= -805879757;
assign addr[5464]= -662153826;
assign addr[5465]= -515068990;
assign addr[5466]= -365371365;
assign addr[5467]= -213820322;
assign addr[5468]= -61184634;
assign addr[5469]= 91761426;
assign addr[5470]= 244242007;
assign addr[5471]= 395483624;
assign addr[5472]= 544719071;
assign addr[5473]= 691191324;
assign addr[5474]= 834157373;
assign addr[5475]= 972891995;
assign addr[5476]= 1106691431;
assign addr[5477]= 1234876957;
assign addr[5478]= 1356798326;
assign addr[5479]= 1471837070;
assign addr[5480]= 1579409630;
assign addr[5481]= 1678970324;
assign addr[5482]= 1770014111;
assign addr[5483]= 1852079154;
assign addr[5484]= 1924749160;
assign addr[5485]= 1987655498;
assign addr[5486]= 2040479063;
assign addr[5487]= 2082951896;
assign addr[5488]= 2114858546;
assign addr[5489]= 2136037160;
assign addr[5490]= 2146380306;
assign addr[5491]= 2145835515;
assign addr[5492]= 2134405552;
assign addr[5493]= 2112148396;
assign addr[5494]= 2079176953;
assign addr[5495]= 2035658475;
assign addr[5496]= 1981813720;
assign addr[5497]= 1917915825;
assign addr[5498]= 1844288924;
assign addr[5499]= 1761306505;
assign addr[5500]= 1669389513;
assign addr[5501]= 1569004214;
assign addr[5502]= 1460659832;
assign addr[5503]= 1344905966;
assign addr[5504]= 1222329801;
assign addr[5505]= 1093553126;
assign addr[5506]= 959229189;
assign addr[5507]= 820039373;
assign addr[5508]= 676689746;
assign addr[5509]= 529907477;
assign addr[5510]= 380437148;
assign addr[5511]= 229036977;
assign addr[5512]= 76474970;
assign addr[5513]= -76474970;
assign addr[5514]= -229036977;
assign addr[5515]= -380437148;
assign addr[5516]= -529907477;
assign addr[5517]= -676689746;
assign addr[5518]= -820039373;
assign addr[5519]= -959229189;
assign addr[5520]= -1093553126;
assign addr[5521]= -1222329801;
assign addr[5522]= -1344905966;
assign addr[5523]= -1460659832;
assign addr[5524]= -1569004214;
assign addr[5525]= -1669389513;
assign addr[5526]= -1761306505;
assign addr[5527]= -1844288924;
assign addr[5528]= -1917915825;
assign addr[5529]= -1981813720;
assign addr[5530]= -2035658475;
assign addr[5531]= -2079176953;
assign addr[5532]= -2112148396;
assign addr[5533]= -2134405552;
assign addr[5534]= -2145835515;
assign addr[5535]= -2146380306;
assign addr[5536]= -2136037160;
assign addr[5537]= -2114858546;
assign addr[5538]= -2082951896;
assign addr[5539]= -2040479063;
assign addr[5540]= -1987655498;
assign addr[5541]= -1924749160;
assign addr[5542]= -1852079154;
assign addr[5543]= -1770014111;
assign addr[5544]= -1678970324;
assign addr[5545]= -1579409630;
assign addr[5546]= -1471837070;
assign addr[5547]= -1356798326;
assign addr[5548]= -1234876957;
assign addr[5549]= -1106691431;
assign addr[5550]= -972891995;
assign addr[5551]= -834157373;
assign addr[5552]= -691191324;
assign addr[5553]= -544719071;
assign addr[5554]= -395483624;
assign addr[5555]= -244242007;
assign addr[5556]= -91761426;
assign addr[5557]= 61184634;
assign addr[5558]= 213820322;
assign addr[5559]= 365371365;
assign addr[5560]= 515068990;
assign addr[5561]= 662153826;
assign addr[5562]= 805879757;
assign addr[5563]= 945517704;
assign addr[5564]= 1080359326;
assign addr[5565]= 1209720613;
assign addr[5566]= 1332945355;
assign addr[5567]= 1449408469;
assign addr[5568]= 1558519173;
assign addr[5569]= 1659723983;
assign addr[5570]= 1752509516;
assign addr[5571]= 1836405100;
assign addr[5572]= 1910985158;
assign addr[5573]= 1975871368;
assign addr[5574]= 2030734582;
assign addr[5575]= 2075296495;
assign addr[5576]= 2109331059;
assign addr[5577]= 2132665626;
assign addr[5578]= 2145181827;
assign addr[5579]= 2146816171;
assign addr[5580]= 2137560369;
assign addr[5581]= 2117461370;
assign addr[5582]= 2086621133;
assign addr[5583]= 2045196100;
assign addr[5584]= 1993396407;
assign addr[5585]= 1931484818;
assign addr[5586]= 1859775393;
assign addr[5587]= 1778631892;
assign addr[5588]= 1688465931;
assign addr[5589]= 1589734894;
assign addr[5590]= 1482939614;
assign addr[5591]= 1368621831;
assign addr[5592]= 1247361445;
assign addr[5593]= 1119773573;
assign addr[5594]= 986505429;
assign addr[5595]= 848233042;
assign addr[5596]= 705657826;
assign addr[5597]= 559503022;
assign addr[5598]= 410510029;
assign addr[5599]= 259434643;
assign addr[5600]= 107043224;
assign addr[5601]= -45891193;
assign addr[5602]= -198592817;
assign addr[5603]= -350287041;
assign addr[5604]= -500204365;
assign addr[5605]= -647584304;
assign addr[5606]= -791679244;
assign addr[5607]= -931758235;
assign addr[5608]= -1067110699;
assign addr[5609]= -1197050035;
assign addr[5610]= -1320917099;
assign addr[5611]= -1438083551;
assign addr[5612]= -1547955041;
assign addr[5613]= -1649974225;
assign addr[5614]= -1743623590;
assign addr[5615]= -1828428082;
assign addr[5616]= -1903957513;
assign addr[5617]= -1969828744;
assign addr[5618]= -2025707632;
assign addr[5619]= -2071310720;
assign addr[5620]= -2106406677;
assign addr[5621]= -2130817471;
assign addr[5622]= -2144419275;
assign addr[5623]= -2147143090;
assign addr[5624]= -2138975100;
assign addr[5625]= -2119956737;
assign addr[5626]= -2090184478;
assign addr[5627]= -2049809346;
assign addr[5628]= -1999036154;
assign addr[5629]= -1938122457;
assign addr[5630]= -1867377253;
assign addr[5631]= -1787159411;
assign addr[5632]= -1697875851;
assign addr[5633]= -1599979481;
assign addr[5634]= -1493966902;
assign addr[5635]= -1380375881;
assign addr[5636]= -1259782632;
assign addr[5637]= -1132798888;
assign addr[5638]= -1000068799;
assign addr[5639]= -862265664;
assign addr[5640]= -720088517;
assign addr[5641]= -574258580;
assign addr[5642]= -425515602;
assign addr[5643]= -274614114;
assign addr[5644]= -122319591;
assign addr[5645]= 30595422;
assign addr[5646]= 183355234;
assign addr[5647]= 335184940;
assign addr[5648]= 485314355;
assign addr[5649]= 632981917;
assign addr[5650]= 777438554;
assign addr[5651]= 917951481;
assign addr[5652]= 1053807919;
assign addr[5653]= 1184318708;
assign addr[5654]= 1308821808;
assign addr[5655]= 1426685652;
assign addr[5656]= 1537312353;
assign addr[5657]= 1640140734;
assign addr[5658]= 1734649179;
assign addr[5659]= 1820358275;
assign addr[5660]= 1896833245;
assign addr[5661]= 1963686155;
assign addr[5662]= 2020577882;
assign addr[5663]= 2067219829;
assign addr[5664]= 2103375398;
assign addr[5665]= 2128861181;
assign addr[5666]= 2143547897;
assign addr[5667]= 2147361045;
assign addr[5668]= 2140281282;
assign addr[5669]= 2122344521;
assign addr[5670]= 2093641749;
assign addr[5671]= 2054318569;
assign addr[5672]= 2004574453;
assign addr[5673]= 1944661739;
assign addr[5674]= 1874884346;
assign addr[5675]= 1795596234;
assign addr[5676]= 1707199606;
assign addr[5677]= 1610142873;
assign addr[5678]= 1504918373;
assign addr[5679]= 1392059879;
assign addr[5680]= 1272139887;
assign addr[5681]= 1145766716;
assign addr[5682]= 1013581418;
assign addr[5683]= 876254528;
assign addr[5684]= 734482665;
assign addr[5685]= 588984994;
assign addr[5686]= 440499581;
assign addr[5687]= 289779648;
assign addr[5688]= 137589750;
assign addr[5689]= -15298099;
assign addr[5690]= -168108346;
assign addr[5691]= -320065829;
assign addr[5692]= -470399716;
assign addr[5693]= -618347408;
assign addr[5694]= -763158411;
assign addr[5695]= -904098143;
assign addr[5696]= -1040451659;
assign addr[5697]= -1171527280;
assign addr[5698]= -1296660098;
assign addr[5699]= -1415215352;
assign addr[5700]= -1526591649;
assign addr[5701]= -1630224009;
assign addr[5702]= -1725586737;
assign addr[5703]= -1812196087;
assign addr[5704]= -1889612716;
assign addr[5705]= -1957443913;
assign addr[5706]= -2015345591;
assign addr[5707]= -2063024031;
assign addr[5708]= -2100237377;
assign addr[5709]= -2126796855;
assign addr[5710]= -2142567738;
assign addr[5711]= -2147470025;
assign addr[5712]= -2141478848;
assign addr[5713]= -2124624598;
assign addr[5714]= -2096992772;
assign addr[5715]= -2058723538;
assign addr[5716]= -2010011024;
assign addr[5717]= -1951102334;
assign addr[5718]= -1882296293;
assign addr[5719]= -1803941934;
assign addr[5720]= -1716436725;
assign addr[5721]= -1620224553;
assign addr[5722]= -1515793473;
assign addr[5723]= -1403673233;
assign addr[5724]= -1284432584;
assign addr[5725]= -1158676398;
assign addr[5726]= -1027042599;
assign addr[5727]= -890198924;
assign addr[5728]= -748839539;
assign addr[5729]= -603681519;
assign addr[5730]= -455461206;
assign addr[5731]= -304930476;
assign addr[5732]= -152852926;
assign addr[5733]= 0;
assign addr[5734]= 152852926;
assign addr[5735]= 304930476;
assign addr[5736]= 455461206;
assign addr[5737]= 603681519;
assign addr[5738]= 748839539;
assign addr[5739]= 890198924;
assign addr[5740]= 1027042599;
assign addr[5741]= 1158676398;
assign addr[5742]= 1284432584;
assign addr[5743]= 1403673233;
assign addr[5744]= 1515793473;
assign addr[5745]= 1620224553;
assign addr[5746]= 1716436725;
assign addr[5747]= 1803941934;
assign addr[5748]= 1882296293;
assign addr[5749]= 1951102334;
assign addr[5750]= 2010011024;
assign addr[5751]= 2058723538;
assign addr[5752]= 2096992772;
assign addr[5753]= 2124624598;
assign addr[5754]= 2141478848;
assign addr[5755]= 2147470025;
assign addr[5756]= 2142567738;
assign addr[5757]= 2126796855;
assign addr[5758]= 2100237377;
assign addr[5759]= 2063024031;
assign addr[5760]= 2015345591;
assign addr[5761]= 1957443913;
assign addr[5762]= 1889612716;
assign addr[5763]= 1812196087;
assign addr[5764]= 1725586737;
assign addr[5765]= 1630224009;
assign addr[5766]= 1526591649;
assign addr[5767]= 1415215352;
assign addr[5768]= 1296660098;
assign addr[5769]= 1171527280;
assign addr[5770]= 1040451659;
assign addr[5771]= 904098143;
assign addr[5772]= 763158411;
assign addr[5773]= 618347408;
assign addr[5774]= 470399716;
assign addr[5775]= 320065829;
assign addr[5776]= 168108346;
assign addr[5777]= 15298099;
assign addr[5778]= -137589750;
assign addr[5779]= -289779648;
assign addr[5780]= -440499581;
assign addr[5781]= -588984994;
assign addr[5782]= -734482665;
assign addr[5783]= -876254528;
assign addr[5784]= -1013581418;
assign addr[5785]= -1145766716;
assign addr[5786]= -1272139887;
assign addr[5787]= -1392059879;
assign addr[5788]= -1504918373;
assign addr[5789]= -1610142873;
assign addr[5790]= -1707199606;
assign addr[5791]= -1795596234;
assign addr[5792]= -1874884346;
assign addr[5793]= -1944661739;
assign addr[5794]= -2004574453;
assign addr[5795]= -2054318569;
assign addr[5796]= -2093641749;
assign addr[5797]= -2122344521;
assign addr[5798]= -2140281282;
assign addr[5799]= -2147361045;
assign addr[5800]= -2143547897;
assign addr[5801]= -2128861181;
assign addr[5802]= -2103375398;
assign addr[5803]= -2067219829;
assign addr[5804]= -2020577882;
assign addr[5805]= -1963686155;
assign addr[5806]= -1896833245;
assign addr[5807]= -1820358275;
assign addr[5808]= -1734649179;
assign addr[5809]= -1640140734;
assign addr[5810]= -1537312353;
assign addr[5811]= -1426685652;
assign addr[5812]= -1308821808;
assign addr[5813]= -1184318708;
assign addr[5814]= -1053807919;
assign addr[5815]= -917951481;
assign addr[5816]= -777438554;
assign addr[5817]= -632981917;
assign addr[5818]= -485314355;
assign addr[5819]= -335184940;
assign addr[5820]= -183355234;
assign addr[5821]= -30595422;
assign addr[5822]= 122319591;
assign addr[5823]= 274614114;
assign addr[5824]= 425515602;
assign addr[5825]= 574258580;
assign addr[5826]= 720088517;
assign addr[5827]= 862265664;
assign addr[5828]= 1000068799;
assign addr[5829]= 1132798888;
assign addr[5830]= 1259782632;
assign addr[5831]= 1380375881;
assign addr[5832]= 1493966902;
assign addr[5833]= 1599979481;
assign addr[5834]= 1697875851;
assign addr[5835]= 1787159411;
assign addr[5836]= 1867377253;
assign addr[5837]= 1938122457;
assign addr[5838]= 1999036154;
assign addr[5839]= 2049809346;
assign addr[5840]= 2090184478;
assign addr[5841]= 2119956737;
assign addr[5842]= 2138975100;
assign addr[5843]= 2147143090;
assign addr[5844]= 2144419275;
assign addr[5845]= 2130817471;
assign addr[5846]= 2106406677;
assign addr[5847]= 2071310720;
assign addr[5848]= 2025707632;
assign addr[5849]= 1969828744;
assign addr[5850]= 1903957513;
assign addr[5851]= 1828428082;
assign addr[5852]= 1743623590;
assign addr[5853]= 1649974225;
assign addr[5854]= 1547955041;
assign addr[5855]= 1438083551;
assign addr[5856]= 1320917099;
assign addr[5857]= 1197050035;
assign addr[5858]= 1067110699;
assign addr[5859]= 931758235;
assign addr[5860]= 791679244;
assign addr[5861]= 647584304;
assign addr[5862]= 500204365;
assign addr[5863]= 350287041;
assign addr[5864]= 198592817;
assign addr[5865]= 45891193;
assign addr[5866]= -107043224;
assign addr[5867]= -259434643;
assign addr[5868]= -410510029;
assign addr[5869]= -559503022;
assign addr[5870]= -705657826;
assign addr[5871]= -848233042;
assign addr[5872]= -986505429;
assign addr[5873]= -1119773573;
assign addr[5874]= -1247361445;
assign addr[5875]= -1368621831;
assign addr[5876]= -1482939614;
assign addr[5877]= -1589734894;
assign addr[5878]= -1688465931;
assign addr[5879]= -1778631892;
assign addr[5880]= -1859775393;
assign addr[5881]= -1931484818;
assign addr[5882]= -1993396407;
assign addr[5883]= -2045196100;
assign addr[5884]= -2086621133;
assign addr[5885]= -2117461370;
assign addr[5886]= -2137560369;
assign addr[5887]= -2146816171;
assign addr[5888]= -2145181827;
assign addr[5889]= -2132665626;
assign addr[5890]= -2109331059;
assign addr[5891]= -2075296495;
assign addr[5892]= -2030734582;
assign addr[5893]= -1975871368;
assign addr[5894]= -1910985158;
assign addr[5895]= -1836405100;
assign addr[5896]= -1752509516;
assign addr[5897]= -1659723983;
assign addr[5898]= -1558519173;
assign addr[5899]= -1449408469;
assign addr[5900]= -1332945355;
assign addr[5901]= -1209720613;
assign addr[5902]= -1080359326;
assign addr[5903]= -945517704;
assign addr[5904]= -805879757;
assign addr[5905]= -662153826;
assign addr[5906]= -515068990;
assign addr[5907]= -365371365;
assign addr[5908]= -213820322;
assign addr[5909]= -61184634;
assign addr[5910]= 91761426;
assign addr[5911]= 244242007;
assign addr[5912]= 395483624;
assign addr[5913]= 544719071;
assign addr[5914]= 691191324;
assign addr[5915]= 834157373;
assign addr[5916]= 972891995;
assign addr[5917]= 1106691431;
assign addr[5918]= 1234876957;
assign addr[5919]= 1356798326;
assign addr[5920]= 1471837070;
assign addr[5921]= 1579409630;
assign addr[5922]= 1678970324;
assign addr[5923]= 1770014111;
assign addr[5924]= 1852079154;
assign addr[5925]= 1924749160;
assign addr[5926]= 1987655498;
assign addr[5927]= 2040479063;
assign addr[5928]= 2082951896;
assign addr[5929]= 2114858546;
assign addr[5930]= 2136037160;
assign addr[5931]= 2146380306;
assign addr[5932]= 2145835515;
assign addr[5933]= 2134405552;
assign addr[5934]= 2112148396;
assign addr[5935]= 2079176953;
assign addr[5936]= 2035658475;
assign addr[5937]= 1981813720;
assign addr[5938]= 1917915825;
assign addr[5939]= 1844288924;
assign addr[5940]= 1761306505;
assign addr[5941]= 1669389513;
assign addr[5942]= 1569004214;
assign addr[5943]= 1460659832;
assign addr[5944]= 1344905966;
assign addr[5945]= 1222329801;
assign addr[5946]= 1093553126;
assign addr[5947]= 959229189;
assign addr[5948]= 820039373;
assign addr[5949]= 676689746;
assign addr[5950]= 529907477;
assign addr[5951]= 380437148;
assign addr[5952]= 229036977;
assign addr[5953]= 76474970;
assign addr[5954]= -76474970;
assign addr[5955]= -229036977;
assign addr[5956]= -380437148;
assign addr[5957]= -529907477;
assign addr[5958]= -676689746;
assign addr[5959]= -820039373;
assign addr[5960]= -959229189;
assign addr[5961]= -1093553126;
assign addr[5962]= -1222329801;
assign addr[5963]= -1344905966;
assign addr[5964]= -1460659832;
assign addr[5965]= -1569004214;
assign addr[5966]= -1669389513;
assign addr[5967]= -1761306505;
assign addr[5968]= -1844288924;
assign addr[5969]= -1917915825;
assign addr[5970]= -1981813720;
assign addr[5971]= -2035658475;
assign addr[5972]= -2079176953;
assign addr[5973]= -2112148396;
assign addr[5974]= -2134405552;
assign addr[5975]= -2145835515;
assign addr[5976]= -2146380306;
assign addr[5977]= -2136037160;
assign addr[5978]= -2114858546;
assign addr[5979]= -2082951896;
assign addr[5980]= -2040479063;
assign addr[5981]= -1987655498;
assign addr[5982]= -1924749160;
assign addr[5983]= -1852079154;
assign addr[5984]= -1770014111;
assign addr[5985]= -1678970324;
assign addr[5986]= -1579409630;
assign addr[5987]= -1471837070;
assign addr[5988]= -1356798326;
assign addr[5989]= -1234876957;
assign addr[5990]= -1106691431;
assign addr[5991]= -972891995;
assign addr[5992]= -834157373;
assign addr[5993]= -691191324;
assign addr[5994]= -544719071;
assign addr[5995]= -395483624;
assign addr[5996]= -244242007;
assign addr[5997]= -91761426;
assign addr[5998]= 61184634;
assign addr[5999]= 213820322;
assign addr[6000]= 365371365;
assign addr[6001]= 515068990;
assign addr[6002]= 662153826;
assign addr[6003]= 805879757;
assign addr[6004]= 945517704;
assign addr[6005]= 1080359326;
assign addr[6006]= 1209720613;
assign addr[6007]= 1332945355;
assign addr[6008]= 1449408469;
assign addr[6009]= 1558519173;
assign addr[6010]= 1659723983;
assign addr[6011]= 1752509516;
assign addr[6012]= 1836405100;
assign addr[6013]= 1910985158;
assign addr[6014]= 1975871368;
assign addr[6015]= 2030734582;
assign addr[6016]= 2075296495;
assign addr[6017]= 2109331059;
assign addr[6018]= 2132665626;
assign addr[6019]= 2145181827;
assign addr[6020]= 2146816171;
assign addr[6021]= 2137560369;
assign addr[6022]= 2117461370;
assign addr[6023]= 2086621133;
assign addr[6024]= 2045196100;
assign addr[6025]= 1993396407;
assign addr[6026]= 1931484818;
assign addr[6027]= 1859775393;
assign addr[6028]= 1778631892;
assign addr[6029]= 1688465931;
assign addr[6030]= 1589734894;
assign addr[6031]= 1482939614;
assign addr[6032]= 1368621831;
assign addr[6033]= 1247361445;
assign addr[6034]= 1119773573;
assign addr[6035]= 986505429;
assign addr[6036]= 848233042;
assign addr[6037]= 705657826;
assign addr[6038]= 559503022;
assign addr[6039]= 410510029;
assign addr[6040]= 259434643;
assign addr[6041]= 107043224;
assign addr[6042]= -45891193;
assign addr[6043]= -198592817;
assign addr[6044]= -350287041;
assign addr[6045]= -500204365;
assign addr[6046]= -647584304;
assign addr[6047]= -791679244;
assign addr[6048]= -931758235;
assign addr[6049]= -1067110699;
assign addr[6050]= -1197050035;
assign addr[6051]= -1320917099;
assign addr[6052]= -1438083551;
assign addr[6053]= -1547955041;
assign addr[6054]= -1649974225;
assign addr[6055]= -1743623590;
assign addr[6056]= -1828428082;
assign addr[6057]= -1903957513;
assign addr[6058]= -1969828744;
assign addr[6059]= -2025707632;
assign addr[6060]= -2071310720;
assign addr[6061]= -2106406677;
assign addr[6062]= -2130817471;
assign addr[6063]= -2144419275;
assign addr[6064]= -2147143090;
assign addr[6065]= -2138975100;
assign addr[6066]= -2119956737;
assign addr[6067]= -2090184478;
assign addr[6068]= -2049809346;
assign addr[6069]= -1999036154;
assign addr[6070]= -1938122457;
assign addr[6071]= -1867377253;
assign addr[6072]= -1787159411;
assign addr[6073]= -1697875851;
assign addr[6074]= -1599979481;
assign addr[6075]= -1493966902;
assign addr[6076]= -1380375881;
assign addr[6077]= -1259782632;
assign addr[6078]= -1132798888;
assign addr[6079]= -1000068799;
assign addr[6080]= -862265664;
assign addr[6081]= -720088517;
assign addr[6082]= -574258580;
assign addr[6083]= -425515602;
assign addr[6084]= -274614114;
assign addr[6085]= -122319591;
assign addr[6086]= 30595422;
assign addr[6087]= 183355234;
assign addr[6088]= 335184940;
assign addr[6089]= 485314355;
assign addr[6090]= 632981917;
assign addr[6091]= 777438554;
assign addr[6092]= 917951481;
assign addr[6093]= 1053807919;
assign addr[6094]= 1184318708;
assign addr[6095]= 1308821808;
assign addr[6096]= 1426685652;
assign addr[6097]= 1537312353;
assign addr[6098]= 1640140734;
assign addr[6099]= 1734649179;
assign addr[6100]= 1820358275;
assign addr[6101]= 1896833245;
assign addr[6102]= 1963686155;
assign addr[6103]= 2020577882;
assign addr[6104]= 2067219829;
assign addr[6105]= 2103375398;
assign addr[6106]= 2128861181;
assign addr[6107]= 2143547897;
assign addr[6108]= 2147361045;
assign addr[6109]= 2140281282;
assign addr[6110]= 2122344521;
assign addr[6111]= 2093641749;
assign addr[6112]= 2054318569;
assign addr[6113]= 2004574453;
assign addr[6114]= 1944661739;
assign addr[6115]= 1874884346;
assign addr[6116]= 1795596234;
assign addr[6117]= 1707199606;
assign addr[6118]= 1610142873;
assign addr[6119]= 1504918373;
assign addr[6120]= 1392059879;
assign addr[6121]= 1272139887;
assign addr[6122]= 1145766716;
assign addr[6123]= 1013581418;
assign addr[6124]= 876254528;
assign addr[6125]= 734482665;
assign addr[6126]= 588984994;
assign addr[6127]= 440499581;
assign addr[6128]= 289779648;
assign addr[6129]= 137589750;
assign addr[6130]= -15298099;
assign addr[6131]= -168108346;
assign addr[6132]= -320065829;
assign addr[6133]= -470399716;
assign addr[6134]= -618347408;
assign addr[6135]= -763158411;
assign addr[6136]= -904098143;
assign addr[6137]= -1040451659;
assign addr[6138]= -1171527280;
assign addr[6139]= -1296660098;
assign addr[6140]= -1415215352;
assign addr[6141]= -1526591649;
assign addr[6142]= -1630224009;
assign addr[6143]= -1725586737;
assign addr[6144]= -1812196087;
assign addr[6145]= -1889612716;
assign addr[6146]= -1957443913;
assign addr[6147]= -2015345591;
assign addr[6148]= -2063024031;
assign addr[6149]= -2100237377;
assign addr[6150]= -2126796855;
assign addr[6151]= -2142567738;
assign addr[6152]= -2147470025;
assign addr[6153]= -2141478848;
assign addr[6154]= -2124624598;
assign addr[6155]= -2096992772;
assign addr[6156]= -2058723538;
assign addr[6157]= -2010011024;
assign addr[6158]= -1951102334;
assign addr[6159]= -1882296293;
assign addr[6160]= -1803941934;
assign addr[6161]= -1716436725;
assign addr[6162]= -1620224553;
assign addr[6163]= -1515793473;
assign addr[6164]= -1403673233;
assign addr[6165]= -1284432584;
assign addr[6166]= -1158676398;
assign addr[6167]= -1027042599;
assign addr[6168]= -890198924;
assign addr[6169]= -748839539;
assign addr[6170]= -603681519;
assign addr[6171]= -455461206;
assign addr[6172]= -304930476;
assign addr[6173]= -152852926;
assign addr[6174]= 0;
assign addr[6175]= 152852926;
assign addr[6176]= 304930476;
assign addr[6177]= 455461206;
assign addr[6178]= 603681519;
assign addr[6179]= 748839539;
assign addr[6180]= 890198924;
assign addr[6181]= 1027042599;
assign addr[6182]= 1158676398;
assign addr[6183]= 1284432584;
assign addr[6184]= 1403673233;
assign addr[6185]= 1515793473;
assign addr[6186]= 1620224553;
assign addr[6187]= 1716436725;
assign addr[6188]= 1803941934;
assign addr[6189]= 1882296293;
assign addr[6190]= 1951102334;
assign addr[6191]= 2010011024;
assign addr[6192]= 2058723538;
assign addr[6193]= 2096992772;
assign addr[6194]= 2124624598;
assign addr[6195]= 2141478848;
assign addr[6196]= 2147470025;
assign addr[6197]= 2142567738;
assign addr[6198]= 2126796855;
assign addr[6199]= 2100237377;
assign addr[6200]= 2063024031;
assign addr[6201]= 2015345591;
assign addr[6202]= 1957443913;
assign addr[6203]= 1889612716;
assign addr[6204]= 1812196087;
assign addr[6205]= 1725586737;
assign addr[6206]= 1630224009;
assign addr[6207]= 1526591649;
assign addr[6208]= 1415215352;
assign addr[6209]= 1296660098;
assign addr[6210]= 1171527280;
assign addr[6211]= 1040451659;
assign addr[6212]= 904098143;
assign addr[6213]= 763158411;
assign addr[6214]= 618347408;
assign addr[6215]= 470399716;
assign addr[6216]= 320065829;
assign addr[6217]= 168108346;
assign addr[6218]= 15298099;
assign addr[6219]= -137589750;
assign addr[6220]= -289779648;
assign addr[6221]= -440499581;
assign addr[6222]= -588984994;
assign addr[6223]= -734482665;
assign addr[6224]= -876254528;
assign addr[6225]= -1013581418;
assign addr[6226]= -1145766716;
assign addr[6227]= -1272139887;
assign addr[6228]= -1392059879;
assign addr[6229]= -1504918373;
assign addr[6230]= -1610142873;
assign addr[6231]= -1707199606;
assign addr[6232]= -1795596234;
assign addr[6233]= -1874884346;
assign addr[6234]= -1944661739;
assign addr[6235]= -2004574453;
assign addr[6236]= -2054318569;
assign addr[6237]= -2093641749;
assign addr[6238]= -2122344521;
assign addr[6239]= -2140281282;
assign addr[6240]= -2147361045;
assign addr[6241]= -2143547897;
assign addr[6242]= -2128861181;
assign addr[6243]= -2103375398;
assign addr[6244]= -2067219829;
assign addr[6245]= -2020577882;
assign addr[6246]= -1963686155;
assign addr[6247]= -1896833245;
assign addr[6248]= -1820358275;
assign addr[6249]= -1734649179;
assign addr[6250]= -1640140734;
assign addr[6251]= -1537312353;
assign addr[6252]= -1426685652;
assign addr[6253]= -1308821808;
assign addr[6254]= -1184318708;
assign addr[6255]= -1053807919;
assign addr[6256]= -917951481;
assign addr[6257]= -777438554;
assign addr[6258]= -632981917;
assign addr[6259]= -485314355;
assign addr[6260]= -335184940;
assign addr[6261]= -183355234;
assign addr[6262]= -30595422;
assign addr[6263]= 122319591;
assign addr[6264]= 274614114;
assign addr[6265]= 425515602;
assign addr[6266]= 574258580;
assign addr[6267]= 720088517;
assign addr[6268]= 862265664;
assign addr[6269]= 1000068799;
assign addr[6270]= 1132798888;
assign addr[6271]= 1259782632;
assign addr[6272]= 1380375881;
assign addr[6273]= 1493966902;
assign addr[6274]= 1599979481;
assign addr[6275]= 1697875851;
assign addr[6276]= 1787159411;
assign addr[6277]= 1867377253;
assign addr[6278]= 1938122457;
assign addr[6279]= 1999036154;
assign addr[6280]= 2049809346;
assign addr[6281]= 2090184478;
assign addr[6282]= 2119956737;
assign addr[6283]= 2138975100;
assign addr[6284]= 2147143090;
assign addr[6285]= 2144419275;
assign addr[6286]= 2130817471;
assign addr[6287]= 2106406677;
assign addr[6288]= 2071310720;
assign addr[6289]= 2025707632;
assign addr[6290]= 1969828744;
assign addr[6291]= 1903957513;
assign addr[6292]= 1828428082;
assign addr[6293]= 1743623590;
assign addr[6294]= 1649974225;
assign addr[6295]= 1547955041;
assign addr[6296]= 1438083551;
assign addr[6297]= 1320917099;
assign addr[6298]= 1197050035;
assign addr[6299]= 1067110699;
assign addr[6300]= 931758235;
assign addr[6301]= 791679244;
assign addr[6302]= 647584304;
assign addr[6303]= 500204365;
assign addr[6304]= 350287041;
assign addr[6305]= 198592817;
assign addr[6306]= 45891193;
assign addr[6307]= -107043224;
assign addr[6308]= -259434643;
assign addr[6309]= -410510029;
assign addr[6310]= -559503022;
assign addr[6311]= -705657826;
assign addr[6312]= -848233042;
assign addr[6313]= -986505429;
assign addr[6314]= -1119773573;
assign addr[6315]= -1247361445;
assign addr[6316]= -1368621831;
assign addr[6317]= -1482939614;
assign addr[6318]= -1589734894;
assign addr[6319]= -1688465931;
assign addr[6320]= -1778631892;
assign addr[6321]= -1859775393;
assign addr[6322]= -1931484818;
assign addr[6323]= -1993396407;
assign addr[6324]= -2045196100;
assign addr[6325]= -2086621133;
assign addr[6326]= -2117461370;
assign addr[6327]= -2137560369;
assign addr[6328]= -2146816171;
assign addr[6329]= -2145181827;
assign addr[6330]= -2132665626;
assign addr[6331]= -2109331059;
assign addr[6332]= -2075296495;
assign addr[6333]= -2030734582;
assign addr[6334]= -1975871368;
assign addr[6335]= -1910985158;
assign addr[6336]= -1836405100;
assign addr[6337]= -1752509516;
assign addr[6338]= -1659723983;
assign addr[6339]= -1558519173;
assign addr[6340]= -1449408469;
assign addr[6341]= -1332945355;
assign addr[6342]= -1209720613;
assign addr[6343]= -1080359326;
assign addr[6344]= -945517704;
assign addr[6345]= -805879757;
assign addr[6346]= -662153826;
assign addr[6347]= -515068990;
assign addr[6348]= -365371365;
assign addr[6349]= -213820322;
assign addr[6350]= -61184634;
assign addr[6351]= 91761426;
assign addr[6352]= 244242007;
assign addr[6353]= 395483624;
assign addr[6354]= 544719071;
assign addr[6355]= 691191324;
assign addr[6356]= 834157373;
assign addr[6357]= 972891995;
assign addr[6358]= 1106691431;
assign addr[6359]= 1234876957;
assign addr[6360]= 1356798326;
assign addr[6361]= 1471837070;
assign addr[6362]= 1579409630;
assign addr[6363]= 1678970324;
assign addr[6364]= 1770014111;
assign addr[6365]= 1852079154;
assign addr[6366]= 1924749160;
assign addr[6367]= 1987655498;
assign addr[6368]= 2040479063;
assign addr[6369]= 2082951896;
assign addr[6370]= 2114858546;
assign addr[6371]= 2136037160;
assign addr[6372]= 2146380306;
assign addr[6373]= 2145835515;
assign addr[6374]= 2134405552;
assign addr[6375]= 2112148396;
assign addr[6376]= 2079176953;
assign addr[6377]= 2035658475;
assign addr[6378]= 1981813720;
assign addr[6379]= 1917915825;
assign addr[6380]= 1844288924;
assign addr[6381]= 1761306505;
assign addr[6382]= 1669389513;
assign addr[6383]= 1569004214;
assign addr[6384]= 1460659832;
assign addr[6385]= 1344905966;
assign addr[6386]= 1222329801;
assign addr[6387]= 1093553126;
assign addr[6388]= 959229189;
assign addr[6389]= 820039373;
assign addr[6390]= 676689746;
assign addr[6391]= 529907477;
assign addr[6392]= 380437148;
assign addr[6393]= 229036977;
assign addr[6394]= 76474970;
assign addr[6395]= -76474970;
assign addr[6396]= -229036977;
assign addr[6397]= -380437148;
assign addr[6398]= -529907477;
assign addr[6399]= -676689746;
assign addr[6400]= -820039373;
assign addr[6401]= -959229189;
assign addr[6402]= -1093553126;
assign addr[6403]= -1222329801;
assign addr[6404]= -1344905966;
assign addr[6405]= -1460659832;
assign addr[6406]= -1569004214;
assign addr[6407]= -1669389513;
assign addr[6408]= -1761306505;
assign addr[6409]= -1844288924;
assign addr[6410]= -1917915825;
assign addr[6411]= -1981813720;
assign addr[6412]= -2035658475;
assign addr[6413]= -2079176953;
assign addr[6414]= -2112148396;
assign addr[6415]= -2134405552;
assign addr[6416]= -2145835515;
assign addr[6417]= -2146380306;
assign addr[6418]= -2136037160;
assign addr[6419]= -2114858546;
assign addr[6420]= -2082951896;
assign addr[6421]= -2040479063;
assign addr[6422]= -1987655498;
assign addr[6423]= -1924749160;
assign addr[6424]= -1852079154;
assign addr[6425]= -1770014111;
assign addr[6426]= -1678970324;
assign addr[6427]= -1579409630;
assign addr[6428]= -1471837070;
assign addr[6429]= -1356798326;
assign addr[6430]= -1234876957;
assign addr[6431]= -1106691431;
assign addr[6432]= -972891995;
assign addr[6433]= -834157373;
assign addr[6434]= -691191324;
assign addr[6435]= -544719071;
assign addr[6436]= -395483624;
assign addr[6437]= -244242007;
assign addr[6438]= -91761426;
assign addr[6439]= 61184634;
assign addr[6440]= 213820322;
assign addr[6441]= 365371365;
assign addr[6442]= 515068990;
assign addr[6443]= 662153826;
assign addr[6444]= 805879757;
assign addr[6445]= 945517704;
assign addr[6446]= 1080359326;
assign addr[6447]= 1209720613;
assign addr[6448]= 1332945355;
assign addr[6449]= 1449408469;
assign addr[6450]= 1558519173;
assign addr[6451]= 1659723983;
assign addr[6452]= 1752509516;
assign addr[6453]= 1836405100;
assign addr[6454]= 1910985158;
assign addr[6455]= 1975871368;
assign addr[6456]= 2030734582;
assign addr[6457]= 2075296495;
assign addr[6458]= 2109331059;
assign addr[6459]= 2132665626;
assign addr[6460]= 2145181827;
assign addr[6461]= 2146816171;
assign addr[6462]= 2137560369;
assign addr[6463]= 2117461370;
assign addr[6464]= 2086621133;
assign addr[6465]= 2045196100;
assign addr[6466]= 1993396407;
assign addr[6467]= 1931484818;
assign addr[6468]= 1859775393;
assign addr[6469]= 1778631892;
assign addr[6470]= 1688465931;
assign addr[6471]= 1589734894;
assign addr[6472]= 1482939614;
assign addr[6473]= 1368621831;
assign addr[6474]= 1247361445;
assign addr[6475]= 1119773573;
assign addr[6476]= 986505429;
assign addr[6477]= 848233042;
assign addr[6478]= 705657826;
assign addr[6479]= 559503022;
assign addr[6480]= 410510029;
assign addr[6481]= 259434643;
assign addr[6482]= 107043224;
assign addr[6483]= -45891193;
assign addr[6484]= -198592817;
assign addr[6485]= -350287041;
assign addr[6486]= -500204365;
assign addr[6487]= -647584304;
assign addr[6488]= -791679244;
assign addr[6489]= -931758235;
assign addr[6490]= -1067110699;
assign addr[6491]= -1197050035;
assign addr[6492]= -1320917099;
assign addr[6493]= -1438083551;
assign addr[6494]= -1547955041;
assign addr[6495]= -1649974225;
assign addr[6496]= -1743623590;
assign addr[6497]= -1828428082;
assign addr[6498]= -1903957513;
assign addr[6499]= -1969828744;
assign addr[6500]= -2025707632;
assign addr[6501]= -2071310720;
assign addr[6502]= -2106406677;
assign addr[6503]= -2130817471;
assign addr[6504]= -2144419275;
assign addr[6505]= -2147143090;
assign addr[6506]= -2138975100;
assign addr[6507]= -2119956737;
assign addr[6508]= -2090184478;
assign addr[6509]= -2049809346;
assign addr[6510]= -1999036154;
assign addr[6511]= -1938122457;
assign addr[6512]= -1867377253;
assign addr[6513]= -1787159411;
assign addr[6514]= -1697875851;
assign addr[6515]= -1599979481;
assign addr[6516]= -1493966902;
assign addr[6517]= -1380375881;
assign addr[6518]= -1259782632;
assign addr[6519]= -1132798888;
assign addr[6520]= -1000068799;
assign addr[6521]= -862265664;
assign addr[6522]= -720088517;
assign addr[6523]= -574258580;
assign addr[6524]= -425515602;
assign addr[6525]= -274614114;
assign addr[6526]= -122319591;
assign addr[6527]= 30595422;
assign addr[6528]= 183355234;
assign addr[6529]= 335184940;
assign addr[6530]= 485314355;
assign addr[6531]= 632981917;
assign addr[6532]= 777438554;
assign addr[6533]= 917951481;
assign addr[6534]= 1053807919;
assign addr[6535]= 1184318708;
assign addr[6536]= 1308821808;
assign addr[6537]= 1426685652;
assign addr[6538]= 1537312353;
assign addr[6539]= 1640140734;
assign addr[6540]= 1734649179;
assign addr[6541]= 1820358275;
assign addr[6542]= 1896833245;
assign addr[6543]= 1963686155;
assign addr[6544]= 2020577882;
assign addr[6545]= 2067219829;
assign addr[6546]= 2103375398;
assign addr[6547]= 2128861181;
assign addr[6548]= 2143547897;
assign addr[6549]= 2147361045;
assign addr[6550]= 2140281282;
assign addr[6551]= 2122344521;
assign addr[6552]= 2093641749;
assign addr[6553]= 2054318569;
assign addr[6554]= 2004574453;
assign addr[6555]= 1944661739;
assign addr[6556]= 1874884346;
assign addr[6557]= 1795596234;
assign addr[6558]= 1707199606;
assign addr[6559]= 1610142873;
assign addr[6560]= 1504918373;
assign addr[6561]= 1392059879;
assign addr[6562]= 1272139887;
assign addr[6563]= 1145766716;
assign addr[6564]= 1013581418;
assign addr[6565]= 876254528;
assign addr[6566]= 734482665;
assign addr[6567]= 588984994;
assign addr[6568]= 440499581;
assign addr[6569]= 289779648;
assign addr[6570]= 137589750;
assign addr[6571]= -15298099;
assign addr[6572]= -168108346;
assign addr[6573]= -320065829;
assign addr[6574]= -470399716;
assign addr[6575]= -618347408;
assign addr[6576]= -763158411;
assign addr[6577]= -904098143;
assign addr[6578]= -1040451659;
assign addr[6579]= -1171527280;
assign addr[6580]= -1296660098;
assign addr[6581]= -1415215352;
assign addr[6582]= -1526591649;
assign addr[6583]= -1630224009;
assign addr[6584]= -1725586737;
assign addr[6585]= -1812196087;
assign addr[6586]= -1889612716;
assign addr[6587]= -1957443913;
assign addr[6588]= -2015345591;
assign addr[6589]= -2063024031;
assign addr[6590]= -2100237377;
assign addr[6591]= -2126796855;
assign addr[6592]= -2142567738;
assign addr[6593]= -2147470025;
assign addr[6594]= -2141478848;
assign addr[6595]= -2124624598;
assign addr[6596]= -2096992772;
assign addr[6597]= -2058723538;
assign addr[6598]= -2010011024;
assign addr[6599]= -1951102334;
assign addr[6600]= -1882296293;
assign addr[6601]= -1803941934;
assign addr[6602]= -1716436725;
assign addr[6603]= -1620224553;
assign addr[6604]= -1515793473;
assign addr[6605]= -1403673233;
assign addr[6606]= -1284432584;
assign addr[6607]= -1158676398;
assign addr[6608]= -1027042599;
assign addr[6609]= -890198924;
assign addr[6610]= -748839539;
assign addr[6611]= -603681519;
assign addr[6612]= -455461206;
assign addr[6613]= -304930476;
assign addr[6614]= -152852926;
assign addr[6615]= 0;
assign addr[6616]= 152852926;
assign addr[6617]= 304930476;
assign addr[6618]= 455461206;
assign addr[6619]= 603681519;
assign addr[6620]= 748839539;
assign addr[6621]= 890198924;
assign addr[6622]= 1027042599;
assign addr[6623]= 1158676398;
assign addr[6624]= 1284432584;
assign addr[6625]= 1403673233;
assign addr[6626]= 1515793473;
assign addr[6627]= 1620224553;
assign addr[6628]= 1716436725;
assign addr[6629]= 1803941934;
assign addr[6630]= 1882296293;
assign addr[6631]= 1951102334;
assign addr[6632]= 2010011024;
assign addr[6633]= 2058723538;
assign addr[6634]= 2096992772;
assign addr[6635]= 2124624598;
assign addr[6636]= 2141478848;
assign addr[6637]= 2147470025;
assign addr[6638]= 2142567738;
assign addr[6639]= 2126796855;
assign addr[6640]= 2100237377;
assign addr[6641]= 2063024031;
assign addr[6642]= 2015345591;
assign addr[6643]= 1957443913;
assign addr[6644]= 1889612716;
assign addr[6645]= 1812196087;
assign addr[6646]= 1725586737;
assign addr[6647]= 1630224009;
assign addr[6648]= 1526591649;
assign addr[6649]= 1415215352;
assign addr[6650]= 1296660098;
assign addr[6651]= 1171527280;
assign addr[6652]= 1040451659;
assign addr[6653]= 904098143;
assign addr[6654]= 763158411;
assign addr[6655]= 618347408;
assign addr[6656]= 470399716;
assign addr[6657]= 320065829;
assign addr[6658]= 168108346;
assign addr[6659]= 15298099;
assign addr[6660]= -137589750;
assign addr[6661]= -289779648;
assign addr[6662]= -440499581;
assign addr[6663]= -588984994;
assign addr[6664]= -734482665;
assign addr[6665]= -876254528;
assign addr[6666]= -1013581418;
assign addr[6667]= -1145766716;
assign addr[6668]= -1272139887;
assign addr[6669]= -1392059879;
assign addr[6670]= -1504918373;
assign addr[6671]= -1610142873;
assign addr[6672]= -1707199606;
assign addr[6673]= -1795596234;
assign addr[6674]= -1874884346;
assign addr[6675]= -1944661739;
assign addr[6676]= -2004574453;
assign addr[6677]= -2054318569;
assign addr[6678]= -2093641749;
assign addr[6679]= -2122344521;
assign addr[6680]= -2140281282;
assign addr[6681]= -2147361045;
assign addr[6682]= -2143547897;
assign addr[6683]= -2128861181;
assign addr[6684]= -2103375398;
assign addr[6685]= -2067219829;
assign addr[6686]= -2020577882;
assign addr[6687]= -1963686155;
assign addr[6688]= -1896833245;
assign addr[6689]= -1820358275;
assign addr[6690]= -1734649179;
assign addr[6691]= -1640140734;
assign addr[6692]= -1537312353;
assign addr[6693]= -1426685652;
assign addr[6694]= -1308821808;
assign addr[6695]= -1184318708;
assign addr[6696]= -1053807919;
assign addr[6697]= -917951481;
assign addr[6698]= -777438554;
assign addr[6699]= -632981917;
assign addr[6700]= -485314355;
assign addr[6701]= -335184940;
assign addr[6702]= -183355234;
assign addr[6703]= -30595422;
assign addr[6704]= 122319591;
assign addr[6705]= 274614114;
assign addr[6706]= 425515602;
assign addr[6707]= 574258580;
assign addr[6708]= 720088517;
assign addr[6709]= 862265664;
assign addr[6710]= 1000068799;
assign addr[6711]= 1132798888;
assign addr[6712]= 1259782632;
assign addr[6713]= 1380375881;
assign addr[6714]= 1493966902;
assign addr[6715]= 1599979481;
assign addr[6716]= 1697875851;
assign addr[6717]= 1787159411;
assign addr[6718]= 1867377253;
assign addr[6719]= 1938122457;
assign addr[6720]= 1999036154;
assign addr[6721]= 2049809346;
assign addr[6722]= 2090184478;
assign addr[6723]= 2119956737;
assign addr[6724]= 2138975100;
assign addr[6725]= 2147143090;
assign addr[6726]= 2144419275;
assign addr[6727]= 2130817471;
assign addr[6728]= 2106406677;
assign addr[6729]= 2071310720;
assign addr[6730]= 2025707632;
assign addr[6731]= 1969828744;
assign addr[6732]= 1903957513;
assign addr[6733]= 1828428082;
assign addr[6734]= 1743623590;
assign addr[6735]= 1649974225;
assign addr[6736]= 1547955041;
assign addr[6737]= 1438083551;
assign addr[6738]= 1320917099;
assign addr[6739]= 1197050035;
assign addr[6740]= 1067110699;
assign addr[6741]= 931758235;
assign addr[6742]= 791679244;
assign addr[6743]= 647584304;
assign addr[6744]= 500204365;
assign addr[6745]= 350287041;
assign addr[6746]= 198592817;
assign addr[6747]= 45891193;
assign addr[6748]= -107043224;
assign addr[6749]= -259434643;
assign addr[6750]= -410510029;
assign addr[6751]= -559503022;
assign addr[6752]= -705657826;
assign addr[6753]= -848233042;
assign addr[6754]= -986505429;
assign addr[6755]= -1119773573;
assign addr[6756]= -1247361445;
assign addr[6757]= -1368621831;
assign addr[6758]= -1482939614;
assign addr[6759]= -1589734894;
assign addr[6760]= -1688465931;
assign addr[6761]= -1778631892;
assign addr[6762]= -1859775393;
assign addr[6763]= -1931484818;
assign addr[6764]= -1993396407;
assign addr[6765]= -2045196100;
assign addr[6766]= -2086621133;
assign addr[6767]= -2117461370;
assign addr[6768]= -2137560369;
assign addr[6769]= -2146816171;
assign addr[6770]= -2145181827;
assign addr[6771]= -2132665626;
assign addr[6772]= -2109331059;
assign addr[6773]= -2075296495;
assign addr[6774]= -2030734582;
assign addr[6775]= -1975871368;
assign addr[6776]= -1910985158;
assign addr[6777]= -1836405100;
assign addr[6778]= -1752509516;
assign addr[6779]= -1659723983;
assign addr[6780]= -1558519173;
assign addr[6781]= -1449408469;
assign addr[6782]= -1332945355;
assign addr[6783]= -1209720613;
assign addr[6784]= -1080359326;
assign addr[6785]= -945517704;
assign addr[6786]= -805879757;
assign addr[6787]= -662153826;
assign addr[6788]= -515068990;
assign addr[6789]= -365371365;
assign addr[6790]= -213820322;
assign addr[6791]= -61184634;
assign addr[6792]= 91761426;
assign addr[6793]= 244242007;
assign addr[6794]= 395483624;
assign addr[6795]= 544719071;
assign addr[6796]= 691191324;
assign addr[6797]= 834157373;
assign addr[6798]= 972891995;
assign addr[6799]= 1106691431;
assign addr[6800]= 1234876957;
assign addr[6801]= 1356798326;
assign addr[6802]= 1471837070;
assign addr[6803]= 1579409630;
assign addr[6804]= 1678970324;
assign addr[6805]= 1770014111;
assign addr[6806]= 1852079154;
assign addr[6807]= 1924749160;
assign addr[6808]= 1987655498;
assign addr[6809]= 2040479063;
assign addr[6810]= 2082951896;
assign addr[6811]= 2114858546;
assign addr[6812]= 2136037160;
assign addr[6813]= 2146380306;
assign addr[6814]= 2145835515;
assign addr[6815]= 2134405552;
assign addr[6816]= 2112148396;
assign addr[6817]= 2079176953;
assign addr[6818]= 2035658475;
assign addr[6819]= 1981813720;
assign addr[6820]= 1917915825;
assign addr[6821]= 1844288924;
assign addr[6822]= 1761306505;
assign addr[6823]= 1669389513;
assign addr[6824]= 1569004214;
assign addr[6825]= 1460659832;
assign addr[6826]= 1344905966;
assign addr[6827]= 1222329801;
assign addr[6828]= 1093553126;
assign addr[6829]= 959229189;
assign addr[6830]= 820039373;
assign addr[6831]= 676689746;
assign addr[6832]= 529907477;
assign addr[6833]= 380437148;
assign addr[6834]= 229036977;
assign addr[6835]= 76474970;
assign addr[6836]= -76474970;
assign addr[6837]= -229036977;
assign addr[6838]= -380437148;
assign addr[6839]= -529907477;
assign addr[6840]= -676689746;
assign addr[6841]= -820039373;
assign addr[6842]= -959229189;
assign addr[6843]= -1093553126;
assign addr[6844]= -1222329801;
assign addr[6845]= -1344905966;
assign addr[6846]= -1460659832;
assign addr[6847]= -1569004214;
assign addr[6848]= -1669389513;
assign addr[6849]= -1761306505;
assign addr[6850]= -1844288924;
assign addr[6851]= -1917915825;
assign addr[6852]= -1981813720;
assign addr[6853]= -2035658475;
assign addr[6854]= -2079176953;
assign addr[6855]= -2112148396;
assign addr[6856]= -2134405552;
assign addr[6857]= -2145835515;
assign addr[6858]= -2146380306;
assign addr[6859]= -2136037160;
assign addr[6860]= -2114858546;
assign addr[6861]= -2082951896;
assign addr[6862]= -2040479063;
assign addr[6863]= -1987655498;
assign addr[6864]= -1924749160;
assign addr[6865]= -1852079154;
assign addr[6866]= -1770014111;
assign addr[6867]= -1678970324;
assign addr[6868]= -1579409630;
assign addr[6869]= -1471837070;
assign addr[6870]= -1356798326;
assign addr[6871]= -1234876957;
assign addr[6872]= -1106691431;
assign addr[6873]= -972891995;
assign addr[6874]= -834157373;
assign addr[6875]= -691191324;
assign addr[6876]= -544719071;
assign addr[6877]= -395483624;
assign addr[6878]= -244242007;
assign addr[6879]= -91761426;
assign addr[6880]= 61184634;
assign addr[6881]= 213820322;
assign addr[6882]= 365371365;
assign addr[6883]= 515068990;
assign addr[6884]= 662153826;
assign addr[6885]= 805879757;
assign addr[6886]= 945517704;
assign addr[6887]= 1080359326;
assign addr[6888]= 1209720613;
assign addr[6889]= 1332945355;
assign addr[6890]= 1449408469;
assign addr[6891]= 1558519173;
assign addr[6892]= 1659723983;
assign addr[6893]= 1752509516;
assign addr[6894]= 1836405100;
assign addr[6895]= 1910985158;
assign addr[6896]= 1975871368;
assign addr[6897]= 2030734582;
assign addr[6898]= 2075296495;
assign addr[6899]= 2109331059;
assign addr[6900]= 2132665626;
assign addr[6901]= 2145181827;
assign addr[6902]= 2146816171;
assign addr[6903]= 2137560369;
assign addr[6904]= 2117461370;
assign addr[6905]= 2086621133;
assign addr[6906]= 2045196100;
assign addr[6907]= 1993396407;
assign addr[6908]= 1931484818;
assign addr[6909]= 1859775393;
assign addr[6910]= 1778631892;
assign addr[6911]= 1688465931;
assign addr[6912]= 1589734894;
assign addr[6913]= 1482939614;
assign addr[6914]= 1368621831;
assign addr[6915]= 1247361445;
assign addr[6916]= 1119773573;
assign addr[6917]= 986505429;
assign addr[6918]= 848233042;
assign addr[6919]= 705657826;
assign addr[6920]= 559503022;
assign addr[6921]= 410510029;
assign addr[6922]= 259434643;
assign addr[6923]= 107043224;
assign addr[6924]= -45891193;
assign addr[6925]= -198592817;
assign addr[6926]= -350287041;
assign addr[6927]= -500204365;
assign addr[6928]= -647584304;
assign addr[6929]= -791679244;
assign addr[6930]= -931758235;
assign addr[6931]= -1067110699;
assign addr[6932]= -1197050035;
assign addr[6933]= -1320917099;
assign addr[6934]= -1438083551;
assign addr[6935]= -1547955041;
assign addr[6936]= -1649974225;
assign addr[6937]= -1743623590;
assign addr[6938]= -1828428082;
assign addr[6939]= -1903957513;
assign addr[6940]= -1969828744;
assign addr[6941]= -2025707632;
assign addr[6942]= -2071310720;
assign addr[6943]= -2106406677;
assign addr[6944]= -2130817471;
assign addr[6945]= -2144419275;
assign addr[6946]= -2147143090;
assign addr[6947]= -2138975100;
assign addr[6948]= -2119956737;
assign addr[6949]= -2090184478;
assign addr[6950]= -2049809346;
assign addr[6951]= -1999036154;
assign addr[6952]= -1938122457;
assign addr[6953]= -1867377253;
assign addr[6954]= -1787159411;
assign addr[6955]= -1697875851;
assign addr[6956]= -1599979481;
assign addr[6957]= -1493966902;
assign addr[6958]= -1380375881;
assign addr[6959]= -1259782632;
assign addr[6960]= -1132798888;
assign addr[6961]= -1000068799;
assign addr[6962]= -862265664;
assign addr[6963]= -720088517;
assign addr[6964]= -574258580;
assign addr[6965]= -425515602;
assign addr[6966]= -274614114;
assign addr[6967]= -122319591;
assign addr[6968]= 30595422;
assign addr[6969]= 183355234;
assign addr[6970]= 335184940;
assign addr[6971]= 485314355;
assign addr[6972]= 632981917;
assign addr[6973]= 777438554;
assign addr[6974]= 917951481;
assign addr[6975]= 1053807919;
assign addr[6976]= 1184318708;
assign addr[6977]= 1308821808;
assign addr[6978]= 1426685652;
assign addr[6979]= 1537312353;
assign addr[6980]= 1640140734;
assign addr[6981]= 1734649179;
assign addr[6982]= 1820358275;
assign addr[6983]= 1896833245;
assign addr[6984]= 1963686155;
assign addr[6985]= 2020577882;
assign addr[6986]= 2067219829;
assign addr[6987]= 2103375398;
assign addr[6988]= 2128861181;
assign addr[6989]= 2143547897;
assign addr[6990]= 2147361045;
assign addr[6991]= 2140281282;
assign addr[6992]= 2122344521;
assign addr[6993]= 2093641749;
assign addr[6994]= 2054318569;
assign addr[6995]= 2004574453;
assign addr[6996]= 1944661739;
assign addr[6997]= 1874884346;
assign addr[6998]= 1795596234;
assign addr[6999]= 1707199606;
assign addr[7000]= 1610142873;
assign addr[7001]= 1504918373;
assign addr[7002]= 1392059879;
assign addr[7003]= 1272139887;
assign addr[7004]= 1145766716;
assign addr[7005]= 1013581418;
assign addr[7006]= 876254528;
assign addr[7007]= 734482665;
assign addr[7008]= 588984994;
assign addr[7009]= 440499581;
assign addr[7010]= 289779648;
assign addr[7011]= 137589750;
assign addr[7012]= -15298099;
assign addr[7013]= -168108346;
assign addr[7014]= -320065829;
assign addr[7015]= -470399716;
assign addr[7016]= -618347408;
assign addr[7017]= -763158411;
assign addr[7018]= -904098143;
assign addr[7019]= -1040451659;
assign addr[7020]= -1171527280;
assign addr[7021]= -1296660098;
assign addr[7022]= -1415215352;
assign addr[7023]= -1526591649;
assign addr[7024]= -1630224009;
assign addr[7025]= -1725586737;
assign addr[7026]= -1812196087;
assign addr[7027]= -1889612716;
assign addr[7028]= -1957443913;
assign addr[7029]= -2015345591;
assign addr[7030]= -2063024031;
assign addr[7031]= -2100237377;
assign addr[7032]= -2126796855;
assign addr[7033]= -2142567738;
assign addr[7034]= -2147470025;
assign addr[7035]= -2141478848;
assign addr[7036]= -2124624598;
assign addr[7037]= -2096992772;
assign addr[7038]= -2058723538;
assign addr[7039]= -2010011024;
assign addr[7040]= -1951102334;
assign addr[7041]= -1882296293;
assign addr[7042]= -1803941934;
assign addr[7043]= -1716436725;
assign addr[7044]= -1620224553;
assign addr[7045]= -1515793473;
assign addr[7046]= -1403673233;
assign addr[7047]= -1284432584;
assign addr[7048]= -1158676398;
assign addr[7049]= -1027042599;
assign addr[7050]= -890198924;
assign addr[7051]= -748839539;
assign addr[7052]= -603681519;
assign addr[7053]= -455461206;
assign addr[7054]= -304930476;
assign addr[7055]= -152852926;
assign addr[7056]= 0;
assign addr[7057]= 152852926;
assign addr[7058]= 304930476;
assign addr[7059]= 455461206;
assign addr[7060]= 603681519;
assign addr[7061]= 748839539;
assign addr[7062]= 890198924;
assign addr[7063]= 1027042599;
assign addr[7064]= 1158676398;
assign addr[7065]= 1284432584;
assign addr[7066]= 1403673233;
assign addr[7067]= 1515793473;
assign addr[7068]= 1620224553;
assign addr[7069]= 1716436725;
assign addr[7070]= 1803941934;
assign addr[7071]= 1882296293;
assign addr[7072]= 1951102334;
assign addr[7073]= 2010011024;
assign addr[7074]= 2058723538;
assign addr[7075]= 2096992772;
assign addr[7076]= 2124624598;
assign addr[7077]= 2141478848;
assign addr[7078]= 2147470025;
assign addr[7079]= 2142567738;
assign addr[7080]= 2126796855;
assign addr[7081]= 2100237377;
assign addr[7082]= 2063024031;
assign addr[7083]= 2015345591;
assign addr[7084]= 1957443913;
assign addr[7085]= 1889612716;
assign addr[7086]= 1812196087;
assign addr[7087]= 1725586737;
assign addr[7088]= 1630224009;
assign addr[7089]= 1526591649;
assign addr[7090]= 1415215352;
assign addr[7091]= 1296660098;
assign addr[7092]= 1171527280;
assign addr[7093]= 1040451659;
assign addr[7094]= 904098143;
assign addr[7095]= 763158411;
assign addr[7096]= 618347408;
assign addr[7097]= 470399716;
assign addr[7098]= 320065829;
assign addr[7099]= 168108346;
assign addr[7100]= 15298099;
assign addr[7101]= -137589750;
assign addr[7102]= -289779648;
assign addr[7103]= -440499581;
assign addr[7104]= -588984994;
assign addr[7105]= -734482665;
assign addr[7106]= -876254528;
assign addr[7107]= -1013581418;
assign addr[7108]= -1145766716;
assign addr[7109]= -1272139887;
assign addr[7110]= -1392059879;
assign addr[7111]= -1504918373;
assign addr[7112]= -1610142873;
assign addr[7113]= -1707199606;
assign addr[7114]= -1795596234;
assign addr[7115]= -1874884346;
assign addr[7116]= -1944661739;
assign addr[7117]= -2004574453;
assign addr[7118]= -2054318569;
assign addr[7119]= -2093641749;
assign addr[7120]= -2122344521;
assign addr[7121]= -2140281282;
assign addr[7122]= -2147361045;
assign addr[7123]= -2143547897;
assign addr[7124]= -2128861181;
assign addr[7125]= -2103375398;
assign addr[7126]= -2067219829;
assign addr[7127]= -2020577882;
assign addr[7128]= -1963686155;
assign addr[7129]= -1896833245;
assign addr[7130]= -1820358275;
assign addr[7131]= -1734649179;
assign addr[7132]= -1640140734;
assign addr[7133]= -1537312353;
assign addr[7134]= -1426685652;
assign addr[7135]= -1308821808;
assign addr[7136]= -1184318708;
assign addr[7137]= -1053807919;
assign addr[7138]= -917951481;
assign addr[7139]= -777438554;
assign addr[7140]= -632981917;
assign addr[7141]= -485314355;
assign addr[7142]= -335184940;
assign addr[7143]= -183355234;
assign addr[7144]= -30595422;
assign addr[7145]= 122319591;
assign addr[7146]= 274614114;
assign addr[7147]= 425515602;
assign addr[7148]= 574258580;
assign addr[7149]= 720088517;
assign addr[7150]= 862265664;
assign addr[7151]= 1000068799;
assign addr[7152]= 1132798888;
assign addr[7153]= 1259782632;
assign addr[7154]= 1380375881;
assign addr[7155]= 1493966902;
assign addr[7156]= 1599979481;
assign addr[7157]= 1697875851;
assign addr[7158]= 1787159411;
assign addr[7159]= 1867377253;
assign addr[7160]= 1938122457;
assign addr[7161]= 1999036154;
assign addr[7162]= 2049809346;
assign addr[7163]= 2090184478;
assign addr[7164]= 2119956737;
assign addr[7165]= 2138975100;
assign addr[7166]= 2147143090;
assign addr[7167]= 2144419275;
assign addr[7168]= 2130817471;
assign addr[7169]= 2106406677;
assign addr[7170]= 2071310720;
assign addr[7171]= 2025707632;
assign addr[7172]= 1969828744;
assign addr[7173]= 1903957513;
assign addr[7174]= 1828428082;
assign addr[7175]= 1743623590;
assign addr[7176]= 1649974225;
assign addr[7177]= 1547955041;
assign addr[7178]= 1438083551;
assign addr[7179]= 1320917099;
assign addr[7180]= 1197050035;
assign addr[7181]= 1067110699;
assign addr[7182]= 931758235;
assign addr[7183]= 791679244;
assign addr[7184]= 647584304;
assign addr[7185]= 500204365;
assign addr[7186]= 350287041;
assign addr[7187]= 198592817;
assign addr[7188]= 45891193;
assign addr[7189]= -107043224;
assign addr[7190]= -259434643;
assign addr[7191]= -410510029;
assign addr[7192]= -559503022;
assign addr[7193]= -705657826;
assign addr[7194]= -848233042;
assign addr[7195]= -986505429;
assign addr[7196]= -1119773573;
assign addr[7197]= -1247361445;
assign addr[7198]= -1368621831;
assign addr[7199]= -1482939614;
assign addr[7200]= -1589734894;
assign addr[7201]= -1688465931;
assign addr[7202]= -1778631892;
assign addr[7203]= -1859775393;
assign addr[7204]= -1931484818;
assign addr[7205]= -1993396407;
assign addr[7206]= -2045196100;
assign addr[7207]= -2086621133;
assign addr[7208]= -2117461370;
assign addr[7209]= -2137560369;
assign addr[7210]= -2146816171;
assign addr[7211]= -2145181827;
assign addr[7212]= -2132665626;
assign addr[7213]= -2109331059;
assign addr[7214]= -2075296495;
assign addr[7215]= -2030734582;
assign addr[7216]= -1975871368;
assign addr[7217]= -1910985158;
assign addr[7218]= -1836405100;
assign addr[7219]= -1752509516;
assign addr[7220]= -1659723983;
assign addr[7221]= -1558519173;
assign addr[7222]= -1449408469;
assign addr[7223]= -1332945355;
assign addr[7224]= -1209720613;
assign addr[7225]= -1080359326;
assign addr[7226]= -945517704;
assign addr[7227]= -805879757;
assign addr[7228]= -662153826;
assign addr[7229]= -515068990;
assign addr[7230]= -365371365;
assign addr[7231]= -213820322;
assign addr[7232]= -61184634;
assign addr[7233]= 91761426;
assign addr[7234]= 244242007;
assign addr[7235]= 395483624;
assign addr[7236]= 544719071;
assign addr[7237]= 691191324;
assign addr[7238]= 834157373;
assign addr[7239]= 972891995;
assign addr[7240]= 1106691431;
assign addr[7241]= 1234876957;
assign addr[7242]= 1356798326;
assign addr[7243]= 1471837070;
assign addr[7244]= 1579409630;
assign addr[7245]= 1678970324;
assign addr[7246]= 1770014111;
assign addr[7247]= 1852079154;
assign addr[7248]= 1924749160;
assign addr[7249]= 1987655498;
assign addr[7250]= 2040479063;
assign addr[7251]= 2082951896;
assign addr[7252]= 2114858546;
assign addr[7253]= 2136037160;
assign addr[7254]= 2146380306;
assign addr[7255]= 2145835515;
assign addr[7256]= 2134405552;
assign addr[7257]= 2112148396;
assign addr[7258]= 2079176953;
assign addr[7259]= 2035658475;
assign addr[7260]= 1981813720;
assign addr[7261]= 1917915825;
assign addr[7262]= 1844288924;
assign addr[7263]= 1761306505;
assign addr[7264]= 1669389513;
assign addr[7265]= 1569004214;
assign addr[7266]= 1460659832;
assign addr[7267]= 1344905966;
assign addr[7268]= 1222329801;
assign addr[7269]= 1093553126;
assign addr[7270]= 959229189;
assign addr[7271]= 820039373;
assign addr[7272]= 676689746;
assign addr[7273]= 529907477;
assign addr[7274]= 380437148;
assign addr[7275]= 229036977;
assign addr[7276]= 76474970;
assign addr[7277]= -76474970;
assign addr[7278]= -229036977;
assign addr[7279]= -380437148;
assign addr[7280]= -529907477;
assign addr[7281]= -676689746;
assign addr[7282]= -820039373;
assign addr[7283]= -959229189;
assign addr[7284]= -1093553126;
assign addr[7285]= -1222329801;
assign addr[7286]= -1344905966;
assign addr[7287]= -1460659832;
assign addr[7288]= -1569004214;
assign addr[7289]= -1669389513;
assign addr[7290]= -1761306505;
assign addr[7291]= -1844288924;
assign addr[7292]= -1917915825;
assign addr[7293]= -1981813720;
assign addr[7294]= -2035658475;
assign addr[7295]= -2079176953;
assign addr[7296]= -2112148396;
assign addr[7297]= -2134405552;
assign addr[7298]= -2145835515;
assign addr[7299]= -2146380306;
assign addr[7300]= -2136037160;
assign addr[7301]= -2114858546;
assign addr[7302]= -2082951896;
assign addr[7303]= -2040479063;
assign addr[7304]= -1987655498;
assign addr[7305]= -1924749160;
assign addr[7306]= -1852079154;
assign addr[7307]= -1770014111;
assign addr[7308]= -1678970324;
assign addr[7309]= -1579409630;
assign addr[7310]= -1471837070;
assign addr[7311]= -1356798326;
assign addr[7312]= -1234876957;
assign addr[7313]= -1106691431;
assign addr[7314]= -972891995;
assign addr[7315]= -834157373;
assign addr[7316]= -691191324;
assign addr[7317]= -544719071;
assign addr[7318]= -395483624;
assign addr[7319]= -244242007;
assign addr[7320]= -91761426;
assign addr[7321]= 61184634;
assign addr[7322]= 213820322;
assign addr[7323]= 365371365;
assign addr[7324]= 515068990;
assign addr[7325]= 662153826;
assign addr[7326]= 805879757;
assign addr[7327]= 945517704;
assign addr[7328]= 1080359326;
assign addr[7329]= 1209720613;
assign addr[7330]= 1332945355;
assign addr[7331]= 1449408469;
assign addr[7332]= 1558519173;
assign addr[7333]= 1659723983;
assign addr[7334]= 1752509516;
assign addr[7335]= 1836405100;
assign addr[7336]= 1910985158;
assign addr[7337]= 1975871368;
assign addr[7338]= 2030734582;
assign addr[7339]= 2075296495;
assign addr[7340]= 2109331059;
assign addr[7341]= 2132665626;
assign addr[7342]= 2145181827;
assign addr[7343]= 2146816171;
assign addr[7344]= 2137560369;
assign addr[7345]= 2117461370;
assign addr[7346]= 2086621133;
assign addr[7347]= 2045196100;
assign addr[7348]= 1993396407;
assign addr[7349]= 1931484818;
assign addr[7350]= 1859775393;
assign addr[7351]= 1778631892;
assign addr[7352]= 1688465931;
assign addr[7353]= 1589734894;
assign addr[7354]= 1482939614;
assign addr[7355]= 1368621831;
assign addr[7356]= 1247361445;
assign addr[7357]= 1119773573;
assign addr[7358]= 986505429;
assign addr[7359]= 848233042;
assign addr[7360]= 705657826;
assign addr[7361]= 559503022;
assign addr[7362]= 410510029;
assign addr[7363]= 259434643;
assign addr[7364]= 107043224;
assign addr[7365]= -45891193;
assign addr[7366]= -198592817;
assign addr[7367]= -350287041;
assign addr[7368]= -500204365;
assign addr[7369]= -647584304;
assign addr[7370]= -791679244;
assign addr[7371]= -931758235;
assign addr[7372]= -1067110699;
assign addr[7373]= -1197050035;
assign addr[7374]= -1320917099;
assign addr[7375]= -1438083551;
assign addr[7376]= -1547955041;
assign addr[7377]= -1649974225;
assign addr[7378]= -1743623590;
assign addr[7379]= -1828428082;
assign addr[7380]= -1903957513;
assign addr[7381]= -1969828744;
assign addr[7382]= -2025707632;
assign addr[7383]= -2071310720;
assign addr[7384]= -2106406677;
assign addr[7385]= -2130817471;
assign addr[7386]= -2144419275;
assign addr[7387]= -2147143090;
assign addr[7388]= -2138975100;
assign addr[7389]= -2119956737;
assign addr[7390]= -2090184478;
assign addr[7391]= -2049809346;
assign addr[7392]= -1999036154;
assign addr[7393]= -1938122457;
assign addr[7394]= -1867377253;
assign addr[7395]= -1787159411;
assign addr[7396]= -1697875851;
assign addr[7397]= -1599979481;
assign addr[7398]= -1493966902;
assign addr[7399]= -1380375881;
assign addr[7400]= -1259782632;
assign addr[7401]= -1132798888;
assign addr[7402]= -1000068799;
assign addr[7403]= -862265664;
assign addr[7404]= -720088517;
assign addr[7405]= -574258580;
assign addr[7406]= -425515602;
assign addr[7407]= -274614114;
assign addr[7408]= -122319591;
assign addr[7409]= 30595422;
assign addr[7410]= 183355234;
assign addr[7411]= 335184940;
assign addr[7412]= 485314355;
assign addr[7413]= 632981917;
assign addr[7414]= 777438554;
assign addr[7415]= 917951481;
assign addr[7416]= 1053807919;
assign addr[7417]= 1184318708;
assign addr[7418]= 1308821808;
assign addr[7419]= 1426685652;
assign addr[7420]= 1537312353;
assign addr[7421]= 1640140734;
assign addr[7422]= 1734649179;
assign addr[7423]= 1820358275;
assign addr[7424]= 1896833245;
assign addr[7425]= 1963686155;
assign addr[7426]= 2020577882;
assign addr[7427]= 2067219829;
assign addr[7428]= 2103375398;
assign addr[7429]= 2128861181;
assign addr[7430]= 2143547897;
assign addr[7431]= 2147361045;
assign addr[7432]= 2140281282;
assign addr[7433]= 2122344521;
assign addr[7434]= 2093641749;
assign addr[7435]= 2054318569;
assign addr[7436]= 2004574453;
assign addr[7437]= 1944661739;
assign addr[7438]= 1874884346;
assign addr[7439]= 1795596234;
assign addr[7440]= 1707199606;
assign addr[7441]= 1610142873;
assign addr[7442]= 1504918373;
assign addr[7443]= 1392059879;
assign addr[7444]= 1272139887;
assign addr[7445]= 1145766716;
assign addr[7446]= 1013581418;
assign addr[7447]= 876254528;
assign addr[7448]= 734482665;
assign addr[7449]= 588984994;
assign addr[7450]= 440499581;
assign addr[7451]= 289779648;
assign addr[7452]= 137589750;
assign addr[7453]= -15298099;
assign addr[7454]= -168108346;
assign addr[7455]= -320065829;
assign addr[7456]= -470399716;
assign addr[7457]= -618347408;
assign addr[7458]= -763158411;
assign addr[7459]= -904098143;
assign addr[7460]= -1040451659;
assign addr[7461]= -1171527280;
assign addr[7462]= -1296660098;
assign addr[7463]= -1415215352;
assign addr[7464]= -1526591649;
assign addr[7465]= -1630224009;
assign addr[7466]= -1725586737;
assign addr[7467]= -1812196087;
assign addr[7468]= -1889612716;
assign addr[7469]= -1957443913;
assign addr[7470]= -2015345591;
assign addr[7471]= -2063024031;
assign addr[7472]= -2100237377;
assign addr[7473]= -2126796855;
assign addr[7474]= -2142567738;
assign addr[7475]= -2147470025;
assign addr[7476]= -2141478848;
assign addr[7477]= -2124624598;
assign addr[7478]= -2096992772;
assign addr[7479]= -2058723538;
assign addr[7480]= -2010011024;
assign addr[7481]= -1951102334;
assign addr[7482]= -1882296293;
assign addr[7483]= -1803941934;
assign addr[7484]= -1716436725;
assign addr[7485]= -1620224553;
assign addr[7486]= -1515793473;
assign addr[7487]= -1403673233;
assign addr[7488]= -1284432584;
assign addr[7489]= -1158676398;
assign addr[7490]= -1027042599;
assign addr[7491]= -890198924;
assign addr[7492]= -748839539;
assign addr[7493]= -603681519;
assign addr[7494]= -455461206;
assign addr[7495]= -304930476;
assign addr[7496]= -152852926;
assign addr[7497]= 0;
assign addr[7498]= 152852926;
assign addr[7499]= 304930476;
assign addr[7500]= 455461206;
assign addr[7501]= 603681519;
assign addr[7502]= 748839539;
assign addr[7503]= 890198924;
assign addr[7504]= 1027042599;
assign addr[7505]= 1158676398;
assign addr[7506]= 1284432584;
assign addr[7507]= 1403673233;
assign addr[7508]= 1515793473;
assign addr[7509]= 1620224553;
assign addr[7510]= 1716436725;
assign addr[7511]= 1803941934;
assign addr[7512]= 1882296293;
assign addr[7513]= 1951102334;
assign addr[7514]= 2010011024;
assign addr[7515]= 2058723538;
assign addr[7516]= 2096992772;
assign addr[7517]= 2124624598;
assign addr[7518]= 2141478848;
assign addr[7519]= 2147470025;
assign addr[7520]= 2142567738;
assign addr[7521]= 2126796855;
assign addr[7522]= 2100237377;
assign addr[7523]= 2063024031;
assign addr[7524]= 2015345591;
assign addr[7525]= 1957443913;
assign addr[7526]= 1889612716;
assign addr[7527]= 1812196087;
assign addr[7528]= 1725586737;
assign addr[7529]= 1630224009;
assign addr[7530]= 1526591649;
assign addr[7531]= 1415215352;
assign addr[7532]= 1296660098;
assign addr[7533]= 1171527280;
assign addr[7534]= 1040451659;
assign addr[7535]= 904098143;
assign addr[7536]= 763158411;
assign addr[7537]= 618347408;
assign addr[7538]= 470399716;
assign addr[7539]= 320065829;
assign addr[7540]= 168108346;
assign addr[7541]= 15298099;
assign addr[7542]= -137589750;
assign addr[7543]= -289779648;
assign addr[7544]= -440499581;
assign addr[7545]= -588984994;
assign addr[7546]= -734482665;
assign addr[7547]= -876254528;
assign addr[7548]= -1013581418;
assign addr[7549]= -1145766716;
assign addr[7550]= -1272139887;
assign addr[7551]= -1392059879;
assign addr[7552]= -1504918373;
assign addr[7553]= -1610142873;
assign addr[7554]= -1707199606;
assign addr[7555]= -1795596234;
assign addr[7556]= -1874884346;
assign addr[7557]= -1944661739;
assign addr[7558]= -2004574453;
assign addr[7559]= -2054318569;
assign addr[7560]= -2093641749;
assign addr[7561]= -2122344521;
assign addr[7562]= -2140281282;
assign addr[7563]= -2147361045;
assign addr[7564]= -2143547897;
assign addr[7565]= -2128861181;
assign addr[7566]= -2103375398;
assign addr[7567]= -2067219829;
assign addr[7568]= -2020577882;
assign addr[7569]= -1963686155;
assign addr[7570]= -1896833245;
assign addr[7571]= -1820358275;
assign addr[7572]= -1734649179;
assign addr[7573]= -1640140734;
assign addr[7574]= -1537312353;
assign addr[7575]= -1426685652;
assign addr[7576]= -1308821808;
assign addr[7577]= -1184318708;
assign addr[7578]= -1053807919;
assign addr[7579]= -917951481;
assign addr[7580]= -777438554;
assign addr[7581]= -632981917;
assign addr[7582]= -485314355;
assign addr[7583]= -335184940;
assign addr[7584]= -183355234;
assign addr[7585]= -30595422;
assign addr[7586]= 122319591;
assign addr[7587]= 274614114;
assign addr[7588]= 425515602;
assign addr[7589]= 574258580;
assign addr[7590]= 720088517;
assign addr[7591]= 862265664;
assign addr[7592]= 1000068799;
assign addr[7593]= 1132798888;
assign addr[7594]= 1259782632;
assign addr[7595]= 1380375881;
assign addr[7596]= 1493966902;
assign addr[7597]= 1599979481;
assign addr[7598]= 1697875851;
assign addr[7599]= 1787159411;
assign addr[7600]= 1867377253;
assign addr[7601]= 1938122457;
assign addr[7602]= 1999036154;
assign addr[7603]= 2049809346;
assign addr[7604]= 2090184478;
assign addr[7605]= 2119956737;
assign addr[7606]= 2138975100;
assign addr[7607]= 2147143090;
assign addr[7608]= 2144419275;
assign addr[7609]= 2130817471;
assign addr[7610]= 2106406677;
assign addr[7611]= 2071310720;
assign addr[7612]= 2025707632;
assign addr[7613]= 1969828744;
assign addr[7614]= 1903957513;
assign addr[7615]= 1828428082;
assign addr[7616]= 1743623590;
assign addr[7617]= 1649974225;
assign addr[7618]= 1547955041;
assign addr[7619]= 1438083551;
assign addr[7620]= 1320917099;
assign addr[7621]= 1197050035;
assign addr[7622]= 1067110699;
assign addr[7623]= 931758235;
assign addr[7624]= 791679244;
assign addr[7625]= 647584304;
assign addr[7626]= 500204365;
assign addr[7627]= 350287041;
assign addr[7628]= 198592817;
assign addr[7629]= 45891193;
assign addr[7630]= -107043224;
assign addr[7631]= -259434643;
assign addr[7632]= -410510029;
assign addr[7633]= -559503022;
assign addr[7634]= -705657826;
assign addr[7635]= -848233042;
assign addr[7636]= -986505429;
assign addr[7637]= -1119773573;
assign addr[7638]= -1247361445;
assign addr[7639]= -1368621831;
assign addr[7640]= -1482939614;
assign addr[7641]= -1589734894;
assign addr[7642]= -1688465931;
assign addr[7643]= -1778631892;
assign addr[7644]= -1859775393;
assign addr[7645]= -1931484818;
assign addr[7646]= -1993396407;
assign addr[7647]= -2045196100;
assign addr[7648]= -2086621133;
assign addr[7649]= -2117461370;
assign addr[7650]= -2137560369;
assign addr[7651]= -2146816171;
assign addr[7652]= -2145181827;
assign addr[7653]= -2132665626;
assign addr[7654]= -2109331059;
assign addr[7655]= -2075296495;
assign addr[7656]= -2030734582;
assign addr[7657]= -1975871368;
assign addr[7658]= -1910985158;
assign addr[7659]= -1836405100;
assign addr[7660]= -1752509516;
assign addr[7661]= -1659723983;
assign addr[7662]= -1558519173;
assign addr[7663]= -1449408469;
assign addr[7664]= -1332945355;
assign addr[7665]= -1209720613;
assign addr[7666]= -1080359326;
assign addr[7667]= -945517704;
assign addr[7668]= -805879757;
assign addr[7669]= -662153826;
assign addr[7670]= -515068990;
assign addr[7671]= -365371365;
assign addr[7672]= -213820322;
assign addr[7673]= -61184634;
assign addr[7674]= 91761426;
assign addr[7675]= 244242007;
assign addr[7676]= 395483624;
assign addr[7677]= 544719071;
assign addr[7678]= 691191324;
assign addr[7679]= 834157373;
assign addr[7680]= 972891995;
assign addr[7681]= 1106691431;
assign addr[7682]= 1234876957;
assign addr[7683]= 1356798326;
assign addr[7684]= 1471837070;
assign addr[7685]= 1579409630;
assign addr[7686]= 1678970324;
assign addr[7687]= 1770014111;
assign addr[7688]= 1852079154;
assign addr[7689]= 1924749160;
assign addr[7690]= 1987655498;
assign addr[7691]= 2040479063;
assign addr[7692]= 2082951896;
assign addr[7693]= 2114858546;
assign addr[7694]= 2136037160;
assign addr[7695]= 2146380306;
assign addr[7696]= 2145835515;
assign addr[7697]= 2134405552;
assign addr[7698]= 2112148396;
assign addr[7699]= 2079176953;
assign addr[7700]= 2035658475;
assign addr[7701]= 1981813720;
assign addr[7702]= 1917915825;
assign addr[7703]= 1844288924;
assign addr[7704]= 1761306505;
assign addr[7705]= 1669389513;
assign addr[7706]= 1569004214;
assign addr[7707]= 1460659832;
assign addr[7708]= 1344905966;
assign addr[7709]= 1222329801;
assign addr[7710]= 1093553126;
assign addr[7711]= 959229189;
assign addr[7712]= 820039373;
assign addr[7713]= 676689746;
assign addr[7714]= 529907477;
assign addr[7715]= 380437148;
assign addr[7716]= 229036977;
assign addr[7717]= 76474970;
assign addr[7718]= -76474970;
assign addr[7719]= -229036977;
assign addr[7720]= -380437148;
assign addr[7721]= -529907477;
assign addr[7722]= -676689746;
assign addr[7723]= -820039373;
assign addr[7724]= -959229189;
assign addr[7725]= -1093553126;
assign addr[7726]= -1222329801;
assign addr[7727]= -1344905966;
assign addr[7728]= -1460659832;
assign addr[7729]= -1569004214;
assign addr[7730]= -1669389513;
assign addr[7731]= -1761306505;
assign addr[7732]= -1844288924;
assign addr[7733]= -1917915825;
assign addr[7734]= -1981813720;
assign addr[7735]= -2035658475;
assign addr[7736]= -2079176953;
assign addr[7737]= -2112148396;
assign addr[7738]= -2134405552;
assign addr[7739]= -2145835515;
assign addr[7740]= -2146380306;
assign addr[7741]= -2136037160;
assign addr[7742]= -2114858546;
assign addr[7743]= -2082951896;
assign addr[7744]= -2040479063;
assign addr[7745]= -1987655498;
assign addr[7746]= -1924749160;
assign addr[7747]= -1852079154;
assign addr[7748]= -1770014111;
assign addr[7749]= -1678970324;
assign addr[7750]= -1579409630;
assign addr[7751]= -1471837070;
assign addr[7752]= -1356798326;
assign addr[7753]= -1234876957;
assign addr[7754]= -1106691431;
assign addr[7755]= -972891995;
assign addr[7756]= -834157373;
assign addr[7757]= -691191324;
assign addr[7758]= -544719071;
assign addr[7759]= -395483624;
assign addr[7760]= -244242007;
assign addr[7761]= -91761426;
assign addr[7762]= 61184634;
assign addr[7763]= 213820322;
assign addr[7764]= 365371365;
assign addr[7765]= 515068990;
assign addr[7766]= 662153826;
assign addr[7767]= 805879757;
assign addr[7768]= 945517704;
assign addr[7769]= 1080359326;
assign addr[7770]= 1209720613;
assign addr[7771]= 1332945355;
assign addr[7772]= 1449408469;
assign addr[7773]= 1558519173;
assign addr[7774]= 1659723983;
assign addr[7775]= 1752509516;
assign addr[7776]= 1836405100;
assign addr[7777]= 1910985158;
assign addr[7778]= 1975871368;
assign addr[7779]= 2030734582;
assign addr[7780]= 2075296495;
assign addr[7781]= 2109331059;
assign addr[7782]= 2132665626;
assign addr[7783]= 2145181827;
assign addr[7784]= 2146816171;
assign addr[7785]= 2137560369;
assign addr[7786]= 2117461370;
assign addr[7787]= 2086621133;
assign addr[7788]= 2045196100;
assign addr[7789]= 1993396407;
assign addr[7790]= 1931484818;
assign addr[7791]= 1859775393;
assign addr[7792]= 1778631892;
assign addr[7793]= 1688465931;
assign addr[7794]= 1589734894;
assign addr[7795]= 1482939614;
assign addr[7796]= 1368621831;
assign addr[7797]= 1247361445;
assign addr[7798]= 1119773573;
assign addr[7799]= 986505429;
assign addr[7800]= 848233042;
assign addr[7801]= 705657826;
assign addr[7802]= 559503022;
assign addr[7803]= 410510029;
assign addr[7804]= 259434643;
assign addr[7805]= 107043224;
assign addr[7806]= -45891193;
assign addr[7807]= -198592817;
assign addr[7808]= -350287041;
assign addr[7809]= -500204365;
assign addr[7810]= -647584304;
assign addr[7811]= -791679244;
assign addr[7812]= -931758235;
assign addr[7813]= -1067110699;
assign addr[7814]= -1197050035;
assign addr[7815]= -1320917099;
assign addr[7816]= -1438083551;
assign addr[7817]= -1547955041;
assign addr[7818]= -1649974225;
assign addr[7819]= -1743623590;
assign addr[7820]= -1828428082;
assign addr[7821]= -1903957513;
assign addr[7822]= -1969828744;
assign addr[7823]= -2025707632;
assign addr[7824]= -2071310720;
assign addr[7825]= -2106406677;
assign addr[7826]= -2130817471;
assign addr[7827]= -2144419275;
assign addr[7828]= -2147143090;
assign addr[7829]= -2138975100;
assign addr[7830]= -2119956737;
assign addr[7831]= -2090184478;
assign addr[7832]= -2049809346;
assign addr[7833]= -1999036154;
assign addr[7834]= -1938122457;
assign addr[7835]= -1867377253;
assign addr[7836]= -1787159411;
assign addr[7837]= -1697875851;
assign addr[7838]= -1599979481;
assign addr[7839]= -1493966902;
assign addr[7840]= -1380375881;
assign addr[7841]= -1259782632;
assign addr[7842]= -1132798888;
assign addr[7843]= -1000068799;
assign addr[7844]= -862265664;
assign addr[7845]= -720088517;
assign addr[7846]= -574258580;
assign addr[7847]= -425515602;
assign addr[7848]= -274614114;
assign addr[7849]= -122319591;
assign addr[7850]= 30595422;
assign addr[7851]= 183355234;
assign addr[7852]= 335184940;
assign addr[7853]= 485314355;
assign addr[7854]= 632981917;
assign addr[7855]= 777438554;
assign addr[7856]= 917951481;
assign addr[7857]= 1053807919;
assign addr[7858]= 1184318708;
assign addr[7859]= 1308821808;
assign addr[7860]= 1426685652;
assign addr[7861]= 1537312353;
assign addr[7862]= 1640140734;
assign addr[7863]= 1734649179;
assign addr[7864]= 1820358275;
assign addr[7865]= 1896833245;
assign addr[7866]= 1963686155;
assign addr[7867]= 2020577882;
assign addr[7868]= 2067219829;
assign addr[7869]= 2103375398;
assign addr[7870]= 2128861181;
assign addr[7871]= 2143547897;
assign addr[7872]= 2147361045;
assign addr[7873]= 2140281282;
assign addr[7874]= 2122344521;
assign addr[7875]= 2093641749;
assign addr[7876]= 2054318569;
assign addr[7877]= 2004574453;
assign addr[7878]= 1944661739;
assign addr[7879]= 1874884346;
assign addr[7880]= 1795596234;
assign addr[7881]= 1707199606;
assign addr[7882]= 1610142873;
assign addr[7883]= 1504918373;
assign addr[7884]= 1392059879;
assign addr[7885]= 1272139887;
assign addr[7886]= 1145766716;
assign addr[7887]= 1013581418;
assign addr[7888]= 876254528;
assign addr[7889]= 734482665;
assign addr[7890]= 588984994;
assign addr[7891]= 440499581;
assign addr[7892]= 289779648;
assign addr[7893]= 137589750;
assign addr[7894]= -15298099;
assign addr[7895]= -168108346;
assign addr[7896]= -320065829;
assign addr[7897]= -470399716;
assign addr[7898]= -618347408;
assign addr[7899]= -763158411;
assign addr[7900]= -904098143;
assign addr[7901]= -1040451659;
assign addr[7902]= -1171527280;
assign addr[7903]= -1296660098;
assign addr[7904]= -1415215352;
assign addr[7905]= -1526591649;
assign addr[7906]= -1630224009;
assign addr[7907]= -1725586737;
assign addr[7908]= -1812196087;
assign addr[7909]= -1889612716;
assign addr[7910]= -1957443913;
assign addr[7911]= -2015345591;
assign addr[7912]= -2063024031;
assign addr[7913]= -2100237377;
assign addr[7914]= -2126796855;
assign addr[7915]= -2142567738;
assign addr[7916]= -2147470025;
assign addr[7917]= -2141478848;
assign addr[7918]= -2124624598;
assign addr[7919]= -2096992772;
assign addr[7920]= -2058723538;
assign addr[7921]= -2010011024;
assign addr[7922]= -1951102334;
assign addr[7923]= -1882296293;
assign addr[7924]= -1803941934;
assign addr[7925]= -1716436725;
assign addr[7926]= -1620224553;
assign addr[7927]= -1515793473;
assign addr[7928]= -1403673233;
assign addr[7929]= -1284432584;
assign addr[7930]= -1158676398;
assign addr[7931]= -1027042599;
assign addr[7932]= -890198924;
assign addr[7933]= -748839539;
assign addr[7934]= -603681519;
assign addr[7935]= -455461206;
assign addr[7936]= -304930476;
assign addr[7937]= -152852926;
assign addr[7938]= 0;
assign addr[7939]= 152852926;
assign addr[7940]= 304930476;
assign addr[7941]= 455461206;
assign addr[7942]= 603681519;
assign addr[7943]= 748839539;
assign addr[7944]= 890198924;
assign addr[7945]= 1027042599;
assign addr[7946]= 1158676398;
assign addr[7947]= 1284432584;
assign addr[7948]= 1403673233;
assign addr[7949]= 1515793473;
assign addr[7950]= 1620224553;
assign addr[7951]= 1716436725;
assign addr[7952]= 1803941934;
assign addr[7953]= 1882296293;
assign addr[7954]= 1951102334;
assign addr[7955]= 2010011024;
assign addr[7956]= 2058723538;
assign addr[7957]= 2096992772;
assign addr[7958]= 2124624598;
assign addr[7959]= 2141478848;
assign addr[7960]= 2147470025;
assign addr[7961]= 2142567738;
assign addr[7962]= 2126796855;
assign addr[7963]= 2100237377;
assign addr[7964]= 2063024031;
assign addr[7965]= 2015345591;
assign addr[7966]= 1957443913;
assign addr[7967]= 1889612716;
assign addr[7968]= 1812196087;
assign addr[7969]= 1725586737;
assign addr[7970]= 1630224009;
assign addr[7971]= 1526591649;
assign addr[7972]= 1415215352;
assign addr[7973]= 1296660098;
assign addr[7974]= 1171527280;
assign addr[7975]= 1040451659;
assign addr[7976]= 904098143;
assign addr[7977]= 763158411;
assign addr[7978]= 618347408;
assign addr[7979]= 470399716;
assign addr[7980]= 320065829;
assign addr[7981]= 168108346;
assign addr[7982]= 15298099;
assign addr[7983]= -137589750;
assign addr[7984]= -289779648;
assign addr[7985]= -440499581;
assign addr[7986]= -588984994;
assign addr[7987]= -734482665;
assign addr[7988]= -876254528;
assign addr[7989]= -1013581418;
assign addr[7990]= -1145766716;
assign addr[7991]= -1272139887;
assign addr[7992]= -1392059879;
assign addr[7993]= -1504918373;
assign addr[7994]= -1610142873;
assign addr[7995]= -1707199606;
assign addr[7996]= -1795596234;
assign addr[7997]= -1874884346;
assign addr[7998]= -1944661739;
assign addr[7999]= -2004574453;
assign addr[8000]= -2054318569;
assign addr[8001]= -2093641749;
assign addr[8002]= -2122344521;
assign addr[8003]= -2140281282;
assign addr[8004]= -2147361045;
assign addr[8005]= -2143547897;
assign addr[8006]= -2128861181;
assign addr[8007]= -2103375398;
assign addr[8008]= -2067219829;
assign addr[8009]= -2020577882;
assign addr[8010]= -1963686155;
assign addr[8011]= -1896833245;
assign addr[8012]= -1820358275;
assign addr[8013]= -1734649179;
assign addr[8014]= -1640140734;
assign addr[8015]= -1537312353;
assign addr[8016]= -1426685652;
assign addr[8017]= -1308821808;
assign addr[8018]= -1184318708;
assign addr[8019]= -1053807919;
assign addr[8020]= -917951481;
assign addr[8021]= -777438554;
assign addr[8022]= -632981917;
assign addr[8023]= -485314355;
assign addr[8024]= -335184940;
assign addr[8025]= -183355234;
assign addr[8026]= -30595422;
assign addr[8027]= 122319591;
assign addr[8028]= 274614114;
assign addr[8029]= 425515602;
assign addr[8030]= 574258580;
assign addr[8031]= 720088517;
assign addr[8032]= 862265664;
assign addr[8033]= 1000068799;
assign addr[8034]= 1132798888;
assign addr[8035]= 1259782632;
assign addr[8036]= 1380375881;
assign addr[8037]= 1493966902;
assign addr[8038]= 1599979481;
assign addr[8039]= 1697875851;
assign addr[8040]= 1787159411;
assign addr[8041]= 1867377253;
assign addr[8042]= 1938122457;
assign addr[8043]= 1999036154;
assign addr[8044]= 2049809346;
assign addr[8045]= 2090184478;
assign addr[8046]= 2119956737;
assign addr[8047]= 2138975100;
assign addr[8048]= 2147143090;
assign addr[8049]= 2144419275;
assign addr[8050]= 2130817471;
assign addr[8051]= 2106406677;
assign addr[8052]= 2071310720;
assign addr[8053]= 2025707632;
assign addr[8054]= 1969828744;
assign addr[8055]= 1903957513;
assign addr[8056]= 1828428082;
assign addr[8057]= 1743623590;
assign addr[8058]= 1649974225;
assign addr[8059]= 1547955041;
assign addr[8060]= 1438083551;
assign addr[8061]= 1320917099;
assign addr[8062]= 1197050035;
assign addr[8063]= 1067110699;
assign addr[8064]= 931758235;
assign addr[8065]= 791679244;
assign addr[8066]= 647584304;
assign addr[8067]= 500204365;
assign addr[8068]= 350287041;
assign addr[8069]= 198592817;
assign addr[8070]= 45891193;
assign addr[8071]= -107043224;
assign addr[8072]= -259434643;
assign addr[8073]= -410510029;
assign addr[8074]= -559503022;
assign addr[8075]= -705657826;
assign addr[8076]= -848233042;
assign addr[8077]= -986505429;
assign addr[8078]= -1119773573;
assign addr[8079]= -1247361445;
assign addr[8080]= -1368621831;
assign addr[8081]= -1482939614;
assign addr[8082]= -1589734894;
assign addr[8083]= -1688465931;
assign addr[8084]= -1778631892;
assign addr[8085]= -1859775393;
assign addr[8086]= -1931484818;
assign addr[8087]= -1993396407;
assign addr[8088]= -2045196100;
assign addr[8089]= -2086621133;
assign addr[8090]= -2117461370;
assign addr[8091]= -2137560369;
assign addr[8092]= -2146816171;
assign addr[8093]= -2145181827;
assign addr[8094]= -2132665626;
assign addr[8095]= -2109331059;
assign addr[8096]= -2075296495;
assign addr[8097]= -2030734582;
assign addr[8098]= -1975871368;
assign addr[8099]= -1910985158;
assign addr[8100]= -1836405100;
assign addr[8101]= -1752509516;
assign addr[8102]= -1659723983;
assign addr[8103]= -1558519173;
assign addr[8104]= -1449408469;
assign addr[8105]= -1332945355;
assign addr[8106]= -1209720613;
assign addr[8107]= -1080359326;
assign addr[8108]= -945517704;
assign addr[8109]= -805879757;
assign addr[8110]= -662153826;
assign addr[8111]= -515068990;
assign addr[8112]= -365371365;
assign addr[8113]= -213820322;
assign addr[8114]= -61184634;
assign addr[8115]= 91761426;
assign addr[8116]= 244242007;
assign addr[8117]= 395483624;
assign addr[8118]= 544719071;
assign addr[8119]= 691191324;
assign addr[8120]= 834157373;
assign addr[8121]= 972891995;
assign addr[8122]= 1106691431;
assign addr[8123]= 1234876957;
assign addr[8124]= 1356798326;
assign addr[8125]= 1471837070;
assign addr[8126]= 1579409630;
assign addr[8127]= 1678970324;
assign addr[8128]= 1770014111;
assign addr[8129]= 1852079154;
assign addr[8130]= 1924749160;
assign addr[8131]= 1987655498;
assign addr[8132]= 2040479063;
assign addr[8133]= 2082951896;
assign addr[8134]= 2114858546;
assign addr[8135]= 2136037160;
assign addr[8136]= 2146380306;
assign addr[8137]= 2145835515;
assign addr[8138]= 2134405552;
assign addr[8139]= 2112148396;
assign addr[8140]= 2079176953;
assign addr[8141]= 2035658475;
assign addr[8142]= 1981813720;
assign addr[8143]= 1917915825;
assign addr[8144]= 1844288924;
assign addr[8145]= 1761306505;
assign addr[8146]= 1669389513;
assign addr[8147]= 1569004214;
assign addr[8148]= 1460659832;
assign addr[8149]= 1344905966;
assign addr[8150]= 1222329801;
assign addr[8151]= 1093553126;
assign addr[8152]= 959229189;
assign addr[8153]= 820039373;
assign addr[8154]= 676689746;
assign addr[8155]= 529907477;
assign addr[8156]= 380437148;
assign addr[8157]= 229036977;
assign addr[8158]= 76474970;
assign addr[8159]= -76474970;
assign addr[8160]= -229036977;
assign addr[8161]= -380437148;
assign addr[8162]= -529907477;
assign addr[8163]= -676689746;
assign addr[8164]= -820039373;
assign addr[8165]= -959229189;
assign addr[8166]= -1093553126;
assign addr[8167]= -1222329801;
assign addr[8168]= -1344905966;
assign addr[8169]= -1460659832;
assign addr[8170]= -1569004214;
assign addr[8171]= -1669389513;
assign addr[8172]= -1761306505;
assign addr[8173]= -1844288924;
assign addr[8174]= -1917915825;
assign addr[8175]= -1981813720;
assign addr[8176]= -2035658475;
assign addr[8177]= -2079176953;
assign addr[8178]= -2112148396;
assign addr[8179]= -2134405552;
assign addr[8180]= -2145835515;
assign addr[8181]= -2146380306;
assign addr[8182]= -2136037160;
assign addr[8183]= -2114858546;
assign addr[8184]= -2082951896;
assign addr[8185]= -2040479063;
assign addr[8186]= -1987655498;
assign addr[8187]= -1924749160;
assign addr[8188]= -1852079154;
assign addr[8189]= -1770014111;
assign addr[8190]= -1678970324;
assign addr[8191]= -1579409630;
assign addr[8192]= -1471837070;
assign addr[8193]= -1356798326;
assign addr[8194]= -1234876957;
assign addr[8195]= -1106691431;
assign addr[8196]= -972891995;
assign addr[8197]= -834157373;
assign addr[8198]= -691191324;
assign addr[8199]= -544719071;
assign addr[8200]= -395483624;
assign addr[8201]= -244242007;
assign addr[8202]= -91761426;
assign addr[8203]= 61184634;
assign addr[8204]= 213820322;
assign addr[8205]= 365371365;
assign addr[8206]= 515068990;
assign addr[8207]= 662153826;
assign addr[8208]= 805879757;
assign addr[8209]= 945517704;
assign addr[8210]= 1080359326;
assign addr[8211]= 1209720613;
assign addr[8212]= 1332945355;
assign addr[8213]= 1449408469;
assign addr[8214]= 1558519173;
assign addr[8215]= 1659723983;
assign addr[8216]= 1752509516;
assign addr[8217]= 1836405100;
assign addr[8218]= 1910985158;
assign addr[8219]= 1975871368;
assign addr[8220]= 2030734582;
assign addr[8221]= 2075296495;
assign addr[8222]= 2109331059;
assign addr[8223]= 2132665626;
assign addr[8224]= 2145181827;
assign addr[8225]= 2146816171;
assign addr[8226]= 2137560369;
assign addr[8227]= 2117461370;
assign addr[8228]= 2086621133;
assign addr[8229]= 2045196100;
assign addr[8230]= 1993396407;
assign addr[8231]= 1931484818;
assign addr[8232]= 1859775393;
assign addr[8233]= 1778631892;
assign addr[8234]= 1688465931;
assign addr[8235]= 1589734894;
assign addr[8236]= 1482939614;
assign addr[8237]= 1368621831;
assign addr[8238]= 1247361445;
assign addr[8239]= 1119773573;
assign addr[8240]= 986505429;
assign addr[8241]= 848233042;
assign addr[8242]= 705657826;
assign addr[8243]= 559503022;
assign addr[8244]= 410510029;
assign addr[8245]= 259434643;
assign addr[8246]= 107043224;
assign addr[8247]= -45891193;
assign addr[8248]= -198592817;
assign addr[8249]= -350287041;
assign addr[8250]= -500204365;
assign addr[8251]= -647584304;
assign addr[8252]= -791679244;
assign addr[8253]= -931758235;
assign addr[8254]= -1067110699;
assign addr[8255]= -1197050035;
assign addr[8256]= -1320917099;
assign addr[8257]= -1438083551;
assign addr[8258]= -1547955041;
assign addr[8259]= -1649974225;
assign addr[8260]= -1743623590;
assign addr[8261]= -1828428082;
assign addr[8262]= -1903957513;
assign addr[8263]= -1969828744;
assign addr[8264]= -2025707632;
assign addr[8265]= -2071310720;
assign addr[8266]= -2106406677;
assign addr[8267]= -2130817471;
assign addr[8268]= -2144419275;
assign addr[8269]= -2147143090;
assign addr[8270]= -2138975100;
assign addr[8271]= -2119956737;
assign addr[8272]= -2090184478;
assign addr[8273]= -2049809346;
assign addr[8274]= -1999036154;
assign addr[8275]= -1938122457;
assign addr[8276]= -1867377253;
assign addr[8277]= -1787159411;
assign addr[8278]= -1697875851;
assign addr[8279]= -1599979481;
assign addr[8280]= -1493966902;
assign addr[8281]= -1380375881;
assign addr[8282]= -1259782632;
assign addr[8283]= -1132798888;
assign addr[8284]= -1000068799;
assign addr[8285]= -862265664;
assign addr[8286]= -720088517;
assign addr[8287]= -574258580;
assign addr[8288]= -425515602;
assign addr[8289]= -274614114;
assign addr[8290]= -122319591;
assign addr[8291]= 30595422;
assign addr[8292]= 183355234;
assign addr[8293]= 335184940;
assign addr[8294]= 485314355;
assign addr[8295]= 632981917;
assign addr[8296]= 777438554;
assign addr[8297]= 917951481;
assign addr[8298]= 1053807919;
assign addr[8299]= 1184318708;
assign addr[8300]= 1308821808;
assign addr[8301]= 1426685652;
assign addr[8302]= 1537312353;
assign addr[8303]= 1640140734;
assign addr[8304]= 1734649179;
assign addr[8305]= 1820358275;
assign addr[8306]= 1896833245;
assign addr[8307]= 1963686155;
assign addr[8308]= 2020577882;
assign addr[8309]= 2067219829;
assign addr[8310]= 2103375398;
assign addr[8311]= 2128861181;
assign addr[8312]= 2143547897;
assign addr[8313]= 2147361045;
assign addr[8314]= 2140281282;
assign addr[8315]= 2122344521;
assign addr[8316]= 2093641749;
assign addr[8317]= 2054318569;
assign addr[8318]= 2004574453;
assign addr[8319]= 1944661739;
assign addr[8320]= 1874884346;
assign addr[8321]= 1795596234;
assign addr[8322]= 1707199606;
assign addr[8323]= 1610142873;
assign addr[8324]= 1504918373;
assign addr[8325]= 1392059879;
assign addr[8326]= 1272139887;
assign addr[8327]= 1145766716;
assign addr[8328]= 1013581418;
assign addr[8329]= 876254528;
assign addr[8330]= 734482665;
assign addr[8331]= 588984994;
assign addr[8332]= 440499581;
assign addr[8333]= 289779648;
assign addr[8334]= 137589750;
assign addr[8335]= -15298099;
assign addr[8336]= -168108346;
assign addr[8337]= -320065829;
assign addr[8338]= -470399716;
assign addr[8339]= -618347408;
assign addr[8340]= -763158411;
assign addr[8341]= -904098143;
assign addr[8342]= -1040451659;
assign addr[8343]= -1171527280;
assign addr[8344]= -1296660098;
assign addr[8345]= -1415215352;
assign addr[8346]= -1526591649;
assign addr[8347]= -1630224009;
assign addr[8348]= -1725586737;
assign addr[8349]= -1812196087;
assign addr[8350]= -1889612716;
assign addr[8351]= -1957443913;
assign addr[8352]= -2015345591;
assign addr[8353]= -2063024031;
assign addr[8354]= -2100237377;
assign addr[8355]= -2126796855;
assign addr[8356]= -2142567738;
assign addr[8357]= -2147470025;
assign addr[8358]= -2141478848;
assign addr[8359]= -2124624598;
assign addr[8360]= -2096992772;
assign addr[8361]= -2058723538;
assign addr[8362]= -2010011024;
assign addr[8363]= -1951102334;
assign addr[8364]= -1882296293;
assign addr[8365]= -1803941934;
assign addr[8366]= -1716436725;
assign addr[8367]= -1620224553;
assign addr[8368]= -1515793473;
assign addr[8369]= -1403673233;
assign addr[8370]= -1284432584;
assign addr[8371]= -1158676398;
assign addr[8372]= -1027042599;
assign addr[8373]= -890198924;
assign addr[8374]= -748839539;
assign addr[8375]= -603681519;
assign addr[8376]= -455461206;
assign addr[8377]= -304930476;
assign addr[8378]= -152852926;
assign addr[8379]= 0;
assign addr[8380]= 152852926;
assign addr[8381]= 304930476;
assign addr[8382]= 455461206;
assign addr[8383]= 603681519;
assign addr[8384]= 748839539;
assign addr[8385]= 890198924;
assign addr[8386]= 1027042599;
assign addr[8387]= 1158676398;
assign addr[8388]= 1284432584;
assign addr[8389]= 1403673233;
assign addr[8390]= 1515793473;
assign addr[8391]= 1620224553;
assign addr[8392]= 1716436725;
assign addr[8393]= 1803941934;
assign addr[8394]= 1882296293;
assign addr[8395]= 1951102334;
assign addr[8396]= 2010011024;
assign addr[8397]= 2058723538;
assign addr[8398]= 2096992772;
assign addr[8399]= 2124624598;
assign addr[8400]= 2141478848;
assign addr[8401]= 2147470025;
assign addr[8402]= 2142567738;
assign addr[8403]= 2126796855;
assign addr[8404]= 2100237377;
assign addr[8405]= 2063024031;
assign addr[8406]= 2015345591;
assign addr[8407]= 1957443913;
assign addr[8408]= 1889612716;
assign addr[8409]= 1812196087;
assign addr[8410]= 1725586737;
assign addr[8411]= 1630224009;
assign addr[8412]= 1526591649;
assign addr[8413]= 1415215352;
assign addr[8414]= 1296660098;
assign addr[8415]= 1171527280;
assign addr[8416]= 1040451659;
assign addr[8417]= 904098143;
assign addr[8418]= 763158411;
assign addr[8419]= 618347408;
assign addr[8420]= 470399716;
assign addr[8421]= 320065829;
assign addr[8422]= 168108346;
assign addr[8423]= 15298099;
assign addr[8424]= -137589750;
assign addr[8425]= -289779648;
assign addr[8426]= -440499581;
assign addr[8427]= -588984994;
assign addr[8428]= -734482665;
assign addr[8429]= -876254528;
assign addr[8430]= -1013581418;
assign addr[8431]= -1145766716;
assign addr[8432]= -1272139887;
assign addr[8433]= -1392059879;
assign addr[8434]= -1504918373;
assign addr[8435]= -1610142873;
assign addr[8436]= -1707199606;
assign addr[8437]= -1795596234;
assign addr[8438]= -1874884346;
assign addr[8439]= -1944661739;
assign addr[8440]= -2004574453;
assign addr[8441]= -2054318569;
assign addr[8442]= -2093641749;
assign addr[8443]= -2122344521;
assign addr[8444]= -2140281282;
assign addr[8445]= -2147361045;
assign addr[8446]= -2143547897;
assign addr[8447]= -2128861181;
assign addr[8448]= -2103375398;
assign addr[8449]= -2067219829;
assign addr[8450]= -2020577882;
assign addr[8451]= -1963686155;
assign addr[8452]= -1896833245;
assign addr[8453]= -1820358275;
assign addr[8454]= -1734649179;
assign addr[8455]= -1640140734;
assign addr[8456]= -1537312353;
assign addr[8457]= -1426685652;
assign addr[8458]= -1308821808;
assign addr[8459]= -1184318708;
assign addr[8460]= -1053807919;
assign addr[8461]= -917951481;
assign addr[8462]= -777438554;
assign addr[8463]= -632981917;
assign addr[8464]= -485314355;
assign addr[8465]= -335184940;
assign addr[8466]= -183355234;
assign addr[8467]= -30595422;
assign addr[8468]= 122319591;
assign addr[8469]= 274614114;
assign addr[8470]= 425515602;
assign addr[8471]= 574258580;
assign addr[8472]= 720088517;
assign addr[8473]= 862265664;
assign addr[8474]= 1000068799;
assign addr[8475]= 1132798888;
assign addr[8476]= 1259782632;
assign addr[8477]= 1380375881;
assign addr[8478]= 1493966902;
assign addr[8479]= 1599979481;
assign addr[8480]= 1697875851;
assign addr[8481]= 1787159411;
assign addr[8482]= 1867377253;
assign addr[8483]= 1938122457;
assign addr[8484]= 1999036154;
assign addr[8485]= 2049809346;
assign addr[8486]= 2090184478;
assign addr[8487]= 2119956737;
assign addr[8488]= 2138975100;
assign addr[8489]= 2147143090;
assign addr[8490]= 2144419275;
assign addr[8491]= 2130817471;
assign addr[8492]= 2106406677;
assign addr[8493]= 2071310720;
assign addr[8494]= 2025707632;
assign addr[8495]= 1969828744;
assign addr[8496]= 1903957513;
assign addr[8497]= 1828428082;
assign addr[8498]= 1743623590;
assign addr[8499]= 1649974225;
assign addr[8500]= 1547955041;
assign addr[8501]= 1438083551;
assign addr[8502]= 1320917099;
assign addr[8503]= 1197050035;
assign addr[8504]= 1067110699;
assign addr[8505]= 931758235;
assign addr[8506]= 791679244;
assign addr[8507]= 647584304;
assign addr[8508]= 500204365;
assign addr[8509]= 350287041;
assign addr[8510]= 198592817;
assign addr[8511]= 45891193;
assign addr[8512]= -107043224;
assign addr[8513]= -259434643;
assign addr[8514]= -410510029;
assign addr[8515]= -559503022;
assign addr[8516]= -705657826;
assign addr[8517]= -848233042;
assign addr[8518]= -986505429;
assign addr[8519]= -1119773573;
assign addr[8520]= -1247361445;
assign addr[8521]= -1368621831;
assign addr[8522]= -1482939614;
assign addr[8523]= -1589734894;
assign addr[8524]= -1688465931;
assign addr[8525]= -1778631892;
assign addr[8526]= -1859775393;
assign addr[8527]= -1931484818;
assign addr[8528]= -1993396407;
assign addr[8529]= -2045196100;
assign addr[8530]= -2086621133;
assign addr[8531]= -2117461370;
assign addr[8532]= -2137560369;
assign addr[8533]= -2146816171;
assign addr[8534]= -2145181827;
assign addr[8535]= -2132665626;
assign addr[8536]= -2109331059;
assign addr[8537]= -2075296495;
assign addr[8538]= -2030734582;
assign addr[8539]= -1975871368;
assign addr[8540]= -1910985158;
assign addr[8541]= -1836405100;
assign addr[8542]= -1752509516;
assign addr[8543]= -1659723983;
assign addr[8544]= -1558519173;
assign addr[8545]= -1449408469;
assign addr[8546]= -1332945355;
assign addr[8547]= -1209720613;
assign addr[8548]= -1080359326;
assign addr[8549]= -945517704;
assign addr[8550]= -805879757;
assign addr[8551]= -662153826;
assign addr[8552]= -515068990;
assign addr[8553]= -365371365;
assign addr[8554]= -213820322;
assign addr[8555]= -61184634;
assign addr[8556]= 91761426;
assign addr[8557]= 244242007;
assign addr[8558]= 395483624;
assign addr[8559]= 544719071;
assign addr[8560]= 691191324;
assign addr[8561]= 834157373;
assign addr[8562]= 972891995;
assign addr[8563]= 1106691431;
assign addr[8564]= 1234876957;
assign addr[8565]= 1356798326;
assign addr[8566]= 1471837070;
assign addr[8567]= 1579409630;
assign addr[8568]= 1678970324;
assign addr[8569]= 1770014111;
assign addr[8570]= 1852079154;
assign addr[8571]= 1924749160;
assign addr[8572]= 1987655498;
assign addr[8573]= 2040479063;
assign addr[8574]= 2082951896;
assign addr[8575]= 2114858546;
assign addr[8576]= 2136037160;
assign addr[8577]= 2146380306;
assign addr[8578]= 2145835515;
assign addr[8579]= 2134405552;
assign addr[8580]= 2112148396;
assign addr[8581]= 2079176953;
assign addr[8582]= 2035658475;
assign addr[8583]= 1981813720;
assign addr[8584]= 1917915825;
assign addr[8585]= 1844288924;
assign addr[8586]= 1761306505;
assign addr[8587]= 1669389513;
assign addr[8588]= 1569004214;
assign addr[8589]= 1460659832;
assign addr[8590]= 1344905966;
assign addr[8591]= 1222329801;
assign addr[8592]= 1093553126;
assign addr[8593]= 959229189;
assign addr[8594]= 820039373;
assign addr[8595]= 676689746;
assign addr[8596]= 529907477;
assign addr[8597]= 380437148;
assign addr[8598]= 229036977;
assign addr[8599]= 76474970;
assign addr[8600]= -76474970;
assign addr[8601]= -229036977;
assign addr[8602]= -380437148;
assign addr[8603]= -529907477;
assign addr[8604]= -676689746;
assign addr[8605]= -820039373;
assign addr[8606]= -959229189;
assign addr[8607]= -1093553126;
assign addr[8608]= -1222329801;
assign addr[8609]= -1344905966;
assign addr[8610]= -1460659832;
assign addr[8611]= -1569004214;
assign addr[8612]= -1669389513;
assign addr[8613]= -1761306505;
assign addr[8614]= -1844288924;
assign addr[8615]= -1917915825;
assign addr[8616]= -1981813720;
assign addr[8617]= -2035658475;
assign addr[8618]= -2079176953;
assign addr[8619]= -2112148396;
assign addr[8620]= -2134405552;
assign addr[8621]= -2145835515;
assign addr[8622]= -2146380306;
assign addr[8623]= -2136037160;
assign addr[8624]= -2114858546;
assign addr[8625]= -2082951896;
assign addr[8626]= -2040479063;
assign addr[8627]= -1987655498;
assign addr[8628]= -1924749160;
assign addr[8629]= -1852079154;
assign addr[8630]= -1770014111;
assign addr[8631]= -1678970324;
assign addr[8632]= -1579409630;
assign addr[8633]= -1471837070;
assign addr[8634]= -1356798326;
assign addr[8635]= -1234876957;
assign addr[8636]= -1106691431;
assign addr[8637]= -972891995;
assign addr[8638]= -834157373;
assign addr[8639]= -691191324;
assign addr[8640]= -544719071;
assign addr[8641]= -395483624;
assign addr[8642]= -244242007;
assign addr[8643]= -91761426;
assign addr[8644]= 61184634;
assign addr[8645]= 213820322;
assign addr[8646]= 365371365;
assign addr[8647]= 515068990;
assign addr[8648]= 662153826;
assign addr[8649]= 805879757;
assign addr[8650]= 945517704;
assign addr[8651]= 1080359326;
assign addr[8652]= 1209720613;
assign addr[8653]= 1332945355;
assign addr[8654]= 1449408469;
assign addr[8655]= 1558519173;
assign addr[8656]= 1659723983;
assign addr[8657]= 1752509516;
assign addr[8658]= 1836405100;
assign addr[8659]= 1910985158;
assign addr[8660]= 1975871368;
assign addr[8661]= 2030734582;
assign addr[8662]= 2075296495;
assign addr[8663]= 2109331059;
assign addr[8664]= 2132665626;
assign addr[8665]= 2145181827;
assign addr[8666]= 2146816171;
assign addr[8667]= 2137560369;
assign addr[8668]= 2117461370;
assign addr[8669]= 2086621133;
assign addr[8670]= 2045196100;
assign addr[8671]= 1993396407;
assign addr[8672]= 1931484818;
assign addr[8673]= 1859775393;
assign addr[8674]= 1778631892;
assign addr[8675]= 1688465931;
assign addr[8676]= 1589734894;
assign addr[8677]= 1482939614;
assign addr[8678]= 1368621831;
assign addr[8679]= 1247361445;
assign addr[8680]= 1119773573;
assign addr[8681]= 986505429;
assign addr[8682]= 848233042;
assign addr[8683]= 705657826;
assign addr[8684]= 559503022;
assign addr[8685]= 410510029;
assign addr[8686]= 259434643;
assign addr[8687]= 107043224;
assign addr[8688]= -45891193;
assign addr[8689]= -198592817;
assign addr[8690]= -350287041;
assign addr[8691]= -500204365;
assign addr[8692]= -647584304;
assign addr[8693]= -791679244;
assign addr[8694]= -931758235;
assign addr[8695]= -1067110699;
assign addr[8696]= -1197050035;
assign addr[8697]= -1320917099;
assign addr[8698]= -1438083551;
assign addr[8699]= -1547955041;
assign addr[8700]= -1649974225;
assign addr[8701]= -1743623590;
assign addr[8702]= -1828428082;
assign addr[8703]= -1903957513;
assign addr[8704]= -1969828744;
assign addr[8705]= -2025707632;
assign addr[8706]= -2071310720;
assign addr[8707]= -2106406677;
assign addr[8708]= -2130817471;
assign addr[8709]= -2144419275;
assign addr[8710]= -2147143090;
assign addr[8711]= -2138975100;
assign addr[8712]= -2119956737;
assign addr[8713]= -2090184478;
assign addr[8714]= -2049809346;
assign addr[8715]= -1999036154;
assign addr[8716]= -1938122457;
assign addr[8717]= -1867377253;
assign addr[8718]= -1787159411;
assign addr[8719]= -1697875851;
assign addr[8720]= -1599979481;
assign addr[8721]= -1493966902;
assign addr[8722]= -1380375881;
assign addr[8723]= -1259782632;
assign addr[8724]= -1132798888;
assign addr[8725]= -1000068799;
assign addr[8726]= -862265664;
assign addr[8727]= -720088517;
assign addr[8728]= -574258580;
assign addr[8729]= -425515602;
assign addr[8730]= -274614114;
assign addr[8731]= -122319591;
assign addr[8732]= 30595422;
assign addr[8733]= 183355234;
assign addr[8734]= 335184940;
assign addr[8735]= 485314355;
assign addr[8736]= 632981917;
assign addr[8737]= 777438554;
assign addr[8738]= 917951481;
assign addr[8739]= 1053807919;
assign addr[8740]= 1184318708;
assign addr[8741]= 1308821808;
assign addr[8742]= 1426685652;
assign addr[8743]= 1537312353;
assign addr[8744]= 1640140734;
assign addr[8745]= 1734649179;
assign addr[8746]= 1820358275;
assign addr[8747]= 1896833245;
assign addr[8748]= 1963686155;
assign addr[8749]= 2020577882;
assign addr[8750]= 2067219829;
assign addr[8751]= 2103375398;
assign addr[8752]= 2128861181;
assign addr[8753]= 2143547897;
assign addr[8754]= 2147361045;
assign addr[8755]= 2140281282;
assign addr[8756]= 2122344521;
assign addr[8757]= 2093641749;
assign addr[8758]= 2054318569;
assign addr[8759]= 2004574453;
assign addr[8760]= 1944661739;
assign addr[8761]= 1874884346;
assign addr[8762]= 1795596234;
assign addr[8763]= 1707199606;
assign addr[8764]= 1610142873;
assign addr[8765]= 1504918373;
assign addr[8766]= 1392059879;
assign addr[8767]= 1272139887;
assign addr[8768]= 1145766716;
assign addr[8769]= 1013581418;
assign addr[8770]= 876254528;
assign addr[8771]= 734482665;
assign addr[8772]= 588984994;
assign addr[8773]= 440499581;
assign addr[8774]= 289779648;
assign addr[8775]= 137589750;
assign addr[8776]= -15298099;
assign addr[8777]= -168108346;
assign addr[8778]= -320065829;
assign addr[8779]= -470399716;
assign addr[8780]= -618347408;
assign addr[8781]= -763158411;
assign addr[8782]= -904098143;
assign addr[8783]= -1040451659;
assign addr[8784]= -1171527280;
assign addr[8785]= -1296660098;
assign addr[8786]= -1415215352;
assign addr[8787]= -1526591649;
assign addr[8788]= -1630224009;
assign addr[8789]= -1725586737;
assign addr[8790]= -1812196087;
assign addr[8791]= -1889612716;
assign addr[8792]= -1957443913;
assign addr[8793]= -2015345591;
assign addr[8794]= -2063024031;
assign addr[8795]= -2100237377;
assign addr[8796]= -2126796855;
assign addr[8797]= -2142567738;
assign addr[8798]= -2147470025;
assign addr[8799]= -2141478848;
assign addr[8800]= -2124624598;
assign addr[8801]= -2096992772;
assign addr[8802]= -2058723538;
assign addr[8803]= -2010011024;
assign addr[8804]= -1951102334;
assign addr[8805]= -1882296293;
assign addr[8806]= -1803941934;
assign addr[8807]= -1716436725;
assign addr[8808]= -1620224553;
assign addr[8809]= -1515793473;
assign addr[8810]= -1403673233;
assign addr[8811]= -1284432584;
assign addr[8812]= -1158676398;
assign addr[8813]= -1027042599;
assign addr[8814]= -890198924;
assign addr[8815]= -748839539;
assign addr[8816]= -603681519;
assign addr[8817]= -455461206;
assign addr[8818]= -304930476;
assign addr[8819]= -152852926;
assign addr[8820]= 0;
assign addr[8821]= 152852926;
assign addr[8822]= 304930476;
assign addr[8823]= 455461206;
assign addr[8824]= 603681519;
assign addr[8825]= 748839539;
assign addr[8826]= 890198924;
assign addr[8827]= 1027042599;
assign addr[8828]= 1158676398;
assign addr[8829]= 1284432584;
assign addr[8830]= 1403673233;
assign addr[8831]= 1515793473;
assign addr[8832]= 1620224553;
assign addr[8833]= 1716436725;
assign addr[8834]= 1803941934;
assign addr[8835]= 1882296293;
assign addr[8836]= 1951102334;
assign addr[8837]= 2010011024;
assign addr[8838]= 2058723538;
assign addr[8839]= 2096992772;
assign addr[8840]= 2124624598;
assign addr[8841]= 2141478848;
assign addr[8842]= 2147470025;
assign addr[8843]= 2142567738;
assign addr[8844]= 2126796855;
assign addr[8845]= 2100237377;
assign addr[8846]= 2063024031;
assign addr[8847]= 2015345591;
assign addr[8848]= 1957443913;
assign addr[8849]= 1889612716;
assign addr[8850]= 1812196087;
assign addr[8851]= 1725586737;
assign addr[8852]= 1630224009;
assign addr[8853]= 1526591649;
assign addr[8854]= 1415215352;
assign addr[8855]= 1296660098;
assign addr[8856]= 1171527280;
assign addr[8857]= 1040451659;
assign addr[8858]= 904098143;
assign addr[8859]= 763158411;
assign addr[8860]= 618347408;
assign addr[8861]= 470399716;
assign addr[8862]= 320065829;
assign addr[8863]= 168108346;
assign addr[8864]= 15298099;
assign addr[8865]= -137589750;
assign addr[8866]= -289779648;
assign addr[8867]= -440499581;
assign addr[8868]= -588984994;
assign addr[8869]= -734482665;
assign addr[8870]= -876254528;
assign addr[8871]= -1013581418;
assign addr[8872]= -1145766716;
assign addr[8873]= -1272139887;
assign addr[8874]= -1392059879;
assign addr[8875]= -1504918373;
assign addr[8876]= -1610142873;
assign addr[8877]= -1707199606;
assign addr[8878]= -1795596234;
assign addr[8879]= -1874884346;
assign addr[8880]= -1944661739;
assign addr[8881]= -2004574453;
assign addr[8882]= -2054318569;
assign addr[8883]= -2093641749;
assign addr[8884]= -2122344521;
assign addr[8885]= -2140281282;
assign addr[8886]= -2147361045;
assign addr[8887]= -2143547897;
assign addr[8888]= -2128861181;
assign addr[8889]= -2103375398;
assign addr[8890]= -2067219829;
assign addr[8891]= -2020577882;
assign addr[8892]= -1963686155;
assign addr[8893]= -1896833245;
assign addr[8894]= -1820358275;
assign addr[8895]= -1734649179;
assign addr[8896]= -1640140734;
assign addr[8897]= -1537312353;
assign addr[8898]= -1426685652;
assign addr[8899]= -1308821808;
assign addr[8900]= -1184318708;
assign addr[8901]= -1053807919;
assign addr[8902]= -917951481;
assign addr[8903]= -777438554;
assign addr[8904]= -632981917;
assign addr[8905]= -485314355;
assign addr[8906]= -335184940;
assign addr[8907]= -183355234;
assign addr[8908]= -30595422;
assign addr[8909]= 122319591;
assign addr[8910]= 274614114;
assign addr[8911]= 425515602;
assign addr[8912]= 574258580;
assign addr[8913]= 720088517;
assign addr[8914]= 862265664;
assign addr[8915]= 1000068799;
assign addr[8916]= 1132798888;
assign addr[8917]= 1259782632;
assign addr[8918]= 1380375881;
assign addr[8919]= 1493966902;
assign addr[8920]= 1599979481;
assign addr[8921]= 1697875851;
assign addr[8922]= 1787159411;
assign addr[8923]= 1867377253;
assign addr[8924]= 1938122457;
assign addr[8925]= 1999036154;
assign addr[8926]= 2049809346;
assign addr[8927]= 2090184478;
assign addr[8928]= 2119956737;
assign addr[8929]= 2138975100;
assign addr[8930]= 2147143090;
assign addr[8931]= 2144419275;
assign addr[8932]= 2130817471;
assign addr[8933]= 2106406677;
assign addr[8934]= 2071310720;
assign addr[8935]= 2025707632;
assign addr[8936]= 1969828744;
assign addr[8937]= 1903957513;
assign addr[8938]= 1828428082;
assign addr[8939]= 1743623590;
assign addr[8940]= 1649974225;
assign addr[8941]= 1547955041;
assign addr[8942]= 1438083551;
assign addr[8943]= 1320917099;
assign addr[8944]= 1197050035;
assign addr[8945]= 1067110699;
assign addr[8946]= 931758235;
assign addr[8947]= 791679244;
assign addr[8948]= 647584304;
assign addr[8949]= 500204365;
assign addr[8950]= 350287041;
assign addr[8951]= 198592817;
assign addr[8952]= 45891193;
assign addr[8953]= -107043224;
assign addr[8954]= -259434643;
assign addr[8955]= -410510029;
assign addr[8956]= -559503022;
assign addr[8957]= -705657826;
assign addr[8958]= -848233042;
assign addr[8959]= -986505429;
assign addr[8960]= -1119773573;
assign addr[8961]= -1247361445;
assign addr[8962]= -1368621831;
assign addr[8963]= -1482939614;
assign addr[8964]= -1589734894;
assign addr[8965]= -1688465931;
assign addr[8966]= -1778631892;
assign addr[8967]= -1859775393;
assign addr[8968]= -1931484818;
assign addr[8969]= -1993396407;
assign addr[8970]= -2045196100;
assign addr[8971]= -2086621133;
assign addr[8972]= -2117461370;
assign addr[8973]= -2137560369;
assign addr[8974]= -2146816171;
assign addr[8975]= -2145181827;
assign addr[8976]= -2132665626;
assign addr[8977]= -2109331059;
assign addr[8978]= -2075296495;
assign addr[8979]= -2030734582;
assign addr[8980]= -1975871368;
assign addr[8981]= -1910985158;
assign addr[8982]= -1836405100;
assign addr[8983]= -1752509516;
assign addr[8984]= -1659723983;
assign addr[8985]= -1558519173;
assign addr[8986]= -1449408469;
assign addr[8987]= -1332945355;
assign addr[8988]= -1209720613;
assign addr[8989]= -1080359326;
assign addr[8990]= -945517704;
assign addr[8991]= -805879757;
assign addr[8992]= -662153826;
assign addr[8993]= -515068990;
assign addr[8994]= -365371365;
assign addr[8995]= -213820322;
assign addr[8996]= -61184634;
assign addr[8997]= 91761426;
assign addr[8998]= 244242007;
assign addr[8999]= 395483624;
assign addr[9000]= 544719071;
assign addr[9001]= 691191324;
assign addr[9002]= 834157373;
assign addr[9003]= 972891995;
assign addr[9004]= 1106691431;
assign addr[9005]= 1234876957;
assign addr[9006]= 1356798326;
assign addr[9007]= 1471837070;
assign addr[9008]= 1579409630;
assign addr[9009]= 1678970324;
assign addr[9010]= 1770014111;
assign addr[9011]= 1852079154;
assign addr[9012]= 1924749160;
assign addr[9013]= 1987655498;
assign addr[9014]= 2040479063;
assign addr[9015]= 2082951896;
assign addr[9016]= 2114858546;
assign addr[9017]= 2136037160;
assign addr[9018]= 2146380306;
assign addr[9019]= 2145835515;
assign addr[9020]= 2134405552;
assign addr[9021]= 2112148396;
assign addr[9022]= 2079176953;
assign addr[9023]= 2035658475;
assign addr[9024]= 1981813720;
assign addr[9025]= 1917915825;
assign addr[9026]= 1844288924;
assign addr[9027]= 1761306505;
assign addr[9028]= 1669389513;
assign addr[9029]= 1569004214;
assign addr[9030]= 1460659832;
assign addr[9031]= 1344905966;
assign addr[9032]= 1222329801;
assign addr[9033]= 1093553126;
assign addr[9034]= 959229189;
assign addr[9035]= 820039373;
assign addr[9036]= 676689746;
assign addr[9037]= 529907477;
assign addr[9038]= 380437148;
assign addr[9039]= 229036977;
assign addr[9040]= 76474970;
assign addr[9041]= -76474970;
assign addr[9042]= -229036977;
assign addr[9043]= -380437148;
assign addr[9044]= -529907477;
assign addr[9045]= -676689746;
assign addr[9046]= -820039373;
assign addr[9047]= -959229189;
assign addr[9048]= -1093553126;
assign addr[9049]= -1222329801;
assign addr[9050]= -1344905966;
assign addr[9051]= -1460659832;
assign addr[9052]= -1569004214;
assign addr[9053]= -1669389513;
assign addr[9054]= -1761306505;
assign addr[9055]= -1844288924;
assign addr[9056]= -1917915825;
assign addr[9057]= -1981813720;
assign addr[9058]= -2035658475;
assign addr[9059]= -2079176953;
assign addr[9060]= -2112148396;
assign addr[9061]= -2134405552;
assign addr[9062]= -2145835515;
assign addr[9063]= -2146380306;
assign addr[9064]= -2136037160;
assign addr[9065]= -2114858546;
assign addr[9066]= -2082951896;
assign addr[9067]= -2040479063;
assign addr[9068]= -1987655498;
assign addr[9069]= -1924749160;
assign addr[9070]= -1852079154;
assign addr[9071]= -1770014111;
assign addr[9072]= -1678970324;
assign addr[9073]= -1579409630;
assign addr[9074]= -1471837070;
assign addr[9075]= -1356798326;
assign addr[9076]= -1234876957;
assign addr[9077]= -1106691431;
assign addr[9078]= -972891995;
assign addr[9079]= -834157373;
assign addr[9080]= -691191324;
assign addr[9081]= -544719071;
assign addr[9082]= -395483624;
assign addr[9083]= -244242007;
assign addr[9084]= -91761426;
assign addr[9085]= 61184634;
assign addr[9086]= 213820322;
assign addr[9087]= 365371365;
assign addr[9088]= 515068990;
assign addr[9089]= 662153826;
assign addr[9090]= 805879757;
assign addr[9091]= 945517704;
assign addr[9092]= 1080359326;
assign addr[9093]= 1209720613;
assign addr[9094]= 1332945355;
assign addr[9095]= 1449408469;
assign addr[9096]= 1558519173;
assign addr[9097]= 1659723983;
assign addr[9098]= 1752509516;
assign addr[9099]= 1836405100;
assign addr[9100]= 1910985158;
assign addr[9101]= 1975871368;
assign addr[9102]= 2030734582;
assign addr[9103]= 2075296495;
assign addr[9104]= 2109331059;
assign addr[9105]= 2132665626;
assign addr[9106]= 2145181827;
assign addr[9107]= 2146816171;
assign addr[9108]= 2137560369;
assign addr[9109]= 2117461370;
assign addr[9110]= 2086621133;
assign addr[9111]= 2045196100;
assign addr[9112]= 1993396407;
assign addr[9113]= 1931484818;
assign addr[9114]= 1859775393;
assign addr[9115]= 1778631892;
assign addr[9116]= 1688465931;
assign addr[9117]= 1589734894;
assign addr[9118]= 1482939614;
assign addr[9119]= 1368621831;
assign addr[9120]= 1247361445;
assign addr[9121]= 1119773573;
assign addr[9122]= 986505429;
assign addr[9123]= 848233042;
assign addr[9124]= 705657826;
assign addr[9125]= 559503022;
assign addr[9126]= 410510029;
assign addr[9127]= 259434643;
assign addr[9128]= 107043224;
assign addr[9129]= -45891193;
assign addr[9130]= -198592817;
assign addr[9131]= -350287041;
assign addr[9132]= -500204365;
assign addr[9133]= -647584304;
assign addr[9134]= -791679244;
assign addr[9135]= -931758235;
assign addr[9136]= -1067110699;
assign addr[9137]= -1197050035;
assign addr[9138]= -1320917099;
assign addr[9139]= -1438083551;
assign addr[9140]= -1547955041;
assign addr[9141]= -1649974225;
assign addr[9142]= -1743623590;
assign addr[9143]= -1828428082;
assign addr[9144]= -1903957513;
assign addr[9145]= -1969828744;
assign addr[9146]= -2025707632;
assign addr[9147]= -2071310720;
assign addr[9148]= -2106406677;
assign addr[9149]= -2130817471;
assign addr[9150]= -2144419275;
assign addr[9151]= -2147143090;
assign addr[9152]= -2138975100;
assign addr[9153]= -2119956737;
assign addr[9154]= -2090184478;
assign addr[9155]= -2049809346;
assign addr[9156]= -1999036154;
assign addr[9157]= -1938122457;
assign addr[9158]= -1867377253;
assign addr[9159]= -1787159411;
assign addr[9160]= -1697875851;
assign addr[9161]= -1599979481;
assign addr[9162]= -1493966902;
assign addr[9163]= -1380375881;
assign addr[9164]= -1259782632;
assign addr[9165]= -1132798888;
assign addr[9166]= -1000068799;
assign addr[9167]= -862265664;
assign addr[9168]= -720088517;
assign addr[9169]= -574258580;
assign addr[9170]= -425515602;
assign addr[9171]= -274614114;
assign addr[9172]= -122319591;
assign addr[9173]= 30595422;
assign addr[9174]= 183355234;
assign addr[9175]= 335184940;
assign addr[9176]= 485314355;
assign addr[9177]= 632981917;
assign addr[9178]= 777438554;
assign addr[9179]= 917951481;
assign addr[9180]= 1053807919;
assign addr[9181]= 1184318708;
assign addr[9182]= 1308821808;
assign addr[9183]= 1426685652;
assign addr[9184]= 1537312353;
assign addr[9185]= 1640140734;
assign addr[9186]= 1734649179;
assign addr[9187]= 1820358275;
assign addr[9188]= 1896833245;
assign addr[9189]= 1963686155;
assign addr[9190]= 2020577882;
assign addr[9191]= 2067219829;
assign addr[9192]= 2103375398;
assign addr[9193]= 2128861181;
assign addr[9194]= 2143547897;
assign addr[9195]= 2147361045;
assign addr[9196]= 2140281282;
assign addr[9197]= 2122344521;
assign addr[9198]= 2093641749;
assign addr[9199]= 2054318569;
assign addr[9200]= 2004574453;
assign addr[9201]= 1944661739;
assign addr[9202]= 1874884346;
assign addr[9203]= 1795596234;
assign addr[9204]= 1707199606;
assign addr[9205]= 1610142873;
assign addr[9206]= 1504918373;
assign addr[9207]= 1392059879;
assign addr[9208]= 1272139887;
assign addr[9209]= 1145766716;
assign addr[9210]= 1013581418;
assign addr[9211]= 876254528;
assign addr[9212]= 734482665;
assign addr[9213]= 588984994;
assign addr[9214]= 440499581;
assign addr[9215]= 289779648;
assign addr[9216]= 137589750;
assign addr[9217]= -15298099;
assign addr[9218]= -168108346;
assign addr[9219]= -320065829;
assign addr[9220]= -470399716;
assign addr[9221]= -618347408;
assign addr[9222]= -763158411;
assign addr[9223]= -904098143;
assign addr[9224]= -1040451659;
assign addr[9225]= -1171527280;
assign addr[9226]= -1296660098;
assign addr[9227]= -1415215352;
assign addr[9228]= -1526591649;
assign addr[9229]= -1630224009;
assign addr[9230]= -1725586737;
assign addr[9231]= -1812196087;
assign addr[9232]= -1889612716;
assign addr[9233]= -1957443913;
assign addr[9234]= -2015345591;
assign addr[9235]= -2063024031;
assign addr[9236]= -2100237377;
assign addr[9237]= -2126796855;
assign addr[9238]= -2142567738;
assign addr[9239]= -2147470025;
assign addr[9240]= -2141478848;
assign addr[9241]= -2124624598;
assign addr[9242]= -2096992772;
assign addr[9243]= -2058723538;
assign addr[9244]= -2010011024;
assign addr[9245]= -1951102334;
assign addr[9246]= -1882296293;
assign addr[9247]= -1803941934;
assign addr[9248]= -1716436725;
assign addr[9249]= -1620224553;
assign addr[9250]= -1515793473;
assign addr[9251]= -1403673233;
assign addr[9252]= -1284432584;
assign addr[9253]= -1158676398;
assign addr[9254]= -1027042599;
assign addr[9255]= -890198924;
assign addr[9256]= -748839539;
assign addr[9257]= -603681519;
assign addr[9258]= -455461206;
assign addr[9259]= -304930476;
assign addr[9260]= -152852926;
assign addr[9261]= 0;
assign addr[9262]= 152852926;
assign addr[9263]= 304930476;
assign addr[9264]= 455461206;
assign addr[9265]= 603681519;
assign addr[9266]= 748839539;
assign addr[9267]= 890198924;
assign addr[9268]= 1027042599;
assign addr[9269]= 1158676398;
assign addr[9270]= 1284432584;
assign addr[9271]= 1403673233;
assign addr[9272]= 1515793473;
assign addr[9273]= 1620224553;
assign addr[9274]= 1716436725;
assign addr[9275]= 1803941934;
assign addr[9276]= 1882296293;
assign addr[9277]= 1951102334;
assign addr[9278]= 2010011024;
assign addr[9279]= 2058723538;
assign addr[9280]= 2096992772;
assign addr[9281]= 2124624598;
assign addr[9282]= 2141478848;
assign addr[9283]= 2147470025;
assign addr[9284]= 2142567738;
assign addr[9285]= 2126796855;
assign addr[9286]= 2100237377;
assign addr[9287]= 2063024031;
assign addr[9288]= 2015345591;
assign addr[9289]= 1957443913;
assign addr[9290]= 1889612716;
assign addr[9291]= 1812196087;
assign addr[9292]= 1725586737;
assign addr[9293]= 1630224009;
assign addr[9294]= 1526591649;
assign addr[9295]= 1415215352;
assign addr[9296]= 1296660098;
assign addr[9297]= 1171527280;
assign addr[9298]= 1040451659;
assign addr[9299]= 904098143;
assign addr[9300]= 763158411;
assign addr[9301]= 618347408;
assign addr[9302]= 470399716;
assign addr[9303]= 320065829;
assign addr[9304]= 168108346;
assign addr[9305]= 15298099;
assign addr[9306]= -137589750;
assign addr[9307]= -289779648;
assign addr[9308]= -440499581;
assign addr[9309]= -588984994;
assign addr[9310]= -734482665;
assign addr[9311]= -876254528;
assign addr[9312]= -1013581418;
assign addr[9313]= -1145766716;
assign addr[9314]= -1272139887;
assign addr[9315]= -1392059879;
assign addr[9316]= -1504918373;
assign addr[9317]= -1610142873;
assign addr[9318]= -1707199606;
assign addr[9319]= -1795596234;
assign addr[9320]= -1874884346;
assign addr[9321]= -1944661739;
assign addr[9322]= -2004574453;
assign addr[9323]= -2054318569;
assign addr[9324]= -2093641749;
assign addr[9325]= -2122344521;
assign addr[9326]= -2140281282;
assign addr[9327]= -2147361045;
assign addr[9328]= -2143547897;
assign addr[9329]= -2128861181;
assign addr[9330]= -2103375398;
assign addr[9331]= -2067219829;
assign addr[9332]= -2020577882;
assign addr[9333]= -1963686155;
assign addr[9334]= -1896833245;
assign addr[9335]= -1820358275;
assign addr[9336]= -1734649179;
assign addr[9337]= -1640140734;
assign addr[9338]= -1537312353;
assign addr[9339]= -1426685652;
assign addr[9340]= -1308821808;
assign addr[9341]= -1184318708;
assign addr[9342]= -1053807919;
assign addr[9343]= -917951481;
assign addr[9344]= -777438554;
assign addr[9345]= -632981917;
assign addr[9346]= -485314355;
assign addr[9347]= -335184940;
assign addr[9348]= -183355234;
assign addr[9349]= -30595422;
assign addr[9350]= 122319591;
assign addr[9351]= 274614114;
assign addr[9352]= 425515602;
assign addr[9353]= 574258580;
assign addr[9354]= 720088517;
assign addr[9355]= 862265664;
assign addr[9356]= 1000068799;
assign addr[9357]= 1132798888;
assign addr[9358]= 1259782632;
assign addr[9359]= 1380375881;
assign addr[9360]= 1493966902;
assign addr[9361]= 1599979481;
assign addr[9362]= 1697875851;
assign addr[9363]= 1787159411;
assign addr[9364]= 1867377253;
assign addr[9365]= 1938122457;
assign addr[9366]= 1999036154;
assign addr[9367]= 2049809346;
assign addr[9368]= 2090184478;
assign addr[9369]= 2119956737;
assign addr[9370]= 2138975100;
assign addr[9371]= 2147143090;
assign addr[9372]= 2144419275;
assign addr[9373]= 2130817471;
assign addr[9374]= 2106406677;
assign addr[9375]= 2071310720;
assign addr[9376]= 2025707632;
assign addr[9377]= 1969828744;
assign addr[9378]= 1903957513;
assign addr[9379]= 1828428082;
assign addr[9380]= 1743623590;
assign addr[9381]= 1649974225;
assign addr[9382]= 1547955041;
assign addr[9383]= 1438083551;
assign addr[9384]= 1320917099;
assign addr[9385]= 1197050035;
assign addr[9386]= 1067110699;
assign addr[9387]= 931758235;
assign addr[9388]= 791679244;
assign addr[9389]= 647584304;
assign addr[9390]= 500204365;
assign addr[9391]= 350287041;
assign addr[9392]= 198592817;
assign addr[9393]= 45891193;
assign addr[9394]= -107043224;
assign addr[9395]= -259434643;
assign addr[9396]= -410510029;
assign addr[9397]= -559503022;
assign addr[9398]= -705657826;
assign addr[9399]= -848233042;
assign addr[9400]= -986505429;
assign addr[9401]= -1119773573;
assign addr[9402]= -1247361445;
assign addr[9403]= -1368621831;
assign addr[9404]= -1482939614;
assign addr[9405]= -1589734894;
assign addr[9406]= -1688465931;
assign addr[9407]= -1778631892;
assign addr[9408]= -1859775393;
assign addr[9409]= -1931484818;
assign addr[9410]= -1993396407;
assign addr[9411]= -2045196100;
assign addr[9412]= -2086621133;
assign addr[9413]= -2117461370;
assign addr[9414]= -2137560369;
assign addr[9415]= -2146816171;
assign addr[9416]= -2145181827;
assign addr[9417]= -2132665626;
assign addr[9418]= -2109331059;
assign addr[9419]= -2075296495;
assign addr[9420]= -2030734582;
assign addr[9421]= -1975871368;
assign addr[9422]= -1910985158;
assign addr[9423]= -1836405100;
assign addr[9424]= -1752509516;
assign addr[9425]= -1659723983;
assign addr[9426]= -1558519173;
assign addr[9427]= -1449408469;
assign addr[9428]= -1332945355;
assign addr[9429]= -1209720613;
assign addr[9430]= -1080359326;
assign addr[9431]= -945517704;
assign addr[9432]= -805879757;
assign addr[9433]= -662153826;
assign addr[9434]= -515068990;
assign addr[9435]= -365371365;
assign addr[9436]= -213820322;
assign addr[9437]= -61184634;
assign addr[9438]= 91761426;
assign addr[9439]= 244242007;
assign addr[9440]= 395483624;
assign addr[9441]= 544719071;
assign addr[9442]= 691191324;
assign addr[9443]= 834157373;
assign addr[9444]= 972891995;
assign addr[9445]= 1106691431;
assign addr[9446]= 1234876957;
assign addr[9447]= 1356798326;
assign addr[9448]= 1471837070;
assign addr[9449]= 1579409630;
assign addr[9450]= 1678970324;
assign addr[9451]= 1770014111;
assign addr[9452]= 1852079154;
assign addr[9453]= 1924749160;
assign addr[9454]= 1987655498;
assign addr[9455]= 2040479063;
assign addr[9456]= 2082951896;
assign addr[9457]= 2114858546;
assign addr[9458]= 2136037160;
assign addr[9459]= 2146380306;
assign addr[9460]= 2145835515;
assign addr[9461]= 2134405552;
assign addr[9462]= 2112148396;
assign addr[9463]= 2079176953;
assign addr[9464]= 2035658475;
assign addr[9465]= 1981813720;
assign addr[9466]= 1917915825;
assign addr[9467]= 1844288924;
assign addr[9468]= 1761306505;
assign addr[9469]= 1669389513;
assign addr[9470]= 1569004214;
assign addr[9471]= 1460659832;
assign addr[9472]= 1344905966;
assign addr[9473]= 1222329801;
assign addr[9474]= 1093553126;
assign addr[9475]= 959229189;
assign addr[9476]= 820039373;
assign addr[9477]= 676689746;
assign addr[9478]= 529907477;
assign addr[9479]= 380437148;
assign addr[9480]= 229036977;
assign addr[9481]= 76474970;
assign addr[9482]= -76474970;
assign addr[9483]= -229036977;
assign addr[9484]= -380437148;
assign addr[9485]= -529907477;
assign addr[9486]= -676689746;
assign addr[9487]= -820039373;
assign addr[9488]= -959229189;
assign addr[9489]= -1093553126;
assign addr[9490]= -1222329801;
assign addr[9491]= -1344905966;
assign addr[9492]= -1460659832;
assign addr[9493]= -1569004214;
assign addr[9494]= -1669389513;
assign addr[9495]= -1761306505;
assign addr[9496]= -1844288924;
assign addr[9497]= -1917915825;
assign addr[9498]= -1981813720;
assign addr[9499]= -2035658475;
assign addr[9500]= -2079176953;
assign addr[9501]= -2112148396;
assign addr[9502]= -2134405552;
assign addr[9503]= -2145835515;
assign addr[9504]= -2146380306;
assign addr[9505]= -2136037160;
assign addr[9506]= -2114858546;
assign addr[9507]= -2082951896;
assign addr[9508]= -2040479063;
assign addr[9509]= -1987655498;
assign addr[9510]= -1924749160;
assign addr[9511]= -1852079154;
assign addr[9512]= -1770014111;
assign addr[9513]= -1678970324;
assign addr[9514]= -1579409630;
assign addr[9515]= -1471837070;
assign addr[9516]= -1356798326;
assign addr[9517]= -1234876957;
assign addr[9518]= -1106691431;
assign addr[9519]= -972891995;
assign addr[9520]= -834157373;
assign addr[9521]= -691191324;
assign addr[9522]= -544719071;
assign addr[9523]= -395483624;
assign addr[9524]= -244242007;
assign addr[9525]= -91761426;
assign addr[9526]= 61184634;
assign addr[9527]= 213820322;
assign addr[9528]= 365371365;
assign addr[9529]= 515068990;
assign addr[9530]= 662153826;
assign addr[9531]= 805879757;
assign addr[9532]= 945517704;
assign addr[9533]= 1080359326;
assign addr[9534]= 1209720613;
assign addr[9535]= 1332945355;
assign addr[9536]= 1449408469;
assign addr[9537]= 1558519173;
assign addr[9538]= 1659723983;
assign addr[9539]= 1752509516;
assign addr[9540]= 1836405100;
assign addr[9541]= 1910985158;
assign addr[9542]= 1975871368;
assign addr[9543]= 2030734582;
assign addr[9544]= 2075296495;
assign addr[9545]= 2109331059;
assign addr[9546]= 2132665626;
assign addr[9547]= 2145181827;
assign addr[9548]= 2146816171;
assign addr[9549]= 2137560369;
assign addr[9550]= 2117461370;
assign addr[9551]= 2086621133;
assign addr[9552]= 2045196100;
assign addr[9553]= 1993396407;
assign addr[9554]= 1931484818;
assign addr[9555]= 1859775393;
assign addr[9556]= 1778631892;
assign addr[9557]= 1688465931;
assign addr[9558]= 1589734894;
assign addr[9559]= 1482939614;
assign addr[9560]= 1368621831;
assign addr[9561]= 1247361445;
assign addr[9562]= 1119773573;
assign addr[9563]= 986505429;
assign addr[9564]= 848233042;
assign addr[9565]= 705657826;
assign addr[9566]= 559503022;
assign addr[9567]= 410510029;
assign addr[9568]= 259434643;
assign addr[9569]= 107043224;
assign addr[9570]= -45891193;
assign addr[9571]= -198592817;
assign addr[9572]= -350287041;
assign addr[9573]= -500204365;
assign addr[9574]= -647584304;
assign addr[9575]= -791679244;
assign addr[9576]= -931758235;
assign addr[9577]= -1067110699;
assign addr[9578]= -1197050035;
assign addr[9579]= -1320917099;
assign addr[9580]= -1438083551;
assign addr[9581]= -1547955041;
assign addr[9582]= -1649974225;
assign addr[9583]= -1743623590;
assign addr[9584]= -1828428082;
assign addr[9585]= -1903957513;
assign addr[9586]= -1969828744;
assign addr[9587]= -2025707632;
assign addr[9588]= -2071310720;
assign addr[9589]= -2106406677;
assign addr[9590]= -2130817471;
assign addr[9591]= -2144419275;
assign addr[9592]= -2147143090;
assign addr[9593]= -2138975100;
assign addr[9594]= -2119956737;
assign addr[9595]= -2090184478;
assign addr[9596]= -2049809346;
assign addr[9597]= -1999036154;
assign addr[9598]= -1938122457;
assign addr[9599]= -1867377253;
assign addr[9600]= -1787159411;
assign addr[9601]= -1697875851;
assign addr[9602]= -1599979481;
assign addr[9603]= -1493966902;
assign addr[9604]= -1380375881;
assign addr[9605]= -1259782632;
assign addr[9606]= -1132798888;
assign addr[9607]= -1000068799;
assign addr[9608]= -862265664;
assign addr[9609]= -720088517;
assign addr[9610]= -574258580;
assign addr[9611]= -425515602;
assign addr[9612]= -274614114;
assign addr[9613]= -122319591;
assign addr[9614]= 30595422;
assign addr[9615]= 183355234;
assign addr[9616]= 335184940;
assign addr[9617]= 485314355;
assign addr[9618]= 632981917;
assign addr[9619]= 777438554;
assign addr[9620]= 917951481;
assign addr[9621]= 1053807919;
assign addr[9622]= 1184318708;
assign addr[9623]= 1308821808;
assign addr[9624]= 1426685652;
assign addr[9625]= 1537312353;
assign addr[9626]= 1640140734;
assign addr[9627]= 1734649179;
assign addr[9628]= 1820358275;
assign addr[9629]= 1896833245;
assign addr[9630]= 1963686155;
assign addr[9631]= 2020577882;
assign addr[9632]= 2067219829;
assign addr[9633]= 2103375398;
assign addr[9634]= 2128861181;
assign addr[9635]= 2143547897;
assign addr[9636]= 2147361045;
assign addr[9637]= 2140281282;
assign addr[9638]= 2122344521;
assign addr[9639]= 2093641749;
assign addr[9640]= 2054318569;
assign addr[9641]= 2004574453;
assign addr[9642]= 1944661739;
assign addr[9643]= 1874884346;
assign addr[9644]= 1795596234;
assign addr[9645]= 1707199606;
assign addr[9646]= 1610142873;
assign addr[9647]= 1504918373;
assign addr[9648]= 1392059879;
assign addr[9649]= 1272139887;
assign addr[9650]= 1145766716;
assign addr[9651]= 1013581418;
assign addr[9652]= 876254528;
assign addr[9653]= 734482665;
assign addr[9654]= 588984994;
assign addr[9655]= 440499581;
assign addr[9656]= 289779648;
assign addr[9657]= 137589750;
assign addr[9658]= -15298099;
assign addr[9659]= -168108346;
assign addr[9660]= -320065829;
assign addr[9661]= -470399716;
assign addr[9662]= -618347408;
assign addr[9663]= -763158411;
assign addr[9664]= -904098143;
assign addr[9665]= -1040451659;
assign addr[9666]= -1171527280;
assign addr[9667]= -1296660098;
assign addr[9668]= -1415215352;
assign addr[9669]= -1526591649;
assign addr[9670]= -1630224009;
assign addr[9671]= -1725586737;
assign addr[9672]= -1812196087;
assign addr[9673]= -1889612716;
assign addr[9674]= -1957443913;
assign addr[9675]= -2015345591;
assign addr[9676]= -2063024031;
assign addr[9677]= -2100237377;
assign addr[9678]= -2126796855;
assign addr[9679]= -2142567738;
assign addr[9680]= -2147470025;
assign addr[9681]= -2141478848;
assign addr[9682]= -2124624598;
assign addr[9683]= -2096992772;
assign addr[9684]= -2058723538;
assign addr[9685]= -2010011024;
assign addr[9686]= -1951102334;
assign addr[9687]= -1882296293;
assign addr[9688]= -1803941934;
assign addr[9689]= -1716436725;
assign addr[9690]= -1620224553;
assign addr[9691]= -1515793473;
assign addr[9692]= -1403673233;
assign addr[9693]= -1284432584;
assign addr[9694]= -1158676398;
assign addr[9695]= -1027042599;
assign addr[9696]= -890198924;
assign addr[9697]= -748839539;
assign addr[9698]= -603681519;
assign addr[9699]= -455461206;
assign addr[9700]= -304930476;
assign addr[9701]= -152852926;
assign addr[9702]= 0;
assign addr[9703]= 152852926;
assign addr[9704]= 304930476;
assign addr[9705]= 455461206;
assign addr[9706]= 603681519;
assign addr[9707]= 748839539;
assign addr[9708]= 890198924;
assign addr[9709]= 1027042599;
assign addr[9710]= 1158676398;
assign addr[9711]= 1284432584;
assign addr[9712]= 1403673233;
assign addr[9713]= 1515793473;
assign addr[9714]= 1620224553;
assign addr[9715]= 1716436725;
assign addr[9716]= 1803941934;
assign addr[9717]= 1882296293;
assign addr[9718]= 1951102334;
assign addr[9719]= 2010011024;
assign addr[9720]= 2058723538;
assign addr[9721]= 2096992772;
assign addr[9722]= 2124624598;
assign addr[9723]= 2141478848;
assign addr[9724]= 2147470025;
assign addr[9725]= 2142567738;
assign addr[9726]= 2126796855;
assign addr[9727]= 2100237377;
assign addr[9728]= 2063024031;
assign addr[9729]= 2015345591;
assign addr[9730]= 1957443913;
assign addr[9731]= 1889612716;
assign addr[9732]= 1812196087;
assign addr[9733]= 1725586737;
assign addr[9734]= 1630224009;
assign addr[9735]= 1526591649;
assign addr[9736]= 1415215352;
assign addr[9737]= 1296660098;
assign addr[9738]= 1171527280;
assign addr[9739]= 1040451659;
assign addr[9740]= 904098143;
assign addr[9741]= 763158411;
assign addr[9742]= 618347408;
assign addr[9743]= 470399716;
assign addr[9744]= 320065829;
assign addr[9745]= 168108346;
assign addr[9746]= 15298099;
assign addr[9747]= -137589750;
assign addr[9748]= -289779648;
assign addr[9749]= -440499581;
assign addr[9750]= -588984994;
assign addr[9751]= -734482665;
assign addr[9752]= -876254528;
assign addr[9753]= -1013581418;
assign addr[9754]= -1145766716;
assign addr[9755]= -1272139887;
assign addr[9756]= -1392059879;
assign addr[9757]= -1504918373;
assign addr[9758]= -1610142873;
assign addr[9759]= -1707199606;
assign addr[9760]= -1795596234;
assign addr[9761]= -1874884346;
assign addr[9762]= -1944661739;
assign addr[9763]= -2004574453;
assign addr[9764]= -2054318569;
assign addr[9765]= -2093641749;
assign addr[9766]= -2122344521;
assign addr[9767]= -2140281282;
assign addr[9768]= -2147361045;
assign addr[9769]= -2143547897;
assign addr[9770]= -2128861181;
assign addr[9771]= -2103375398;
assign addr[9772]= -2067219829;
assign addr[9773]= -2020577882;
assign addr[9774]= -1963686155;
assign addr[9775]= -1896833245;
assign addr[9776]= -1820358275;
assign addr[9777]= -1734649179;
assign addr[9778]= -1640140734;
assign addr[9779]= -1537312353;
assign addr[9780]= -1426685652;
assign addr[9781]= -1308821808;
assign addr[9782]= -1184318708;
assign addr[9783]= -1053807919;
assign addr[9784]= -917951481;
assign addr[9785]= -777438554;
assign addr[9786]= -632981917;
assign addr[9787]= -485314355;
assign addr[9788]= -335184940;
assign addr[9789]= -183355234;
assign addr[9790]= -30595422;
assign addr[9791]= 122319591;
assign addr[9792]= 274614114;
assign addr[9793]= 425515602;
assign addr[9794]= 574258580;
assign addr[9795]= 720088517;
assign addr[9796]= 862265664;
assign addr[9797]= 1000068799;
assign addr[9798]= 1132798888;
assign addr[9799]= 1259782632;
assign addr[9800]= 1380375881;
assign addr[9801]= 1493966902;
assign addr[9802]= 1599979481;
assign addr[9803]= 1697875851;
assign addr[9804]= 1787159411;
assign addr[9805]= 1867377253;
assign addr[9806]= 1938122457;
assign addr[9807]= 1999036154;
assign addr[9808]= 2049809346;
assign addr[9809]= 2090184478;
assign addr[9810]= 2119956737;
assign addr[9811]= 2138975100;
assign addr[9812]= 2147143090;
assign addr[9813]= 2144419275;
assign addr[9814]= 2130817471;
assign addr[9815]= 2106406677;
assign addr[9816]= 2071310720;
assign addr[9817]= 2025707632;
assign addr[9818]= 1969828744;
assign addr[9819]= 1903957513;
assign addr[9820]= 1828428082;
assign addr[9821]= 1743623590;
assign addr[9822]= 1649974225;
assign addr[9823]= 1547955041;
assign addr[9824]= 1438083551;
assign addr[9825]= 1320917099;
assign addr[9826]= 1197050035;
assign addr[9827]= 1067110699;
assign addr[9828]= 931758235;
assign addr[9829]= 791679244;
assign addr[9830]= 647584304;
assign addr[9831]= 500204365;
assign addr[9832]= 350287041;
assign addr[9833]= 198592817;
assign addr[9834]= 45891193;
assign addr[9835]= -107043224;
assign addr[9836]= -259434643;
assign addr[9837]= -410510029;
assign addr[9838]= -559503022;
assign addr[9839]= -705657826;
assign addr[9840]= -848233042;
assign addr[9841]= -986505429;
assign addr[9842]= -1119773573;
assign addr[9843]= -1247361445;
assign addr[9844]= -1368621831;
assign addr[9845]= -1482939614;
assign addr[9846]= -1589734894;
assign addr[9847]= -1688465931;
assign addr[9848]= -1778631892;
assign addr[9849]= -1859775393;
assign addr[9850]= -1931484818;
assign addr[9851]= -1993396407;
assign addr[9852]= -2045196100;
assign addr[9853]= -2086621133;
assign addr[9854]= -2117461370;
assign addr[9855]= -2137560369;
assign addr[9856]= -2146816171;
assign addr[9857]= -2145181827;
assign addr[9858]= -2132665626;
assign addr[9859]= -2109331059;
assign addr[9860]= -2075296495;
assign addr[9861]= -2030734582;
assign addr[9862]= -1975871368;
assign addr[9863]= -1910985158;
assign addr[9864]= -1836405100;
assign addr[9865]= -1752509516;
assign addr[9866]= -1659723983;
assign addr[9867]= -1558519173;
assign addr[9868]= -1449408469;
assign addr[9869]= -1332945355;
assign addr[9870]= -1209720613;
assign addr[9871]= -1080359326;
assign addr[9872]= -945517704;
assign addr[9873]= -805879757;
assign addr[9874]= -662153826;
assign addr[9875]= -515068990;
assign addr[9876]= -365371365;
assign addr[9877]= -213820322;
assign addr[9878]= -61184634;
assign addr[9879]= 91761426;
assign addr[9880]= 244242007;
assign addr[9881]= 395483624;
assign addr[9882]= 544719071;
assign addr[9883]= 691191324;
assign addr[9884]= 834157373;
assign addr[9885]= 972891995;
assign addr[9886]= 1106691431;
assign addr[9887]= 1234876957;
assign addr[9888]= 1356798326;
assign addr[9889]= 1471837070;
assign addr[9890]= 1579409630;
assign addr[9891]= 1678970324;
assign addr[9892]= 1770014111;
assign addr[9893]= 1852079154;
assign addr[9894]= 1924749160;
assign addr[9895]= 1987655498;
assign addr[9896]= 2040479063;
assign addr[9897]= 2082951896;
assign addr[9898]= 2114858546;
assign addr[9899]= 2136037160;
assign addr[9900]= 2146380306;
assign addr[9901]= 2145835515;
assign addr[9902]= 2134405552;
assign addr[9903]= 2112148396;
assign addr[9904]= 2079176953;
assign addr[9905]= 2035658475;
assign addr[9906]= 1981813720;
assign addr[9907]= 1917915825;
assign addr[9908]= 1844288924;
assign addr[9909]= 1761306505;
assign addr[9910]= 1669389513;
assign addr[9911]= 1569004214;
assign addr[9912]= 1460659832;
assign addr[9913]= 1344905966;
assign addr[9914]= 1222329801;
assign addr[9915]= 1093553126;
assign addr[9916]= 959229189;
assign addr[9917]= 820039373;
assign addr[9918]= 676689746;
assign addr[9919]= 529907477;
assign addr[9920]= 380437148;
assign addr[9921]= 229036977;
assign addr[9922]= 76474970;
assign addr[9923]= -76474970;
assign addr[9924]= -229036977;
assign addr[9925]= -380437148;
assign addr[9926]= -529907477;
assign addr[9927]= -676689746;
assign addr[9928]= -820039373;
assign addr[9929]= -959229189;
assign addr[9930]= -1093553126;
assign addr[9931]= -1222329801;
assign addr[9932]= -1344905966;
assign addr[9933]= -1460659832;
assign addr[9934]= -1569004214;
assign addr[9935]= -1669389513;
assign addr[9936]= -1761306505;
assign addr[9937]= -1844288924;
assign addr[9938]= -1917915825;
assign addr[9939]= -1981813720;
assign addr[9940]= -2035658475;
assign addr[9941]= -2079176953;
assign addr[9942]= -2112148396;
assign addr[9943]= -2134405552;
assign addr[9944]= -2145835515;
assign addr[9945]= -2146380306;
assign addr[9946]= -2136037160;
assign addr[9947]= -2114858546;
assign addr[9948]= -2082951896;
assign addr[9949]= -2040479063;
assign addr[9950]= -1987655498;
assign addr[9951]= -1924749160;
assign addr[9952]= -1852079154;
assign addr[9953]= -1770014111;
assign addr[9954]= -1678970324;
assign addr[9955]= -1579409630;
assign addr[9956]= -1471837070;
assign addr[9957]= -1356798326;
assign addr[9958]= -1234876957;
assign addr[9959]= -1106691431;
assign addr[9960]= -972891995;
assign addr[9961]= -834157373;
assign addr[9962]= -691191324;
assign addr[9963]= -544719071;
assign addr[9964]= -395483624;
assign addr[9965]= -244242007;
assign addr[9966]= -91761426;
assign addr[9967]= 61184634;
assign addr[9968]= 213820322;
assign addr[9969]= 365371365;
assign addr[9970]= 515068990;
assign addr[9971]= 662153826;
assign addr[9972]= 805879757;
assign addr[9973]= 945517704;
assign addr[9974]= 1080359326;
assign addr[9975]= 1209720613;
assign addr[9976]= 1332945355;
assign addr[9977]= 1449408469;
assign addr[9978]= 1558519173;
assign addr[9979]= 1659723983;
assign addr[9980]= 1752509516;
assign addr[9981]= 1836405100;
assign addr[9982]= 1910985158;
assign addr[9983]= 1975871368;
assign addr[9984]= 2030734582;
assign addr[9985]= 2075296495;
assign addr[9986]= 2109331059;
assign addr[9987]= 2132665626;
assign addr[9988]= 2145181827;
assign addr[9989]= 2146816171;
assign addr[9990]= 2137560369;
assign addr[9991]= 2117461370;
assign addr[9992]= 2086621133;
assign addr[9993]= 2045196100;
assign addr[9994]= 1993396407;
assign addr[9995]= 1931484818;
assign addr[9996]= 1859775393;
assign addr[9997]= 1778631892;
assign addr[9998]= 1688465931;
assign addr[9999]= 1589734894;
assign addr[10000]= 1482939614;
assign addr[10001]= 1368621831;
assign addr[10002]= 1247361445;
assign addr[10003]= 1119773573;
assign addr[10004]= 986505429;
assign addr[10005]= 848233042;
assign addr[10006]= 705657826;
assign addr[10007]= 559503022;
assign addr[10008]= 410510029;
assign addr[10009]= 259434643;
assign addr[10010]= 107043224;
assign addr[10011]= -45891193;
assign addr[10012]= -198592817;
assign addr[10013]= -350287041;
assign addr[10014]= -500204365;
assign addr[10015]= -647584304;
assign addr[10016]= -791679244;
assign addr[10017]= -931758235;
assign addr[10018]= -1067110699;
assign addr[10019]= -1197050035;
assign addr[10020]= -1320917099;
assign addr[10021]= -1438083551;
assign addr[10022]= -1547955041;
assign addr[10023]= -1649974225;
assign addr[10024]= -1743623590;
assign addr[10025]= -1828428082;
assign addr[10026]= -1903957513;
assign addr[10027]= -1969828744;
assign addr[10028]= -2025707632;
assign addr[10029]= -2071310720;
assign addr[10030]= -2106406677;
assign addr[10031]= -2130817471;
assign addr[10032]= -2144419275;
assign addr[10033]= -2147143090;
assign addr[10034]= -2138975100;
assign addr[10035]= -2119956737;
assign addr[10036]= -2090184478;
assign addr[10037]= -2049809346;
assign addr[10038]= -1999036154;
assign addr[10039]= -1938122457;
assign addr[10040]= -1867377253;
assign addr[10041]= -1787159411;
assign addr[10042]= -1697875851;
assign addr[10043]= -1599979481;
assign addr[10044]= -1493966902;
assign addr[10045]= -1380375881;
assign addr[10046]= -1259782632;
assign addr[10047]= -1132798888;
assign addr[10048]= -1000068799;
assign addr[10049]= -862265664;
assign addr[10050]= -720088517;
assign addr[10051]= -574258580;
assign addr[10052]= -425515602;
assign addr[10053]= -274614114;
assign addr[10054]= -122319591;
assign addr[10055]= 30595422;
assign addr[10056]= 183355234;
assign addr[10057]= 335184940;
assign addr[10058]= 485314355;
assign addr[10059]= 632981917;
assign addr[10060]= 777438554;
assign addr[10061]= 917951481;
assign addr[10062]= 1053807919;
assign addr[10063]= 1184318708;
assign addr[10064]= 1308821808;
assign addr[10065]= 1426685652;
assign addr[10066]= 1537312353;
assign addr[10067]= 1640140734;
assign addr[10068]= 1734649179;
assign addr[10069]= 1820358275;
assign addr[10070]= 1896833245;
assign addr[10071]= 1963686155;
assign addr[10072]= 2020577882;
assign addr[10073]= 2067219829;
assign addr[10074]= 2103375398;
assign addr[10075]= 2128861181;
assign addr[10076]= 2143547897;
assign addr[10077]= 2147361045;
assign addr[10078]= 2140281282;
assign addr[10079]= 2122344521;
assign addr[10080]= 2093641749;
assign addr[10081]= 2054318569;
assign addr[10082]= 2004574453;
assign addr[10083]= 1944661739;
assign addr[10084]= 1874884346;
assign addr[10085]= 1795596234;
assign addr[10086]= 1707199606;
assign addr[10087]= 1610142873;
assign addr[10088]= 1504918373;
assign addr[10089]= 1392059879;
assign addr[10090]= 1272139887;
assign addr[10091]= 1145766716;
assign addr[10092]= 1013581418;
assign addr[10093]= 876254528;
assign addr[10094]= 734482665;
assign addr[10095]= 588984994;
assign addr[10096]= 440499581;
assign addr[10097]= 289779648;
assign addr[10098]= 137589750;
assign addr[10099]= -15298099;
assign addr[10100]= -168108346;
assign addr[10101]= -320065829;
assign addr[10102]= -470399716;
assign addr[10103]= -618347408;
assign addr[10104]= -763158411;
assign addr[10105]= -904098143;
assign addr[10106]= -1040451659;
assign addr[10107]= -1171527280;
assign addr[10108]= -1296660098;
assign addr[10109]= -1415215352;
assign addr[10110]= -1526591649;
assign addr[10111]= -1630224009;
assign addr[10112]= -1725586737;
assign addr[10113]= -1812196087;
assign addr[10114]= -1889612716;
assign addr[10115]= -1957443913;
assign addr[10116]= -2015345591;
assign addr[10117]= -2063024031;
assign addr[10118]= -2100237377;
assign addr[10119]= -2126796855;
assign addr[10120]= -2142567738;
assign addr[10121]= -2147470025;
assign addr[10122]= -2141478848;
assign addr[10123]= -2124624598;
assign addr[10124]= -2096992772;
assign addr[10125]= -2058723538;
assign addr[10126]= -2010011024;
assign addr[10127]= -1951102334;
assign addr[10128]= -1882296293;
assign addr[10129]= -1803941934;
assign addr[10130]= -1716436725;
assign addr[10131]= -1620224553;
assign addr[10132]= -1515793473;
assign addr[10133]= -1403673233;
assign addr[10134]= -1284432584;
assign addr[10135]= -1158676398;
assign addr[10136]= -1027042599;
assign addr[10137]= -890198924;
assign addr[10138]= -748839539;
assign addr[10139]= -603681519;
assign addr[10140]= -455461206;
assign addr[10141]= -304930476;
assign addr[10142]= -152852926;
assign addr[10143]= 0;
assign addr[10144]= 152852926;
assign addr[10145]= 304930476;
assign addr[10146]= 455461206;
assign addr[10147]= 603681519;
assign addr[10148]= 748839539;
assign addr[10149]= 890198924;
assign addr[10150]= 1027042599;
assign addr[10151]= 1158676398;
assign addr[10152]= 1284432584;
assign addr[10153]= 1403673233;
assign addr[10154]= 1515793473;
assign addr[10155]= 1620224553;
assign addr[10156]= 1716436725;
assign addr[10157]= 1803941934;
assign addr[10158]= 1882296293;
assign addr[10159]= 1951102334;
assign addr[10160]= 2010011024;
assign addr[10161]= 2058723538;
assign addr[10162]= 2096992772;
assign addr[10163]= 2124624598;
assign addr[10164]= 2141478848;
assign addr[10165]= 2147470025;
assign addr[10166]= 2142567738;
assign addr[10167]= 2126796855;
assign addr[10168]= 2100237377;
assign addr[10169]= 2063024031;
assign addr[10170]= 2015345591;
assign addr[10171]= 1957443913;
assign addr[10172]= 1889612716;
assign addr[10173]= 1812196087;
assign addr[10174]= 1725586737;
assign addr[10175]= 1630224009;
assign addr[10176]= 1526591649;
assign addr[10177]= 1415215352;
assign addr[10178]= 1296660098;
assign addr[10179]= 1171527280;
assign addr[10180]= 1040451659;
assign addr[10181]= 904098143;
assign addr[10182]= 763158411;
assign addr[10183]= 618347408;
assign addr[10184]= 470399716;
assign addr[10185]= 320065829;
assign addr[10186]= 168108346;
assign addr[10187]= 15298099;
assign addr[10188]= -137589750;
assign addr[10189]= -289779648;
assign addr[10190]= -440499581;
assign addr[10191]= -588984994;
assign addr[10192]= -734482665;
assign addr[10193]= -876254528;
assign addr[10194]= -1013581418;
assign addr[10195]= -1145766716;
assign addr[10196]= -1272139887;
assign addr[10197]= -1392059879;
assign addr[10198]= -1504918373;
assign addr[10199]= -1610142873;
assign addr[10200]= -1707199606;
assign addr[10201]= -1795596234;
assign addr[10202]= -1874884346;
assign addr[10203]= -1944661739;
assign addr[10204]= -2004574453;
assign addr[10205]= -2054318569;
assign addr[10206]= -2093641749;
assign addr[10207]= -2122344521;
assign addr[10208]= -2140281282;
assign addr[10209]= -2147361045;
assign addr[10210]= -2143547897;
assign addr[10211]= -2128861181;
assign addr[10212]= -2103375398;
assign addr[10213]= -2067219829;
assign addr[10214]= -2020577882;
assign addr[10215]= -1963686155;
assign addr[10216]= -1896833245;
assign addr[10217]= -1820358275;
assign addr[10218]= -1734649179;
assign addr[10219]= -1640140734;
assign addr[10220]= -1537312353;
assign addr[10221]= -1426685652;
assign addr[10222]= -1308821808;
assign addr[10223]= -1184318708;
assign addr[10224]= -1053807919;
assign addr[10225]= -917951481;
assign addr[10226]= -777438554;
assign addr[10227]= -632981917;
assign addr[10228]= -485314355;
assign addr[10229]= -335184940;
assign addr[10230]= -183355234;
assign addr[10231]= -30595422;
assign addr[10232]= 122319591;
assign addr[10233]= 274614114;
assign addr[10234]= 425515602;
assign addr[10235]= 574258580;
assign addr[10236]= 720088517;
assign addr[10237]= 862265664;
assign addr[10238]= 1000068799;
assign addr[10239]= 1132798888;
assign addr[10240]= 1259782632;
assign addr[10241]= 1380375881;
assign addr[10242]= 1493966902;
assign addr[10243]= 1599979481;
assign addr[10244]= 1697875851;
assign addr[10245]= 1787159411;
assign addr[10246]= 1867377253;
assign addr[10247]= 1938122457;
assign addr[10248]= 1999036154;
assign addr[10249]= 2049809346;
assign addr[10250]= 2090184478;
assign addr[10251]= 2119956737;
assign addr[10252]= 2138975100;
assign addr[10253]= 2147143090;
assign addr[10254]= 2144419275;
assign addr[10255]= 2130817471;
assign addr[10256]= 2106406677;
assign addr[10257]= 2071310720;
assign addr[10258]= 2025707632;
assign addr[10259]= 1969828744;
assign addr[10260]= 1903957513;
assign addr[10261]= 1828428082;
assign addr[10262]= 1743623590;
assign addr[10263]= 1649974225;
assign addr[10264]= 1547955041;
assign addr[10265]= 1438083551;
assign addr[10266]= 1320917099;
assign addr[10267]= 1197050035;
assign addr[10268]= 1067110699;
assign addr[10269]= 931758235;
assign addr[10270]= 791679244;
assign addr[10271]= 647584304;
assign addr[10272]= 500204365;
assign addr[10273]= 350287041;
assign addr[10274]= 198592817;
assign addr[10275]= 45891193;
assign addr[10276]= -107043224;
assign addr[10277]= -259434643;
assign addr[10278]= -410510029;
assign addr[10279]= -559503022;
assign addr[10280]= -705657826;
assign addr[10281]= -848233042;
assign addr[10282]= -986505429;
assign addr[10283]= -1119773573;
assign addr[10284]= -1247361445;
assign addr[10285]= -1368621831;
assign addr[10286]= -1482939614;
assign addr[10287]= -1589734894;
assign addr[10288]= -1688465931;
assign addr[10289]= -1778631892;
assign addr[10290]= -1859775393;
assign addr[10291]= -1931484818;
assign addr[10292]= -1993396407;
assign addr[10293]= -2045196100;
assign addr[10294]= -2086621133;
assign addr[10295]= -2117461370;
assign addr[10296]= -2137560369;
assign addr[10297]= -2146816171;
assign addr[10298]= -2145181827;
assign addr[10299]= -2132665626;
assign addr[10300]= -2109331059;
assign addr[10301]= -2075296495;
assign addr[10302]= -2030734582;
assign addr[10303]= -1975871368;
assign addr[10304]= -1910985158;
assign addr[10305]= -1836405100;
assign addr[10306]= -1752509516;
assign addr[10307]= -1659723983;
assign addr[10308]= -1558519173;
assign addr[10309]= -1449408469;
assign addr[10310]= -1332945355;
assign addr[10311]= -1209720613;
assign addr[10312]= -1080359326;
assign addr[10313]= -945517704;
assign addr[10314]= -805879757;
assign addr[10315]= -662153826;
assign addr[10316]= -515068990;
assign addr[10317]= -365371365;
assign addr[10318]= -213820322;
assign addr[10319]= -61184634;
assign addr[10320]= 91761426;
assign addr[10321]= 244242007;
assign addr[10322]= 395483624;
assign addr[10323]= 544719071;
assign addr[10324]= 691191324;
assign addr[10325]= 834157373;
assign addr[10326]= 972891995;
assign addr[10327]= 1106691431;
assign addr[10328]= 1234876957;
assign addr[10329]= 1356798326;
assign addr[10330]= 1471837070;
assign addr[10331]= 1579409630;
assign addr[10332]= 1678970324;
assign addr[10333]= 1770014111;
assign addr[10334]= 1852079154;
assign addr[10335]= 1924749160;
assign addr[10336]= 1987655498;
assign addr[10337]= 2040479063;
assign addr[10338]= 2082951896;
assign addr[10339]= 2114858546;
assign addr[10340]= 2136037160;
assign addr[10341]= 2146380306;
assign addr[10342]= 2145835515;
assign addr[10343]= 2134405552;
assign addr[10344]= 2112148396;
assign addr[10345]= 2079176953;
assign addr[10346]= 2035658475;
assign addr[10347]= 1981813720;
assign addr[10348]= 1917915825;
assign addr[10349]= 1844288924;
assign addr[10350]= 1761306505;
assign addr[10351]= 1669389513;
assign addr[10352]= 1569004214;
assign addr[10353]= 1460659832;
assign addr[10354]= 1344905966;
assign addr[10355]= 1222329801;
assign addr[10356]= 1093553126;
assign addr[10357]= 959229189;
assign addr[10358]= 820039373;
assign addr[10359]= 676689746;
assign addr[10360]= 529907477;
assign addr[10361]= 380437148;
assign addr[10362]= 229036977;
assign addr[10363]= 76474970;
assign addr[10364]= -76474970;
assign addr[10365]= -229036977;
assign addr[10366]= -380437148;
assign addr[10367]= -529907477;
assign addr[10368]= -676689746;
assign addr[10369]= -820039373;
assign addr[10370]= -959229189;
assign addr[10371]= -1093553126;
assign addr[10372]= -1222329801;
assign addr[10373]= -1344905966;
assign addr[10374]= -1460659832;
assign addr[10375]= -1569004214;
assign addr[10376]= -1669389513;
assign addr[10377]= -1761306505;
assign addr[10378]= -1844288924;
assign addr[10379]= -1917915825;
assign addr[10380]= -1981813720;
assign addr[10381]= -2035658475;
assign addr[10382]= -2079176953;
assign addr[10383]= -2112148396;
assign addr[10384]= -2134405552;
assign addr[10385]= -2145835515;
assign addr[10386]= -2146380306;
assign addr[10387]= -2136037160;
assign addr[10388]= -2114858546;
assign addr[10389]= -2082951896;
assign addr[10390]= -2040479063;
assign addr[10391]= -1987655498;
assign addr[10392]= -1924749160;
assign addr[10393]= -1852079154;
assign addr[10394]= -1770014111;
assign addr[10395]= -1678970324;
assign addr[10396]= -1579409630;
assign addr[10397]= -1471837070;
assign addr[10398]= -1356798326;
assign addr[10399]= -1234876957;
assign addr[10400]= -1106691431;
assign addr[10401]= -972891995;
assign addr[10402]= -834157373;
assign addr[10403]= -691191324;
assign addr[10404]= -544719071;
assign addr[10405]= -395483624;
assign addr[10406]= -244242007;
assign addr[10407]= -91761426;
assign addr[10408]= 61184634;
assign addr[10409]= 213820322;
assign addr[10410]= 365371365;
assign addr[10411]= 515068990;
assign addr[10412]= 662153826;
assign addr[10413]= 805879757;
assign addr[10414]= 945517704;
assign addr[10415]= 1080359326;
assign addr[10416]= 1209720613;
assign addr[10417]= 1332945355;
assign addr[10418]= 1449408469;
assign addr[10419]= 1558519173;
assign addr[10420]= 1659723983;
assign addr[10421]= 1752509516;
assign addr[10422]= 1836405100;
assign addr[10423]= 1910985158;
assign addr[10424]= 1975871368;
assign addr[10425]= 2030734582;
assign addr[10426]= 2075296495;
assign addr[10427]= 2109331059;
assign addr[10428]= 2132665626;
assign addr[10429]= 2145181827;
assign addr[10430]= 2146816171;
assign addr[10431]= 2137560369;
assign addr[10432]= 2117461370;
assign addr[10433]= 2086621133;
assign addr[10434]= 2045196100;
assign addr[10435]= 1993396407;
assign addr[10436]= 1931484818;
assign addr[10437]= 1859775393;
assign addr[10438]= 1778631892;
assign addr[10439]= 1688465931;
assign addr[10440]= 1589734894;
assign addr[10441]= 1482939614;
assign addr[10442]= 1368621831;
assign addr[10443]= 1247361445;
assign addr[10444]= 1119773573;
assign addr[10445]= 986505429;
assign addr[10446]= 848233042;
assign addr[10447]= 705657826;
assign addr[10448]= 559503022;
assign addr[10449]= 410510029;
assign addr[10450]= 259434643;
assign addr[10451]= 107043224;
assign addr[10452]= -45891193;
assign addr[10453]= -198592817;
assign addr[10454]= -350287041;
assign addr[10455]= -500204365;
assign addr[10456]= -647584304;
assign addr[10457]= -791679244;
assign addr[10458]= -931758235;
assign addr[10459]= -1067110699;
assign addr[10460]= -1197050035;
assign addr[10461]= -1320917099;
assign addr[10462]= -1438083551;
assign addr[10463]= -1547955041;
assign addr[10464]= -1649974225;
assign addr[10465]= -1743623590;
assign addr[10466]= -1828428082;
assign addr[10467]= -1903957513;
assign addr[10468]= -1969828744;
assign addr[10469]= -2025707632;
assign addr[10470]= -2071310720;
assign addr[10471]= -2106406677;
assign addr[10472]= -2130817471;
assign addr[10473]= -2144419275;
assign addr[10474]= -2147143090;
assign addr[10475]= -2138975100;
assign addr[10476]= -2119956737;
assign addr[10477]= -2090184478;
assign addr[10478]= -2049809346;
assign addr[10479]= -1999036154;
assign addr[10480]= -1938122457;
assign addr[10481]= -1867377253;
assign addr[10482]= -1787159411;
assign addr[10483]= -1697875851;
assign addr[10484]= -1599979481;
assign addr[10485]= -1493966902;
assign addr[10486]= -1380375881;
assign addr[10487]= -1259782632;
assign addr[10488]= -1132798888;
assign addr[10489]= -1000068799;
assign addr[10490]= -862265664;
assign addr[10491]= -720088517;
assign addr[10492]= -574258580;
assign addr[10493]= -425515602;
assign addr[10494]= -274614114;
assign addr[10495]= -122319591;
assign addr[10496]= 30595422;
assign addr[10497]= 183355234;
assign addr[10498]= 335184940;
assign addr[10499]= 485314355;
assign addr[10500]= 632981917;
assign addr[10501]= 777438554;
assign addr[10502]= 917951481;
assign addr[10503]= 1053807919;
assign addr[10504]= 1184318708;
assign addr[10505]= 1308821808;
assign addr[10506]= 1426685652;
assign addr[10507]= 1537312353;
assign addr[10508]= 1640140734;
assign addr[10509]= 1734649179;
assign addr[10510]= 1820358275;
assign addr[10511]= 1896833245;
assign addr[10512]= 1963686155;
assign addr[10513]= 2020577882;
assign addr[10514]= 2067219829;
assign addr[10515]= 2103375398;
assign addr[10516]= 2128861181;
assign addr[10517]= 2143547897;
assign addr[10518]= 2147361045;
assign addr[10519]= 2140281282;
assign addr[10520]= 2122344521;
assign addr[10521]= 2093641749;
assign addr[10522]= 2054318569;
assign addr[10523]= 2004574453;
assign addr[10524]= 1944661739;
assign addr[10525]= 1874884346;
assign addr[10526]= 1795596234;
assign addr[10527]= 1707199606;
assign addr[10528]= 1610142873;
assign addr[10529]= 1504918373;
assign addr[10530]= 1392059879;
assign addr[10531]= 1272139887;
assign addr[10532]= 1145766716;
assign addr[10533]= 1013581418;
assign addr[10534]= 876254528;
assign addr[10535]= 734482665;
assign addr[10536]= 588984994;
assign addr[10537]= 440499581;
assign addr[10538]= 289779648;
assign addr[10539]= 137589750;
assign addr[10540]= -15298099;
assign addr[10541]= -168108346;
assign addr[10542]= -320065829;
assign addr[10543]= -470399716;
assign addr[10544]= -618347408;
assign addr[10545]= -763158411;
assign addr[10546]= -904098143;
assign addr[10547]= -1040451659;
assign addr[10548]= -1171527280;
assign addr[10549]= -1296660098;
assign addr[10550]= -1415215352;
assign addr[10551]= -1526591649;
assign addr[10552]= -1630224009;
assign addr[10553]= -1725586737;
assign addr[10554]= -1812196087;
assign addr[10555]= -1889612716;
assign addr[10556]= -1957443913;
assign addr[10557]= -2015345591;
assign addr[10558]= -2063024031;
assign addr[10559]= -2100237377;
assign addr[10560]= -2126796855;
assign addr[10561]= -2142567738;
assign addr[10562]= -2147470025;
assign addr[10563]= -2141478848;
assign addr[10564]= -2124624598;
assign addr[10565]= -2096992772;
assign addr[10566]= -2058723538;
assign addr[10567]= -2010011024;
assign addr[10568]= -1951102334;
assign addr[10569]= -1882296293;
assign addr[10570]= -1803941934;
assign addr[10571]= -1716436725;
assign addr[10572]= -1620224553;
assign addr[10573]= -1515793473;
assign addr[10574]= -1403673233;
assign addr[10575]= -1284432584;
assign addr[10576]= -1158676398;
assign addr[10577]= -1027042599;
assign addr[10578]= -890198924;
assign addr[10579]= -748839539;
assign addr[10580]= -603681519;
assign addr[10581]= -455461206;
assign addr[10582]= -304930476;
assign addr[10583]= -152852926;
assign addr[10584]= 0;
assign addr[10585]= 152852926;
assign addr[10586]= 304930476;
assign addr[10587]= 455461206;
assign addr[10588]= 603681519;
assign addr[10589]= 748839539;
assign addr[10590]= 890198924;
assign addr[10591]= 1027042599;
assign addr[10592]= 1158676398;
assign addr[10593]= 1284432584;
assign addr[10594]= 1403673233;
assign addr[10595]= 1515793473;
assign addr[10596]= 1620224553;
assign addr[10597]= 1716436725;
assign addr[10598]= 1803941934;
assign addr[10599]= 1882296293;
assign addr[10600]= 1951102334;
assign addr[10601]= 2010011024;
assign addr[10602]= 2058723538;
assign addr[10603]= 2096992772;
assign addr[10604]= 2124624598;
assign addr[10605]= 2141478848;
assign addr[10606]= 2147470025;
assign addr[10607]= 2142567738;
assign addr[10608]= 2126796855;
assign addr[10609]= 2100237377;
assign addr[10610]= 2063024031;
assign addr[10611]= 2015345591;
assign addr[10612]= 1957443913;
assign addr[10613]= 1889612716;
assign addr[10614]= 1812196087;
assign addr[10615]= 1725586737;
assign addr[10616]= 1630224009;
assign addr[10617]= 1526591649;
assign addr[10618]= 1415215352;
assign addr[10619]= 1296660098;
assign addr[10620]= 1171527280;
assign addr[10621]= 1040451659;
assign addr[10622]= 904098143;
assign addr[10623]= 763158411;
assign addr[10624]= 618347408;
assign addr[10625]= 470399716;
assign addr[10626]= 320065829;
assign addr[10627]= 168108346;
assign addr[10628]= 15298099;
assign addr[10629]= -137589750;
assign addr[10630]= -289779648;
assign addr[10631]= -440499581;
assign addr[10632]= -588984994;
assign addr[10633]= -734482665;
assign addr[10634]= -876254528;
assign addr[10635]= -1013581418;
assign addr[10636]= -1145766716;
assign addr[10637]= -1272139887;
assign addr[10638]= -1392059879;
assign addr[10639]= -1504918373;
assign addr[10640]= -1610142873;
assign addr[10641]= -1707199606;
assign addr[10642]= -1795596234;
assign addr[10643]= -1874884346;
assign addr[10644]= -1944661739;
assign addr[10645]= -2004574453;
assign addr[10646]= -2054318569;
assign addr[10647]= -2093641749;
assign addr[10648]= -2122344521;
assign addr[10649]= -2140281282;
assign addr[10650]= -2147361045;
assign addr[10651]= -2143547897;
assign addr[10652]= -2128861181;
assign addr[10653]= -2103375398;
assign addr[10654]= -2067219829;
assign addr[10655]= -2020577882;
assign addr[10656]= -1963686155;
assign addr[10657]= -1896833245;
assign addr[10658]= -1820358275;
assign addr[10659]= -1734649179;
assign addr[10660]= -1640140734;
assign addr[10661]= -1537312353;
assign addr[10662]= -1426685652;
assign addr[10663]= -1308821808;
assign addr[10664]= -1184318708;
assign addr[10665]= -1053807919;
assign addr[10666]= -917951481;
assign addr[10667]= -777438554;
assign addr[10668]= -632981917;
assign addr[10669]= -485314355;
assign addr[10670]= -335184940;
assign addr[10671]= -183355234;
assign addr[10672]= -30595422;
assign addr[10673]= 122319591;
assign addr[10674]= 274614114;
assign addr[10675]= 425515602;
assign addr[10676]= 574258580;
assign addr[10677]= 720088517;
assign addr[10678]= 862265664;
assign addr[10679]= 1000068799;
assign addr[10680]= 1132798888;
assign addr[10681]= 1259782632;
assign addr[10682]= 1380375881;
assign addr[10683]= 1493966902;
assign addr[10684]= 1599979481;
assign addr[10685]= 1697875851;
assign addr[10686]= 1787159411;
assign addr[10687]= 1867377253;
assign addr[10688]= 1938122457;
assign addr[10689]= 1999036154;
assign addr[10690]= 2049809346;
assign addr[10691]= 2090184478;
assign addr[10692]= 2119956737;
assign addr[10693]= 2138975100;
assign addr[10694]= 2147143090;
assign addr[10695]= 2144419275;
assign addr[10696]= 2130817471;
assign addr[10697]= 2106406677;
assign addr[10698]= 2071310720;
assign addr[10699]= 2025707632;
assign addr[10700]= 1969828744;
assign addr[10701]= 1903957513;
assign addr[10702]= 1828428082;
assign addr[10703]= 1743623590;
assign addr[10704]= 1649974225;
assign addr[10705]= 1547955041;
assign addr[10706]= 1438083551;
assign addr[10707]= 1320917099;
assign addr[10708]= 1197050035;
assign addr[10709]= 1067110699;
assign addr[10710]= 931758235;
assign addr[10711]= 791679244;
assign addr[10712]= 647584304;
assign addr[10713]= 500204365;
assign addr[10714]= 350287041;
assign addr[10715]= 198592817;
assign addr[10716]= 45891193;
assign addr[10717]= -107043224;
assign addr[10718]= -259434643;
assign addr[10719]= -410510029;
assign addr[10720]= -559503022;
assign addr[10721]= -705657826;
assign addr[10722]= -848233042;
assign addr[10723]= -986505429;
assign addr[10724]= -1119773573;
assign addr[10725]= -1247361445;
assign addr[10726]= -1368621831;
assign addr[10727]= -1482939614;
assign addr[10728]= -1589734894;
assign addr[10729]= -1688465931;
assign addr[10730]= -1778631892;
assign addr[10731]= -1859775393;
assign addr[10732]= -1931484818;
assign addr[10733]= -1993396407;
assign addr[10734]= -2045196100;
assign addr[10735]= -2086621133;
assign addr[10736]= -2117461370;
assign addr[10737]= -2137560369;
assign addr[10738]= -2146816171;
assign addr[10739]= -2145181827;
assign addr[10740]= -2132665626;
assign addr[10741]= -2109331059;
assign addr[10742]= -2075296495;
assign addr[10743]= -2030734582;
assign addr[10744]= -1975871368;
assign addr[10745]= -1910985158;
assign addr[10746]= -1836405100;
assign addr[10747]= -1752509516;
assign addr[10748]= -1659723983;
assign addr[10749]= -1558519173;
assign addr[10750]= -1449408469;
assign addr[10751]= -1332945355;
assign addr[10752]= -1209720613;
assign addr[10753]= -1080359326;
assign addr[10754]= -945517704;
assign addr[10755]= -805879757;
assign addr[10756]= -662153826;
assign addr[10757]= -515068990;
assign addr[10758]= -365371365;
assign addr[10759]= -213820322;
assign addr[10760]= -61184634;
assign addr[10761]= 91761426;
assign addr[10762]= 244242007;
assign addr[10763]= 395483624;
assign addr[10764]= 544719071;
assign addr[10765]= 691191324;
assign addr[10766]= 834157373;
assign addr[10767]= 972891995;
assign addr[10768]= 1106691431;
assign addr[10769]= 1234876957;
assign addr[10770]= 1356798326;
assign addr[10771]= 1471837070;
assign addr[10772]= 1579409630;
assign addr[10773]= 1678970324;
assign addr[10774]= 1770014111;
assign addr[10775]= 1852079154;
assign addr[10776]= 1924749160;
assign addr[10777]= 1987655498;
assign addr[10778]= 2040479063;
assign addr[10779]= 2082951896;
assign addr[10780]= 2114858546;
assign addr[10781]= 2136037160;
assign addr[10782]= 2146380306;
assign addr[10783]= 2145835515;
assign addr[10784]= 2134405552;
assign addr[10785]= 2112148396;
assign addr[10786]= 2079176953;
assign addr[10787]= 2035658475;
assign addr[10788]= 1981813720;
assign addr[10789]= 1917915825;
assign addr[10790]= 1844288924;
assign addr[10791]= 1761306505;
assign addr[10792]= 1669389513;
assign addr[10793]= 1569004214;
assign addr[10794]= 1460659832;
assign addr[10795]= 1344905966;
assign addr[10796]= 1222329801;
assign addr[10797]= 1093553126;
assign addr[10798]= 959229189;
assign addr[10799]= 820039373;
assign addr[10800]= 676689746;
assign addr[10801]= 529907477;
assign addr[10802]= 380437148;
assign addr[10803]= 229036977;
assign addr[10804]= 76474970;
assign addr[10805]= -76474970;
assign addr[10806]= -229036977;
assign addr[10807]= -380437148;
assign addr[10808]= -529907477;
assign addr[10809]= -676689746;
assign addr[10810]= -820039373;
assign addr[10811]= -959229189;
assign addr[10812]= -1093553126;
assign addr[10813]= -1222329801;
assign addr[10814]= -1344905966;
assign addr[10815]= -1460659832;
assign addr[10816]= -1569004214;
assign addr[10817]= -1669389513;
assign addr[10818]= -1761306505;
assign addr[10819]= -1844288924;
assign addr[10820]= -1917915825;
assign addr[10821]= -1981813720;
assign addr[10822]= -2035658475;
assign addr[10823]= -2079176953;
assign addr[10824]= -2112148396;
assign addr[10825]= -2134405552;
assign addr[10826]= -2145835515;
assign addr[10827]= -2146380306;
assign addr[10828]= -2136037160;
assign addr[10829]= -2114858546;
assign addr[10830]= -2082951896;
assign addr[10831]= -2040479063;
assign addr[10832]= -1987655498;
assign addr[10833]= -1924749160;
assign addr[10834]= -1852079154;
assign addr[10835]= -1770014111;
assign addr[10836]= -1678970324;
assign addr[10837]= -1579409630;
assign addr[10838]= -1471837070;
assign addr[10839]= -1356798326;
assign addr[10840]= -1234876957;
assign addr[10841]= -1106691431;
assign addr[10842]= -972891995;
assign addr[10843]= -834157373;
assign addr[10844]= -691191324;
assign addr[10845]= -544719071;
assign addr[10846]= -395483624;
assign addr[10847]= -244242007;
assign addr[10848]= -91761426;
assign addr[10849]= 61184634;
assign addr[10850]= 213820322;
assign addr[10851]= 365371365;
assign addr[10852]= 515068990;
assign addr[10853]= 662153826;
assign addr[10854]= 805879757;
assign addr[10855]= 945517704;
assign addr[10856]= 1080359326;
assign addr[10857]= 1209720613;
assign addr[10858]= 1332945355;
assign addr[10859]= 1449408469;
assign addr[10860]= 1558519173;
assign addr[10861]= 1659723983;
assign addr[10862]= 1752509516;
assign addr[10863]= 1836405100;
assign addr[10864]= 1910985158;
assign addr[10865]= 1975871368;
assign addr[10866]= 2030734582;
assign addr[10867]= 2075296495;
assign addr[10868]= 2109331059;
assign addr[10869]= 2132665626;
assign addr[10870]= 2145181827;
assign addr[10871]= 2146816171;
assign addr[10872]= 2137560369;
assign addr[10873]= 2117461370;
assign addr[10874]= 2086621133;
assign addr[10875]= 2045196100;
assign addr[10876]= 1993396407;
assign addr[10877]= 1931484818;
assign addr[10878]= 1859775393;
assign addr[10879]= 1778631892;
assign addr[10880]= 1688465931;
assign addr[10881]= 1589734894;
assign addr[10882]= 1482939614;
assign addr[10883]= 1368621831;
assign addr[10884]= 1247361445;
assign addr[10885]= 1119773573;
assign addr[10886]= 986505429;
assign addr[10887]= 848233042;
assign addr[10888]= 705657826;
assign addr[10889]= 559503022;
assign addr[10890]= 410510029;
assign addr[10891]= 259434643;
assign addr[10892]= 107043224;
assign addr[10893]= -45891193;
assign addr[10894]= -198592817;
assign addr[10895]= -350287041;
assign addr[10896]= -500204365;
assign addr[10897]= -647584304;
assign addr[10898]= -791679244;
assign addr[10899]= -931758235;
assign addr[10900]= -1067110699;
assign addr[10901]= -1197050035;
assign addr[10902]= -1320917099;
assign addr[10903]= -1438083551;
assign addr[10904]= -1547955041;
assign addr[10905]= -1649974225;
assign addr[10906]= -1743623590;
assign addr[10907]= -1828428082;
assign addr[10908]= -1903957513;
assign addr[10909]= -1969828744;
assign addr[10910]= -2025707632;
assign addr[10911]= -2071310720;
assign addr[10912]= -2106406677;
assign addr[10913]= -2130817471;
assign addr[10914]= -2144419275;
assign addr[10915]= -2147143090;
assign addr[10916]= -2138975100;
assign addr[10917]= -2119956737;
assign addr[10918]= -2090184478;
assign addr[10919]= -2049809346;
assign addr[10920]= -1999036154;
assign addr[10921]= -1938122457;
assign addr[10922]= -1867377253;
assign addr[10923]= -1787159411;
assign addr[10924]= -1697875851;
assign addr[10925]= -1599979481;
assign addr[10926]= -1493966902;
assign addr[10927]= -1380375881;
assign addr[10928]= -1259782632;
assign addr[10929]= -1132798888;
assign addr[10930]= -1000068799;
assign addr[10931]= -862265664;
assign addr[10932]= -720088517;
assign addr[10933]= -574258580;
assign addr[10934]= -425515602;
assign addr[10935]= -274614114;
assign addr[10936]= -122319591;
assign addr[10937]= 30595422;
assign addr[10938]= 183355234;
assign addr[10939]= 335184940;
assign addr[10940]= 485314355;
assign addr[10941]= 632981917;
assign addr[10942]= 777438554;
assign addr[10943]= 917951481;
assign addr[10944]= 1053807919;
assign addr[10945]= 1184318708;
assign addr[10946]= 1308821808;
assign addr[10947]= 1426685652;
assign addr[10948]= 1537312353;
assign addr[10949]= 1640140734;
assign addr[10950]= 1734649179;
assign addr[10951]= 1820358275;
assign addr[10952]= 1896833245;
assign addr[10953]= 1963686155;
assign addr[10954]= 2020577882;
assign addr[10955]= 2067219829;
assign addr[10956]= 2103375398;
assign addr[10957]= 2128861181;
assign addr[10958]= 2143547897;
assign addr[10959]= 2147361045;
assign addr[10960]= 2140281282;
assign addr[10961]= 2122344521;
assign addr[10962]= 2093641749;
assign addr[10963]= 2054318569;
assign addr[10964]= 2004574453;
assign addr[10965]= 1944661739;
assign addr[10966]= 1874884346;
assign addr[10967]= 1795596234;
assign addr[10968]= 1707199606;
assign addr[10969]= 1610142873;
assign addr[10970]= 1504918373;
assign addr[10971]= 1392059879;
assign addr[10972]= 1272139887;
assign addr[10973]= 1145766716;
assign addr[10974]= 1013581418;
assign addr[10975]= 876254528;
assign addr[10976]= 734482665;
assign addr[10977]= 588984994;
assign addr[10978]= 440499581;
assign addr[10979]= 289779648;
assign addr[10980]= 137589750;
assign addr[10981]= -15298099;
assign addr[10982]= -168108346;
assign addr[10983]= -320065829;
assign addr[10984]= -470399716;
assign addr[10985]= -618347408;
assign addr[10986]= -763158411;
assign addr[10987]= -904098143;
assign addr[10988]= -1040451659;
assign addr[10989]= -1171527280;
assign addr[10990]= -1296660098;
assign addr[10991]= -1415215352;
assign addr[10992]= -1526591649;
assign addr[10993]= -1630224009;
assign addr[10994]= -1725586737;
assign addr[10995]= -1812196087;
assign addr[10996]= -1889612716;
assign addr[10997]= -1957443913;
assign addr[10998]= -2015345591;
assign addr[10999]= -2063024031;
assign addr[11000]= -2100237377;
assign addr[11001]= -2126796855;
assign addr[11002]= -2142567738;
assign addr[11003]= -2147470025;
assign addr[11004]= -2141478848;
assign addr[11005]= -2124624598;
assign addr[11006]= -2096992772;
assign addr[11007]= -2058723538;
assign addr[11008]= -2010011024;
assign addr[11009]= -1951102334;
assign addr[11010]= -1882296293;
assign addr[11011]= -1803941934;
assign addr[11012]= -1716436725;
assign addr[11013]= -1620224553;
assign addr[11014]= -1515793473;
assign addr[11015]= -1403673233;
assign addr[11016]= -1284432584;
assign addr[11017]= -1158676398;
assign addr[11018]= -1027042599;
assign addr[11019]= -890198924;
assign addr[11020]= -748839539;
assign addr[11021]= -603681519;
assign addr[11022]= -455461206;
assign addr[11023]= -304930476;
assign addr[11024]= -152852926;
assign addr[11025]= 0;
assign addr[11026]= 152852926;
assign addr[11027]= 304930476;
assign addr[11028]= 455461206;
assign addr[11029]= 603681519;
assign addr[11030]= 748839539;
assign addr[11031]= 890198924;
assign addr[11032]= 1027042599;
assign addr[11033]= 1158676398;
assign addr[11034]= 1284432584;
assign addr[11035]= 1403673233;
assign addr[11036]= 1515793473;
assign addr[11037]= 1620224553;
assign addr[11038]= 1716436725;
assign addr[11039]= 1803941934;
assign addr[11040]= 1882296293;
assign addr[11041]= 1951102334;
assign addr[11042]= 2010011024;
assign addr[11043]= 2058723538;
assign addr[11044]= 2096992772;
assign addr[11045]= 2124624598;
assign addr[11046]= 2141478848;
assign addr[11047]= 2147470025;
assign addr[11048]= 2142567738;
assign addr[11049]= 2126796855;
assign addr[11050]= 2100237377;
assign addr[11051]= 2063024031;
assign addr[11052]= 2015345591;
assign addr[11053]= 1957443913;
assign addr[11054]= 1889612716;
assign addr[11055]= 1812196087;
assign addr[11056]= 1725586737;
assign addr[11057]= 1630224009;
assign addr[11058]= 1526591649;
assign addr[11059]= 1415215352;
assign addr[11060]= 1296660098;
assign addr[11061]= 1171527280;
assign addr[11062]= 1040451659;
assign addr[11063]= 904098143;
assign addr[11064]= 763158411;
assign addr[11065]= 618347408;
assign addr[11066]= 470399716;
assign addr[11067]= 320065829;
assign addr[11068]= 168108346;
assign addr[11069]= 15298099;
assign addr[11070]= -137589750;
assign addr[11071]= -289779648;
assign addr[11072]= -440499581;
assign addr[11073]= -588984994;
assign addr[11074]= -734482665;
assign addr[11075]= -876254528;
assign addr[11076]= -1013581418;
assign addr[11077]= -1145766716;
assign addr[11078]= -1272139887;
assign addr[11079]= -1392059879;
assign addr[11080]= -1504918373;
assign addr[11081]= -1610142873;
assign addr[11082]= -1707199606;
assign addr[11083]= -1795596234;
assign addr[11084]= -1874884346;
assign addr[11085]= -1944661739;
assign addr[11086]= -2004574453;
assign addr[11087]= -2054318569;
assign addr[11088]= -2093641749;
assign addr[11089]= -2122344521;
assign addr[11090]= -2140281282;
assign addr[11091]= -2147361045;
assign addr[11092]= -2143547897;
assign addr[11093]= -2128861181;
assign addr[11094]= -2103375398;
assign addr[11095]= -2067219829;
assign addr[11096]= -2020577882;
assign addr[11097]= -1963686155;
assign addr[11098]= -1896833245;
assign addr[11099]= -1820358275;
assign addr[11100]= -1734649179;
assign addr[11101]= -1640140734;
assign addr[11102]= -1537312353;
assign addr[11103]= -1426685652;
assign addr[11104]= -1308821808;
assign addr[11105]= -1184318708;
assign addr[11106]= -1053807919;
assign addr[11107]= -917951481;
assign addr[11108]= -777438554;
assign addr[11109]= -632981917;
assign addr[11110]= -485314355;
assign addr[11111]= -335184940;
assign addr[11112]= -183355234;
assign addr[11113]= -30595422;
assign addr[11114]= 122319591;
assign addr[11115]= 274614114;
assign addr[11116]= 425515602;
assign addr[11117]= 574258580;
assign addr[11118]= 720088517;
assign addr[11119]= 862265664;
assign addr[11120]= 1000068799;
assign addr[11121]= 1132798888;
assign addr[11122]= 1259782632;
assign addr[11123]= 1380375881;
assign addr[11124]= 1493966902;
assign addr[11125]= 1599979481;
assign addr[11126]= 1697875851;
assign addr[11127]= 1787159411;
assign addr[11128]= 1867377253;
assign addr[11129]= 1938122457;
assign addr[11130]= 1999036154;
assign addr[11131]= 2049809346;
assign addr[11132]= 2090184478;
assign addr[11133]= 2119956737;
assign addr[11134]= 2138975100;
assign addr[11135]= 2147143090;
assign addr[11136]= 2144419275;
assign addr[11137]= 2130817471;
assign addr[11138]= 2106406677;
assign addr[11139]= 2071310720;
assign addr[11140]= 2025707632;
assign addr[11141]= 1969828744;
assign addr[11142]= 1903957513;
assign addr[11143]= 1828428082;
assign addr[11144]= 1743623590;
assign addr[11145]= 1649974225;
assign addr[11146]= 1547955041;
assign addr[11147]= 1438083551;
assign addr[11148]= 1320917099;
assign addr[11149]= 1197050035;
assign addr[11150]= 1067110699;
assign addr[11151]= 931758235;
assign addr[11152]= 791679244;
assign addr[11153]= 647584304;
assign addr[11154]= 500204365;
assign addr[11155]= 350287041;
assign addr[11156]= 198592817;
assign addr[11157]= 45891193;
assign addr[11158]= -107043224;
assign addr[11159]= -259434643;
assign addr[11160]= -410510029;
assign addr[11161]= -559503022;
assign addr[11162]= -705657826;
assign addr[11163]= -848233042;
assign addr[11164]= -986505429;
assign addr[11165]= -1119773573;
assign addr[11166]= -1247361445;
assign addr[11167]= -1368621831;
assign addr[11168]= -1482939614;
assign addr[11169]= -1589734894;
assign addr[11170]= -1688465931;
assign addr[11171]= -1778631892;
assign addr[11172]= -1859775393;
assign addr[11173]= -1931484818;
assign addr[11174]= -1993396407;
assign addr[11175]= -2045196100;
assign addr[11176]= -2086621133;
assign addr[11177]= -2117461370;
assign addr[11178]= -2137560369;
assign addr[11179]= -2146816171;
assign addr[11180]= -2145181827;
assign addr[11181]= -2132665626;
assign addr[11182]= -2109331059;
assign addr[11183]= -2075296495;
assign addr[11184]= -2030734582;
assign addr[11185]= -1975871368;
assign addr[11186]= -1910985158;
assign addr[11187]= -1836405100;
assign addr[11188]= -1752509516;
assign addr[11189]= -1659723983;
assign addr[11190]= -1558519173;
assign addr[11191]= -1449408469;
assign addr[11192]= -1332945355;
assign addr[11193]= -1209720613;
assign addr[11194]= -1080359326;
assign addr[11195]= -945517704;
assign addr[11196]= -805879757;
assign addr[11197]= -662153826;
assign addr[11198]= -515068990;
assign addr[11199]= -365371365;
assign addr[11200]= -213820322;
assign addr[11201]= -61184634;
assign addr[11202]= 91761426;
assign addr[11203]= 244242007;
assign addr[11204]= 395483624;
assign addr[11205]= 544719071;
assign addr[11206]= 691191324;
assign addr[11207]= 834157373;
assign addr[11208]= 972891995;
assign addr[11209]= 1106691431;
assign addr[11210]= 1234876957;
assign addr[11211]= 1356798326;
assign addr[11212]= 1471837070;
assign addr[11213]= 1579409630;
assign addr[11214]= 1678970324;
assign addr[11215]= 1770014111;
assign addr[11216]= 1852079154;
assign addr[11217]= 1924749160;
assign addr[11218]= 1987655498;
assign addr[11219]= 2040479063;
assign addr[11220]= 2082951896;
assign addr[11221]= 2114858546;
assign addr[11222]= 2136037160;
assign addr[11223]= 2146380306;
assign addr[11224]= 2145835515;
assign addr[11225]= 2134405552;
assign addr[11226]= 2112148396;
assign addr[11227]= 2079176953;
assign addr[11228]= 2035658475;
assign addr[11229]= 1981813720;
assign addr[11230]= 1917915825;
assign addr[11231]= 1844288924;
assign addr[11232]= 1761306505;
assign addr[11233]= 1669389513;
assign addr[11234]= 1569004214;
assign addr[11235]= 1460659832;
assign addr[11236]= 1344905966;
assign addr[11237]= 1222329801;
assign addr[11238]= 1093553126;
assign addr[11239]= 959229189;
assign addr[11240]= 820039373;
assign addr[11241]= 676689746;
assign addr[11242]= 529907477;
assign addr[11243]= 380437148;
assign addr[11244]= 229036977;
assign addr[11245]= 76474970;
assign addr[11246]= -76474970;
assign addr[11247]= -229036977;
assign addr[11248]= -380437148;
assign addr[11249]= -529907477;
assign addr[11250]= -676689746;
assign addr[11251]= -820039373;
assign addr[11252]= -959229189;
assign addr[11253]= -1093553126;
assign addr[11254]= -1222329801;
assign addr[11255]= -1344905966;
assign addr[11256]= -1460659832;
assign addr[11257]= -1569004214;
assign addr[11258]= -1669389513;
assign addr[11259]= -1761306505;
assign addr[11260]= -1844288924;
assign addr[11261]= -1917915825;
assign addr[11262]= -1981813720;
assign addr[11263]= -2035658475;
assign addr[11264]= -2079176953;
assign addr[11265]= -2112148396;
assign addr[11266]= -2134405552;
assign addr[11267]= -2145835515;
assign addr[11268]= -2146380306;
assign addr[11269]= -2136037160;
assign addr[11270]= -2114858546;
assign addr[11271]= -2082951896;
assign addr[11272]= -2040479063;
assign addr[11273]= -1987655498;
assign addr[11274]= -1924749160;
assign addr[11275]= -1852079154;
assign addr[11276]= -1770014111;
assign addr[11277]= -1678970324;
assign addr[11278]= -1579409630;
assign addr[11279]= -1471837070;
assign addr[11280]= -1356798326;
assign addr[11281]= -1234876957;
assign addr[11282]= -1106691431;
assign addr[11283]= -972891995;
assign addr[11284]= -834157373;
assign addr[11285]= -691191324;
assign addr[11286]= -544719071;
assign addr[11287]= -395483624;
assign addr[11288]= -244242007;
assign addr[11289]= -91761426;
assign addr[11290]= 61184634;
assign addr[11291]= 213820322;
assign addr[11292]= 365371365;
assign addr[11293]= 515068990;
assign addr[11294]= 662153826;
assign addr[11295]= 805879757;
assign addr[11296]= 945517704;
assign addr[11297]= 1080359326;
assign addr[11298]= 1209720613;
assign addr[11299]= 1332945355;
assign addr[11300]= 1449408469;
assign addr[11301]= 1558519173;
assign addr[11302]= 1659723983;
assign addr[11303]= 1752509516;
assign addr[11304]= 1836405100;
assign addr[11305]= 1910985158;
assign addr[11306]= 1975871368;
assign addr[11307]= 2030734582;
assign addr[11308]= 2075296495;
assign addr[11309]= 2109331059;
assign addr[11310]= 2132665626;
assign addr[11311]= 2145181827;
assign addr[11312]= 2146816171;
assign addr[11313]= 2137560369;
assign addr[11314]= 2117461370;
assign addr[11315]= 2086621133;
assign addr[11316]= 2045196100;
assign addr[11317]= 1993396407;
assign addr[11318]= 1931484818;
assign addr[11319]= 1859775393;
assign addr[11320]= 1778631892;
assign addr[11321]= 1688465931;
assign addr[11322]= 1589734894;
assign addr[11323]= 1482939614;
assign addr[11324]= 1368621831;
assign addr[11325]= 1247361445;
assign addr[11326]= 1119773573;
assign addr[11327]= 986505429;
assign addr[11328]= 848233042;
assign addr[11329]= 705657826;
assign addr[11330]= 559503022;
assign addr[11331]= 410510029;
assign addr[11332]= 259434643;
assign addr[11333]= 107043224;
assign addr[11334]= -45891193;
assign addr[11335]= -198592817;
assign addr[11336]= -350287041;
assign addr[11337]= -500204365;
assign addr[11338]= -647584304;
assign addr[11339]= -791679244;
assign addr[11340]= -931758235;
assign addr[11341]= -1067110699;
assign addr[11342]= -1197050035;
assign addr[11343]= -1320917099;
assign addr[11344]= -1438083551;
assign addr[11345]= -1547955041;
assign addr[11346]= -1649974225;
assign addr[11347]= -1743623590;
assign addr[11348]= -1828428082;
assign addr[11349]= -1903957513;
assign addr[11350]= -1969828744;
assign addr[11351]= -2025707632;
assign addr[11352]= -2071310720;
assign addr[11353]= -2106406677;
assign addr[11354]= -2130817471;
assign addr[11355]= -2144419275;
assign addr[11356]= -2147143090;
assign addr[11357]= -2138975100;
assign addr[11358]= -2119956737;
assign addr[11359]= -2090184478;
assign addr[11360]= -2049809346;
assign addr[11361]= -1999036154;
assign addr[11362]= -1938122457;
assign addr[11363]= -1867377253;
assign addr[11364]= -1787159411;
assign addr[11365]= -1697875851;
assign addr[11366]= -1599979481;
assign addr[11367]= -1493966902;
assign addr[11368]= -1380375881;
assign addr[11369]= -1259782632;
assign addr[11370]= -1132798888;
assign addr[11371]= -1000068799;
assign addr[11372]= -862265664;
assign addr[11373]= -720088517;
assign addr[11374]= -574258580;
assign addr[11375]= -425515602;
assign addr[11376]= -274614114;
assign addr[11377]= -122319591;
assign addr[11378]= 30595422;
assign addr[11379]= 183355234;
assign addr[11380]= 335184940;
assign addr[11381]= 485314355;
assign addr[11382]= 632981917;
assign addr[11383]= 777438554;
assign addr[11384]= 917951481;
assign addr[11385]= 1053807919;
assign addr[11386]= 1184318708;
assign addr[11387]= 1308821808;
assign addr[11388]= 1426685652;
assign addr[11389]= 1537312353;
assign addr[11390]= 1640140734;
assign addr[11391]= 1734649179;
assign addr[11392]= 1820358275;
assign addr[11393]= 1896833245;
assign addr[11394]= 1963686155;
assign addr[11395]= 2020577882;
assign addr[11396]= 2067219829;
assign addr[11397]= 2103375398;
assign addr[11398]= 2128861181;
assign addr[11399]= 2143547897;
assign addr[11400]= 2147361045;
assign addr[11401]= 2140281282;
assign addr[11402]= 2122344521;
assign addr[11403]= 2093641749;
assign addr[11404]= 2054318569;
assign addr[11405]= 2004574453;
assign addr[11406]= 1944661739;
assign addr[11407]= 1874884346;
assign addr[11408]= 1795596234;
assign addr[11409]= 1707199606;
assign addr[11410]= 1610142873;
assign addr[11411]= 1504918373;
assign addr[11412]= 1392059879;
assign addr[11413]= 1272139887;
assign addr[11414]= 1145766716;
assign addr[11415]= 1013581418;
assign addr[11416]= 876254528;
assign addr[11417]= 734482665;
assign addr[11418]= 588984994;
assign addr[11419]= 440499581;
assign addr[11420]= 289779648;
assign addr[11421]= 137589750;
assign addr[11422]= -15298099;
assign addr[11423]= -168108346;
assign addr[11424]= -320065829;
assign addr[11425]= -470399716;
assign addr[11426]= -618347408;
assign addr[11427]= -763158411;
assign addr[11428]= -904098143;
assign addr[11429]= -1040451659;
assign addr[11430]= -1171527280;
assign addr[11431]= -1296660098;
assign addr[11432]= -1415215352;
assign addr[11433]= -1526591649;
assign addr[11434]= -1630224009;
assign addr[11435]= -1725586737;
assign addr[11436]= -1812196087;
assign addr[11437]= -1889612716;
assign addr[11438]= -1957443913;
assign addr[11439]= -2015345591;
assign addr[11440]= -2063024031;
assign addr[11441]= -2100237377;
assign addr[11442]= -2126796855;
assign addr[11443]= -2142567738;
assign addr[11444]= -2147470025;
assign addr[11445]= -2141478848;
assign addr[11446]= -2124624598;
assign addr[11447]= -2096992772;
assign addr[11448]= -2058723538;
assign addr[11449]= -2010011024;
assign addr[11450]= -1951102334;
assign addr[11451]= -1882296293;
assign addr[11452]= -1803941934;
assign addr[11453]= -1716436725;
assign addr[11454]= -1620224553;
assign addr[11455]= -1515793473;
assign addr[11456]= -1403673233;
assign addr[11457]= -1284432584;
assign addr[11458]= -1158676398;
assign addr[11459]= -1027042599;
assign addr[11460]= -890198924;
assign addr[11461]= -748839539;
assign addr[11462]= -603681519;
assign addr[11463]= -455461206;
assign addr[11464]= -304930476;
assign addr[11465]= -152852926;
assign addr[11466]= 0;
assign addr[11467]= 152852926;
assign addr[11468]= 304930476;
assign addr[11469]= 455461206;
assign addr[11470]= 603681519;
assign addr[11471]= 748839539;
assign addr[11472]= 890198924;
assign addr[11473]= 1027042599;
assign addr[11474]= 1158676398;
assign addr[11475]= 1284432584;
assign addr[11476]= 1403673233;
assign addr[11477]= 1515793473;
assign addr[11478]= 1620224553;
assign addr[11479]= 1716436725;
assign addr[11480]= 1803941934;
assign addr[11481]= 1882296293;
assign addr[11482]= 1951102334;
assign addr[11483]= 2010011024;
assign addr[11484]= 2058723538;
assign addr[11485]= 2096992772;
assign addr[11486]= 2124624598;
assign addr[11487]= 2141478848;
assign addr[11488]= 2147470025;
assign addr[11489]= 2142567738;
assign addr[11490]= 2126796855;
assign addr[11491]= 2100237377;
assign addr[11492]= 2063024031;
assign addr[11493]= 2015345591;
assign addr[11494]= 1957443913;
assign addr[11495]= 1889612716;
assign addr[11496]= 1812196087;
assign addr[11497]= 1725586737;
assign addr[11498]= 1630224009;
assign addr[11499]= 1526591649;
assign addr[11500]= 1415215352;
assign addr[11501]= 1296660098;
assign addr[11502]= 1171527280;
assign addr[11503]= 1040451659;
assign addr[11504]= 904098143;
assign addr[11505]= 763158411;
assign addr[11506]= 618347408;
assign addr[11507]= 470399716;
assign addr[11508]= 320065829;
assign addr[11509]= 168108346;
assign addr[11510]= 15298099;
assign addr[11511]= -137589750;
assign addr[11512]= -289779648;
assign addr[11513]= -440499581;
assign addr[11514]= -588984994;
assign addr[11515]= -734482665;
assign addr[11516]= -876254528;
assign addr[11517]= -1013581418;
assign addr[11518]= -1145766716;
assign addr[11519]= -1272139887;
assign addr[11520]= -1392059879;
assign addr[11521]= -1504918373;
assign addr[11522]= -1610142873;
assign addr[11523]= -1707199606;
assign addr[11524]= -1795596234;
assign addr[11525]= -1874884346;
assign addr[11526]= -1944661739;
assign addr[11527]= -2004574453;
assign addr[11528]= -2054318569;
assign addr[11529]= -2093641749;
assign addr[11530]= -2122344521;
assign addr[11531]= -2140281282;
assign addr[11532]= -2147361045;
assign addr[11533]= -2143547897;
assign addr[11534]= -2128861181;
assign addr[11535]= -2103375398;
assign addr[11536]= -2067219829;
assign addr[11537]= -2020577882;
assign addr[11538]= -1963686155;
assign addr[11539]= -1896833245;
assign addr[11540]= -1820358275;
assign addr[11541]= -1734649179;
assign addr[11542]= -1640140734;
assign addr[11543]= -1537312353;
assign addr[11544]= -1426685652;
assign addr[11545]= -1308821808;
assign addr[11546]= -1184318708;
assign addr[11547]= -1053807919;
assign addr[11548]= -917951481;
assign addr[11549]= -777438554;
assign addr[11550]= -632981917;
assign addr[11551]= -485314355;
assign addr[11552]= -335184940;
assign addr[11553]= -183355234;
assign addr[11554]= -30595422;
assign addr[11555]= 122319591;
assign addr[11556]= 274614114;
assign addr[11557]= 425515602;
assign addr[11558]= 574258580;
assign addr[11559]= 720088517;
assign addr[11560]= 862265664;
assign addr[11561]= 1000068799;
assign addr[11562]= 1132798888;
assign addr[11563]= 1259782632;
assign addr[11564]= 1380375881;
assign addr[11565]= 1493966902;
assign addr[11566]= 1599979481;
assign addr[11567]= 1697875851;
assign addr[11568]= 1787159411;
assign addr[11569]= 1867377253;
assign addr[11570]= 1938122457;
assign addr[11571]= 1999036154;
assign addr[11572]= 2049809346;
assign addr[11573]= 2090184478;
assign addr[11574]= 2119956737;
assign addr[11575]= 2138975100;
assign addr[11576]= 2147143090;
assign addr[11577]= 2144419275;
assign addr[11578]= 2130817471;
assign addr[11579]= 2106406677;
assign addr[11580]= 2071310720;
assign addr[11581]= 2025707632;
assign addr[11582]= 1969828744;
assign addr[11583]= 1903957513;
assign addr[11584]= 1828428082;
assign addr[11585]= 1743623590;
assign addr[11586]= 1649974225;
assign addr[11587]= 1547955041;
assign addr[11588]= 1438083551;
assign addr[11589]= 1320917099;
assign addr[11590]= 1197050035;
assign addr[11591]= 1067110699;
assign addr[11592]= 931758235;
assign addr[11593]= 791679244;
assign addr[11594]= 647584304;
assign addr[11595]= 500204365;
assign addr[11596]= 350287041;
assign addr[11597]= 198592817;
assign addr[11598]= 45891193;
assign addr[11599]= -107043224;
assign addr[11600]= -259434643;
assign addr[11601]= -410510029;
assign addr[11602]= -559503022;
assign addr[11603]= -705657826;
assign addr[11604]= -848233042;
assign addr[11605]= -986505429;
assign addr[11606]= -1119773573;
assign addr[11607]= -1247361445;
assign addr[11608]= -1368621831;
assign addr[11609]= -1482939614;
assign addr[11610]= -1589734894;
assign addr[11611]= -1688465931;
assign addr[11612]= -1778631892;
assign addr[11613]= -1859775393;
assign addr[11614]= -1931484818;
assign addr[11615]= -1993396407;
assign addr[11616]= -2045196100;
assign addr[11617]= -2086621133;
assign addr[11618]= -2117461370;
assign addr[11619]= -2137560369;
assign addr[11620]= -2146816171;
assign addr[11621]= -2145181827;
assign addr[11622]= -2132665626;
assign addr[11623]= -2109331059;
assign addr[11624]= -2075296495;
assign addr[11625]= -2030734582;
assign addr[11626]= -1975871368;
assign addr[11627]= -1910985158;
assign addr[11628]= -1836405100;
assign addr[11629]= -1752509516;
assign addr[11630]= -1659723983;
assign addr[11631]= -1558519173;
assign addr[11632]= -1449408469;
assign addr[11633]= -1332945355;
assign addr[11634]= -1209720613;
assign addr[11635]= -1080359326;
assign addr[11636]= -945517704;
assign addr[11637]= -805879757;
assign addr[11638]= -662153826;
assign addr[11639]= -515068990;
assign addr[11640]= -365371365;
assign addr[11641]= -213820322;
assign addr[11642]= -61184634;
assign addr[11643]= 91761426;
assign addr[11644]= 244242007;
assign addr[11645]= 395483624;
assign addr[11646]= 544719071;
assign addr[11647]= 691191324;
assign addr[11648]= 834157373;
assign addr[11649]= 972891995;
assign addr[11650]= 1106691431;
assign addr[11651]= 1234876957;
assign addr[11652]= 1356798326;
assign addr[11653]= 1471837070;
assign addr[11654]= 1579409630;
assign addr[11655]= 1678970324;
assign addr[11656]= 1770014111;
assign addr[11657]= 1852079154;
assign addr[11658]= 1924749160;
assign addr[11659]= 1987655498;
assign addr[11660]= 2040479063;
assign addr[11661]= 2082951896;
assign addr[11662]= 2114858546;
assign addr[11663]= 2136037160;
assign addr[11664]= 2146380306;
assign addr[11665]= 2145835515;
assign addr[11666]= 2134405552;
assign addr[11667]= 2112148396;
assign addr[11668]= 2079176953;
assign addr[11669]= 2035658475;
assign addr[11670]= 1981813720;
assign addr[11671]= 1917915825;
assign addr[11672]= 1844288924;
assign addr[11673]= 1761306505;
assign addr[11674]= 1669389513;
assign addr[11675]= 1569004214;
assign addr[11676]= 1460659832;
assign addr[11677]= 1344905966;
assign addr[11678]= 1222329801;
assign addr[11679]= 1093553126;
assign addr[11680]= 959229189;
assign addr[11681]= 820039373;
assign addr[11682]= 676689746;
assign addr[11683]= 529907477;
assign addr[11684]= 380437148;
assign addr[11685]= 229036977;
assign addr[11686]= 76474970;
assign addr[11687]= -76474970;
assign addr[11688]= -229036977;
assign addr[11689]= -380437148;
assign addr[11690]= -529907477;
assign addr[11691]= -676689746;
assign addr[11692]= -820039373;
assign addr[11693]= -959229189;
assign addr[11694]= -1093553126;
assign addr[11695]= -1222329801;
assign addr[11696]= -1344905966;
assign addr[11697]= -1460659832;
assign addr[11698]= -1569004214;
assign addr[11699]= -1669389513;
assign addr[11700]= -1761306505;
assign addr[11701]= -1844288924;
assign addr[11702]= -1917915825;
assign addr[11703]= -1981813720;
assign addr[11704]= -2035658475;
assign addr[11705]= -2079176953;
assign addr[11706]= -2112148396;
assign addr[11707]= -2134405552;
assign addr[11708]= -2145835515;
assign addr[11709]= -2146380306;
assign addr[11710]= -2136037160;
assign addr[11711]= -2114858546;
assign addr[11712]= -2082951896;
assign addr[11713]= -2040479063;
assign addr[11714]= -1987655498;
assign addr[11715]= -1924749160;
assign addr[11716]= -1852079154;
assign addr[11717]= -1770014111;
assign addr[11718]= -1678970324;
assign addr[11719]= -1579409630;
assign addr[11720]= -1471837070;
assign addr[11721]= -1356798326;
assign addr[11722]= -1234876957;
assign addr[11723]= -1106691431;
assign addr[11724]= -972891995;
assign addr[11725]= -834157373;
assign addr[11726]= -691191324;
assign addr[11727]= -544719071;
assign addr[11728]= -395483624;
assign addr[11729]= -244242007;
assign addr[11730]= -91761426;
assign addr[11731]= 61184634;
assign addr[11732]= 213820322;
assign addr[11733]= 365371365;
assign addr[11734]= 515068990;
assign addr[11735]= 662153826;
assign addr[11736]= 805879757;
assign addr[11737]= 945517704;
assign addr[11738]= 1080359326;
assign addr[11739]= 1209720613;
assign addr[11740]= 1332945355;
assign addr[11741]= 1449408469;
assign addr[11742]= 1558519173;
assign addr[11743]= 1659723983;
assign addr[11744]= 1752509516;
assign addr[11745]= 1836405100;
assign addr[11746]= 1910985158;
assign addr[11747]= 1975871368;
assign addr[11748]= 2030734582;
assign addr[11749]= 2075296495;
assign addr[11750]= 2109331059;
assign addr[11751]= 2132665626;
assign addr[11752]= 2145181827;
assign addr[11753]= 2146816171;
assign addr[11754]= 2137560369;
assign addr[11755]= 2117461370;
assign addr[11756]= 2086621133;
assign addr[11757]= 2045196100;
assign addr[11758]= 1993396407;
assign addr[11759]= 1931484818;
assign addr[11760]= 1859775393;
assign addr[11761]= 1778631892;
assign addr[11762]= 1688465931;
assign addr[11763]= 1589734894;
assign addr[11764]= 1482939614;
assign addr[11765]= 1368621831;
assign addr[11766]= 1247361445;
assign addr[11767]= 1119773573;
assign addr[11768]= 986505429;
assign addr[11769]= 848233042;
assign addr[11770]= 705657826;
assign addr[11771]= 559503022;
assign addr[11772]= 410510029;
assign addr[11773]= 259434643;
assign addr[11774]= 107043224;
assign addr[11775]= -45891193;
assign addr[11776]= -198592817;
assign addr[11777]= -350287041;
assign addr[11778]= -500204365;
assign addr[11779]= -647584304;
assign addr[11780]= -791679244;
assign addr[11781]= -931758235;
assign addr[11782]= -1067110699;
assign addr[11783]= -1197050035;
assign addr[11784]= -1320917099;
assign addr[11785]= -1438083551;
assign addr[11786]= -1547955041;
assign addr[11787]= -1649974225;
assign addr[11788]= -1743623590;
assign addr[11789]= -1828428082;
assign addr[11790]= -1903957513;
assign addr[11791]= -1969828744;
assign addr[11792]= -2025707632;
assign addr[11793]= -2071310720;
assign addr[11794]= -2106406677;
assign addr[11795]= -2130817471;
assign addr[11796]= -2144419275;
assign addr[11797]= -2147143090;
assign addr[11798]= -2138975100;
assign addr[11799]= -2119956737;
assign addr[11800]= -2090184478;
assign addr[11801]= -2049809346;
assign addr[11802]= -1999036154;
assign addr[11803]= -1938122457;
assign addr[11804]= -1867377253;
assign addr[11805]= -1787159411;
assign addr[11806]= -1697875851;
assign addr[11807]= -1599979481;
assign addr[11808]= -1493966902;
assign addr[11809]= -1380375881;
assign addr[11810]= -1259782632;
assign addr[11811]= -1132798888;
assign addr[11812]= -1000068799;
assign addr[11813]= -862265664;
assign addr[11814]= -720088517;
assign addr[11815]= -574258580;
assign addr[11816]= -425515602;
assign addr[11817]= -274614114;
assign addr[11818]= -122319591;
assign addr[11819]= 30595422;
assign addr[11820]= 183355234;
assign addr[11821]= 335184940;
assign addr[11822]= 485314355;
assign addr[11823]= 632981917;
assign addr[11824]= 777438554;
assign addr[11825]= 917951481;
assign addr[11826]= 1053807919;
assign addr[11827]= 1184318708;
assign addr[11828]= 1308821808;
assign addr[11829]= 1426685652;
assign addr[11830]= 1537312353;
assign addr[11831]= 1640140734;
assign addr[11832]= 1734649179;
assign addr[11833]= 1820358275;
assign addr[11834]= 1896833245;
assign addr[11835]= 1963686155;
assign addr[11836]= 2020577882;
assign addr[11837]= 2067219829;
assign addr[11838]= 2103375398;
assign addr[11839]= 2128861181;
assign addr[11840]= 2143547897;
assign addr[11841]= 2147361045;
assign addr[11842]= 2140281282;
assign addr[11843]= 2122344521;
assign addr[11844]= 2093641749;
assign addr[11845]= 2054318569;
assign addr[11846]= 2004574453;
assign addr[11847]= 1944661739;
assign addr[11848]= 1874884346;
assign addr[11849]= 1795596234;
assign addr[11850]= 1707199606;
assign addr[11851]= 1610142873;
assign addr[11852]= 1504918373;
assign addr[11853]= 1392059879;
assign addr[11854]= 1272139887;
assign addr[11855]= 1145766716;
assign addr[11856]= 1013581418;
assign addr[11857]= 876254528;
assign addr[11858]= 734482665;
assign addr[11859]= 588984994;
assign addr[11860]= 440499581;
assign addr[11861]= 289779648;
assign addr[11862]= 137589750;
assign addr[11863]= -15298099;
assign addr[11864]= -168108346;
assign addr[11865]= -320065829;
assign addr[11866]= -470399716;
assign addr[11867]= -618347408;
assign addr[11868]= -763158411;
assign addr[11869]= -904098143;
assign addr[11870]= -1040451659;
assign addr[11871]= -1171527280;
assign addr[11872]= -1296660098;
assign addr[11873]= -1415215352;
assign addr[11874]= -1526591649;
assign addr[11875]= -1630224009;
assign addr[11876]= -1725586737;
assign addr[11877]= -1812196087;
assign addr[11878]= -1889612716;
assign addr[11879]= -1957443913;
assign addr[11880]= -2015345591;
assign addr[11881]= -2063024031;
assign addr[11882]= -2100237377;
assign addr[11883]= -2126796855;
assign addr[11884]= -2142567738;
assign addr[11885]= -2147470025;
assign addr[11886]= -2141478848;
assign addr[11887]= -2124624598;
assign addr[11888]= -2096992772;
assign addr[11889]= -2058723538;
assign addr[11890]= -2010011024;
assign addr[11891]= -1951102334;
assign addr[11892]= -1882296293;
assign addr[11893]= -1803941934;
assign addr[11894]= -1716436725;
assign addr[11895]= -1620224553;
assign addr[11896]= -1515793473;
assign addr[11897]= -1403673233;
assign addr[11898]= -1284432584;
assign addr[11899]= -1158676398;
assign addr[11900]= -1027042599;
assign addr[11901]= -890198924;
assign addr[11902]= -748839539;
assign addr[11903]= -603681519;
assign addr[11904]= -455461206;
assign addr[11905]= -304930476;
assign addr[11906]= -152852926;
assign addr[11907]= 0;
assign addr[11908]= 152852926;
assign addr[11909]= 304930476;
assign addr[11910]= 455461206;
assign addr[11911]= 603681519;
assign addr[11912]= 748839539;
assign addr[11913]= 890198924;
assign addr[11914]= 1027042599;
assign addr[11915]= 1158676398;
assign addr[11916]= 1284432584;
assign addr[11917]= 1403673233;
assign addr[11918]= 1515793473;
assign addr[11919]= 1620224553;
assign addr[11920]= 1716436725;
assign addr[11921]= 1803941934;
assign addr[11922]= 1882296293;
assign addr[11923]= 1951102334;
assign addr[11924]= 2010011024;
assign addr[11925]= 2058723538;
assign addr[11926]= 2096992772;
assign addr[11927]= 2124624598;
assign addr[11928]= 2141478848;
assign addr[11929]= 2147470025;
assign addr[11930]= 2142567738;
assign addr[11931]= 2126796855;
assign addr[11932]= 2100237377;
assign addr[11933]= 2063024031;
assign addr[11934]= 2015345591;
assign addr[11935]= 1957443913;
assign addr[11936]= 1889612716;
assign addr[11937]= 1812196087;
assign addr[11938]= 1725586737;
assign addr[11939]= 1630224009;
assign addr[11940]= 1526591649;
assign addr[11941]= 1415215352;
assign addr[11942]= 1296660098;
assign addr[11943]= 1171527280;
assign addr[11944]= 1040451659;
assign addr[11945]= 904098143;
assign addr[11946]= 763158411;
assign addr[11947]= 618347408;
assign addr[11948]= 470399716;
assign addr[11949]= 320065829;
assign addr[11950]= 168108346;
assign addr[11951]= 15298099;
assign addr[11952]= -137589750;
assign addr[11953]= -289779648;
assign addr[11954]= -440499581;
assign addr[11955]= -588984994;
assign addr[11956]= -734482665;
assign addr[11957]= -876254528;
assign addr[11958]= -1013581418;
assign addr[11959]= -1145766716;
assign addr[11960]= -1272139887;
assign addr[11961]= -1392059879;
assign addr[11962]= -1504918373;
assign addr[11963]= -1610142873;
assign addr[11964]= -1707199606;
assign addr[11965]= -1795596234;
assign addr[11966]= -1874884346;
assign addr[11967]= -1944661739;
assign addr[11968]= -2004574453;
assign addr[11969]= -2054318569;
assign addr[11970]= -2093641749;
assign addr[11971]= -2122344521;
assign addr[11972]= -2140281282;
assign addr[11973]= -2147361045;
assign addr[11974]= -2143547897;
assign addr[11975]= -2128861181;
assign addr[11976]= -2103375398;
assign addr[11977]= -2067219829;
assign addr[11978]= -2020577882;
assign addr[11979]= -1963686155;
assign addr[11980]= -1896833245;
assign addr[11981]= -1820358275;
assign addr[11982]= -1734649179;
assign addr[11983]= -1640140734;
assign addr[11984]= -1537312353;
assign addr[11985]= -1426685652;
assign addr[11986]= -1308821808;
assign addr[11987]= -1184318708;
assign addr[11988]= -1053807919;
assign addr[11989]= -917951481;
assign addr[11990]= -777438554;
assign addr[11991]= -632981917;
assign addr[11992]= -485314355;
assign addr[11993]= -335184940;
assign addr[11994]= -183355234;
assign addr[11995]= -30595422;
assign addr[11996]= 122319591;
assign addr[11997]= 274614114;
assign addr[11998]= 425515602;
assign addr[11999]= 574258580;
assign addr[12000]= 720088517;
assign addr[12001]= 862265664;
assign addr[12002]= 1000068799;
assign addr[12003]= 1132798888;
assign addr[12004]= 1259782632;
assign addr[12005]= 1380375881;
assign addr[12006]= 1493966902;
assign addr[12007]= 1599979481;
assign addr[12008]= 1697875851;
assign addr[12009]= 1787159411;
assign addr[12010]= 1867377253;
assign addr[12011]= 1938122457;
assign addr[12012]= 1999036154;
assign addr[12013]= 2049809346;
assign addr[12014]= 2090184478;
assign addr[12015]= 2119956737;
assign addr[12016]= 2138975100;
assign addr[12017]= 2147143090;
assign addr[12018]= 2144419275;
assign addr[12019]= 2130817471;
assign addr[12020]= 2106406677;
assign addr[12021]= 2071310720;
assign addr[12022]= 2025707632;
assign addr[12023]= 1969828744;
assign addr[12024]= 1903957513;
assign addr[12025]= 1828428082;
assign addr[12026]= 1743623590;
assign addr[12027]= 1649974225;
assign addr[12028]= 1547955041;
assign addr[12029]= 1438083551;
assign addr[12030]= 1320917099;
assign addr[12031]= 1197050035;
assign addr[12032]= 1067110699;
assign addr[12033]= 931758235;
assign addr[12034]= 791679244;
assign addr[12035]= 647584304;
assign addr[12036]= 500204365;
assign addr[12037]= 350287041;
assign addr[12038]= 198592817;
assign addr[12039]= 45891193;
assign addr[12040]= -107043224;
assign addr[12041]= -259434643;
assign addr[12042]= -410510029;
assign addr[12043]= -559503022;
assign addr[12044]= -705657826;
assign addr[12045]= -848233042;
assign addr[12046]= -986505429;
assign addr[12047]= -1119773573;
assign addr[12048]= -1247361445;
assign addr[12049]= -1368621831;
assign addr[12050]= -1482939614;
assign addr[12051]= -1589734894;
assign addr[12052]= -1688465931;
assign addr[12053]= -1778631892;
assign addr[12054]= -1859775393;
assign addr[12055]= -1931484818;
assign addr[12056]= -1993396407;
assign addr[12057]= -2045196100;
assign addr[12058]= -2086621133;
assign addr[12059]= -2117461370;
assign addr[12060]= -2137560369;
assign addr[12061]= -2146816171;
assign addr[12062]= -2145181827;
assign addr[12063]= -2132665626;
assign addr[12064]= -2109331059;
assign addr[12065]= -2075296495;
assign addr[12066]= -2030734582;
assign addr[12067]= -1975871368;
assign addr[12068]= -1910985158;
assign addr[12069]= -1836405100;
assign addr[12070]= -1752509516;
assign addr[12071]= -1659723983;
assign addr[12072]= -1558519173;
assign addr[12073]= -1449408469;
assign addr[12074]= -1332945355;
assign addr[12075]= -1209720613;
assign addr[12076]= -1080359326;
assign addr[12077]= -945517704;
assign addr[12078]= -805879757;
assign addr[12079]= -662153826;
assign addr[12080]= -515068990;
assign addr[12081]= -365371365;
assign addr[12082]= -213820322;
assign addr[12083]= -61184634;
assign addr[12084]= 91761426;
assign addr[12085]= 244242007;
assign addr[12086]= 395483624;
assign addr[12087]= 544719071;
assign addr[12088]= 691191324;
assign addr[12089]= 834157373;
assign addr[12090]= 972891995;
assign addr[12091]= 1106691431;
assign addr[12092]= 1234876957;
assign addr[12093]= 1356798326;
assign addr[12094]= 1471837070;
assign addr[12095]= 1579409630;
assign addr[12096]= 1678970324;
assign addr[12097]= 1770014111;
assign addr[12098]= 1852079154;
assign addr[12099]= 1924749160;
assign addr[12100]= 1987655498;
assign addr[12101]= 2040479063;
assign addr[12102]= 2082951896;
assign addr[12103]= 2114858546;
assign addr[12104]= 2136037160;
assign addr[12105]= 2146380306;
assign addr[12106]= 2145835515;
assign addr[12107]= 2134405552;
assign addr[12108]= 2112148396;
assign addr[12109]= 2079176953;
assign addr[12110]= 2035658475;
assign addr[12111]= 1981813720;
assign addr[12112]= 1917915825;
assign addr[12113]= 1844288924;
assign addr[12114]= 1761306505;
assign addr[12115]= 1669389513;
assign addr[12116]= 1569004214;
assign addr[12117]= 1460659832;
assign addr[12118]= 1344905966;
assign addr[12119]= 1222329801;
assign addr[12120]= 1093553126;
assign addr[12121]= 959229189;
assign addr[12122]= 820039373;
assign addr[12123]= 676689746;
assign addr[12124]= 529907477;
assign addr[12125]= 380437148;
assign addr[12126]= 229036977;
assign addr[12127]= 76474970;
assign addr[12128]= -76474970;
assign addr[12129]= -229036977;
assign addr[12130]= -380437148;
assign addr[12131]= -529907477;
assign addr[12132]= -676689746;
assign addr[12133]= -820039373;
assign addr[12134]= -959229189;
assign addr[12135]= -1093553126;
assign addr[12136]= -1222329801;
assign addr[12137]= -1344905966;
assign addr[12138]= -1460659832;
assign addr[12139]= -1569004214;
assign addr[12140]= -1669389513;
assign addr[12141]= -1761306505;
assign addr[12142]= -1844288924;
assign addr[12143]= -1917915825;
assign addr[12144]= -1981813720;
assign addr[12145]= -2035658475;
assign addr[12146]= -2079176953;
assign addr[12147]= -2112148396;
assign addr[12148]= -2134405552;
assign addr[12149]= -2145835515;
assign addr[12150]= -2146380306;
assign addr[12151]= -2136037160;
assign addr[12152]= -2114858546;
assign addr[12153]= -2082951896;
assign addr[12154]= -2040479063;
assign addr[12155]= -1987655498;
assign addr[12156]= -1924749160;
assign addr[12157]= -1852079154;
assign addr[12158]= -1770014111;
assign addr[12159]= -1678970324;
assign addr[12160]= -1579409630;
assign addr[12161]= -1471837070;
assign addr[12162]= -1356798326;
assign addr[12163]= -1234876957;
assign addr[12164]= -1106691431;
assign addr[12165]= -972891995;
assign addr[12166]= -834157373;
assign addr[12167]= -691191324;
assign addr[12168]= -544719071;
assign addr[12169]= -395483624;
assign addr[12170]= -244242007;
assign addr[12171]= -91761426;
assign addr[12172]= 61184634;
assign addr[12173]= 213820322;
assign addr[12174]= 365371365;
assign addr[12175]= 515068990;
assign addr[12176]= 662153826;
assign addr[12177]= 805879757;
assign addr[12178]= 945517704;
assign addr[12179]= 1080359326;
assign addr[12180]= 1209720613;
assign addr[12181]= 1332945355;
assign addr[12182]= 1449408469;
assign addr[12183]= 1558519173;
assign addr[12184]= 1659723983;
assign addr[12185]= 1752509516;
assign addr[12186]= 1836405100;
assign addr[12187]= 1910985158;
assign addr[12188]= 1975871368;
assign addr[12189]= 2030734582;
assign addr[12190]= 2075296495;
assign addr[12191]= 2109331059;
assign addr[12192]= 2132665626;
assign addr[12193]= 2145181827;
assign addr[12194]= 2146816171;
assign addr[12195]= 2137560369;
assign addr[12196]= 2117461370;
assign addr[12197]= 2086621133;
assign addr[12198]= 2045196100;
assign addr[12199]= 1993396407;
assign addr[12200]= 1931484818;
assign addr[12201]= 1859775393;
assign addr[12202]= 1778631892;
assign addr[12203]= 1688465931;
assign addr[12204]= 1589734894;
assign addr[12205]= 1482939614;
assign addr[12206]= 1368621831;
assign addr[12207]= 1247361445;
assign addr[12208]= 1119773573;
assign addr[12209]= 986505429;
assign addr[12210]= 848233042;
assign addr[12211]= 705657826;
assign addr[12212]= 559503022;
assign addr[12213]= 410510029;
assign addr[12214]= 259434643;
assign addr[12215]= 107043224;
assign addr[12216]= -45891193;
assign addr[12217]= -198592817;
assign addr[12218]= -350287041;
assign addr[12219]= -500204365;
assign addr[12220]= -647584304;
assign addr[12221]= -791679244;
assign addr[12222]= -931758235;
assign addr[12223]= -1067110699;
assign addr[12224]= -1197050035;
assign addr[12225]= -1320917099;
assign addr[12226]= -1438083551;
assign addr[12227]= -1547955041;
assign addr[12228]= -1649974225;
assign addr[12229]= -1743623590;
assign addr[12230]= -1828428082;
assign addr[12231]= -1903957513;
assign addr[12232]= -1969828744;
assign addr[12233]= -2025707632;
assign addr[12234]= -2071310720;
assign addr[12235]= -2106406677;
assign addr[12236]= -2130817471;
assign addr[12237]= -2144419275;
assign addr[12238]= -2147143090;
assign addr[12239]= -2138975100;
assign addr[12240]= -2119956737;
assign addr[12241]= -2090184478;
assign addr[12242]= -2049809346;
assign addr[12243]= -1999036154;
assign addr[12244]= -1938122457;
assign addr[12245]= -1867377253;
assign addr[12246]= -1787159411;
assign addr[12247]= -1697875851;
assign addr[12248]= -1599979481;
assign addr[12249]= -1493966902;
assign addr[12250]= -1380375881;
assign addr[12251]= -1259782632;
assign addr[12252]= -1132798888;
assign addr[12253]= -1000068799;
assign addr[12254]= -862265664;
assign addr[12255]= -720088517;
assign addr[12256]= -574258580;
assign addr[12257]= -425515602;
assign addr[12258]= -274614114;
assign addr[12259]= -122319591;
assign addr[12260]= 30595422;
assign addr[12261]= 183355234;
assign addr[12262]= 335184940;
assign addr[12263]= 485314355;
assign addr[12264]= 632981917;
assign addr[12265]= 777438554;
assign addr[12266]= 917951481;
assign addr[12267]= 1053807919;
assign addr[12268]= 1184318708;
assign addr[12269]= 1308821808;
assign addr[12270]= 1426685652;
assign addr[12271]= 1537312353;
assign addr[12272]= 1640140734;
assign addr[12273]= 1734649179;
assign addr[12274]= 1820358275;
assign addr[12275]= 1896833245;
assign addr[12276]= 1963686155;
assign addr[12277]= 2020577882;
assign addr[12278]= 2067219829;
assign addr[12279]= 2103375398;
assign addr[12280]= 2128861181;
assign addr[12281]= 2143547897;
assign addr[12282]= 2147361045;
assign addr[12283]= 2140281282;
assign addr[12284]= 2122344521;
assign addr[12285]= 2093641749;
assign addr[12286]= 2054318569;
assign addr[12287]= 2004574453;
assign addr[12288]= 1944661739;
assign addr[12289]= 1874884346;
assign addr[12290]= 1795596234;
assign addr[12291]= 1707199606;
assign addr[12292]= 1610142873;
assign addr[12293]= 1504918373;
assign addr[12294]= 1392059879;
assign addr[12295]= 1272139887;
assign addr[12296]= 1145766716;
assign addr[12297]= 1013581418;
assign addr[12298]= 876254528;
assign addr[12299]= 734482665;
assign addr[12300]= 588984994;
assign addr[12301]= 440499581;
assign addr[12302]= 289779648;
assign addr[12303]= 137589750;
assign addr[12304]= -15298099;
assign addr[12305]= -168108346;
assign addr[12306]= -320065829;
assign addr[12307]= -470399716;
assign addr[12308]= -618347408;
assign addr[12309]= -763158411;
assign addr[12310]= -904098143;
assign addr[12311]= -1040451659;
assign addr[12312]= -1171527280;
assign addr[12313]= -1296660098;
assign addr[12314]= -1415215352;
assign addr[12315]= -1526591649;
assign addr[12316]= -1630224009;
assign addr[12317]= -1725586737;
assign addr[12318]= -1812196087;
assign addr[12319]= -1889612716;
assign addr[12320]= -1957443913;
assign addr[12321]= -2015345591;
assign addr[12322]= -2063024031;
assign addr[12323]= -2100237377;
assign addr[12324]= -2126796855;
assign addr[12325]= -2142567738;
assign addr[12326]= -2147470025;
assign addr[12327]= -2141478848;
assign addr[12328]= -2124624598;
assign addr[12329]= -2096992772;
assign addr[12330]= -2058723538;
assign addr[12331]= -2010011024;
assign addr[12332]= -1951102334;
assign addr[12333]= -1882296293;
assign addr[12334]= -1803941934;
assign addr[12335]= -1716436725;
assign addr[12336]= -1620224553;
assign addr[12337]= -1515793473;
assign addr[12338]= -1403673233;
assign addr[12339]= -1284432584;
assign addr[12340]= -1158676398;
assign addr[12341]= -1027042599;
assign addr[12342]= -890198924;
assign addr[12343]= -748839539;
assign addr[12344]= -603681519;
assign addr[12345]= -455461206;
assign addr[12346]= -304930476;
assign addr[12347]= -152852926;
assign addr[12348]= 0;
assign addr[12349]= 152852926;
assign addr[12350]= 304930476;
assign addr[12351]= 455461206;
assign addr[12352]= 603681519;
assign addr[12353]= 748839539;
assign addr[12354]= 890198924;
assign addr[12355]= 1027042599;
assign addr[12356]= 1158676398;
assign addr[12357]= 1284432584;
assign addr[12358]= 1403673233;
assign addr[12359]= 1515793473;
assign addr[12360]= 1620224553;
assign addr[12361]= 1716436725;
assign addr[12362]= 1803941934;
assign addr[12363]= 1882296293;
assign addr[12364]= 1951102334;
assign addr[12365]= 2010011024;
assign addr[12366]= 2058723538;
assign addr[12367]= 2096992772;
assign addr[12368]= 2124624598;
assign addr[12369]= 2141478848;
assign addr[12370]= 2147470025;
assign addr[12371]= 2142567738;
assign addr[12372]= 2126796855;
assign addr[12373]= 2100237377;
assign addr[12374]= 2063024031;
assign addr[12375]= 2015345591;
assign addr[12376]= 1957443913;
assign addr[12377]= 1889612716;
assign addr[12378]= 1812196087;
assign addr[12379]= 1725586737;
assign addr[12380]= 1630224009;
assign addr[12381]= 1526591649;
assign addr[12382]= 1415215352;
assign addr[12383]= 1296660098;
assign addr[12384]= 1171527280;
assign addr[12385]= 1040451659;
assign addr[12386]= 904098143;
assign addr[12387]= 763158411;
assign addr[12388]= 618347408;
assign addr[12389]= 470399716;
assign addr[12390]= 320065829;
assign addr[12391]= 168108346;
assign addr[12392]= 15298099;
assign addr[12393]= -137589750;
assign addr[12394]= -289779648;
assign addr[12395]= -440499581;
assign addr[12396]= -588984994;
assign addr[12397]= -734482665;
assign addr[12398]= -876254528;
assign addr[12399]= -1013581418;
assign addr[12400]= -1145766716;
assign addr[12401]= -1272139887;
assign addr[12402]= -1392059879;
assign addr[12403]= -1504918373;
assign addr[12404]= -1610142873;
assign addr[12405]= -1707199606;
assign addr[12406]= -1795596234;
assign addr[12407]= -1874884346;
assign addr[12408]= -1944661739;
assign addr[12409]= -2004574453;
assign addr[12410]= -2054318569;
assign addr[12411]= -2093641749;
assign addr[12412]= -2122344521;
assign addr[12413]= -2140281282;
assign addr[12414]= -2147361045;
assign addr[12415]= -2143547897;
assign addr[12416]= -2128861181;
assign addr[12417]= -2103375398;
assign addr[12418]= -2067219829;
assign addr[12419]= -2020577882;
assign addr[12420]= -1963686155;
assign addr[12421]= -1896833245;
assign addr[12422]= -1820358275;
assign addr[12423]= -1734649179;
assign addr[12424]= -1640140734;
assign addr[12425]= -1537312353;
assign addr[12426]= -1426685652;
assign addr[12427]= -1308821808;
assign addr[12428]= -1184318708;
assign addr[12429]= -1053807919;
assign addr[12430]= -917951481;
assign addr[12431]= -777438554;
assign addr[12432]= -632981917;
assign addr[12433]= -485314355;
assign addr[12434]= -335184940;
assign addr[12435]= -183355234;
assign addr[12436]= -30595422;
assign addr[12437]= 122319591;
assign addr[12438]= 274614114;
assign addr[12439]= 425515602;
assign addr[12440]= 574258580;
assign addr[12441]= 720088517;
assign addr[12442]= 862265664;
assign addr[12443]= 1000068799;
assign addr[12444]= 1132798888;
assign addr[12445]= 1259782632;
assign addr[12446]= 1380375881;
assign addr[12447]= 1493966902;
assign addr[12448]= 1599979481;
assign addr[12449]= 1697875851;
assign addr[12450]= 1787159411;
assign addr[12451]= 1867377253;
assign addr[12452]= 1938122457;
assign addr[12453]= 1999036154;
assign addr[12454]= 2049809346;
assign addr[12455]= 2090184478;
assign addr[12456]= 2119956737;
assign addr[12457]= 2138975100;
assign addr[12458]= 2147143090;
assign addr[12459]= 2144419275;
assign addr[12460]= 2130817471;
assign addr[12461]= 2106406677;
assign addr[12462]= 2071310720;
assign addr[12463]= 2025707632;
assign addr[12464]= 1969828744;
assign addr[12465]= 1903957513;
assign addr[12466]= 1828428082;
assign addr[12467]= 1743623590;
assign addr[12468]= 1649974225;
assign addr[12469]= 1547955041;
assign addr[12470]= 1438083551;
assign addr[12471]= 1320917099;
assign addr[12472]= 1197050035;
assign addr[12473]= 1067110699;
assign addr[12474]= 931758235;
assign addr[12475]= 791679244;
assign addr[12476]= 647584304;
assign addr[12477]= 500204365;
assign addr[12478]= 350287041;
assign addr[12479]= 198592817;
assign addr[12480]= 45891193;
assign addr[12481]= -107043224;
assign addr[12482]= -259434643;
assign addr[12483]= -410510029;
assign addr[12484]= -559503022;
assign addr[12485]= -705657826;
assign addr[12486]= -848233042;
assign addr[12487]= -986505429;
assign addr[12488]= -1119773573;
assign addr[12489]= -1247361445;
assign addr[12490]= -1368621831;
assign addr[12491]= -1482939614;
assign addr[12492]= -1589734894;
assign addr[12493]= -1688465931;
assign addr[12494]= -1778631892;
assign addr[12495]= -1859775393;
assign addr[12496]= -1931484818;
assign addr[12497]= -1993396407;
assign addr[12498]= -2045196100;
assign addr[12499]= -2086621133;
assign addr[12500]= -2117461370;
assign addr[12501]= -2137560369;
assign addr[12502]= -2146816171;
assign addr[12503]= -2145181827;
assign addr[12504]= -2132665626;
assign addr[12505]= -2109331059;
assign addr[12506]= -2075296495;
assign addr[12507]= -2030734582;
assign addr[12508]= -1975871368;
assign addr[12509]= -1910985158;
assign addr[12510]= -1836405100;
assign addr[12511]= -1752509516;
assign addr[12512]= -1659723983;
assign addr[12513]= -1558519173;
assign addr[12514]= -1449408469;
assign addr[12515]= -1332945355;
assign addr[12516]= -1209720613;
assign addr[12517]= -1080359326;
assign addr[12518]= -945517704;
assign addr[12519]= -805879757;
assign addr[12520]= -662153826;
assign addr[12521]= -515068990;
assign addr[12522]= -365371365;
assign addr[12523]= -213820322;
assign addr[12524]= -61184634;
assign addr[12525]= 91761426;
assign addr[12526]= 244242007;
assign addr[12527]= 395483624;
assign addr[12528]= 544719071;
assign addr[12529]= 691191324;
assign addr[12530]= 834157373;
assign addr[12531]= 972891995;
assign addr[12532]= 1106691431;
assign addr[12533]= 1234876957;
assign addr[12534]= 1356798326;
assign addr[12535]= 1471837070;
assign addr[12536]= 1579409630;
assign addr[12537]= 1678970324;
assign addr[12538]= 1770014111;
assign addr[12539]= 1852079154;
assign addr[12540]= 1924749160;
assign addr[12541]= 1987655498;
assign addr[12542]= 2040479063;
assign addr[12543]= 2082951896;
assign addr[12544]= 2114858546;
assign addr[12545]= 2136037160;
assign addr[12546]= 2146380306;
assign addr[12547]= 2145835515;
assign addr[12548]= 2134405552;
assign addr[12549]= 2112148396;
assign addr[12550]= 2079176953;
assign addr[12551]= 2035658475;
assign addr[12552]= 1981813720;
assign addr[12553]= 1917915825;
assign addr[12554]= 1844288924;
assign addr[12555]= 1761306505;
assign addr[12556]= 1669389513;
assign addr[12557]= 1569004214;
assign addr[12558]= 1460659832;
assign addr[12559]= 1344905966;
assign addr[12560]= 1222329801;
assign addr[12561]= 1093553126;
assign addr[12562]= 959229189;
assign addr[12563]= 820039373;
assign addr[12564]= 676689746;
assign addr[12565]= 529907477;
assign addr[12566]= 380437148;
assign addr[12567]= 229036977;
assign addr[12568]= 76474970;
assign addr[12569]= -76474970;
assign addr[12570]= -229036977;
assign addr[12571]= -380437148;
assign addr[12572]= -529907477;
assign addr[12573]= -676689746;
assign addr[12574]= -820039373;
assign addr[12575]= -959229189;
assign addr[12576]= -1093553126;
assign addr[12577]= -1222329801;
assign addr[12578]= -1344905966;
assign addr[12579]= -1460659832;
assign addr[12580]= -1569004214;
assign addr[12581]= -1669389513;
assign addr[12582]= -1761306505;
assign addr[12583]= -1844288924;
assign addr[12584]= -1917915825;
assign addr[12585]= -1981813720;
assign addr[12586]= -2035658475;
assign addr[12587]= -2079176953;
assign addr[12588]= -2112148396;
assign addr[12589]= -2134405552;
assign addr[12590]= -2145835515;
assign addr[12591]= -2146380306;
assign addr[12592]= -2136037160;
assign addr[12593]= -2114858546;
assign addr[12594]= -2082951896;
assign addr[12595]= -2040479063;
assign addr[12596]= -1987655498;
assign addr[12597]= -1924749160;
assign addr[12598]= -1852079154;
assign addr[12599]= -1770014111;
assign addr[12600]= -1678970324;
assign addr[12601]= -1579409630;
assign addr[12602]= -1471837070;
assign addr[12603]= -1356798326;
assign addr[12604]= -1234876957;
assign addr[12605]= -1106691431;
assign addr[12606]= -972891995;
assign addr[12607]= -834157373;
assign addr[12608]= -691191324;
assign addr[12609]= -544719071;
assign addr[12610]= -395483624;
assign addr[12611]= -244242007;
assign addr[12612]= -91761426;
assign addr[12613]= 61184634;
assign addr[12614]= 213820322;
assign addr[12615]= 365371365;
assign addr[12616]= 515068990;
assign addr[12617]= 662153826;
assign addr[12618]= 805879757;
assign addr[12619]= 945517704;
assign addr[12620]= 1080359326;
assign addr[12621]= 1209720613;
assign addr[12622]= 1332945355;
assign addr[12623]= 1449408469;
assign addr[12624]= 1558519173;
assign addr[12625]= 1659723983;
assign addr[12626]= 1752509516;
assign addr[12627]= 1836405100;
assign addr[12628]= 1910985158;
assign addr[12629]= 1975871368;
assign addr[12630]= 2030734582;
assign addr[12631]= 2075296495;
assign addr[12632]= 2109331059;
assign addr[12633]= 2132665626;
assign addr[12634]= 2145181827;
assign addr[12635]= 2146816171;
assign addr[12636]= 2137560369;
assign addr[12637]= 2117461370;
assign addr[12638]= 2086621133;
assign addr[12639]= 2045196100;
assign addr[12640]= 1993396407;
assign addr[12641]= 1931484818;
assign addr[12642]= 1859775393;
assign addr[12643]= 1778631892;
assign addr[12644]= 1688465931;
assign addr[12645]= 1589734894;
assign addr[12646]= 1482939614;
assign addr[12647]= 1368621831;
assign addr[12648]= 1247361445;
assign addr[12649]= 1119773573;
assign addr[12650]= 986505429;
assign addr[12651]= 848233042;
assign addr[12652]= 705657826;
assign addr[12653]= 559503022;
assign addr[12654]= 410510029;
assign addr[12655]= 259434643;
assign addr[12656]= 107043224;
assign addr[12657]= -45891193;
assign addr[12658]= -198592817;
assign addr[12659]= -350287041;
assign addr[12660]= -500204365;
assign addr[12661]= -647584304;
assign addr[12662]= -791679244;
assign addr[12663]= -931758235;
assign addr[12664]= -1067110699;
assign addr[12665]= -1197050035;
assign addr[12666]= -1320917099;
assign addr[12667]= -1438083551;
assign addr[12668]= -1547955041;
assign addr[12669]= -1649974225;
assign addr[12670]= -1743623590;
assign addr[12671]= -1828428082;
assign addr[12672]= -1903957513;
assign addr[12673]= -1969828744;
assign addr[12674]= -2025707632;
assign addr[12675]= -2071310720;
assign addr[12676]= -2106406677;
assign addr[12677]= -2130817471;
assign addr[12678]= -2144419275;
assign addr[12679]= -2147143090;
assign addr[12680]= -2138975100;
assign addr[12681]= -2119956737;
assign addr[12682]= -2090184478;
assign addr[12683]= -2049809346;
assign addr[12684]= -1999036154;
assign addr[12685]= -1938122457;
assign addr[12686]= -1867377253;
assign addr[12687]= -1787159411;
assign addr[12688]= -1697875851;
assign addr[12689]= -1599979481;
assign addr[12690]= -1493966902;
assign addr[12691]= -1380375881;
assign addr[12692]= -1259782632;
assign addr[12693]= -1132798888;
assign addr[12694]= -1000068799;
assign addr[12695]= -862265664;
assign addr[12696]= -720088517;
assign addr[12697]= -574258580;
assign addr[12698]= -425515602;
assign addr[12699]= -274614114;
assign addr[12700]= -122319591;
assign addr[12701]= 30595422;
assign addr[12702]= 183355234;
assign addr[12703]= 335184940;
assign addr[12704]= 485314355;
assign addr[12705]= 632981917;
assign addr[12706]= 777438554;
assign addr[12707]= 917951481;
assign addr[12708]= 1053807919;
assign addr[12709]= 1184318708;
assign addr[12710]= 1308821808;
assign addr[12711]= 1426685652;
assign addr[12712]= 1537312353;
assign addr[12713]= 1640140734;
assign addr[12714]= 1734649179;
assign addr[12715]= 1820358275;
assign addr[12716]= 1896833245;
assign addr[12717]= 1963686155;
assign addr[12718]= 2020577882;
assign addr[12719]= 2067219829;
assign addr[12720]= 2103375398;
assign addr[12721]= 2128861181;
assign addr[12722]= 2143547897;
assign addr[12723]= 2147361045;
assign addr[12724]= 2140281282;
assign addr[12725]= 2122344521;
assign addr[12726]= 2093641749;
assign addr[12727]= 2054318569;
assign addr[12728]= 2004574453;
assign addr[12729]= 1944661739;
assign addr[12730]= 1874884346;
assign addr[12731]= 1795596234;
assign addr[12732]= 1707199606;
assign addr[12733]= 1610142873;
assign addr[12734]= 1504918373;
assign addr[12735]= 1392059879;
assign addr[12736]= 1272139887;
assign addr[12737]= 1145766716;
assign addr[12738]= 1013581418;
assign addr[12739]= 876254528;
assign addr[12740]= 734482665;
assign addr[12741]= 588984994;
assign addr[12742]= 440499581;
assign addr[12743]= 289779648;
assign addr[12744]= 137589750;
assign addr[12745]= -15298099;
assign addr[12746]= -168108346;
assign addr[12747]= -320065829;
assign addr[12748]= -470399716;
assign addr[12749]= -618347408;
assign addr[12750]= -763158411;
assign addr[12751]= -904098143;
assign addr[12752]= -1040451659;
assign addr[12753]= -1171527280;
assign addr[12754]= -1296660098;
assign addr[12755]= -1415215352;
assign addr[12756]= -1526591649;
assign addr[12757]= -1630224009;
assign addr[12758]= -1725586737;
assign addr[12759]= -1812196087;
assign addr[12760]= -1889612716;
assign addr[12761]= -1957443913;
assign addr[12762]= -2015345591;
assign addr[12763]= -2063024031;
assign addr[12764]= -2100237377;
assign addr[12765]= -2126796855;
assign addr[12766]= -2142567738;
assign addr[12767]= -2147470025;
assign addr[12768]= -2141478848;
assign addr[12769]= -2124624598;
assign addr[12770]= -2096992772;
assign addr[12771]= -2058723538;
assign addr[12772]= -2010011024;
assign addr[12773]= -1951102334;
assign addr[12774]= -1882296293;
assign addr[12775]= -1803941934;
assign addr[12776]= -1716436725;
assign addr[12777]= -1620224553;
assign addr[12778]= -1515793473;
assign addr[12779]= -1403673233;
assign addr[12780]= -1284432584;
assign addr[12781]= -1158676398;
assign addr[12782]= -1027042599;
assign addr[12783]= -890198924;
assign addr[12784]= -748839539;
assign addr[12785]= -603681519;
assign addr[12786]= -455461206;
assign addr[12787]= -304930476;
assign addr[12788]= -152852926;
assign addr[12789]= 0;
assign addr[12790]= 152852926;
assign addr[12791]= 304930476;
assign addr[12792]= 455461206;
assign addr[12793]= 603681519;
assign addr[12794]= 748839539;
assign addr[12795]= 890198924;
assign addr[12796]= 1027042599;
assign addr[12797]= 1158676398;
assign addr[12798]= 1284432584;
assign addr[12799]= 1403673233;
assign addr[12800]= 1515793473;
assign addr[12801]= 1620224553;
assign addr[12802]= 1716436725;
assign addr[12803]= 1803941934;
assign addr[12804]= 1882296293;
assign addr[12805]= 1951102334;
assign addr[12806]= 2010011024;
assign addr[12807]= 2058723538;
assign addr[12808]= 2096992772;
assign addr[12809]= 2124624598;
assign addr[12810]= 2141478848;
assign addr[12811]= 2147470025;
assign addr[12812]= 2142567738;
assign addr[12813]= 2126796855;
assign addr[12814]= 2100237377;
assign addr[12815]= 2063024031;
assign addr[12816]= 2015345591;
assign addr[12817]= 1957443913;
assign addr[12818]= 1889612716;
assign addr[12819]= 1812196087;
assign addr[12820]= 1725586737;
assign addr[12821]= 1630224009;
assign addr[12822]= 1526591649;
assign addr[12823]= 1415215352;
assign addr[12824]= 1296660098;
assign addr[12825]= 1171527280;
assign addr[12826]= 1040451659;
assign addr[12827]= 904098143;
assign addr[12828]= 763158411;
assign addr[12829]= 618347408;
assign addr[12830]= 470399716;
assign addr[12831]= 320065829;
assign addr[12832]= 168108346;
assign addr[12833]= 15298099;
assign addr[12834]= -137589750;
assign addr[12835]= -289779648;
assign addr[12836]= -440499581;
assign addr[12837]= -588984994;
assign addr[12838]= -734482665;
assign addr[12839]= -876254528;
assign addr[12840]= -1013581418;
assign addr[12841]= -1145766716;
assign addr[12842]= -1272139887;
assign addr[12843]= -1392059879;
assign addr[12844]= -1504918373;
assign addr[12845]= -1610142873;
assign addr[12846]= -1707199606;
assign addr[12847]= -1795596234;
assign addr[12848]= -1874884346;
assign addr[12849]= -1944661739;
assign addr[12850]= -2004574453;
assign addr[12851]= -2054318569;
assign addr[12852]= -2093641749;
assign addr[12853]= -2122344521;
assign addr[12854]= -2140281282;
assign addr[12855]= -2147361045;
assign addr[12856]= -2143547897;
assign addr[12857]= -2128861181;
assign addr[12858]= -2103375398;
assign addr[12859]= -2067219829;
assign addr[12860]= -2020577882;
assign addr[12861]= -1963686155;
assign addr[12862]= -1896833245;
assign addr[12863]= -1820358275;
assign addr[12864]= -1734649179;
assign addr[12865]= -1640140734;
assign addr[12866]= -1537312353;
assign addr[12867]= -1426685652;
assign addr[12868]= -1308821808;
assign addr[12869]= -1184318708;
assign addr[12870]= -1053807919;
assign addr[12871]= -917951481;
assign addr[12872]= -777438554;
assign addr[12873]= -632981917;
assign addr[12874]= -485314355;
assign addr[12875]= -335184940;
assign addr[12876]= -183355234;
assign addr[12877]= -30595422;
assign addr[12878]= 122319591;
assign addr[12879]= 274614114;
assign addr[12880]= 425515602;
assign addr[12881]= 574258580;
assign addr[12882]= 720088517;
assign addr[12883]= 862265664;
assign addr[12884]= 1000068799;
assign addr[12885]= 1132798888;
assign addr[12886]= 1259782632;
assign addr[12887]= 1380375881;
assign addr[12888]= 1493966902;
assign addr[12889]= 1599979481;
assign addr[12890]= 1697875851;
assign addr[12891]= 1787159411;
assign addr[12892]= 1867377253;
assign addr[12893]= 1938122457;
assign addr[12894]= 1999036154;
assign addr[12895]= 2049809346;
assign addr[12896]= 2090184478;
assign addr[12897]= 2119956737;
assign addr[12898]= 2138975100;
assign addr[12899]= 2147143090;
assign addr[12900]= 2144419275;
assign addr[12901]= 2130817471;
assign addr[12902]= 2106406677;
assign addr[12903]= 2071310720;
assign addr[12904]= 2025707632;
assign addr[12905]= 1969828744;
assign addr[12906]= 1903957513;
assign addr[12907]= 1828428082;
assign addr[12908]= 1743623590;
assign addr[12909]= 1649974225;
assign addr[12910]= 1547955041;
assign addr[12911]= 1438083551;
assign addr[12912]= 1320917099;
assign addr[12913]= 1197050035;
assign addr[12914]= 1067110699;
assign addr[12915]= 931758235;
assign addr[12916]= 791679244;
assign addr[12917]= 647584304;
assign addr[12918]= 500204365;
assign addr[12919]= 350287041;
assign addr[12920]= 198592817;
assign addr[12921]= 45891193;
assign addr[12922]= -107043224;
assign addr[12923]= -259434643;
assign addr[12924]= -410510029;
assign addr[12925]= -559503022;
assign addr[12926]= -705657826;
assign addr[12927]= -848233042;
assign addr[12928]= -986505429;
assign addr[12929]= -1119773573;
assign addr[12930]= -1247361445;
assign addr[12931]= -1368621831;
assign addr[12932]= -1482939614;
assign addr[12933]= -1589734894;
assign addr[12934]= -1688465931;
assign addr[12935]= -1778631892;
assign addr[12936]= -1859775393;
assign addr[12937]= -1931484818;
assign addr[12938]= -1993396407;
assign addr[12939]= -2045196100;
assign addr[12940]= -2086621133;
assign addr[12941]= -2117461370;
assign addr[12942]= -2137560369;
assign addr[12943]= -2146816171;
assign addr[12944]= -2145181827;
assign addr[12945]= -2132665626;
assign addr[12946]= -2109331059;
assign addr[12947]= -2075296495;
assign addr[12948]= -2030734582;
assign addr[12949]= -1975871368;
assign addr[12950]= -1910985158;
assign addr[12951]= -1836405100;
assign addr[12952]= -1752509516;
assign addr[12953]= -1659723983;
assign addr[12954]= -1558519173;
assign addr[12955]= -1449408469;
assign addr[12956]= -1332945355;
assign addr[12957]= -1209720613;
assign addr[12958]= -1080359326;
assign addr[12959]= -945517704;
assign addr[12960]= -805879757;
assign addr[12961]= -662153826;
assign addr[12962]= -515068990;
assign addr[12963]= -365371365;
assign addr[12964]= -213820322;
assign addr[12965]= -61184634;
assign addr[12966]= 91761426;
assign addr[12967]= 244242007;
assign addr[12968]= 395483624;
assign addr[12969]= 544719071;
assign addr[12970]= 691191324;
assign addr[12971]= 834157373;
assign addr[12972]= 972891995;
assign addr[12973]= 1106691431;
assign addr[12974]= 1234876957;
assign addr[12975]= 1356798326;
assign addr[12976]= 1471837070;
assign addr[12977]= 1579409630;
assign addr[12978]= 1678970324;
assign addr[12979]= 1770014111;
assign addr[12980]= 1852079154;
assign addr[12981]= 1924749160;
assign addr[12982]= 1987655498;
assign addr[12983]= 2040479063;
assign addr[12984]= 2082951896;
assign addr[12985]= 2114858546;
assign addr[12986]= 2136037160;
assign addr[12987]= 2146380306;
assign addr[12988]= 2145835515;
assign addr[12989]= 2134405552;
assign addr[12990]= 2112148396;
assign addr[12991]= 2079176953;
assign addr[12992]= 2035658475;
assign addr[12993]= 1981813720;
assign addr[12994]= 1917915825;
assign addr[12995]= 1844288924;
assign addr[12996]= 1761306505;
assign addr[12997]= 1669389513;
assign addr[12998]= 1569004214;
assign addr[12999]= 1460659832;
assign addr[13000]= 1344905966;
assign addr[13001]= 1222329801;
assign addr[13002]= 1093553126;
assign addr[13003]= 959229189;
assign addr[13004]= 820039373;
assign addr[13005]= 676689746;
assign addr[13006]= 529907477;
assign addr[13007]= 380437148;
assign addr[13008]= 229036977;
assign addr[13009]= 76474970;
assign addr[13010]= -76474970;
assign addr[13011]= -229036977;
assign addr[13012]= -380437148;
assign addr[13013]= -529907477;
assign addr[13014]= -676689746;
assign addr[13015]= -820039373;
assign addr[13016]= -959229189;
assign addr[13017]= -1093553126;
assign addr[13018]= -1222329801;
assign addr[13019]= -1344905966;
assign addr[13020]= -1460659832;
assign addr[13021]= -1569004214;
assign addr[13022]= -1669389513;
assign addr[13023]= -1761306505;
assign addr[13024]= -1844288924;
assign addr[13025]= -1917915825;
assign addr[13026]= -1981813720;
assign addr[13027]= -2035658475;
assign addr[13028]= -2079176953;
assign addr[13029]= -2112148396;
assign addr[13030]= -2134405552;
assign addr[13031]= -2145835515;
assign addr[13032]= -2146380306;
assign addr[13033]= -2136037160;
assign addr[13034]= -2114858546;
assign addr[13035]= -2082951896;
assign addr[13036]= -2040479063;
assign addr[13037]= -1987655498;
assign addr[13038]= -1924749160;
assign addr[13039]= -1852079154;
assign addr[13040]= -1770014111;
assign addr[13041]= -1678970324;
assign addr[13042]= -1579409630;
assign addr[13043]= -1471837070;
assign addr[13044]= -1356798326;
assign addr[13045]= -1234876957;
assign addr[13046]= -1106691431;
assign addr[13047]= -972891995;
assign addr[13048]= -834157373;
assign addr[13049]= -691191324;
assign addr[13050]= -544719071;
assign addr[13051]= -395483624;
assign addr[13052]= -244242007;
assign addr[13053]= -91761426;
assign addr[13054]= 61184634;
assign addr[13055]= 213820322;
assign addr[13056]= 365371365;
assign addr[13057]= 515068990;
assign addr[13058]= 662153826;
assign addr[13059]= 805879757;
assign addr[13060]= 945517704;
assign addr[13061]= 1080359326;
assign addr[13062]= 1209720613;
assign addr[13063]= 1332945355;
assign addr[13064]= 1449408469;
assign addr[13065]= 1558519173;
assign addr[13066]= 1659723983;
assign addr[13067]= 1752509516;
assign addr[13068]= 1836405100;
assign addr[13069]= 1910985158;
assign addr[13070]= 1975871368;
assign addr[13071]= 2030734582;
assign addr[13072]= 2075296495;
assign addr[13073]= 2109331059;
assign addr[13074]= 2132665626;
assign addr[13075]= 2145181827;
assign addr[13076]= 2146816171;
assign addr[13077]= 2137560369;
assign addr[13078]= 2117461370;
assign addr[13079]= 2086621133;
assign addr[13080]= 2045196100;
assign addr[13081]= 1993396407;
assign addr[13082]= 1931484818;
assign addr[13083]= 1859775393;
assign addr[13084]= 1778631892;
assign addr[13085]= 1688465931;
assign addr[13086]= 1589734894;
assign addr[13087]= 1482939614;
assign addr[13088]= 1368621831;
assign addr[13089]= 1247361445;
assign addr[13090]= 1119773573;
assign addr[13091]= 986505429;
assign addr[13092]= 848233042;
assign addr[13093]= 705657826;
assign addr[13094]= 559503022;
assign addr[13095]= 410510029;
assign addr[13096]= 259434643;
assign addr[13097]= 107043224;
assign addr[13098]= -45891193;
assign addr[13099]= -198592817;
assign addr[13100]= -350287041;
assign addr[13101]= -500204365;
assign addr[13102]= -647584304;
assign addr[13103]= -791679244;
assign addr[13104]= -931758235;
assign addr[13105]= -1067110699;
assign addr[13106]= -1197050035;
assign addr[13107]= -1320917099;
assign addr[13108]= -1438083551;
assign addr[13109]= -1547955041;
assign addr[13110]= -1649974225;
assign addr[13111]= -1743623590;
assign addr[13112]= -1828428082;
assign addr[13113]= -1903957513;
assign addr[13114]= -1969828744;
assign addr[13115]= -2025707632;
assign addr[13116]= -2071310720;
assign addr[13117]= -2106406677;
assign addr[13118]= -2130817471;
assign addr[13119]= -2144419275;
assign addr[13120]= -2147143090;
assign addr[13121]= -2138975100;
assign addr[13122]= -2119956737;
assign addr[13123]= -2090184478;
assign addr[13124]= -2049809346;
assign addr[13125]= -1999036154;
assign addr[13126]= -1938122457;
assign addr[13127]= -1867377253;
assign addr[13128]= -1787159411;
assign addr[13129]= -1697875851;
assign addr[13130]= -1599979481;
assign addr[13131]= -1493966902;
assign addr[13132]= -1380375881;
assign addr[13133]= -1259782632;
assign addr[13134]= -1132798888;
assign addr[13135]= -1000068799;
assign addr[13136]= -862265664;
assign addr[13137]= -720088517;
assign addr[13138]= -574258580;
assign addr[13139]= -425515602;
assign addr[13140]= -274614114;
assign addr[13141]= -122319591;
assign addr[13142]= 30595422;
assign addr[13143]= 183355234;
assign addr[13144]= 335184940;
assign addr[13145]= 485314355;
assign addr[13146]= 632981917;
assign addr[13147]= 777438554;
assign addr[13148]= 917951481;
assign addr[13149]= 1053807919;
assign addr[13150]= 1184318708;
assign addr[13151]= 1308821808;
assign addr[13152]= 1426685652;
assign addr[13153]= 1537312353;
assign addr[13154]= 1640140734;
assign addr[13155]= 1734649179;
assign addr[13156]= 1820358275;
assign addr[13157]= 1896833245;
assign addr[13158]= 1963686155;
assign addr[13159]= 2020577882;
assign addr[13160]= 2067219829;
assign addr[13161]= 2103375398;
assign addr[13162]= 2128861181;
assign addr[13163]= 2143547897;
assign addr[13164]= 2147361045;
assign addr[13165]= 2140281282;
assign addr[13166]= 2122344521;
assign addr[13167]= 2093641749;
assign addr[13168]= 2054318569;
assign addr[13169]= 2004574453;
assign addr[13170]= 1944661739;
assign addr[13171]= 1874884346;
assign addr[13172]= 1795596234;
assign addr[13173]= 1707199606;
assign addr[13174]= 1610142873;
assign addr[13175]= 1504918373;
assign addr[13176]= 1392059879;
assign addr[13177]= 1272139887;
assign addr[13178]= 1145766716;
assign addr[13179]= 1013581418;
assign addr[13180]= 876254528;
assign addr[13181]= 734482665;
assign addr[13182]= 588984994;
assign addr[13183]= 440499581;
assign addr[13184]= 289779648;
assign addr[13185]= 137589750;
assign addr[13186]= -15298099;
assign addr[13187]= -168108346;
assign addr[13188]= -320065829;
assign addr[13189]= -470399716;
assign addr[13190]= -618347408;
assign addr[13191]= -763158411;
assign addr[13192]= -904098143;
assign addr[13193]= -1040451659;
assign addr[13194]= -1171527280;
assign addr[13195]= -1296660098;
assign addr[13196]= -1415215352;
assign addr[13197]= -1526591649;
assign addr[13198]= -1630224009;
assign addr[13199]= -1725586737;
assign addr[13200]= -1812196087;
assign addr[13201]= -1889612716;
assign addr[13202]= -1957443913;
assign addr[13203]= -2015345591;
assign addr[13204]= -2063024031;
assign addr[13205]= -2100237377;
assign addr[13206]= -2126796855;
assign addr[13207]= -2142567738;
assign addr[13208]= -2147470025;
assign addr[13209]= -2141478848;
assign addr[13210]= -2124624598;
assign addr[13211]= -2096992772;
assign addr[13212]= -2058723538;
assign addr[13213]= -2010011024;
assign addr[13214]= -1951102334;
assign addr[13215]= -1882296293;
assign addr[13216]= -1803941934;
assign addr[13217]= -1716436725;
assign addr[13218]= -1620224553;
assign addr[13219]= -1515793473;
assign addr[13220]= -1403673233;
assign addr[13221]= -1284432584;
assign addr[13222]= -1158676398;
assign addr[13223]= -1027042599;
assign addr[13224]= -890198924;
assign addr[13225]= -748839539;
assign addr[13226]= -603681519;
assign addr[13227]= -455461206;
assign addr[13228]= -304930476;
assign addr[13229]= -152852926;
assign addr[13230]= 0;
assign addr[13231]= 152852926;
assign addr[13232]= 304930476;
assign addr[13233]= 455461206;
assign addr[13234]= 603681519;
assign addr[13235]= 748839539;
assign addr[13236]= 890198924;
assign addr[13237]= 1027042599;
assign addr[13238]= 1158676398;
assign addr[13239]= 1284432584;
assign addr[13240]= 1403673233;
assign addr[13241]= 1515793473;
assign addr[13242]= 1620224553;
assign addr[13243]= 1716436725;
assign addr[13244]= 1803941934;
assign addr[13245]= 1882296293;
assign addr[13246]= 1951102334;
assign addr[13247]= 2010011024;
assign addr[13248]= 2058723538;
assign addr[13249]= 2096992772;
assign addr[13250]= 2124624598;
assign addr[13251]= 2141478848;
assign addr[13252]= 2147470025;
assign addr[13253]= 2142567738;
assign addr[13254]= 2126796855;
assign addr[13255]= 2100237377;
assign addr[13256]= 2063024031;
assign addr[13257]= 2015345591;
assign addr[13258]= 1957443913;
assign addr[13259]= 1889612716;
assign addr[13260]= 1812196087;
assign addr[13261]= 1725586737;
assign addr[13262]= 1630224009;
assign addr[13263]= 1526591649;
assign addr[13264]= 1415215352;
assign addr[13265]= 1296660098;
assign addr[13266]= 1171527280;
assign addr[13267]= 1040451659;
assign addr[13268]= 904098143;
assign addr[13269]= 763158411;
assign addr[13270]= 618347408;
assign addr[13271]= 470399716;
assign addr[13272]= 320065829;
assign addr[13273]= 168108346;
assign addr[13274]= 15298099;
assign addr[13275]= -137589750;
assign addr[13276]= -289779648;
assign addr[13277]= -440499581;
assign addr[13278]= -588984994;
assign addr[13279]= -734482665;
assign addr[13280]= -876254528;
assign addr[13281]= -1013581418;
assign addr[13282]= -1145766716;
assign addr[13283]= -1272139887;
assign addr[13284]= -1392059879;
assign addr[13285]= -1504918373;
assign addr[13286]= -1610142873;
assign addr[13287]= -1707199606;
assign addr[13288]= -1795596234;
assign addr[13289]= -1874884346;
assign addr[13290]= -1944661739;
assign addr[13291]= -2004574453;
assign addr[13292]= -2054318569;
assign addr[13293]= -2093641749;
assign addr[13294]= -2122344521;
assign addr[13295]= -2140281282;
assign addr[13296]= -2147361045;
assign addr[13297]= -2143547897;
assign addr[13298]= -2128861181;
assign addr[13299]= -2103375398;
assign addr[13300]= -2067219829;
assign addr[13301]= -2020577882;
assign addr[13302]= -1963686155;
assign addr[13303]= -1896833245;
assign addr[13304]= -1820358275;
assign addr[13305]= -1734649179;
assign addr[13306]= -1640140734;
assign addr[13307]= -1537312353;
assign addr[13308]= -1426685652;
assign addr[13309]= -1308821808;
assign addr[13310]= -1184318708;
assign addr[13311]= -1053807919;
assign addr[13312]= -917951481;
assign addr[13313]= -777438554;
assign addr[13314]= -632981917;
assign addr[13315]= -485314355;
assign addr[13316]= -335184940;
assign addr[13317]= -183355234;
assign addr[13318]= -30595422;
assign addr[13319]= 122319591;
assign addr[13320]= 274614114;
assign addr[13321]= 425515602;
assign addr[13322]= 574258580;
assign addr[13323]= 720088517;
assign addr[13324]= 862265664;
assign addr[13325]= 1000068799;
assign addr[13326]= 1132798888;
assign addr[13327]= 1259782632;
assign addr[13328]= 1380375881;
assign addr[13329]= 1493966902;
assign addr[13330]= 1599979481;
assign addr[13331]= 1697875851;
assign addr[13332]= 1787159411;
assign addr[13333]= 1867377253;
assign addr[13334]= 1938122457;
assign addr[13335]= 1999036154;
assign addr[13336]= 2049809346;
assign addr[13337]= 2090184478;
assign addr[13338]= 2119956737;
assign addr[13339]= 2138975100;
assign addr[13340]= 2147143090;
assign addr[13341]= 2144419275;
assign addr[13342]= 2130817471;
assign addr[13343]= 2106406677;
assign addr[13344]= 2071310720;
assign addr[13345]= 2025707632;
assign addr[13346]= 1969828744;
assign addr[13347]= 1903957513;
assign addr[13348]= 1828428082;
assign addr[13349]= 1743623590;
assign addr[13350]= 1649974225;
assign addr[13351]= 1547955041;
assign addr[13352]= 1438083551;
assign addr[13353]= 1320917099;
assign addr[13354]= 1197050035;
assign addr[13355]= 1067110699;
assign addr[13356]= 931758235;
assign addr[13357]= 791679244;
assign addr[13358]= 647584304;
assign addr[13359]= 500204365;
assign addr[13360]= 350287041;
assign addr[13361]= 198592817;
assign addr[13362]= 45891193;
assign addr[13363]= -107043224;
assign addr[13364]= -259434643;
assign addr[13365]= -410510029;
assign addr[13366]= -559503022;
assign addr[13367]= -705657826;
assign addr[13368]= -848233042;
assign addr[13369]= -986505429;
assign addr[13370]= -1119773573;
assign addr[13371]= -1247361445;
assign addr[13372]= -1368621831;
assign addr[13373]= -1482939614;
assign addr[13374]= -1589734894;
assign addr[13375]= -1688465931;
assign addr[13376]= -1778631892;
assign addr[13377]= -1859775393;
assign addr[13378]= -1931484818;
assign addr[13379]= -1993396407;
assign addr[13380]= -2045196100;
assign addr[13381]= -2086621133;
assign addr[13382]= -2117461370;
assign addr[13383]= -2137560369;
assign addr[13384]= -2146816171;
assign addr[13385]= -2145181827;
assign addr[13386]= -2132665626;
assign addr[13387]= -2109331059;
assign addr[13388]= -2075296495;
assign addr[13389]= -2030734582;
assign addr[13390]= -1975871368;
assign addr[13391]= -1910985158;
assign addr[13392]= -1836405100;
assign addr[13393]= -1752509516;
assign addr[13394]= -1659723983;
assign addr[13395]= -1558519173;
assign addr[13396]= -1449408469;
assign addr[13397]= -1332945355;
assign addr[13398]= -1209720613;
assign addr[13399]= -1080359326;
assign addr[13400]= -945517704;
assign addr[13401]= -805879757;
assign addr[13402]= -662153826;
assign addr[13403]= -515068990;
assign addr[13404]= -365371365;
assign addr[13405]= -213820322;
assign addr[13406]= -61184634;
assign addr[13407]= 91761426;
assign addr[13408]= 244242007;
assign addr[13409]= 395483624;
assign addr[13410]= 544719071;
assign addr[13411]= 691191324;
assign addr[13412]= 834157373;
assign addr[13413]= 972891995;
assign addr[13414]= 1106691431;
assign addr[13415]= 1234876957;
assign addr[13416]= 1356798326;
assign addr[13417]= 1471837070;
assign addr[13418]= 1579409630;
assign addr[13419]= 1678970324;
assign addr[13420]= 1770014111;
assign addr[13421]= 1852079154;
assign addr[13422]= 1924749160;
assign addr[13423]= 1987655498;
assign addr[13424]= 2040479063;
assign addr[13425]= 2082951896;
assign addr[13426]= 2114858546;
assign addr[13427]= 2136037160;
assign addr[13428]= 2146380306;
assign addr[13429]= 2145835515;
assign addr[13430]= 2134405552;
assign addr[13431]= 2112148396;
assign addr[13432]= 2079176953;
assign addr[13433]= 2035658475;
assign addr[13434]= 1981813720;
assign addr[13435]= 1917915825;
assign addr[13436]= 1844288924;
assign addr[13437]= 1761306505;
assign addr[13438]= 1669389513;
assign addr[13439]= 1569004214;
assign addr[13440]= 1460659832;
assign addr[13441]= 1344905966;
assign addr[13442]= 1222329801;
assign addr[13443]= 1093553126;
assign addr[13444]= 959229189;
assign addr[13445]= 820039373;
assign addr[13446]= 676689746;
assign addr[13447]= 529907477;
assign addr[13448]= 380437148;
assign addr[13449]= 229036977;
assign addr[13450]= 76474970;
assign addr[13451]= -76474970;
assign addr[13452]= -229036977;
assign addr[13453]= -380437148;
assign addr[13454]= -529907477;
assign addr[13455]= -676689746;
assign addr[13456]= -820039373;
assign addr[13457]= -959229189;
assign addr[13458]= -1093553126;
assign addr[13459]= -1222329801;
assign addr[13460]= -1344905966;
assign addr[13461]= -1460659832;
assign addr[13462]= -1569004214;
assign addr[13463]= -1669389513;
assign addr[13464]= -1761306505;
assign addr[13465]= -1844288924;
assign addr[13466]= -1917915825;
assign addr[13467]= -1981813720;
assign addr[13468]= -2035658475;
assign addr[13469]= -2079176953;
assign addr[13470]= -2112148396;
assign addr[13471]= -2134405552;
assign addr[13472]= -2145835515;
assign addr[13473]= -2146380306;
assign addr[13474]= -2136037160;
assign addr[13475]= -2114858546;
assign addr[13476]= -2082951896;
assign addr[13477]= -2040479063;
assign addr[13478]= -1987655498;
assign addr[13479]= -1924749160;
assign addr[13480]= -1852079154;
assign addr[13481]= -1770014111;
assign addr[13482]= -1678970324;
assign addr[13483]= -1579409630;
assign addr[13484]= -1471837070;
assign addr[13485]= -1356798326;
assign addr[13486]= -1234876957;
assign addr[13487]= -1106691431;
assign addr[13488]= -972891995;
assign addr[13489]= -834157373;
assign addr[13490]= -691191324;
assign addr[13491]= -544719071;
assign addr[13492]= -395483624;
assign addr[13493]= -244242007;
assign addr[13494]= -91761426;
assign addr[13495]= 61184634;
assign addr[13496]= 213820322;
assign addr[13497]= 365371365;
assign addr[13498]= 515068990;
assign addr[13499]= 662153826;
assign addr[13500]= 805879757;
assign addr[13501]= 945517704;
assign addr[13502]= 1080359326;
assign addr[13503]= 1209720613;
assign addr[13504]= 1332945355;
assign addr[13505]= 1449408469;
assign addr[13506]= 1558519173;
assign addr[13507]= 1659723983;
assign addr[13508]= 1752509516;
assign addr[13509]= 1836405100;
assign addr[13510]= 1910985158;
assign addr[13511]= 1975871368;
assign addr[13512]= 2030734582;
assign addr[13513]= 2075296495;
assign addr[13514]= 2109331059;
assign addr[13515]= 2132665626;
assign addr[13516]= 2145181827;
assign addr[13517]= 2146816171;
assign addr[13518]= 2137560369;
assign addr[13519]= 2117461370;
assign addr[13520]= 2086621133;
assign addr[13521]= 2045196100;
assign addr[13522]= 1993396407;
assign addr[13523]= 1931484818;
assign addr[13524]= 1859775393;
assign addr[13525]= 1778631892;
assign addr[13526]= 1688465931;
assign addr[13527]= 1589734894;
assign addr[13528]= 1482939614;
assign addr[13529]= 1368621831;
assign addr[13530]= 1247361445;
assign addr[13531]= 1119773573;
assign addr[13532]= 986505429;
assign addr[13533]= 848233042;
assign addr[13534]= 705657826;
assign addr[13535]= 559503022;
assign addr[13536]= 410510029;
assign addr[13537]= 259434643;
assign addr[13538]= 107043224;
assign addr[13539]= -45891193;
assign addr[13540]= -198592817;
assign addr[13541]= -350287041;
assign addr[13542]= -500204365;
assign addr[13543]= -647584304;
assign addr[13544]= -791679244;
assign addr[13545]= -931758235;
assign addr[13546]= -1067110699;
assign addr[13547]= -1197050035;
assign addr[13548]= -1320917099;
assign addr[13549]= -1438083551;
assign addr[13550]= -1547955041;
assign addr[13551]= -1649974225;
assign addr[13552]= -1743623590;
assign addr[13553]= -1828428082;
assign addr[13554]= -1903957513;
assign addr[13555]= -1969828744;
assign addr[13556]= -2025707632;
assign addr[13557]= -2071310720;
assign addr[13558]= -2106406677;
assign addr[13559]= -2130817471;
assign addr[13560]= -2144419275;
assign addr[13561]= -2147143090;
assign addr[13562]= -2138975100;
assign addr[13563]= -2119956737;
assign addr[13564]= -2090184478;
assign addr[13565]= -2049809346;
assign addr[13566]= -1999036154;
assign addr[13567]= -1938122457;
assign addr[13568]= -1867377253;
assign addr[13569]= -1787159411;
assign addr[13570]= -1697875851;
assign addr[13571]= -1599979481;
assign addr[13572]= -1493966902;
assign addr[13573]= -1380375881;
assign addr[13574]= -1259782632;
assign addr[13575]= -1132798888;
assign addr[13576]= -1000068799;
assign addr[13577]= -862265664;
assign addr[13578]= -720088517;
assign addr[13579]= -574258580;
assign addr[13580]= -425515602;
assign addr[13581]= -274614114;
assign addr[13582]= -122319591;
assign addr[13583]= 30595422;
assign addr[13584]= 183355234;
assign addr[13585]= 335184940;
assign addr[13586]= 485314355;
assign addr[13587]= 632981917;
assign addr[13588]= 777438554;
assign addr[13589]= 917951481;
assign addr[13590]= 1053807919;
assign addr[13591]= 1184318708;
assign addr[13592]= 1308821808;
assign addr[13593]= 1426685652;
assign addr[13594]= 1537312353;
assign addr[13595]= 1640140734;
assign addr[13596]= 1734649179;
assign addr[13597]= 1820358275;
assign addr[13598]= 1896833245;
assign addr[13599]= 1963686155;
assign addr[13600]= 2020577882;
assign addr[13601]= 2067219829;
assign addr[13602]= 2103375398;
assign addr[13603]= 2128861181;
assign addr[13604]= 2143547897;
assign addr[13605]= 2147361045;
assign addr[13606]= 2140281282;
assign addr[13607]= 2122344521;
assign addr[13608]= 2093641749;
assign addr[13609]= 2054318569;
assign addr[13610]= 2004574453;
assign addr[13611]= 1944661739;
assign addr[13612]= 1874884346;
assign addr[13613]= 1795596234;
assign addr[13614]= 1707199606;
assign addr[13615]= 1610142873;
assign addr[13616]= 1504918373;
assign addr[13617]= 1392059879;
assign addr[13618]= 1272139887;
assign addr[13619]= 1145766716;
assign addr[13620]= 1013581418;
assign addr[13621]= 876254528;
assign addr[13622]= 734482665;
assign addr[13623]= 588984994;
assign addr[13624]= 440499581;
assign addr[13625]= 289779648;
assign addr[13626]= 137589750;
assign addr[13627]= -15298099;
assign addr[13628]= -168108346;
assign addr[13629]= -320065829;
assign addr[13630]= -470399716;
assign addr[13631]= -618347408;
assign addr[13632]= -763158411;
assign addr[13633]= -904098143;
assign addr[13634]= -1040451659;
assign addr[13635]= -1171527280;
assign addr[13636]= -1296660098;
assign addr[13637]= -1415215352;
assign addr[13638]= -1526591649;
assign addr[13639]= -1630224009;
assign addr[13640]= -1725586737;
assign addr[13641]= -1812196087;
assign addr[13642]= -1889612716;
assign addr[13643]= -1957443913;
assign addr[13644]= -2015345591;
assign addr[13645]= -2063024031;
assign addr[13646]= -2100237377;
assign addr[13647]= -2126796855;
assign addr[13648]= -2142567738;
assign addr[13649]= -2147470025;
assign addr[13650]= -2141478848;
assign addr[13651]= -2124624598;
assign addr[13652]= -2096992772;
assign addr[13653]= -2058723538;
assign addr[13654]= -2010011024;
assign addr[13655]= -1951102334;
assign addr[13656]= -1882296293;
assign addr[13657]= -1803941934;
assign addr[13658]= -1716436725;
assign addr[13659]= -1620224553;
assign addr[13660]= -1515793473;
assign addr[13661]= -1403673233;
assign addr[13662]= -1284432584;
assign addr[13663]= -1158676398;
assign addr[13664]= -1027042599;
assign addr[13665]= -890198924;
assign addr[13666]= -748839539;
assign addr[13667]= -603681519;
assign addr[13668]= -455461206;
assign addr[13669]= -304930476;
assign addr[13670]= -152852926;
assign addr[13671]= 0;
assign addr[13672]= 152852926;
assign addr[13673]= 304930476;
assign addr[13674]= 455461206;
assign addr[13675]= 603681519;
assign addr[13676]= 748839539;
assign addr[13677]= 890198924;
assign addr[13678]= 1027042599;
assign addr[13679]= 1158676398;
assign addr[13680]= 1284432584;
assign addr[13681]= 1403673233;
assign addr[13682]= 1515793473;
assign addr[13683]= 1620224553;
assign addr[13684]= 1716436725;
assign addr[13685]= 1803941934;
assign addr[13686]= 1882296293;
assign addr[13687]= 1951102334;
assign addr[13688]= 2010011024;
assign addr[13689]= 2058723538;
assign addr[13690]= 2096992772;
assign addr[13691]= 2124624598;
assign addr[13692]= 2141478848;
assign addr[13693]= 2147470025;
assign addr[13694]= 2142567738;
assign addr[13695]= 2126796855;
assign addr[13696]= 2100237377;
assign addr[13697]= 2063024031;
assign addr[13698]= 2015345591;
assign addr[13699]= 1957443913;
assign addr[13700]= 1889612716;
assign addr[13701]= 1812196087;
assign addr[13702]= 1725586737;
assign addr[13703]= 1630224009;
assign addr[13704]= 1526591649;
assign addr[13705]= 1415215352;
assign addr[13706]= 1296660098;
assign addr[13707]= 1171527280;
assign addr[13708]= 1040451659;
assign addr[13709]= 904098143;
assign addr[13710]= 763158411;
assign addr[13711]= 618347408;
assign addr[13712]= 470399716;
assign addr[13713]= 320065829;
assign addr[13714]= 168108346;
assign addr[13715]= 15298099;
assign addr[13716]= -137589750;
assign addr[13717]= -289779648;
assign addr[13718]= -440499581;
assign addr[13719]= -588984994;
assign addr[13720]= -734482665;
assign addr[13721]= -876254528;
assign addr[13722]= -1013581418;
assign addr[13723]= -1145766716;
assign addr[13724]= -1272139887;
assign addr[13725]= -1392059879;
assign addr[13726]= -1504918373;
assign addr[13727]= -1610142873;
assign addr[13728]= -1707199606;
assign addr[13729]= -1795596234;
assign addr[13730]= -1874884346;
assign addr[13731]= -1944661739;
assign addr[13732]= -2004574453;
assign addr[13733]= -2054318569;
assign addr[13734]= -2093641749;
assign addr[13735]= -2122344521;
assign addr[13736]= -2140281282;
assign addr[13737]= -2147361045;
assign addr[13738]= -2143547897;
assign addr[13739]= -2128861181;
assign addr[13740]= -2103375398;
assign addr[13741]= -2067219829;
assign addr[13742]= -2020577882;
assign addr[13743]= -1963686155;
assign addr[13744]= -1896833245;
assign addr[13745]= -1820358275;
assign addr[13746]= -1734649179;
assign addr[13747]= -1640140734;
assign addr[13748]= -1537312353;
assign addr[13749]= -1426685652;
assign addr[13750]= -1308821808;
assign addr[13751]= -1184318708;
assign addr[13752]= -1053807919;
assign addr[13753]= -917951481;
assign addr[13754]= -777438554;
assign addr[13755]= -632981917;
assign addr[13756]= -485314355;
assign addr[13757]= -335184940;
assign addr[13758]= -183355234;
assign addr[13759]= -30595422;
assign addr[13760]= 122319591;
assign addr[13761]= 274614114;
assign addr[13762]= 425515602;
assign addr[13763]= 574258580;
assign addr[13764]= 720088517;
assign addr[13765]= 862265664;
assign addr[13766]= 1000068799;
assign addr[13767]= 1132798888;
assign addr[13768]= 1259782632;
assign addr[13769]= 1380375881;
assign addr[13770]= 1493966902;
assign addr[13771]= 1599979481;
assign addr[13772]= 1697875851;
assign addr[13773]= 1787159411;
assign addr[13774]= 1867377253;
assign addr[13775]= 1938122457;
assign addr[13776]= 1999036154;
assign addr[13777]= 2049809346;
assign addr[13778]= 2090184478;
assign addr[13779]= 2119956737;
assign addr[13780]= 2138975100;
assign addr[13781]= 2147143090;
assign addr[13782]= 2144419275;
assign addr[13783]= 2130817471;
assign addr[13784]= 2106406677;
assign addr[13785]= 2071310720;
assign addr[13786]= 2025707632;
assign addr[13787]= 1969828744;
assign addr[13788]= 1903957513;
assign addr[13789]= 1828428082;
assign addr[13790]= 1743623590;
assign addr[13791]= 1649974225;
assign addr[13792]= 1547955041;
assign addr[13793]= 1438083551;
assign addr[13794]= 1320917099;
assign addr[13795]= 1197050035;
assign addr[13796]= 1067110699;
assign addr[13797]= 931758235;
assign addr[13798]= 791679244;
assign addr[13799]= 647584304;
assign addr[13800]= 500204365;
assign addr[13801]= 350287041;
assign addr[13802]= 198592817;
assign addr[13803]= 45891193;
assign addr[13804]= -107043224;
assign addr[13805]= -259434643;
assign addr[13806]= -410510029;
assign addr[13807]= -559503022;
assign addr[13808]= -705657826;
assign addr[13809]= -848233042;
assign addr[13810]= -986505429;
assign addr[13811]= -1119773573;
assign addr[13812]= -1247361445;
assign addr[13813]= -1368621831;
assign addr[13814]= -1482939614;
assign addr[13815]= -1589734894;
assign addr[13816]= -1688465931;
assign addr[13817]= -1778631892;
assign addr[13818]= -1859775393;
assign addr[13819]= -1931484818;
assign addr[13820]= -1993396407;
assign addr[13821]= -2045196100;
assign addr[13822]= -2086621133;
assign addr[13823]= -2117461370;
assign addr[13824]= -2137560369;
assign addr[13825]= -2146816171;
assign addr[13826]= -2145181827;
assign addr[13827]= -2132665626;
assign addr[13828]= -2109331059;
assign addr[13829]= -2075296495;
assign addr[13830]= -2030734582;
assign addr[13831]= -1975871368;
assign addr[13832]= -1910985158;
assign addr[13833]= -1836405100;
assign addr[13834]= -1752509516;
assign addr[13835]= -1659723983;
assign addr[13836]= -1558519173;
assign addr[13837]= -1449408469;
assign addr[13838]= -1332945355;
assign addr[13839]= -1209720613;
assign addr[13840]= -1080359326;
assign addr[13841]= -945517704;
assign addr[13842]= -805879757;
assign addr[13843]= -662153826;
assign addr[13844]= -515068990;
assign addr[13845]= -365371365;
assign addr[13846]= -213820322;
assign addr[13847]= -61184634;
assign addr[13848]= 91761426;
assign addr[13849]= 244242007;
assign addr[13850]= 395483624;
assign addr[13851]= 544719071;
assign addr[13852]= 691191324;
assign addr[13853]= 834157373;
assign addr[13854]= 972891995;
assign addr[13855]= 1106691431;
assign addr[13856]= 1234876957;
assign addr[13857]= 1356798326;
assign addr[13858]= 1471837070;
assign addr[13859]= 1579409630;
assign addr[13860]= 1678970324;
assign addr[13861]= 1770014111;
assign addr[13862]= 1852079154;
assign addr[13863]= 1924749160;
assign addr[13864]= 1987655498;
assign addr[13865]= 2040479063;
assign addr[13866]= 2082951896;
assign addr[13867]= 2114858546;
assign addr[13868]= 2136037160;
assign addr[13869]= 2146380306;
assign addr[13870]= 2145835515;
assign addr[13871]= 2134405552;
assign addr[13872]= 2112148396;
assign addr[13873]= 2079176953;
assign addr[13874]= 2035658475;
assign addr[13875]= 1981813720;
assign addr[13876]= 1917915825;
assign addr[13877]= 1844288924;
assign addr[13878]= 1761306505;
assign addr[13879]= 1669389513;
assign addr[13880]= 1569004214;
assign addr[13881]= 1460659832;
assign addr[13882]= 1344905966;
assign addr[13883]= 1222329801;
assign addr[13884]= 1093553126;
assign addr[13885]= 959229189;
assign addr[13886]= 820039373;
assign addr[13887]= 676689746;
assign addr[13888]= 529907477;
assign addr[13889]= 380437148;
assign addr[13890]= 229036977;
assign addr[13891]= 76474970;
assign addr[13892]= -76474970;
assign addr[13893]= -229036977;
assign addr[13894]= -380437148;
assign addr[13895]= -529907477;
assign addr[13896]= -676689746;
assign addr[13897]= -820039373;
assign addr[13898]= -959229189;
assign addr[13899]= -1093553126;
assign addr[13900]= -1222329801;
assign addr[13901]= -1344905966;
assign addr[13902]= -1460659832;
assign addr[13903]= -1569004214;
assign addr[13904]= -1669389513;
assign addr[13905]= -1761306505;
assign addr[13906]= -1844288924;
assign addr[13907]= -1917915825;
assign addr[13908]= -1981813720;
assign addr[13909]= -2035658475;
assign addr[13910]= -2079176953;
assign addr[13911]= -2112148396;
assign addr[13912]= -2134405552;
assign addr[13913]= -2145835515;
assign addr[13914]= -2146380306;
assign addr[13915]= -2136037160;
assign addr[13916]= -2114858546;
assign addr[13917]= -2082951896;
assign addr[13918]= -2040479063;
assign addr[13919]= -1987655498;
assign addr[13920]= -1924749160;
assign addr[13921]= -1852079154;
assign addr[13922]= -1770014111;
assign addr[13923]= -1678970324;
assign addr[13924]= -1579409630;
assign addr[13925]= -1471837070;
assign addr[13926]= -1356798326;
assign addr[13927]= -1234876957;
assign addr[13928]= -1106691431;
assign addr[13929]= -972891995;
assign addr[13930]= -834157373;
assign addr[13931]= -691191324;
assign addr[13932]= -544719071;
assign addr[13933]= -395483624;
assign addr[13934]= -244242007;
assign addr[13935]= -91761426;
assign addr[13936]= 61184634;
assign addr[13937]= 213820322;
assign addr[13938]= 365371365;
assign addr[13939]= 515068990;
assign addr[13940]= 662153826;
assign addr[13941]= 805879757;
assign addr[13942]= 945517704;
assign addr[13943]= 1080359326;
assign addr[13944]= 1209720613;
assign addr[13945]= 1332945355;
assign addr[13946]= 1449408469;
assign addr[13947]= 1558519173;
assign addr[13948]= 1659723983;
assign addr[13949]= 1752509516;
assign addr[13950]= 1836405100;
assign addr[13951]= 1910985158;
assign addr[13952]= 1975871368;
assign addr[13953]= 2030734582;
assign addr[13954]= 2075296495;
assign addr[13955]= 2109331059;
assign addr[13956]= 2132665626;
assign addr[13957]= 2145181827;
assign addr[13958]= 2146816171;
assign addr[13959]= 2137560369;
assign addr[13960]= 2117461370;
assign addr[13961]= 2086621133;
assign addr[13962]= 2045196100;
assign addr[13963]= 1993396407;
assign addr[13964]= 1931484818;
assign addr[13965]= 1859775393;
assign addr[13966]= 1778631892;
assign addr[13967]= 1688465931;
assign addr[13968]= 1589734894;
assign addr[13969]= 1482939614;
assign addr[13970]= 1368621831;
assign addr[13971]= 1247361445;
assign addr[13972]= 1119773573;
assign addr[13973]= 986505429;
assign addr[13974]= 848233042;
assign addr[13975]= 705657826;
assign addr[13976]= 559503022;
assign addr[13977]= 410510029;
assign addr[13978]= 259434643;
assign addr[13979]= 107043224;
assign addr[13980]= -45891193;
assign addr[13981]= -198592817;
assign addr[13982]= -350287041;
assign addr[13983]= -500204365;
assign addr[13984]= -647584304;
assign addr[13985]= -791679244;
assign addr[13986]= -931758235;
assign addr[13987]= -1067110699;
assign addr[13988]= -1197050035;
assign addr[13989]= -1320917099;
assign addr[13990]= -1438083551;
assign addr[13991]= -1547955041;
assign addr[13992]= -1649974225;
assign addr[13993]= -1743623590;
assign addr[13994]= -1828428082;
assign addr[13995]= -1903957513;
assign addr[13996]= -1969828744;
assign addr[13997]= -2025707632;
assign addr[13998]= -2071310720;
assign addr[13999]= -2106406677;
assign addr[14000]= -2130817471;
assign addr[14001]= -2144419275;
assign addr[14002]= -2147143090;
assign addr[14003]= -2138975100;
assign addr[14004]= -2119956737;
assign addr[14005]= -2090184478;
assign addr[14006]= -2049809346;
assign addr[14007]= -1999036154;
assign addr[14008]= -1938122457;
assign addr[14009]= -1867377253;
assign addr[14010]= -1787159411;
assign addr[14011]= -1697875851;
assign addr[14012]= -1599979481;
assign addr[14013]= -1493966902;
assign addr[14014]= -1380375881;
assign addr[14015]= -1259782632;
assign addr[14016]= -1132798888;
assign addr[14017]= -1000068799;
assign addr[14018]= -862265664;
assign addr[14019]= -720088517;
assign addr[14020]= -574258580;
assign addr[14021]= -425515602;
assign addr[14022]= -274614114;
assign addr[14023]= -122319591;
assign addr[14024]= 30595422;
assign addr[14025]= 183355234;
assign addr[14026]= 335184940;
assign addr[14027]= 485314355;
assign addr[14028]= 632981917;
assign addr[14029]= 777438554;
assign addr[14030]= 917951481;
assign addr[14031]= 1053807919;
assign addr[14032]= 1184318708;
assign addr[14033]= 1308821808;
assign addr[14034]= 1426685652;
assign addr[14035]= 1537312353;
assign addr[14036]= 1640140734;
assign addr[14037]= 1734649179;
assign addr[14038]= 1820358275;
assign addr[14039]= 1896833245;
assign addr[14040]= 1963686155;
assign addr[14041]= 2020577882;
assign addr[14042]= 2067219829;
assign addr[14043]= 2103375398;
assign addr[14044]= 2128861181;
assign addr[14045]= 2143547897;
assign addr[14046]= 2147361045;
assign addr[14047]= 2140281282;
assign addr[14048]= 2122344521;
assign addr[14049]= 2093641749;
assign addr[14050]= 2054318569;
assign addr[14051]= 2004574453;
assign addr[14052]= 1944661739;
assign addr[14053]= 1874884346;
assign addr[14054]= 1795596234;
assign addr[14055]= 1707199606;
assign addr[14056]= 1610142873;
assign addr[14057]= 1504918373;
assign addr[14058]= 1392059879;
assign addr[14059]= 1272139887;
assign addr[14060]= 1145766716;
assign addr[14061]= 1013581418;
assign addr[14062]= 876254528;
assign addr[14063]= 734482665;
assign addr[14064]= 588984994;
assign addr[14065]= 440499581;
assign addr[14066]= 289779648;
assign addr[14067]= 137589750;
assign addr[14068]= -15298099;
assign addr[14069]= -168108346;
assign addr[14070]= -320065829;
assign addr[14071]= -470399716;
assign addr[14072]= -618347408;
assign addr[14073]= -763158411;
assign addr[14074]= -904098143;
assign addr[14075]= -1040451659;
assign addr[14076]= -1171527280;
assign addr[14077]= -1296660098;
assign addr[14078]= -1415215352;
assign addr[14079]= -1526591649;
assign addr[14080]= -1630224009;
assign addr[14081]= -1725586737;
assign addr[14082]= -1812196087;
assign addr[14083]= -1889612716;
assign addr[14084]= -1957443913;
assign addr[14085]= -2015345591;
assign addr[14086]= -2063024031;
assign addr[14087]= -2100237377;
assign addr[14088]= -2126796855;
assign addr[14089]= -2142567738;
assign addr[14090]= -2147470025;
assign addr[14091]= -2141478848;
assign addr[14092]= -2124624598;
assign addr[14093]= -2096992772;
assign addr[14094]= -2058723538;
assign addr[14095]= -2010011024;
assign addr[14096]= -1951102334;
assign addr[14097]= -1882296293;
assign addr[14098]= -1803941934;
assign addr[14099]= -1716436725;
assign addr[14100]= -1620224553;
assign addr[14101]= -1515793473;
assign addr[14102]= -1403673233;
assign addr[14103]= -1284432584;
assign addr[14104]= -1158676398;
assign addr[14105]= -1027042599;
assign addr[14106]= -890198924;
assign addr[14107]= -748839539;
assign addr[14108]= -603681519;
assign addr[14109]= -455461206;
assign addr[14110]= -304930476;
assign addr[14111]= -152852926;
assign addr[14112]= 0;
assign addr[14113]= 152852926;
assign addr[14114]= 304930476;
assign addr[14115]= 455461206;
assign addr[14116]= 603681519;
assign addr[14117]= 748839539;
assign addr[14118]= 890198924;
assign addr[14119]= 1027042599;
assign addr[14120]= 1158676398;
assign addr[14121]= 1284432584;
assign addr[14122]= 1403673233;
assign addr[14123]= 1515793473;
assign addr[14124]= 1620224553;
assign addr[14125]= 1716436725;
assign addr[14126]= 1803941934;
assign addr[14127]= 1882296293;
assign addr[14128]= 1951102334;
assign addr[14129]= 2010011024;
assign addr[14130]= 2058723538;
assign addr[14131]= 2096992772;
assign addr[14132]= 2124624598;
assign addr[14133]= 2141478848;
assign addr[14134]= 2147470025;
assign addr[14135]= 2142567738;
assign addr[14136]= 2126796855;
assign addr[14137]= 2100237377;
assign addr[14138]= 2063024031;
assign addr[14139]= 2015345591;
assign addr[14140]= 1957443913;
assign addr[14141]= 1889612716;
assign addr[14142]= 1812196087;
assign addr[14143]= 1725586737;
assign addr[14144]= 1630224009;
assign addr[14145]= 1526591649;
assign addr[14146]= 1415215352;
assign addr[14147]= 1296660098;
assign addr[14148]= 1171527280;
assign addr[14149]= 1040451659;
assign addr[14150]= 904098143;
assign addr[14151]= 763158411;
assign addr[14152]= 618347408;
assign addr[14153]= 470399716;
assign addr[14154]= 320065829;
assign addr[14155]= 168108346;
assign addr[14156]= 15298099;
assign addr[14157]= -137589750;
assign addr[14158]= -289779648;
assign addr[14159]= -440499581;
assign addr[14160]= -588984994;
assign addr[14161]= -734482665;
assign addr[14162]= -876254528;
assign addr[14163]= -1013581418;
assign addr[14164]= -1145766716;
assign addr[14165]= -1272139887;
assign addr[14166]= -1392059879;
assign addr[14167]= -1504918373;
assign addr[14168]= -1610142873;
assign addr[14169]= -1707199606;
assign addr[14170]= -1795596234;
assign addr[14171]= -1874884346;
assign addr[14172]= -1944661739;
assign addr[14173]= -2004574453;
assign addr[14174]= -2054318569;
assign addr[14175]= -2093641749;
assign addr[14176]= -2122344521;
assign addr[14177]= -2140281282;
assign addr[14178]= -2147361045;
assign addr[14179]= -2143547897;
assign addr[14180]= -2128861181;
assign addr[14181]= -2103375398;
assign addr[14182]= -2067219829;
assign addr[14183]= -2020577882;
assign addr[14184]= -1963686155;
assign addr[14185]= -1896833245;
assign addr[14186]= -1820358275;
assign addr[14187]= -1734649179;
assign addr[14188]= -1640140734;
assign addr[14189]= -1537312353;
assign addr[14190]= -1426685652;
assign addr[14191]= -1308821808;
assign addr[14192]= -1184318708;
assign addr[14193]= -1053807919;
assign addr[14194]= -917951481;
assign addr[14195]= -777438554;
assign addr[14196]= -632981917;
assign addr[14197]= -485314355;
assign addr[14198]= -335184940;
assign addr[14199]= -183355234;
assign addr[14200]= -30595422;
assign addr[14201]= 122319591;
assign addr[14202]= 274614114;
assign addr[14203]= 425515602;
assign addr[14204]= 574258580;
assign addr[14205]= 720088517;
assign addr[14206]= 862265664;
assign addr[14207]= 1000068799;
assign addr[14208]= 1132798888;
assign addr[14209]= 1259782632;
assign addr[14210]= 1380375881;
assign addr[14211]= 1493966902;
assign addr[14212]= 1599979481;
assign addr[14213]= 1697875851;
assign addr[14214]= 1787159411;
assign addr[14215]= 1867377253;
assign addr[14216]= 1938122457;
assign addr[14217]= 1999036154;
assign addr[14218]= 2049809346;
assign addr[14219]= 2090184478;
assign addr[14220]= 2119956737;
assign addr[14221]= 2138975100;
assign addr[14222]= 2147143090;
assign addr[14223]= 2144419275;
assign addr[14224]= 2130817471;
assign addr[14225]= 2106406677;
assign addr[14226]= 2071310720;
assign addr[14227]= 2025707632;
assign addr[14228]= 1969828744;
assign addr[14229]= 1903957513;
assign addr[14230]= 1828428082;
assign addr[14231]= 1743623590;
assign addr[14232]= 1649974225;
assign addr[14233]= 1547955041;
assign addr[14234]= 1438083551;
assign addr[14235]= 1320917099;
assign addr[14236]= 1197050035;
assign addr[14237]= 1067110699;
assign addr[14238]= 931758235;
assign addr[14239]= 791679244;
assign addr[14240]= 647584304;
assign addr[14241]= 500204365;
assign addr[14242]= 350287041;
assign addr[14243]= 198592817;
assign addr[14244]= 45891193;
assign addr[14245]= -107043224;
assign addr[14246]= -259434643;
assign addr[14247]= -410510029;
assign addr[14248]= -559503022;
assign addr[14249]= -705657826;
assign addr[14250]= -848233042;
assign addr[14251]= -986505429;
assign addr[14252]= -1119773573;
assign addr[14253]= -1247361445;
assign addr[14254]= -1368621831;
assign addr[14255]= -1482939614;
assign addr[14256]= -1589734894;
assign addr[14257]= -1688465931;
assign addr[14258]= -1778631892;
assign addr[14259]= -1859775393;
assign addr[14260]= -1931484818;
assign addr[14261]= -1993396407;
assign addr[14262]= -2045196100;
assign addr[14263]= -2086621133;
assign addr[14264]= -2117461370;
assign addr[14265]= -2137560369;
assign addr[14266]= -2146816171;
assign addr[14267]= -2145181827;
assign addr[14268]= -2132665626;
assign addr[14269]= -2109331059;
assign addr[14270]= -2075296495;
assign addr[14271]= -2030734582;
assign addr[14272]= -1975871368;
assign addr[14273]= -1910985158;
assign addr[14274]= -1836405100;
assign addr[14275]= -1752509516;
assign addr[14276]= -1659723983;
assign addr[14277]= -1558519173;
assign addr[14278]= -1449408469;
assign addr[14279]= -1332945355;
assign addr[14280]= -1209720613;
assign addr[14281]= -1080359326;
assign addr[14282]= -945517704;
assign addr[14283]= -805879757;
assign addr[14284]= -662153826;
assign addr[14285]= -515068990;
assign addr[14286]= -365371365;
assign addr[14287]= -213820322;
assign addr[14288]= -61184634;
assign addr[14289]= 91761426;
assign addr[14290]= 244242007;
assign addr[14291]= 395483624;
assign addr[14292]= 544719071;
assign addr[14293]= 691191324;
assign addr[14294]= 834157373;
assign addr[14295]= 972891995;
assign addr[14296]= 1106691431;
assign addr[14297]= 1234876957;
assign addr[14298]= 1356798326;
assign addr[14299]= 1471837070;
assign addr[14300]= 1579409630;
assign addr[14301]= 1678970324;
assign addr[14302]= 1770014111;
assign addr[14303]= 1852079154;
assign addr[14304]= 1924749160;
assign addr[14305]= 1987655498;
assign addr[14306]= 2040479063;
assign addr[14307]= 2082951896;
assign addr[14308]= 2114858546;
assign addr[14309]= 2136037160;
assign addr[14310]= 2146380306;
assign addr[14311]= 2145835515;
assign addr[14312]= 2134405552;
assign addr[14313]= 2112148396;
assign addr[14314]= 2079176953;
assign addr[14315]= 2035658475;
assign addr[14316]= 1981813720;
assign addr[14317]= 1917915825;
assign addr[14318]= 1844288924;
assign addr[14319]= 1761306505;
assign addr[14320]= 1669389513;
assign addr[14321]= 1569004214;
assign addr[14322]= 1460659832;
assign addr[14323]= 1344905966;
assign addr[14324]= 1222329801;
assign addr[14325]= 1093553126;
assign addr[14326]= 959229189;
assign addr[14327]= 820039373;
assign addr[14328]= 676689746;
assign addr[14329]= 529907477;
assign addr[14330]= 380437148;
assign addr[14331]= 229036977;
assign addr[14332]= 76474970;
assign addr[14333]= -76474970;
assign addr[14334]= -229036977;
assign addr[14335]= -380437148;
assign addr[14336]= -529907477;
assign addr[14337]= -676689746;
assign addr[14338]= -820039373;
assign addr[14339]= -959229189;
assign addr[14340]= -1093553126;
assign addr[14341]= -1222329801;
assign addr[14342]= -1344905966;
assign addr[14343]= -1460659832;
assign addr[14344]= -1569004214;
assign addr[14345]= -1669389513;
assign addr[14346]= -1761306505;
assign addr[14347]= -1844288924;
assign addr[14348]= -1917915825;
assign addr[14349]= -1981813720;
assign addr[14350]= -2035658475;
assign addr[14351]= -2079176953;
assign addr[14352]= -2112148396;
assign addr[14353]= -2134405552;
assign addr[14354]= -2145835515;
assign addr[14355]= -2146380306;
assign addr[14356]= -2136037160;
assign addr[14357]= -2114858546;
assign addr[14358]= -2082951896;
assign addr[14359]= -2040479063;
assign addr[14360]= -1987655498;
assign addr[14361]= -1924749160;
assign addr[14362]= -1852079154;
assign addr[14363]= -1770014111;
assign addr[14364]= -1678970324;
assign addr[14365]= -1579409630;
assign addr[14366]= -1471837070;
assign addr[14367]= -1356798326;
assign addr[14368]= -1234876957;
assign addr[14369]= -1106691431;
assign addr[14370]= -972891995;
assign addr[14371]= -834157373;
assign addr[14372]= -691191324;
assign addr[14373]= -544719071;
assign addr[14374]= -395483624;
assign addr[14375]= -244242007;
assign addr[14376]= -91761426;
assign addr[14377]= 61184634;
assign addr[14378]= 213820322;
assign addr[14379]= 365371365;
assign addr[14380]= 515068990;
assign addr[14381]= 662153826;
assign addr[14382]= 805879757;
assign addr[14383]= 945517704;
assign addr[14384]= 1080359326;
assign addr[14385]= 1209720613;
assign addr[14386]= 1332945355;
assign addr[14387]= 1449408469;
assign addr[14388]= 1558519173;
assign addr[14389]= 1659723983;
assign addr[14390]= 1752509516;
assign addr[14391]= 1836405100;
assign addr[14392]= 1910985158;
assign addr[14393]= 1975871368;
assign addr[14394]= 2030734582;
assign addr[14395]= 2075296495;
assign addr[14396]= 2109331059;
assign addr[14397]= 2132665626;
assign addr[14398]= 2145181827;
assign addr[14399]= 2146816171;
assign addr[14400]= 2137560369;
assign addr[14401]= 2117461370;
assign addr[14402]= 2086621133;
assign addr[14403]= 2045196100;
assign addr[14404]= 1993396407;
assign addr[14405]= 1931484818;
assign addr[14406]= 1859775393;
assign addr[14407]= 1778631892;
assign addr[14408]= 1688465931;
assign addr[14409]= 1589734894;
assign addr[14410]= 1482939614;
assign addr[14411]= 1368621831;
assign addr[14412]= 1247361445;
assign addr[14413]= 1119773573;
assign addr[14414]= 986505429;
assign addr[14415]= 848233042;
assign addr[14416]= 705657826;
assign addr[14417]= 559503022;
assign addr[14418]= 410510029;
assign addr[14419]= 259434643;
assign addr[14420]= 107043224;
assign addr[14421]= -45891193;
assign addr[14422]= -198592817;
assign addr[14423]= -350287041;
assign addr[14424]= -500204365;
assign addr[14425]= -647584304;
assign addr[14426]= -791679244;
assign addr[14427]= -931758235;
assign addr[14428]= -1067110699;
assign addr[14429]= -1197050035;
assign addr[14430]= -1320917099;
assign addr[14431]= -1438083551;
assign addr[14432]= -1547955041;
assign addr[14433]= -1649974225;
assign addr[14434]= -1743623590;
assign addr[14435]= -1828428082;
assign addr[14436]= -1903957513;
assign addr[14437]= -1969828744;
assign addr[14438]= -2025707632;
assign addr[14439]= -2071310720;
assign addr[14440]= -2106406677;
assign addr[14441]= -2130817471;
assign addr[14442]= -2144419275;
assign addr[14443]= -2147143090;
assign addr[14444]= -2138975100;
assign addr[14445]= -2119956737;
assign addr[14446]= -2090184478;
assign addr[14447]= -2049809346;
assign addr[14448]= -1999036154;
assign addr[14449]= -1938122457;
assign addr[14450]= -1867377253;
assign addr[14451]= -1787159411;
assign addr[14452]= -1697875851;
assign addr[14453]= -1599979481;
assign addr[14454]= -1493966902;
assign addr[14455]= -1380375881;
assign addr[14456]= -1259782632;
assign addr[14457]= -1132798888;
assign addr[14458]= -1000068799;
assign addr[14459]= -862265664;
assign addr[14460]= -720088517;
assign addr[14461]= -574258580;
assign addr[14462]= -425515602;
assign addr[14463]= -274614114;
assign addr[14464]= -122319591;
assign addr[14465]= 30595422;
assign addr[14466]= 183355234;
assign addr[14467]= 335184940;
assign addr[14468]= 485314355;
assign addr[14469]= 632981917;
assign addr[14470]= 777438554;
assign addr[14471]= 917951481;
assign addr[14472]= 1053807919;
assign addr[14473]= 1184318708;
assign addr[14474]= 1308821808;
assign addr[14475]= 1426685652;
assign addr[14476]= 1537312353;
assign addr[14477]= 1640140734;
assign addr[14478]= 1734649179;
assign addr[14479]= 1820358275;
assign addr[14480]= 1896833245;
assign addr[14481]= 1963686155;
assign addr[14482]= 2020577882;
assign addr[14483]= 2067219829;
assign addr[14484]= 2103375398;
assign addr[14485]= 2128861181;
assign addr[14486]= 2143547897;
assign addr[14487]= 2147361045;
assign addr[14488]= 2140281282;
assign addr[14489]= 2122344521;
assign addr[14490]= 2093641749;
assign addr[14491]= 2054318569;
assign addr[14492]= 2004574453;
assign addr[14493]= 1944661739;
assign addr[14494]= 1874884346;
assign addr[14495]= 1795596234;
assign addr[14496]= 1707199606;
assign addr[14497]= 1610142873;
assign addr[14498]= 1504918373;
assign addr[14499]= 1392059879;
assign addr[14500]= 1272139887;
assign addr[14501]= 1145766716;
assign addr[14502]= 1013581418;
assign addr[14503]= 876254528;
assign addr[14504]= 734482665;
assign addr[14505]= 588984994;
assign addr[14506]= 440499581;
assign addr[14507]= 289779648;
assign addr[14508]= 137589750;
assign addr[14509]= -15298099;
assign addr[14510]= -168108346;
assign addr[14511]= -320065829;
assign addr[14512]= -470399716;
assign addr[14513]= -618347408;
assign addr[14514]= -763158411;
assign addr[14515]= -904098143;
assign addr[14516]= -1040451659;
assign addr[14517]= -1171527280;
assign addr[14518]= -1296660098;
assign addr[14519]= -1415215352;
assign addr[14520]= -1526591649;
assign addr[14521]= -1630224009;
assign addr[14522]= -1725586737;
assign addr[14523]= -1812196087;
assign addr[14524]= -1889612716;
assign addr[14525]= -1957443913;
assign addr[14526]= -2015345591;
assign addr[14527]= -2063024031;
assign addr[14528]= -2100237377;
assign addr[14529]= -2126796855;
assign addr[14530]= -2142567738;
assign addr[14531]= -2147470025;
assign addr[14532]= -2141478848;
assign addr[14533]= -2124624598;
assign addr[14534]= -2096992772;
assign addr[14535]= -2058723538;
assign addr[14536]= -2010011024;
assign addr[14537]= -1951102334;
assign addr[14538]= -1882296293;
assign addr[14539]= -1803941934;
assign addr[14540]= -1716436725;
assign addr[14541]= -1620224553;
assign addr[14542]= -1515793473;
assign addr[14543]= -1403673233;
assign addr[14544]= -1284432584;
assign addr[14545]= -1158676398;
assign addr[14546]= -1027042599;
assign addr[14547]= -890198924;
assign addr[14548]= -748839539;
assign addr[14549]= -603681519;
assign addr[14550]= -455461206;
assign addr[14551]= -304930476;
assign addr[14552]= -152852926;
assign addr[14553]= 0;
assign addr[14554]= 152852926;
assign addr[14555]= 304930476;
assign addr[14556]= 455461206;
assign addr[14557]= 603681519;
assign addr[14558]= 748839539;
assign addr[14559]= 890198924;
assign addr[14560]= 1027042599;
assign addr[14561]= 1158676398;
assign addr[14562]= 1284432584;
assign addr[14563]= 1403673233;
assign addr[14564]= 1515793473;
assign addr[14565]= 1620224553;
assign addr[14566]= 1716436725;
assign addr[14567]= 1803941934;
assign addr[14568]= 1882296293;
assign addr[14569]= 1951102334;
assign addr[14570]= 2010011024;
assign addr[14571]= 2058723538;
assign addr[14572]= 2096992772;
assign addr[14573]= 2124624598;
assign addr[14574]= 2141478848;
assign addr[14575]= 2147470025;
assign addr[14576]= 2142567738;
assign addr[14577]= 2126796855;
assign addr[14578]= 2100237377;
assign addr[14579]= 2063024031;
assign addr[14580]= 2015345591;
assign addr[14581]= 1957443913;
assign addr[14582]= 1889612716;
assign addr[14583]= 1812196087;
assign addr[14584]= 1725586737;
assign addr[14585]= 1630224009;
assign addr[14586]= 1526591649;
assign addr[14587]= 1415215352;
assign addr[14588]= 1296660098;
assign addr[14589]= 1171527280;
assign addr[14590]= 1040451659;
assign addr[14591]= 904098143;
assign addr[14592]= 763158411;
assign addr[14593]= 618347408;
assign addr[14594]= 470399716;
assign addr[14595]= 320065829;
assign addr[14596]= 168108346;
assign addr[14597]= 15298099;
assign addr[14598]= -137589750;
assign addr[14599]= -289779648;
assign addr[14600]= -440499581;
assign addr[14601]= -588984994;
assign addr[14602]= -734482665;
assign addr[14603]= -876254528;
assign addr[14604]= -1013581418;
assign addr[14605]= -1145766716;
assign addr[14606]= -1272139887;
assign addr[14607]= -1392059879;
assign addr[14608]= -1504918373;
assign addr[14609]= -1610142873;
assign addr[14610]= -1707199606;
assign addr[14611]= -1795596234;
assign addr[14612]= -1874884346;
assign addr[14613]= -1944661739;
assign addr[14614]= -2004574453;
assign addr[14615]= -2054318569;
assign addr[14616]= -2093641749;
assign addr[14617]= -2122344521;
assign addr[14618]= -2140281282;
assign addr[14619]= -2147361045;
assign addr[14620]= -2143547897;
assign addr[14621]= -2128861181;
assign addr[14622]= -2103375398;
assign addr[14623]= -2067219829;
assign addr[14624]= -2020577882;
assign addr[14625]= -1963686155;
assign addr[14626]= -1896833245;
assign addr[14627]= -1820358275;
assign addr[14628]= -1734649179;
assign addr[14629]= -1640140734;
assign addr[14630]= -1537312353;
assign addr[14631]= -1426685652;
assign addr[14632]= -1308821808;
assign addr[14633]= -1184318708;
assign addr[14634]= -1053807919;
assign addr[14635]= -917951481;
assign addr[14636]= -777438554;
assign addr[14637]= -632981917;
assign addr[14638]= -485314355;
assign addr[14639]= -335184940;
assign addr[14640]= -183355234;
assign addr[14641]= -30595422;
assign addr[14642]= 122319591;
assign addr[14643]= 274614114;
assign addr[14644]= 425515602;
assign addr[14645]= 574258580;
assign addr[14646]= 720088517;
assign addr[14647]= 862265664;
assign addr[14648]= 1000068799;
assign addr[14649]= 1132798888;
assign addr[14650]= 1259782632;
assign addr[14651]= 1380375881;
assign addr[14652]= 1493966902;
assign addr[14653]= 1599979481;
assign addr[14654]= 1697875851;
assign addr[14655]= 1787159411;
assign addr[14656]= 1867377253;
assign addr[14657]= 1938122457;
assign addr[14658]= 1999036154;
assign addr[14659]= 2049809346;
assign addr[14660]= 2090184478;
assign addr[14661]= 2119956737;
assign addr[14662]= 2138975100;
assign addr[14663]= 2147143090;
assign addr[14664]= 2144419275;
assign addr[14665]= 2130817471;
assign addr[14666]= 2106406677;
assign addr[14667]= 2071310720;
assign addr[14668]= 2025707632;
assign addr[14669]= 1969828744;
assign addr[14670]= 1903957513;
assign addr[14671]= 1828428082;
assign addr[14672]= 1743623590;
assign addr[14673]= 1649974225;
assign addr[14674]= 1547955041;
assign addr[14675]= 1438083551;
assign addr[14676]= 1320917099;
assign addr[14677]= 1197050035;
assign addr[14678]= 1067110699;
assign addr[14679]= 931758235;
assign addr[14680]= 791679244;
assign addr[14681]= 647584304;
assign addr[14682]= 500204365;
assign addr[14683]= 350287041;
assign addr[14684]= 198592817;
assign addr[14685]= 45891193;
assign addr[14686]= -107043224;
assign addr[14687]= -259434643;
assign addr[14688]= -410510029;
assign addr[14689]= -559503022;
assign addr[14690]= -705657826;
assign addr[14691]= -848233042;
assign addr[14692]= -986505429;
assign addr[14693]= -1119773573;
assign addr[14694]= -1247361445;
assign addr[14695]= -1368621831;
assign addr[14696]= -1482939614;
assign addr[14697]= -1589734894;
assign addr[14698]= -1688465931;
assign addr[14699]= -1778631892;
assign addr[14700]= -1859775393;
assign addr[14701]= -1931484818;
assign addr[14702]= -1993396407;
assign addr[14703]= -2045196100;
assign addr[14704]= -2086621133;
assign addr[14705]= -2117461370;
assign addr[14706]= -2137560369;
assign addr[14707]= -2146816171;
assign addr[14708]= -2145181827;
assign addr[14709]= -2132665626;
assign addr[14710]= -2109331059;
assign addr[14711]= -2075296495;
assign addr[14712]= -2030734582;
assign addr[14713]= -1975871368;
assign addr[14714]= -1910985158;
assign addr[14715]= -1836405100;
assign addr[14716]= -1752509516;
assign addr[14717]= -1659723983;
assign addr[14718]= -1558519173;
assign addr[14719]= -1449408469;
assign addr[14720]= -1332945355;
assign addr[14721]= -1209720613;
assign addr[14722]= -1080359326;
assign addr[14723]= -945517704;
assign addr[14724]= -805879757;
assign addr[14725]= -662153826;
assign addr[14726]= -515068990;
assign addr[14727]= -365371365;
assign addr[14728]= -213820322;
assign addr[14729]= -61184634;
assign addr[14730]= 91761426;
assign addr[14731]= 244242007;
assign addr[14732]= 395483624;
assign addr[14733]= 544719071;
assign addr[14734]= 691191324;
assign addr[14735]= 834157373;
assign addr[14736]= 972891995;
assign addr[14737]= 1106691431;
assign addr[14738]= 1234876957;
assign addr[14739]= 1356798326;
assign addr[14740]= 1471837070;
assign addr[14741]= 1579409630;
assign addr[14742]= 1678970324;
assign addr[14743]= 1770014111;
assign addr[14744]= 1852079154;
assign addr[14745]= 1924749160;
assign addr[14746]= 1987655498;
assign addr[14747]= 2040479063;
assign addr[14748]= 2082951896;
assign addr[14749]= 2114858546;
assign addr[14750]= 2136037160;
assign addr[14751]= 2146380306;
assign addr[14752]= 2145835515;
assign addr[14753]= 2134405552;
assign addr[14754]= 2112148396;
assign addr[14755]= 2079176953;
assign addr[14756]= 2035658475;
assign addr[14757]= 1981813720;
assign addr[14758]= 1917915825;
assign addr[14759]= 1844288924;
assign addr[14760]= 1761306505;
assign addr[14761]= 1669389513;
assign addr[14762]= 1569004214;
assign addr[14763]= 1460659832;
assign addr[14764]= 1344905966;
assign addr[14765]= 1222329801;
assign addr[14766]= 1093553126;
assign addr[14767]= 959229189;
assign addr[14768]= 820039373;
assign addr[14769]= 676689746;
assign addr[14770]= 529907477;
assign addr[14771]= 380437148;
assign addr[14772]= 229036977;
assign addr[14773]= 76474970;
assign addr[14774]= -76474970;
assign addr[14775]= -229036977;
assign addr[14776]= -380437148;
assign addr[14777]= -529907477;
assign addr[14778]= -676689746;
assign addr[14779]= -820039373;
assign addr[14780]= -959229189;
assign addr[14781]= -1093553126;
assign addr[14782]= -1222329801;
assign addr[14783]= -1344905966;
assign addr[14784]= -1460659832;
assign addr[14785]= -1569004214;
assign addr[14786]= -1669389513;
assign addr[14787]= -1761306505;
assign addr[14788]= -1844288924;
assign addr[14789]= -1917915825;
assign addr[14790]= -1981813720;
assign addr[14791]= -2035658475;
assign addr[14792]= -2079176953;
assign addr[14793]= -2112148396;
assign addr[14794]= -2134405552;
assign addr[14795]= -2145835515;
assign addr[14796]= -2146380306;
assign addr[14797]= -2136037160;
assign addr[14798]= -2114858546;
assign addr[14799]= -2082951896;
assign addr[14800]= -2040479063;
assign addr[14801]= -1987655498;
assign addr[14802]= -1924749160;
assign addr[14803]= -1852079154;
assign addr[14804]= -1770014111;
assign addr[14805]= -1678970324;
assign addr[14806]= -1579409630;
assign addr[14807]= -1471837070;
assign addr[14808]= -1356798326;
assign addr[14809]= -1234876957;
assign addr[14810]= -1106691431;
assign addr[14811]= -972891995;
assign addr[14812]= -834157373;
assign addr[14813]= -691191324;
assign addr[14814]= -544719071;
assign addr[14815]= -395483624;
assign addr[14816]= -244242007;
assign addr[14817]= -91761426;
assign addr[14818]= 61184634;
assign addr[14819]= 213820322;
assign addr[14820]= 365371365;
assign addr[14821]= 515068990;
assign addr[14822]= 662153826;
assign addr[14823]= 805879757;
assign addr[14824]= 945517704;
assign addr[14825]= 1080359326;
assign addr[14826]= 1209720613;
assign addr[14827]= 1332945355;
assign addr[14828]= 1449408469;
assign addr[14829]= 1558519173;
assign addr[14830]= 1659723983;
assign addr[14831]= 1752509516;
assign addr[14832]= 1836405100;
assign addr[14833]= 1910985158;
assign addr[14834]= 1975871368;
assign addr[14835]= 2030734582;
assign addr[14836]= 2075296495;
assign addr[14837]= 2109331059;
assign addr[14838]= 2132665626;
assign addr[14839]= 2145181827;
assign addr[14840]= 2146816171;
assign addr[14841]= 2137560369;
assign addr[14842]= 2117461370;
assign addr[14843]= 2086621133;
assign addr[14844]= 2045196100;
assign addr[14845]= 1993396407;
assign addr[14846]= 1931484818;
assign addr[14847]= 1859775393;
assign addr[14848]= 1778631892;
assign addr[14849]= 1688465931;
assign addr[14850]= 1589734894;
assign addr[14851]= 1482939614;
assign addr[14852]= 1368621831;
assign addr[14853]= 1247361445;
assign addr[14854]= 1119773573;
assign addr[14855]= 986505429;
assign addr[14856]= 848233042;
assign addr[14857]= 705657826;
assign addr[14858]= 559503022;
assign addr[14859]= 410510029;
assign addr[14860]= 259434643;
assign addr[14861]= 107043224;
assign addr[14862]= -45891193;
assign addr[14863]= -198592817;
assign addr[14864]= -350287041;
assign addr[14865]= -500204365;
assign addr[14866]= -647584304;
assign addr[14867]= -791679244;
assign addr[14868]= -931758235;
assign addr[14869]= -1067110699;
assign addr[14870]= -1197050035;
assign addr[14871]= -1320917099;
assign addr[14872]= -1438083551;
assign addr[14873]= -1547955041;
assign addr[14874]= -1649974225;
assign addr[14875]= -1743623590;
assign addr[14876]= -1828428082;
assign addr[14877]= -1903957513;
assign addr[14878]= -1969828744;
assign addr[14879]= -2025707632;
assign addr[14880]= -2071310720;
assign addr[14881]= -2106406677;
assign addr[14882]= -2130817471;
assign addr[14883]= -2144419275;
assign addr[14884]= -2147143090;
assign addr[14885]= -2138975100;
assign addr[14886]= -2119956737;
assign addr[14887]= -2090184478;
assign addr[14888]= -2049809346;
assign addr[14889]= -1999036154;
assign addr[14890]= -1938122457;
assign addr[14891]= -1867377253;
assign addr[14892]= -1787159411;
assign addr[14893]= -1697875851;
assign addr[14894]= -1599979481;
assign addr[14895]= -1493966902;
assign addr[14896]= -1380375881;
assign addr[14897]= -1259782632;
assign addr[14898]= -1132798888;
assign addr[14899]= -1000068799;
assign addr[14900]= -862265664;
assign addr[14901]= -720088517;
assign addr[14902]= -574258580;
assign addr[14903]= -425515602;
assign addr[14904]= -274614114;
assign addr[14905]= -122319591;
assign addr[14906]= 30595422;
assign addr[14907]= 183355234;
assign addr[14908]= 335184940;
assign addr[14909]= 485314355;
assign addr[14910]= 632981917;
assign addr[14911]= 777438554;
assign addr[14912]= 917951481;
assign addr[14913]= 1053807919;
assign addr[14914]= 1184318708;
assign addr[14915]= 1308821808;
assign addr[14916]= 1426685652;
assign addr[14917]= 1537312353;
assign addr[14918]= 1640140734;
assign addr[14919]= 1734649179;
assign addr[14920]= 1820358275;
assign addr[14921]= 1896833245;
assign addr[14922]= 1963686155;
assign addr[14923]= 2020577882;
assign addr[14924]= 2067219829;
assign addr[14925]= 2103375398;
assign addr[14926]= 2128861181;
assign addr[14927]= 2143547897;
assign addr[14928]= 2147361045;
assign addr[14929]= 2140281282;
assign addr[14930]= 2122344521;
assign addr[14931]= 2093641749;
assign addr[14932]= 2054318569;
assign addr[14933]= 2004574453;
assign addr[14934]= 1944661739;
assign addr[14935]= 1874884346;
assign addr[14936]= 1795596234;
assign addr[14937]= 1707199606;
assign addr[14938]= 1610142873;
assign addr[14939]= 1504918373;
assign addr[14940]= 1392059879;
assign addr[14941]= 1272139887;
assign addr[14942]= 1145766716;
assign addr[14943]= 1013581418;
assign addr[14944]= 876254528;
assign addr[14945]= 734482665;
assign addr[14946]= 588984994;
assign addr[14947]= 440499581;
assign addr[14948]= 289779648;
assign addr[14949]= 137589750;
assign addr[14950]= -15298099;
assign addr[14951]= -168108346;
assign addr[14952]= -320065829;
assign addr[14953]= -470399716;
assign addr[14954]= -618347408;
assign addr[14955]= -763158411;
assign addr[14956]= -904098143;
assign addr[14957]= -1040451659;
assign addr[14958]= -1171527280;
assign addr[14959]= -1296660098;
assign addr[14960]= -1415215352;
assign addr[14961]= -1526591649;
assign addr[14962]= -1630224009;
assign addr[14963]= -1725586737;
assign addr[14964]= -1812196087;
assign addr[14965]= -1889612716;
assign addr[14966]= -1957443913;
assign addr[14967]= -2015345591;
assign addr[14968]= -2063024031;
assign addr[14969]= -2100237377;
assign addr[14970]= -2126796855;
assign addr[14971]= -2142567738;
assign addr[14972]= -2147470025;
assign addr[14973]= -2141478848;
assign addr[14974]= -2124624598;
assign addr[14975]= -2096992772;
assign addr[14976]= -2058723538;
assign addr[14977]= -2010011024;
assign addr[14978]= -1951102334;
assign addr[14979]= -1882296293;
assign addr[14980]= -1803941934;
assign addr[14981]= -1716436725;
assign addr[14982]= -1620224553;
assign addr[14983]= -1515793473;
assign addr[14984]= -1403673233;
assign addr[14985]= -1284432584;
assign addr[14986]= -1158676398;
assign addr[14987]= -1027042599;
assign addr[14988]= -890198924;
assign addr[14989]= -748839539;
assign addr[14990]= -603681519;
assign addr[14991]= -455461206;
assign addr[14992]= -304930476;
assign addr[14993]= -152852926;
assign addr[14994]= 0;
assign addr[14995]= 152852926;
assign addr[14996]= 304930476;
assign addr[14997]= 455461206;
assign addr[14998]= 603681519;
assign addr[14999]= 748839539;
assign addr[15000]= 890198924;
assign addr[15001]= 1027042599;
assign addr[15002]= 1158676398;
assign addr[15003]= 1284432584;
assign addr[15004]= 1403673233;
assign addr[15005]= 1515793473;
assign addr[15006]= 1620224553;
assign addr[15007]= 1716436725;
assign addr[15008]= 1803941934;
assign addr[15009]= 1882296293;
assign addr[15010]= 1951102334;
assign addr[15011]= 2010011024;
assign addr[15012]= 2058723538;
assign addr[15013]= 2096992772;
assign addr[15014]= 2124624598;
assign addr[15015]= 2141478848;
assign addr[15016]= 2147470025;
assign addr[15017]= 2142567738;
assign addr[15018]= 2126796855;
assign addr[15019]= 2100237377;
assign addr[15020]= 2063024031;
assign addr[15021]= 2015345591;
assign addr[15022]= 1957443913;
assign addr[15023]= 1889612716;
assign addr[15024]= 1812196087;
assign addr[15025]= 1725586737;
assign addr[15026]= 1630224009;
assign addr[15027]= 1526591649;
assign addr[15028]= 1415215352;
assign addr[15029]= 1296660098;
assign addr[15030]= 1171527280;
assign addr[15031]= 1040451659;
assign addr[15032]= 904098143;
assign addr[15033]= 763158411;
assign addr[15034]= 618347408;
assign addr[15035]= 470399716;
assign addr[15036]= 320065829;
assign addr[15037]= 168108346;
assign addr[15038]= 15298099;
assign addr[15039]= -137589750;
assign addr[15040]= -289779648;
assign addr[15041]= -440499581;
assign addr[15042]= -588984994;
assign addr[15043]= -734482665;
assign addr[15044]= -876254528;
assign addr[15045]= -1013581418;
assign addr[15046]= -1145766716;
assign addr[15047]= -1272139887;
assign addr[15048]= -1392059879;
assign addr[15049]= -1504918373;
assign addr[15050]= -1610142873;
assign addr[15051]= -1707199606;
assign addr[15052]= -1795596234;
assign addr[15053]= -1874884346;
assign addr[15054]= -1944661739;
assign addr[15055]= -2004574453;
assign addr[15056]= -2054318569;
assign addr[15057]= -2093641749;
assign addr[15058]= -2122344521;
assign addr[15059]= -2140281282;
assign addr[15060]= -2147361045;
assign addr[15061]= -2143547897;
assign addr[15062]= -2128861181;
assign addr[15063]= -2103375398;
assign addr[15064]= -2067219829;
assign addr[15065]= -2020577882;
assign addr[15066]= -1963686155;
assign addr[15067]= -1896833245;
assign addr[15068]= -1820358275;
assign addr[15069]= -1734649179;
assign addr[15070]= -1640140734;
assign addr[15071]= -1537312353;
assign addr[15072]= -1426685652;
assign addr[15073]= -1308821808;
assign addr[15074]= -1184318708;
assign addr[15075]= -1053807919;
assign addr[15076]= -917951481;
assign addr[15077]= -777438554;
assign addr[15078]= -632981917;
assign addr[15079]= -485314355;
assign addr[15080]= -335184940;
assign addr[15081]= -183355234;
assign addr[15082]= -30595422;
assign addr[15083]= 122319591;
assign addr[15084]= 274614114;
assign addr[15085]= 425515602;
assign addr[15086]= 574258580;
assign addr[15087]= 720088517;
assign addr[15088]= 862265664;
assign addr[15089]= 1000068799;
assign addr[15090]= 1132798888;
assign addr[15091]= 1259782632;
assign addr[15092]= 1380375881;
assign addr[15093]= 1493966902;
assign addr[15094]= 1599979481;
assign addr[15095]= 1697875851;
assign addr[15096]= 1787159411;
assign addr[15097]= 1867377253;
assign addr[15098]= 1938122457;
assign addr[15099]= 1999036154;
assign addr[15100]= 2049809346;
assign addr[15101]= 2090184478;
assign addr[15102]= 2119956737;
assign addr[15103]= 2138975100;
assign addr[15104]= 2147143090;
assign addr[15105]= 2144419275;
assign addr[15106]= 2130817471;
assign addr[15107]= 2106406677;
assign addr[15108]= 2071310720;
assign addr[15109]= 2025707632;
assign addr[15110]= 1969828744;
assign addr[15111]= 1903957513;
assign addr[15112]= 1828428082;
assign addr[15113]= 1743623590;
assign addr[15114]= 1649974225;
assign addr[15115]= 1547955041;
assign addr[15116]= 1438083551;
assign addr[15117]= 1320917099;
assign addr[15118]= 1197050035;
assign addr[15119]= 1067110699;
assign addr[15120]= 931758235;
assign addr[15121]= 791679244;
assign addr[15122]= 647584304;
assign addr[15123]= 500204365;
assign addr[15124]= 350287041;
assign addr[15125]= 198592817;
assign addr[15126]= 45891193;
assign addr[15127]= -107043224;
assign addr[15128]= -259434643;
assign addr[15129]= -410510029;
assign addr[15130]= -559503022;
assign addr[15131]= -705657826;
assign addr[15132]= -848233042;
assign addr[15133]= -986505429;
assign addr[15134]= -1119773573;
assign addr[15135]= -1247361445;
assign addr[15136]= -1368621831;
assign addr[15137]= -1482939614;
assign addr[15138]= -1589734894;
assign addr[15139]= -1688465931;
assign addr[15140]= -1778631892;
assign addr[15141]= -1859775393;
assign addr[15142]= -1931484818;
assign addr[15143]= -1993396407;
assign addr[15144]= -2045196100;
assign addr[15145]= -2086621133;
assign addr[15146]= -2117461370;
assign addr[15147]= -2137560369;
assign addr[15148]= -2146816171;
assign addr[15149]= -2145181827;
assign addr[15150]= -2132665626;
assign addr[15151]= -2109331059;
assign addr[15152]= -2075296495;
assign addr[15153]= -2030734582;
assign addr[15154]= -1975871368;
assign addr[15155]= -1910985158;
assign addr[15156]= -1836405100;
assign addr[15157]= -1752509516;
assign addr[15158]= -1659723983;
assign addr[15159]= -1558519173;
assign addr[15160]= -1449408469;
assign addr[15161]= -1332945355;
assign addr[15162]= -1209720613;
assign addr[15163]= -1080359326;
assign addr[15164]= -945517704;
assign addr[15165]= -805879757;
assign addr[15166]= -662153826;
assign addr[15167]= -515068990;
assign addr[15168]= -365371365;
assign addr[15169]= -213820322;
assign addr[15170]= -61184634;
assign addr[15171]= 91761426;
assign addr[15172]= 244242007;
assign addr[15173]= 395483624;
assign addr[15174]= 544719071;
assign addr[15175]= 691191324;
assign addr[15176]= 834157373;
assign addr[15177]= 972891995;
assign addr[15178]= 1106691431;
assign addr[15179]= 1234876957;
assign addr[15180]= 1356798326;
assign addr[15181]= 1471837070;
assign addr[15182]= 1579409630;
assign addr[15183]= 1678970324;
assign addr[15184]= 1770014111;
assign addr[15185]= 1852079154;
assign addr[15186]= 1924749160;
assign addr[15187]= 1987655498;
assign addr[15188]= 2040479063;
assign addr[15189]= 2082951896;
assign addr[15190]= 2114858546;
assign addr[15191]= 2136037160;
assign addr[15192]= 2146380306;
assign addr[15193]= 2145835515;
assign addr[15194]= 2134405552;
assign addr[15195]= 2112148396;
assign addr[15196]= 2079176953;
assign addr[15197]= 2035658475;
assign addr[15198]= 1981813720;
assign addr[15199]= 1917915825;
assign addr[15200]= 1844288924;
assign addr[15201]= 1761306505;
assign addr[15202]= 1669389513;
assign addr[15203]= 1569004214;
assign addr[15204]= 1460659832;
assign addr[15205]= 1344905966;
assign addr[15206]= 1222329801;
assign addr[15207]= 1093553126;
assign addr[15208]= 959229189;
assign addr[15209]= 820039373;
assign addr[15210]= 676689746;
assign addr[15211]= 529907477;
assign addr[15212]= 380437148;
assign addr[15213]= 229036977;
assign addr[15214]= 76474970;
assign addr[15215]= -76474970;
assign addr[15216]= -229036977;
assign addr[15217]= -380437148;
assign addr[15218]= -529907477;
assign addr[15219]= -676689746;
assign addr[15220]= -820039373;
assign addr[15221]= -959229189;
assign addr[15222]= -1093553126;
assign addr[15223]= -1222329801;
assign addr[15224]= -1344905966;
assign addr[15225]= -1460659832;
assign addr[15226]= -1569004214;
assign addr[15227]= -1669389513;
assign addr[15228]= -1761306505;
assign addr[15229]= -1844288924;
assign addr[15230]= -1917915825;
assign addr[15231]= -1981813720;
assign addr[15232]= -2035658475;
assign addr[15233]= -2079176953;
assign addr[15234]= -2112148396;
assign addr[15235]= -2134405552;
assign addr[15236]= -2145835515;
assign addr[15237]= -2146380306;
assign addr[15238]= -2136037160;
assign addr[15239]= -2114858546;
assign addr[15240]= -2082951896;
assign addr[15241]= -2040479063;
assign addr[15242]= -1987655498;
assign addr[15243]= -1924749160;
assign addr[15244]= -1852079154;
assign addr[15245]= -1770014111;
assign addr[15246]= -1678970324;
assign addr[15247]= -1579409630;
assign addr[15248]= -1471837070;
assign addr[15249]= -1356798326;
assign addr[15250]= -1234876957;
assign addr[15251]= -1106691431;
assign addr[15252]= -972891995;
assign addr[15253]= -834157373;
assign addr[15254]= -691191324;
assign addr[15255]= -544719071;
assign addr[15256]= -395483624;
assign addr[15257]= -244242007;
assign addr[15258]= -91761426;
assign addr[15259]= 61184634;
assign addr[15260]= 213820322;
assign addr[15261]= 365371365;
assign addr[15262]= 515068990;
assign addr[15263]= 662153826;
assign addr[15264]= 805879757;
assign addr[15265]= 945517704;
assign addr[15266]= 1080359326;
assign addr[15267]= 1209720613;
assign addr[15268]= 1332945355;
assign addr[15269]= 1449408469;
assign addr[15270]= 1558519173;
assign addr[15271]= 1659723983;
assign addr[15272]= 1752509516;
assign addr[15273]= 1836405100;
assign addr[15274]= 1910985158;
assign addr[15275]= 1975871368;
assign addr[15276]= 2030734582;
assign addr[15277]= 2075296495;
assign addr[15278]= 2109331059;
assign addr[15279]= 2132665626;
assign addr[15280]= 2145181827;
assign addr[15281]= 2146816171;
assign addr[15282]= 2137560369;
assign addr[15283]= 2117461370;
assign addr[15284]= 2086621133;
assign addr[15285]= 2045196100;
assign addr[15286]= 1993396407;
assign addr[15287]= 1931484818;
assign addr[15288]= 1859775393;
assign addr[15289]= 1778631892;
assign addr[15290]= 1688465931;
assign addr[15291]= 1589734894;
assign addr[15292]= 1482939614;
assign addr[15293]= 1368621831;
assign addr[15294]= 1247361445;
assign addr[15295]= 1119773573;
assign addr[15296]= 986505429;
assign addr[15297]= 848233042;
assign addr[15298]= 705657826;
assign addr[15299]= 559503022;
assign addr[15300]= 410510029;
assign addr[15301]= 259434643;
assign addr[15302]= 107043224;
assign addr[15303]= -45891193;
assign addr[15304]= -198592817;
assign addr[15305]= -350287041;
assign addr[15306]= -500204365;
assign addr[15307]= -647584304;
assign addr[15308]= -791679244;
assign addr[15309]= -931758235;
assign addr[15310]= -1067110699;
assign addr[15311]= -1197050035;
assign addr[15312]= -1320917099;
assign addr[15313]= -1438083551;
assign addr[15314]= -1547955041;
assign addr[15315]= -1649974225;
assign addr[15316]= -1743623590;
assign addr[15317]= -1828428082;
assign addr[15318]= -1903957513;
assign addr[15319]= -1969828744;
assign addr[15320]= -2025707632;
assign addr[15321]= -2071310720;
assign addr[15322]= -2106406677;
assign addr[15323]= -2130817471;
assign addr[15324]= -2144419275;
assign addr[15325]= -2147143090;
assign addr[15326]= -2138975100;
assign addr[15327]= -2119956737;
assign addr[15328]= -2090184478;
assign addr[15329]= -2049809346;
assign addr[15330]= -1999036154;
assign addr[15331]= -1938122457;
assign addr[15332]= -1867377253;
assign addr[15333]= -1787159411;
assign addr[15334]= -1697875851;
assign addr[15335]= -1599979481;
assign addr[15336]= -1493966902;
assign addr[15337]= -1380375881;
assign addr[15338]= -1259782632;
assign addr[15339]= -1132798888;
assign addr[15340]= -1000068799;
assign addr[15341]= -862265664;
assign addr[15342]= -720088517;
assign addr[15343]= -574258580;
assign addr[15344]= -425515602;
assign addr[15345]= -274614114;
assign addr[15346]= -122319591;
assign addr[15347]= 30595422;
assign addr[15348]= 183355234;
assign addr[15349]= 335184940;
assign addr[15350]= 485314355;
assign addr[15351]= 632981917;
assign addr[15352]= 777438554;
assign addr[15353]= 917951481;
assign addr[15354]= 1053807919;
assign addr[15355]= 1184318708;
assign addr[15356]= 1308821808;
assign addr[15357]= 1426685652;
assign addr[15358]= 1537312353;
assign addr[15359]= 1640140734;
assign addr[15360]= 1734649179;
assign addr[15361]= 1820358275;
assign addr[15362]= 1896833245;
assign addr[15363]= 1963686155;
assign addr[15364]= 2020577882;
assign addr[15365]= 2067219829;
assign addr[15366]= 2103375398;
assign addr[15367]= 2128861181;
assign addr[15368]= 2143547897;
assign addr[15369]= 2147361045;
assign addr[15370]= 2140281282;
assign addr[15371]= 2122344521;
assign addr[15372]= 2093641749;
assign addr[15373]= 2054318569;
assign addr[15374]= 2004574453;
assign addr[15375]= 1944661739;
assign addr[15376]= 1874884346;
assign addr[15377]= 1795596234;
assign addr[15378]= 1707199606;
assign addr[15379]= 1610142873;
assign addr[15380]= 1504918373;
assign addr[15381]= 1392059879;
assign addr[15382]= 1272139887;
assign addr[15383]= 1145766716;
assign addr[15384]= 1013581418;
assign addr[15385]= 876254528;
assign addr[15386]= 734482665;
assign addr[15387]= 588984994;
assign addr[15388]= 440499581;
assign addr[15389]= 289779648;
assign addr[15390]= 137589750;
assign addr[15391]= -15298099;
assign addr[15392]= -168108346;
assign addr[15393]= -320065829;
assign addr[15394]= -470399716;
assign addr[15395]= -618347408;
assign addr[15396]= -763158411;
assign addr[15397]= -904098143;
assign addr[15398]= -1040451659;
assign addr[15399]= -1171527280;
assign addr[15400]= -1296660098;
assign addr[15401]= -1415215352;
assign addr[15402]= -1526591649;
assign addr[15403]= -1630224009;
assign addr[15404]= -1725586737;
assign addr[15405]= -1812196087;
assign addr[15406]= -1889612716;
assign addr[15407]= -1957443913;
assign addr[15408]= -2015345591;
assign addr[15409]= -2063024031;
assign addr[15410]= -2100237377;
assign addr[15411]= -2126796855;
assign addr[15412]= -2142567738;
assign addr[15413]= -2147470025;
assign addr[15414]= -2141478848;
assign addr[15415]= -2124624598;
assign addr[15416]= -2096992772;
assign addr[15417]= -2058723538;
assign addr[15418]= -2010011024;
assign addr[15419]= -1951102334;
assign addr[15420]= -1882296293;
assign addr[15421]= -1803941934;
assign addr[15422]= -1716436725;
assign addr[15423]= -1620224553;
assign addr[15424]= -1515793473;
assign addr[15425]= -1403673233;
assign addr[15426]= -1284432584;
assign addr[15427]= -1158676398;
assign addr[15428]= -1027042599;
assign addr[15429]= -890198924;
assign addr[15430]= -748839539;
assign addr[15431]= -603681519;
assign addr[15432]= -455461206;
assign addr[15433]= -304930476;
assign addr[15434]= -152852926;
assign addr[15435]= 0;
assign addr[15436]= 152852926;
assign addr[15437]= 304930476;
assign addr[15438]= 455461206;
assign addr[15439]= 603681519;
assign addr[15440]= 748839539;
assign addr[15441]= 890198924;
assign addr[15442]= 1027042599;
assign addr[15443]= 1158676398;
assign addr[15444]= 1284432584;
assign addr[15445]= 1403673233;
assign addr[15446]= 1515793473;
assign addr[15447]= 1620224553;
assign addr[15448]= 1716436725;
assign addr[15449]= 1803941934;
assign addr[15450]= 1882296293;
assign addr[15451]= 1951102334;
assign addr[15452]= 2010011024;
assign addr[15453]= 2058723538;
assign addr[15454]= 2096992772;
assign addr[15455]= 2124624598;
assign addr[15456]= 2141478848;
assign addr[15457]= 2147470025;
assign addr[15458]= 2142567738;
assign addr[15459]= 2126796855;
assign addr[15460]= 2100237377;
assign addr[15461]= 2063024031;
assign addr[15462]= 2015345591;
assign addr[15463]= 1957443913;
assign addr[15464]= 1889612716;
assign addr[15465]= 1812196087;
assign addr[15466]= 1725586737;
assign addr[15467]= 1630224009;
assign addr[15468]= 1526591649;
assign addr[15469]= 1415215352;
assign addr[15470]= 1296660098;
assign addr[15471]= 1171527280;
assign addr[15472]= 1040451659;
assign addr[15473]= 904098143;
assign addr[15474]= 763158411;
assign addr[15475]= 618347408;
assign addr[15476]= 470399716;
assign addr[15477]= 320065829;
assign addr[15478]= 168108346;
assign addr[15479]= 15298099;
assign addr[15480]= -137589750;
assign addr[15481]= -289779648;
assign addr[15482]= -440499581;
assign addr[15483]= -588984994;
assign addr[15484]= -734482665;
assign addr[15485]= -876254528;
assign addr[15486]= -1013581418;
assign addr[15487]= -1145766716;
assign addr[15488]= -1272139887;
assign addr[15489]= -1392059879;
assign addr[15490]= -1504918373;
assign addr[15491]= -1610142873;
assign addr[15492]= -1707199606;
assign addr[15493]= -1795596234;
assign addr[15494]= -1874884346;
assign addr[15495]= -1944661739;
assign addr[15496]= -2004574453;
assign addr[15497]= -2054318569;
assign addr[15498]= -2093641749;
assign addr[15499]= -2122344521;
assign addr[15500]= -2140281282;
assign addr[15501]= -2147361045;
assign addr[15502]= -2143547897;
assign addr[15503]= -2128861181;
assign addr[15504]= -2103375398;
assign addr[15505]= -2067219829;
assign addr[15506]= -2020577882;
assign addr[15507]= -1963686155;
assign addr[15508]= -1896833245;
assign addr[15509]= -1820358275;
assign addr[15510]= -1734649179;
assign addr[15511]= -1640140734;
assign addr[15512]= -1537312353;
assign addr[15513]= -1426685652;
assign addr[15514]= -1308821808;
assign addr[15515]= -1184318708;
assign addr[15516]= -1053807919;
assign addr[15517]= -917951481;
assign addr[15518]= -777438554;
assign addr[15519]= -632981917;
assign addr[15520]= -485314355;
assign addr[15521]= -335184940;
assign addr[15522]= -183355234;
assign addr[15523]= -30595422;
assign addr[15524]= 122319591;
assign addr[15525]= 274614114;
assign addr[15526]= 425515602;
assign addr[15527]= 574258580;
assign addr[15528]= 720088517;
assign addr[15529]= 862265664;
assign addr[15530]= 1000068799;
assign addr[15531]= 1132798888;
assign addr[15532]= 1259782632;
assign addr[15533]= 1380375881;
assign addr[15534]= 1493966902;
assign addr[15535]= 1599979481;
assign addr[15536]= 1697875851;
assign addr[15537]= 1787159411;
assign addr[15538]= 1867377253;
assign addr[15539]= 1938122457;
assign addr[15540]= 1999036154;
assign addr[15541]= 2049809346;
assign addr[15542]= 2090184478;
assign addr[15543]= 2119956737;
assign addr[15544]= 2138975100;
assign addr[15545]= 2147143090;
assign addr[15546]= 2144419275;
assign addr[15547]= 2130817471;
assign addr[15548]= 2106406677;
assign addr[15549]= 2071310720;
assign addr[15550]= 2025707632;
assign addr[15551]= 1969828744;
assign addr[15552]= 1903957513;
assign addr[15553]= 1828428082;
assign addr[15554]= 1743623590;
assign addr[15555]= 1649974225;
assign addr[15556]= 1547955041;
assign addr[15557]= 1438083551;
assign addr[15558]= 1320917099;
assign addr[15559]= 1197050035;
assign addr[15560]= 1067110699;
assign addr[15561]= 931758235;
assign addr[15562]= 791679244;
assign addr[15563]= 647584304;
assign addr[15564]= 500204365;
assign addr[15565]= 350287041;
assign addr[15566]= 198592817;
assign addr[15567]= 45891193;
assign addr[15568]= -107043224;
assign addr[15569]= -259434643;
assign addr[15570]= -410510029;
assign addr[15571]= -559503022;
assign addr[15572]= -705657826;
assign addr[15573]= -848233042;
assign addr[15574]= -986505429;
assign addr[15575]= -1119773573;
assign addr[15576]= -1247361445;
assign addr[15577]= -1368621831;
assign addr[15578]= -1482939614;
assign addr[15579]= -1589734894;
assign addr[15580]= -1688465931;
assign addr[15581]= -1778631892;
assign addr[15582]= -1859775393;
assign addr[15583]= -1931484818;
assign addr[15584]= -1993396407;
assign addr[15585]= -2045196100;
assign addr[15586]= -2086621133;
assign addr[15587]= -2117461370;
assign addr[15588]= -2137560369;
assign addr[15589]= -2146816171;
assign addr[15590]= -2145181827;
assign addr[15591]= -2132665626;
assign addr[15592]= -2109331059;
assign addr[15593]= -2075296495;
assign addr[15594]= -2030734582;
assign addr[15595]= -1975871368;
assign addr[15596]= -1910985158;
assign addr[15597]= -1836405100;
assign addr[15598]= -1752509516;
assign addr[15599]= -1659723983;
assign addr[15600]= -1558519173;
assign addr[15601]= -1449408469;
assign addr[15602]= -1332945355;
assign addr[15603]= -1209720613;
assign addr[15604]= -1080359326;
assign addr[15605]= -945517704;
assign addr[15606]= -805879757;
assign addr[15607]= -662153826;
assign addr[15608]= -515068990;
assign addr[15609]= -365371365;
assign addr[15610]= -213820322;
assign addr[15611]= -61184634;
assign addr[15612]= 91761426;
assign addr[15613]= 244242007;
assign addr[15614]= 395483624;
assign addr[15615]= 544719071;
assign addr[15616]= 691191324;
assign addr[15617]= 834157373;
assign addr[15618]= 972891995;
assign addr[15619]= 1106691431;
assign addr[15620]= 1234876957;
assign addr[15621]= 1356798326;
assign addr[15622]= 1471837070;
assign addr[15623]= 1579409630;
assign addr[15624]= 1678970324;
assign addr[15625]= 1770014111;
assign addr[15626]= 1852079154;
assign addr[15627]= 1924749160;
assign addr[15628]= 1987655498;
assign addr[15629]= 2040479063;
assign addr[15630]= 2082951896;
assign addr[15631]= 2114858546;
assign addr[15632]= 2136037160;
assign addr[15633]= 2146380306;
assign addr[15634]= 2145835515;
assign addr[15635]= 2134405552;
assign addr[15636]= 2112148396;
assign addr[15637]= 2079176953;
assign addr[15638]= 2035658475;
assign addr[15639]= 1981813720;
assign addr[15640]= 1917915825;
assign addr[15641]= 1844288924;
assign addr[15642]= 1761306505;
assign addr[15643]= 1669389513;
assign addr[15644]= 1569004214;
assign addr[15645]= 1460659832;
assign addr[15646]= 1344905966;
assign addr[15647]= 1222329801;
assign addr[15648]= 1093553126;
assign addr[15649]= 959229189;
assign addr[15650]= 820039373;
assign addr[15651]= 676689746;
assign addr[15652]= 529907477;
assign addr[15653]= 380437148;
assign addr[15654]= 229036977;
assign addr[15655]= 76474970;
assign addr[15656]= -76474970;
assign addr[15657]= -229036977;
assign addr[15658]= -380437148;
assign addr[15659]= -529907477;
assign addr[15660]= -676689746;
assign addr[15661]= -820039373;
assign addr[15662]= -959229189;
assign addr[15663]= -1093553126;
assign addr[15664]= -1222329801;
assign addr[15665]= -1344905966;
assign addr[15666]= -1460659832;
assign addr[15667]= -1569004214;
assign addr[15668]= -1669389513;
assign addr[15669]= -1761306505;
assign addr[15670]= -1844288924;
assign addr[15671]= -1917915825;
assign addr[15672]= -1981813720;
assign addr[15673]= -2035658475;
assign addr[15674]= -2079176953;
assign addr[15675]= -2112148396;
assign addr[15676]= -2134405552;
assign addr[15677]= -2145835515;
assign addr[15678]= -2146380306;
assign addr[15679]= -2136037160;
assign addr[15680]= -2114858546;
assign addr[15681]= -2082951896;
assign addr[15682]= -2040479063;
assign addr[15683]= -1987655498;
assign addr[15684]= -1924749160;
assign addr[15685]= -1852079154;
assign addr[15686]= -1770014111;
assign addr[15687]= -1678970324;
assign addr[15688]= -1579409630;
assign addr[15689]= -1471837070;
assign addr[15690]= -1356798326;
assign addr[15691]= -1234876957;
assign addr[15692]= -1106691431;
assign addr[15693]= -972891995;
assign addr[15694]= -834157373;
assign addr[15695]= -691191324;
assign addr[15696]= -544719071;
assign addr[15697]= -395483624;
assign addr[15698]= -244242007;
assign addr[15699]= -91761426;
assign addr[15700]= 61184634;
assign addr[15701]= 213820322;
assign addr[15702]= 365371365;
assign addr[15703]= 515068990;
assign addr[15704]= 662153826;
assign addr[15705]= 805879757;
assign addr[15706]= 945517704;
assign addr[15707]= 1080359326;
assign addr[15708]= 1209720613;
assign addr[15709]= 1332945355;
assign addr[15710]= 1449408469;
assign addr[15711]= 1558519173;
assign addr[15712]= 1659723983;
assign addr[15713]= 1752509516;
assign addr[15714]= 1836405100;
assign addr[15715]= 1910985158;
assign addr[15716]= 1975871368;
assign addr[15717]= 2030734582;
assign addr[15718]= 2075296495;
assign addr[15719]= 2109331059;
assign addr[15720]= 2132665626;
assign addr[15721]= 2145181827;
assign addr[15722]= 2146816171;
assign addr[15723]= 2137560369;
assign addr[15724]= 2117461370;
assign addr[15725]= 2086621133;
assign addr[15726]= 2045196100;
assign addr[15727]= 1993396407;
assign addr[15728]= 1931484818;
assign addr[15729]= 1859775393;
assign addr[15730]= 1778631892;
assign addr[15731]= 1688465931;
assign addr[15732]= 1589734894;
assign addr[15733]= 1482939614;
assign addr[15734]= 1368621831;
assign addr[15735]= 1247361445;
assign addr[15736]= 1119773573;
assign addr[15737]= 986505429;
assign addr[15738]= 848233042;
assign addr[15739]= 705657826;
assign addr[15740]= 559503022;
assign addr[15741]= 410510029;
assign addr[15742]= 259434643;
assign addr[15743]= 107043224;
assign addr[15744]= -45891193;
assign addr[15745]= -198592817;
assign addr[15746]= -350287041;
assign addr[15747]= -500204365;
assign addr[15748]= -647584304;
assign addr[15749]= -791679244;
assign addr[15750]= -931758235;
assign addr[15751]= -1067110699;
assign addr[15752]= -1197050035;
assign addr[15753]= -1320917099;
assign addr[15754]= -1438083551;
assign addr[15755]= -1547955041;
assign addr[15756]= -1649974225;
assign addr[15757]= -1743623590;
assign addr[15758]= -1828428082;
assign addr[15759]= -1903957513;
assign addr[15760]= -1969828744;
assign addr[15761]= -2025707632;
assign addr[15762]= -2071310720;
assign addr[15763]= -2106406677;
assign addr[15764]= -2130817471;
assign addr[15765]= -2144419275;
assign addr[15766]= -2147143090;
assign addr[15767]= -2138975100;
assign addr[15768]= -2119956737;
assign addr[15769]= -2090184478;
assign addr[15770]= -2049809346;
assign addr[15771]= -1999036154;
assign addr[15772]= -1938122457;
assign addr[15773]= -1867377253;
assign addr[15774]= -1787159411;
assign addr[15775]= -1697875851;
assign addr[15776]= -1599979481;
assign addr[15777]= -1493966902;
assign addr[15778]= -1380375881;
assign addr[15779]= -1259782632;
assign addr[15780]= -1132798888;
assign addr[15781]= -1000068799;
assign addr[15782]= -862265664;
assign addr[15783]= -720088517;
assign addr[15784]= -574258580;
assign addr[15785]= -425515602;
assign addr[15786]= -274614114;
assign addr[15787]= -122319591;
assign addr[15788]= 30595422;
assign addr[15789]= 183355234;
assign addr[15790]= 335184940;
assign addr[15791]= 485314355;
assign addr[15792]= 632981917;
assign addr[15793]= 777438554;
assign addr[15794]= 917951481;
assign addr[15795]= 1053807919;
assign addr[15796]= 1184318708;
assign addr[15797]= 1308821808;
assign addr[15798]= 1426685652;
assign addr[15799]= 1537312353;
assign addr[15800]= 1640140734;
assign addr[15801]= 1734649179;
assign addr[15802]= 1820358275;
assign addr[15803]= 1896833245;
assign addr[15804]= 1963686155;
assign addr[15805]= 2020577882;
assign addr[15806]= 2067219829;
assign addr[15807]= 2103375398;
assign addr[15808]= 2128861181;
assign addr[15809]= 2143547897;
assign addr[15810]= 2147361045;
assign addr[15811]= 2140281282;
assign addr[15812]= 2122344521;
assign addr[15813]= 2093641749;
assign addr[15814]= 2054318569;
assign addr[15815]= 2004574453;
assign addr[15816]= 1944661739;
assign addr[15817]= 1874884346;
assign addr[15818]= 1795596234;
assign addr[15819]= 1707199606;
assign addr[15820]= 1610142873;
assign addr[15821]= 1504918373;
assign addr[15822]= 1392059879;
assign addr[15823]= 1272139887;
assign addr[15824]= 1145766716;
assign addr[15825]= 1013581418;
assign addr[15826]= 876254528;
assign addr[15827]= 734482665;
assign addr[15828]= 588984994;
assign addr[15829]= 440499581;
assign addr[15830]= 289779648;
assign addr[15831]= 137589750;
assign addr[15832]= -15298099;
assign addr[15833]= -168108346;
assign addr[15834]= -320065829;
assign addr[15835]= -470399716;
assign addr[15836]= -618347408;
assign addr[15837]= -763158411;
assign addr[15838]= -904098143;
assign addr[15839]= -1040451659;
assign addr[15840]= -1171527280;
assign addr[15841]= -1296660098;
assign addr[15842]= -1415215352;
assign addr[15843]= -1526591649;
assign addr[15844]= -1630224009;
assign addr[15845]= -1725586737;
assign addr[15846]= -1812196087;
assign addr[15847]= -1889612716;
assign addr[15848]= -1957443913;
assign addr[15849]= -2015345591;
assign addr[15850]= -2063024031;
assign addr[15851]= -2100237377;
assign addr[15852]= -2126796855;
assign addr[15853]= -2142567738;
assign addr[15854]= -2147470025;
assign addr[15855]= -2141478848;
assign addr[15856]= -2124624598;
assign addr[15857]= -2096992772;
assign addr[15858]= -2058723538;
assign addr[15859]= -2010011024;
assign addr[15860]= -1951102334;
assign addr[15861]= -1882296293;
assign addr[15862]= -1803941934;
assign addr[15863]= -1716436725;
assign addr[15864]= -1620224553;
assign addr[15865]= -1515793473;
assign addr[15866]= -1403673233;
assign addr[15867]= -1284432584;
assign addr[15868]= -1158676398;
assign addr[15869]= -1027042599;
assign addr[15870]= -890198924;
assign addr[15871]= -748839539;
assign addr[15872]= -603681519;
assign addr[15873]= -455461206;
assign addr[15874]= -304930476;
assign addr[15875]= -152852926;
assign addr[15876]= 0;
assign addr[15877]= 152852926;
assign addr[15878]= 304930476;
assign addr[15879]= 455461206;
assign addr[15880]= 603681519;
assign addr[15881]= 748839539;
assign addr[15882]= 890198924;
assign addr[15883]= 1027042599;
assign addr[15884]= 1158676398;
assign addr[15885]= 1284432584;
assign addr[15886]= 1403673233;
assign addr[15887]= 1515793473;
assign addr[15888]= 1620224553;
assign addr[15889]= 1716436725;
assign addr[15890]= 1803941934;
assign addr[15891]= 1882296293;
assign addr[15892]= 1951102334;
assign addr[15893]= 2010011024;
assign addr[15894]= 2058723538;
assign addr[15895]= 2096992772;
assign addr[15896]= 2124624598;
assign addr[15897]= 2141478848;
assign addr[15898]= 2147470025;
assign addr[15899]= 2142567738;
assign addr[15900]= 2126796855;
assign addr[15901]= 2100237377;
assign addr[15902]= 2063024031;
assign addr[15903]= 2015345591;
assign addr[15904]= 1957443913;
assign addr[15905]= 1889612716;
assign addr[15906]= 1812196087;
assign addr[15907]= 1725586737;
assign addr[15908]= 1630224009;
assign addr[15909]= 1526591649;
assign addr[15910]= 1415215352;
assign addr[15911]= 1296660098;
assign addr[15912]= 1171527280;
assign addr[15913]= 1040451659;
assign addr[15914]= 904098143;
assign addr[15915]= 763158411;
assign addr[15916]= 618347408;
assign addr[15917]= 470399716;
assign addr[15918]= 320065829;
assign addr[15919]= 168108346;
assign addr[15920]= 15298099;
assign addr[15921]= -137589750;
assign addr[15922]= -289779648;
assign addr[15923]= -440499581;
assign addr[15924]= -588984994;
assign addr[15925]= -734482665;
assign addr[15926]= -876254528;
assign addr[15927]= -1013581418;
assign addr[15928]= -1145766716;
assign addr[15929]= -1272139887;
assign addr[15930]= -1392059879;
assign addr[15931]= -1504918373;
assign addr[15932]= -1610142873;
assign addr[15933]= -1707199606;
assign addr[15934]= -1795596234;
assign addr[15935]= -1874884346;
assign addr[15936]= -1944661739;
assign addr[15937]= -2004574453;
assign addr[15938]= -2054318569;
assign addr[15939]= -2093641749;
assign addr[15940]= -2122344521;
assign addr[15941]= -2140281282;
assign addr[15942]= -2147361045;
assign addr[15943]= -2143547897;
assign addr[15944]= -2128861181;
assign addr[15945]= -2103375398;
assign addr[15946]= -2067219829;
assign addr[15947]= -2020577882;
assign addr[15948]= -1963686155;
assign addr[15949]= -1896833245;
assign addr[15950]= -1820358275;
assign addr[15951]= -1734649179;
assign addr[15952]= -1640140734;
assign addr[15953]= -1537312353;
assign addr[15954]= -1426685652;
assign addr[15955]= -1308821808;
assign addr[15956]= -1184318708;
assign addr[15957]= -1053807919;
assign addr[15958]= -917951481;
assign addr[15959]= -777438554;
assign addr[15960]= -632981917;
assign addr[15961]= -485314355;
assign addr[15962]= -335184940;
assign addr[15963]= -183355234;
assign addr[15964]= -30595422;
assign addr[15965]= 122319591;
assign addr[15966]= 274614114;
assign addr[15967]= 425515602;
assign addr[15968]= 574258580;
assign addr[15969]= 720088517;
assign addr[15970]= 862265664;
assign addr[15971]= 1000068799;
assign addr[15972]= 1132798888;
assign addr[15973]= 1259782632;
assign addr[15974]= 1380375881;
assign addr[15975]= 1493966902;
assign addr[15976]= 1599979481;
assign addr[15977]= 1697875851;
assign addr[15978]= 1787159411;
assign addr[15979]= 1867377253;
assign addr[15980]= 1938122457;
assign addr[15981]= 1999036154;
assign addr[15982]= 2049809346;
assign addr[15983]= 2090184478;
assign addr[15984]= 2119956737;
assign addr[15985]= 2138975100;
assign addr[15986]= 2147143090;
assign addr[15987]= 2144419275;
assign addr[15988]= 2130817471;
assign addr[15989]= 2106406677;
assign addr[15990]= 2071310720;
assign addr[15991]= 2025707632;
assign addr[15992]= 1969828744;
assign addr[15993]= 1903957513;
assign addr[15994]= 1828428082;
assign addr[15995]= 1743623590;
assign addr[15996]= 1649974225;
assign addr[15997]= 1547955041;
assign addr[15998]= 1438083551;
assign addr[15999]= 1320917099;
assign addr[16000]= 1197050035;
assign addr[16001]= 1067110699;
assign addr[16002]= 931758235;
assign addr[16003]= 791679244;
assign addr[16004]= 647584304;
assign addr[16005]= 500204365;
assign addr[16006]= 350287041;
assign addr[16007]= 198592817;
assign addr[16008]= 45891193;
assign addr[16009]= -107043224;
assign addr[16010]= -259434643;
assign addr[16011]= -410510029;
assign addr[16012]= -559503022;
assign addr[16013]= -705657826;
assign addr[16014]= -848233042;
assign addr[16015]= -986505429;
assign addr[16016]= -1119773573;
assign addr[16017]= -1247361445;
assign addr[16018]= -1368621831;
assign addr[16019]= -1482939614;
assign addr[16020]= -1589734894;
assign addr[16021]= -1688465931;
assign addr[16022]= -1778631892;
assign addr[16023]= -1859775393;
assign addr[16024]= -1931484818;
assign addr[16025]= -1993396407;
assign addr[16026]= -2045196100;
assign addr[16027]= -2086621133;
assign addr[16028]= -2117461370;
assign addr[16029]= -2137560369;
assign addr[16030]= -2146816171;
assign addr[16031]= -2145181827;
assign addr[16032]= -2132665626;
assign addr[16033]= -2109331059;
assign addr[16034]= -2075296495;
assign addr[16035]= -2030734582;
assign addr[16036]= -1975871368;
assign addr[16037]= -1910985158;
assign addr[16038]= -1836405100;
assign addr[16039]= -1752509516;
assign addr[16040]= -1659723983;
assign addr[16041]= -1558519173;
assign addr[16042]= -1449408469;
assign addr[16043]= -1332945355;
assign addr[16044]= -1209720613;
assign addr[16045]= -1080359326;
assign addr[16046]= -945517704;
assign addr[16047]= -805879757;
assign addr[16048]= -662153826;
assign addr[16049]= -515068990;
assign addr[16050]= -365371365;
assign addr[16051]= -213820322;
assign addr[16052]= -61184634;
assign addr[16053]= 91761426;
assign addr[16054]= 244242007;
assign addr[16055]= 395483624;
assign addr[16056]= 544719071;
assign addr[16057]= 691191324;
assign addr[16058]= 834157373;
assign addr[16059]= 972891995;
assign addr[16060]= 1106691431;
assign addr[16061]= 1234876957;
assign addr[16062]= 1356798326;
assign addr[16063]= 1471837070;
assign addr[16064]= 1579409630;
assign addr[16065]= 1678970324;
assign addr[16066]= 1770014111;
assign addr[16067]= 1852079154;
assign addr[16068]= 1924749160;
assign addr[16069]= 1987655498;
assign addr[16070]= 2040479063;
assign addr[16071]= 2082951896;
assign addr[16072]= 2114858546;
assign addr[16073]= 2136037160;
assign addr[16074]= 2146380306;
assign addr[16075]= 2145835515;
assign addr[16076]= 2134405552;
assign addr[16077]= 2112148396;
assign addr[16078]= 2079176953;
assign addr[16079]= 2035658475;
assign addr[16080]= 1981813720;
assign addr[16081]= 1917915825;
assign addr[16082]= 1844288924;
assign addr[16083]= 1761306505;
assign addr[16084]= 1669389513;
assign addr[16085]= 1569004214;
assign addr[16086]= 1460659832;
assign addr[16087]= 1344905966;
assign addr[16088]= 1222329801;
assign addr[16089]= 1093553126;
assign addr[16090]= 959229189;
assign addr[16091]= 820039373;
assign addr[16092]= 676689746;
assign addr[16093]= 529907477;
assign addr[16094]= 380437148;
assign addr[16095]= 229036977;
assign addr[16096]= 76474970;
assign addr[16097]= -76474970;
assign addr[16098]= -229036977;
assign addr[16099]= -380437148;
assign addr[16100]= -529907477;
assign addr[16101]= -676689746;
assign addr[16102]= -820039373;
assign addr[16103]= -959229189;
assign addr[16104]= -1093553126;
assign addr[16105]= -1222329801;
assign addr[16106]= -1344905966;
assign addr[16107]= -1460659832;
assign addr[16108]= -1569004214;
assign addr[16109]= -1669389513;
assign addr[16110]= -1761306505;
assign addr[16111]= -1844288924;
assign addr[16112]= -1917915825;
assign addr[16113]= -1981813720;
assign addr[16114]= -2035658475;
assign addr[16115]= -2079176953;
assign addr[16116]= -2112148396;
assign addr[16117]= -2134405552;
assign addr[16118]= -2145835515;
assign addr[16119]= -2146380306;
assign addr[16120]= -2136037160;
assign addr[16121]= -2114858546;
assign addr[16122]= -2082951896;
assign addr[16123]= -2040479063;
assign addr[16124]= -1987655498;
assign addr[16125]= -1924749160;
assign addr[16126]= -1852079154;
assign addr[16127]= -1770014111;
assign addr[16128]= -1678970324;
assign addr[16129]= -1579409630;
assign addr[16130]= -1471837070;
assign addr[16131]= -1356798326;
assign addr[16132]= -1234876957;
assign addr[16133]= -1106691431;
assign addr[16134]= -972891995;
assign addr[16135]= -834157373;
assign addr[16136]= -691191324;
assign addr[16137]= -544719071;
assign addr[16138]= -395483624;
assign addr[16139]= -244242007;
assign addr[16140]= -91761426;
assign addr[16141]= 61184634;
assign addr[16142]= 213820322;
assign addr[16143]= 365371365;
assign addr[16144]= 515068990;
assign addr[16145]= 662153826;
assign addr[16146]= 805879757;
assign addr[16147]= 945517704;
assign addr[16148]= 1080359326;
assign addr[16149]= 1209720613;
assign addr[16150]= 1332945355;
assign addr[16151]= 1449408469;
assign addr[16152]= 1558519173;
assign addr[16153]= 1659723983;
assign addr[16154]= 1752509516;
assign addr[16155]= 1836405100;
assign addr[16156]= 1910985158;
assign addr[16157]= 1975871368;
assign addr[16158]= 2030734582;
assign addr[16159]= 2075296495;
assign addr[16160]= 2109331059;
assign addr[16161]= 2132665626;
assign addr[16162]= 2145181827;
assign addr[16163]= 2146816171;
assign addr[16164]= 2137560369;
assign addr[16165]= 2117461370;
assign addr[16166]= 2086621133;
assign addr[16167]= 2045196100;
assign addr[16168]= 1993396407;
assign addr[16169]= 1931484818;
assign addr[16170]= 1859775393;
assign addr[16171]= 1778631892;
assign addr[16172]= 1688465931;
assign addr[16173]= 1589734894;
assign addr[16174]= 1482939614;
assign addr[16175]= 1368621831;
assign addr[16176]= 1247361445;
assign addr[16177]= 1119773573;
assign addr[16178]= 986505429;
assign addr[16179]= 848233042;
assign addr[16180]= 705657826;
assign addr[16181]= 559503022;
assign addr[16182]= 410510029;
assign addr[16183]= 259434643;
assign addr[16184]= 107043224;
assign addr[16185]= -45891193;
assign addr[16186]= -198592817;
assign addr[16187]= -350287041;
assign addr[16188]= -500204365;
assign addr[16189]= -647584304;
assign addr[16190]= -791679244;
assign addr[16191]= -931758235;
assign addr[16192]= -1067110699;
assign addr[16193]= -1197050035;
assign addr[16194]= -1320917099;
assign addr[16195]= -1438083551;
assign addr[16196]= -1547955041;
assign addr[16197]= -1649974225;
assign addr[16198]= -1743623590;
assign addr[16199]= -1828428082;
assign addr[16200]= -1903957513;
assign addr[16201]= -1969828744;
assign addr[16202]= -2025707632;
assign addr[16203]= -2071310720;
assign addr[16204]= -2106406677;
assign addr[16205]= -2130817471;
assign addr[16206]= -2144419275;
assign addr[16207]= -2147143090;
assign addr[16208]= -2138975100;
assign addr[16209]= -2119956737;
assign addr[16210]= -2090184478;
assign addr[16211]= -2049809346;
assign addr[16212]= -1999036154;
assign addr[16213]= -1938122457;
assign addr[16214]= -1867377253;
assign addr[16215]= -1787159411;
assign addr[16216]= -1697875851;
assign addr[16217]= -1599979481;
assign addr[16218]= -1493966902;
assign addr[16219]= -1380375881;
assign addr[16220]= -1259782632;
assign addr[16221]= -1132798888;
assign addr[16222]= -1000068799;
assign addr[16223]= -862265664;
assign addr[16224]= -720088517;
assign addr[16225]= -574258580;
assign addr[16226]= -425515602;
assign addr[16227]= -274614114;
assign addr[16228]= -122319591;
assign addr[16229]= 30595422;
assign addr[16230]= 183355234;
assign addr[16231]= 335184940;
assign addr[16232]= 485314355;
assign addr[16233]= 632981917;
assign addr[16234]= 777438554;
assign addr[16235]= 917951481;
assign addr[16236]= 1053807919;
assign addr[16237]= 1184318708;
assign addr[16238]= 1308821808;
assign addr[16239]= 1426685652;
assign addr[16240]= 1537312353;
assign addr[16241]= 1640140734;
assign addr[16242]= 1734649179;
assign addr[16243]= 1820358275;
assign addr[16244]= 1896833245;
assign addr[16245]= 1963686155;
assign addr[16246]= 2020577882;
assign addr[16247]= 2067219829;
assign addr[16248]= 2103375398;
assign addr[16249]= 2128861181;
assign addr[16250]= 2143547897;
assign addr[16251]= 2147361045;
assign addr[16252]= 2140281282;
assign addr[16253]= 2122344521;
assign addr[16254]= 2093641749;
assign addr[16255]= 2054318569;
assign addr[16256]= 2004574453;
assign addr[16257]= 1944661739;
assign addr[16258]= 1874884346;
assign addr[16259]= 1795596234;
assign addr[16260]= 1707199606;
assign addr[16261]= 1610142873;
assign addr[16262]= 1504918373;
assign addr[16263]= 1392059879;
assign addr[16264]= 1272139887;
assign addr[16265]= 1145766716;
assign addr[16266]= 1013581418;
assign addr[16267]= 876254528;
assign addr[16268]= 734482665;
assign addr[16269]= 588984994;
assign addr[16270]= 440499581;
assign addr[16271]= 289779648;
assign addr[16272]= 137589750;
assign addr[16273]= -15298099;
assign addr[16274]= -168108346;
assign addr[16275]= -320065829;
assign addr[16276]= -470399716;
assign addr[16277]= -618347408;
assign addr[16278]= -763158411;
assign addr[16279]= -904098143;
assign addr[16280]= -1040451659;
assign addr[16281]= -1171527280;
assign addr[16282]= -1296660098;
assign addr[16283]= -1415215352;
assign addr[16284]= -1526591649;
assign addr[16285]= -1630224009;
assign addr[16286]= -1725586737;
assign addr[16287]= -1812196087;
assign addr[16288]= -1889612716;
assign addr[16289]= -1957443913;
assign addr[16290]= -2015345591;
assign addr[16291]= -2063024031;
assign addr[16292]= -2100237377;
assign addr[16293]= -2126796855;
assign addr[16294]= -2142567738;
assign addr[16295]= -2147470025;
assign addr[16296]= -2141478848;
assign addr[16297]= -2124624598;
assign addr[16298]= -2096992772;
assign addr[16299]= -2058723538;
assign addr[16300]= -2010011024;
assign addr[16301]= -1951102334;
assign addr[16302]= -1882296293;
assign addr[16303]= -1803941934;
assign addr[16304]= -1716436725;
assign addr[16305]= -1620224553;
assign addr[16306]= -1515793473;
assign addr[16307]= -1403673233;
assign addr[16308]= -1284432584;
assign addr[16309]= -1158676398;
assign addr[16310]= -1027042599;
assign addr[16311]= -890198924;
assign addr[16312]= -748839539;
assign addr[16313]= -603681519;
assign addr[16314]= -455461206;
assign addr[16315]= -304930476;
assign addr[16316]= -152852926;
assign addr[16317]= 0;
assign addr[16318]= 152852926;
assign addr[16319]= 304930476;
assign addr[16320]= 455461206;
assign addr[16321]= 603681519;
assign addr[16322]= 748839539;
assign addr[16323]= 890198924;
assign addr[16324]= 1027042599;
assign addr[16325]= 1158676398;
assign addr[16326]= 1284432584;
assign addr[16327]= 1403673233;
assign addr[16328]= 1515793473;
assign addr[16329]= 1620224553;
assign addr[16330]= 1716436725;
assign addr[16331]= 1803941934;
assign addr[16332]= 1882296293;
assign addr[16333]= 1951102334;
assign addr[16334]= 2010011024;
assign addr[16335]= 2058723538;
assign addr[16336]= 2096992772;
assign addr[16337]= 2124624598;
assign addr[16338]= 2141478848;
assign addr[16339]= 2147470025;
assign addr[16340]= 2142567738;
assign addr[16341]= 2126796855;
assign addr[16342]= 2100237377;
assign addr[16343]= 2063024031;
assign addr[16344]= 2015345591;
assign addr[16345]= 1957443913;
assign addr[16346]= 1889612716;
assign addr[16347]= 1812196087;
assign addr[16348]= 1725586737;
assign addr[16349]= 1630224009;
assign addr[16350]= 1526591649;
assign addr[16351]= 1415215352;
assign addr[16352]= 1296660098;
assign addr[16353]= 1171527280;
assign addr[16354]= 1040451659;
assign addr[16355]= 904098143;
assign addr[16356]= 763158411;
assign addr[16357]= 618347408;
assign addr[16358]= 470399716;
assign addr[16359]= 320065829;
assign addr[16360]= 168108346;
assign addr[16361]= 15298099;
assign addr[16362]= -137589750;
assign addr[16363]= -289779648;
assign addr[16364]= -440499581;
assign addr[16365]= -588984994;
assign addr[16366]= -734482665;
assign addr[16367]= -876254528;
assign addr[16368]= -1013581418;
assign addr[16369]= -1145766716;
assign addr[16370]= -1272139887;
assign addr[16371]= -1392059879;
assign addr[16372]= -1504918373;
assign addr[16373]= -1610142873;
assign addr[16374]= -1707199606;
assign addr[16375]= -1795596234;
assign addr[16376]= -1874884346;
assign addr[16377]= -1944661739;
assign addr[16378]= -2004574453;
assign addr[16379]= -2054318569;
assign addr[16380]= -2093641749;
assign addr[16381]= -2122344521;
assign addr[16382]= -2140281282;
assign addr[16383]= -2147361045;
assign addr[16384]= -2143547897;
assign addr[16385]= -2128861181;
assign addr[16386]= -2103375398;
assign addr[16387]= -2067219829;
assign addr[16388]= -2020577882;
assign addr[16389]= -1963686155;
assign addr[16390]= -1896833245;
assign addr[16391]= -1820358275;
assign addr[16392]= -1734649179;
assign addr[16393]= -1640140734;
assign addr[16394]= -1537312353;
assign addr[16395]= -1426685652;
assign addr[16396]= -1308821808;
assign addr[16397]= -1184318708;
assign addr[16398]= -1053807919;
assign addr[16399]= -917951481;
assign addr[16400]= -777438554;
assign addr[16401]= -632981917;
assign addr[16402]= -485314355;
assign addr[16403]= -335184940;
assign addr[16404]= -183355234;
assign addr[16405]= -30595422;
assign addr[16406]= 122319591;
assign addr[16407]= 274614114;
assign addr[16408]= 425515602;
assign addr[16409]= 574258580;
assign addr[16410]= 720088517;
assign addr[16411]= 862265664;
assign addr[16412]= 1000068799;
assign addr[16413]= 1132798888;
assign addr[16414]= 1259782632;
assign addr[16415]= 1380375881;
assign addr[16416]= 1493966902;
assign addr[16417]= 1599979481;
assign addr[16418]= 1697875851;
assign addr[16419]= 1787159411;
assign addr[16420]= 1867377253;
assign addr[16421]= 1938122457;
assign addr[16422]= 1999036154;
assign addr[16423]= 2049809346;
assign addr[16424]= 2090184478;
assign addr[16425]= 2119956737;
assign addr[16426]= 2138975100;
assign addr[16427]= 2147143090;
assign addr[16428]= 2144419275;
assign addr[16429]= 2130817471;
assign addr[16430]= 2106406677;
assign addr[16431]= 2071310720;
assign addr[16432]= 2025707632;
assign addr[16433]= 1969828744;
assign addr[16434]= 1903957513;
assign addr[16435]= 1828428082;
assign addr[16436]= 1743623590;
assign addr[16437]= 1649974225;
assign addr[16438]= 1547955041;
assign addr[16439]= 1438083551;
assign addr[16440]= 1320917099;
assign addr[16441]= 1197050035;
assign addr[16442]= 1067110699;
assign addr[16443]= 931758235;
assign addr[16444]= 791679244;
assign addr[16445]= 647584304;
assign addr[16446]= 500204365;
assign addr[16447]= 350287041;
assign addr[16448]= 198592817;
assign addr[16449]= 45891193;
assign addr[16450]= -107043224;
assign addr[16451]= -259434643;
assign addr[16452]= -410510029;
assign addr[16453]= -559503022;
assign addr[16454]= -705657826;
assign addr[16455]= -848233042;
assign addr[16456]= -986505429;
assign addr[16457]= -1119773573;
assign addr[16458]= -1247361445;
assign addr[16459]= -1368621831;
assign addr[16460]= -1482939614;
assign addr[16461]= -1589734894;
assign addr[16462]= -1688465931;
assign addr[16463]= -1778631892;
assign addr[16464]= -1859775393;
assign addr[16465]= -1931484818;
assign addr[16466]= -1993396407;
assign addr[16467]= -2045196100;
assign addr[16468]= -2086621133;
assign addr[16469]= -2117461370;
assign addr[16470]= -2137560369;
assign addr[16471]= -2146816171;
assign addr[16472]= -2145181827;
assign addr[16473]= -2132665626;
assign addr[16474]= -2109331059;
assign addr[16475]= -2075296495;
assign addr[16476]= -2030734582;
assign addr[16477]= -1975871368;
assign addr[16478]= -1910985158;
assign addr[16479]= -1836405100;
assign addr[16480]= -1752509516;
assign addr[16481]= -1659723983;
assign addr[16482]= -1558519173;
assign addr[16483]= -1449408469;
assign addr[16484]= -1332945355;
assign addr[16485]= -1209720613;
assign addr[16486]= -1080359326;
assign addr[16487]= -945517704;
assign addr[16488]= -805879757;
assign addr[16489]= -662153826;
assign addr[16490]= -515068990;
assign addr[16491]= -365371365;
assign addr[16492]= -213820322;
assign addr[16493]= -61184634;
assign addr[16494]= 91761426;
assign addr[16495]= 244242007;
assign addr[16496]= 395483624;
assign addr[16497]= 544719071;
assign addr[16498]= 691191324;
assign addr[16499]= 834157373;
assign addr[16500]= 972891995;
assign addr[16501]= 1106691431;
assign addr[16502]= 1234876957;
assign addr[16503]= 1356798326;
assign addr[16504]= 1471837070;
assign addr[16505]= 1579409630;
assign addr[16506]= 1678970324;
assign addr[16507]= 1770014111;
assign addr[16508]= 1852079154;
assign addr[16509]= 1924749160;
assign addr[16510]= 1987655498;
assign addr[16511]= 2040479063;
assign addr[16512]= 2082951896;
assign addr[16513]= 2114858546;
assign addr[16514]= 2136037160;
assign addr[16515]= 2146380306;
assign addr[16516]= 2145835515;
assign addr[16517]= 2134405552;
assign addr[16518]= 2112148396;
assign addr[16519]= 2079176953;
assign addr[16520]= 2035658475;
assign addr[16521]= 1981813720;
assign addr[16522]= 1917915825;
assign addr[16523]= 1844288924;
assign addr[16524]= 1761306505;
assign addr[16525]= 1669389513;
assign addr[16526]= 1569004214;
assign addr[16527]= 1460659832;
assign addr[16528]= 1344905966;
assign addr[16529]= 1222329801;
assign addr[16530]= 1093553126;
assign addr[16531]= 959229189;
assign addr[16532]= 820039373;
assign addr[16533]= 676689746;
assign addr[16534]= 529907477;
assign addr[16535]= 380437148;
assign addr[16536]= 229036977;
assign addr[16537]= 76474970;
assign addr[16538]= -76474970;
assign addr[16539]= -229036977;
assign addr[16540]= -380437148;
assign addr[16541]= -529907477;
assign addr[16542]= -676689746;
assign addr[16543]= -820039373;
assign addr[16544]= -959229189;
assign addr[16545]= -1093553126;
assign addr[16546]= -1222329801;
assign addr[16547]= -1344905966;
assign addr[16548]= -1460659832;
assign addr[16549]= -1569004214;
assign addr[16550]= -1669389513;
assign addr[16551]= -1761306505;
assign addr[16552]= -1844288924;
assign addr[16553]= -1917915825;
assign addr[16554]= -1981813720;
assign addr[16555]= -2035658475;
assign addr[16556]= -2079176953;
assign addr[16557]= -2112148396;
assign addr[16558]= -2134405552;
assign addr[16559]= -2145835515;
assign addr[16560]= -2146380306;
assign addr[16561]= -2136037160;
assign addr[16562]= -2114858546;
assign addr[16563]= -2082951896;
assign addr[16564]= -2040479063;
assign addr[16565]= -1987655498;
assign addr[16566]= -1924749160;
assign addr[16567]= -1852079154;
assign addr[16568]= -1770014111;
assign addr[16569]= -1678970324;
assign addr[16570]= -1579409630;
assign addr[16571]= -1471837070;
assign addr[16572]= -1356798326;
assign addr[16573]= -1234876957;
assign addr[16574]= -1106691431;
assign addr[16575]= -972891995;
assign addr[16576]= -834157373;
assign addr[16577]= -691191324;
assign addr[16578]= -544719071;
assign addr[16579]= -395483624;
assign addr[16580]= -244242007;
assign addr[16581]= -91761426;
assign addr[16582]= 61184634;
assign addr[16583]= 213820322;
assign addr[16584]= 365371365;
assign addr[16585]= 515068990;
assign addr[16586]= 662153826;
assign addr[16587]= 805879757;
assign addr[16588]= 945517704;
assign addr[16589]= 1080359326;
assign addr[16590]= 1209720613;
assign addr[16591]= 1332945355;
assign addr[16592]= 1449408469;
assign addr[16593]= 1558519173;
assign addr[16594]= 1659723983;
assign addr[16595]= 1752509516;
assign addr[16596]= 1836405100;
assign addr[16597]= 1910985158;
assign addr[16598]= 1975871368;
assign addr[16599]= 2030734582;
assign addr[16600]= 2075296495;
assign addr[16601]= 2109331059;
assign addr[16602]= 2132665626;
assign addr[16603]= 2145181827;
assign addr[16604]= 2146816171;
assign addr[16605]= 2137560369;
assign addr[16606]= 2117461370;
assign addr[16607]= 2086621133;
assign addr[16608]= 2045196100;
assign addr[16609]= 1993396407;
assign addr[16610]= 1931484818;
assign addr[16611]= 1859775393;
assign addr[16612]= 1778631892;
assign addr[16613]= 1688465931;
assign addr[16614]= 1589734894;
assign addr[16615]= 1482939614;
assign addr[16616]= 1368621831;
assign addr[16617]= 1247361445;
assign addr[16618]= 1119773573;
assign addr[16619]= 986505429;
assign addr[16620]= 848233042;
assign addr[16621]= 705657826;
assign addr[16622]= 559503022;
assign addr[16623]= 410510029;
assign addr[16624]= 259434643;
assign addr[16625]= 107043224;
assign addr[16626]= -45891193;
assign addr[16627]= -198592817;
assign addr[16628]= -350287041;
assign addr[16629]= -500204365;
assign addr[16630]= -647584304;
assign addr[16631]= -791679244;
assign addr[16632]= -931758235;
assign addr[16633]= -1067110699;
assign addr[16634]= -1197050035;
assign addr[16635]= -1320917099;
assign addr[16636]= -1438083551;
assign addr[16637]= -1547955041;
assign addr[16638]= -1649974225;
assign addr[16639]= -1743623590;
assign addr[16640]= -1828428082;
assign addr[16641]= -1903957513;
assign addr[16642]= -1969828744;
assign addr[16643]= -2025707632;
assign addr[16644]= -2071310720;
assign addr[16645]= -2106406677;
assign addr[16646]= -2130817471;
assign addr[16647]= -2144419275;
assign addr[16648]= -2147143090;
assign addr[16649]= -2138975100;
assign addr[16650]= -2119956737;
assign addr[16651]= -2090184478;
assign addr[16652]= -2049809346;
assign addr[16653]= -1999036154;
assign addr[16654]= -1938122457;
assign addr[16655]= -1867377253;
assign addr[16656]= -1787159411;
assign addr[16657]= -1697875851;
assign addr[16658]= -1599979481;
assign addr[16659]= -1493966902;
assign addr[16660]= -1380375881;
assign addr[16661]= -1259782632;
assign addr[16662]= -1132798888;
assign addr[16663]= -1000068799;
assign addr[16664]= -862265664;
assign addr[16665]= -720088517;
assign addr[16666]= -574258580;
assign addr[16667]= -425515602;
assign addr[16668]= -274614114;
assign addr[16669]= -122319591;
assign addr[16670]= 30595422;
assign addr[16671]= 183355234;
assign addr[16672]= 335184940;
assign addr[16673]= 485314355;
assign addr[16674]= 632981917;
assign addr[16675]= 777438554;
assign addr[16676]= 917951481;
assign addr[16677]= 1053807919;
assign addr[16678]= 1184318708;
assign addr[16679]= 1308821808;
assign addr[16680]= 1426685652;
assign addr[16681]= 1537312353;
assign addr[16682]= 1640140734;
assign addr[16683]= 1734649179;
assign addr[16684]= 1820358275;
assign addr[16685]= 1896833245;
assign addr[16686]= 1963686155;
assign addr[16687]= 2020577882;
assign addr[16688]= 2067219829;
assign addr[16689]= 2103375398;
assign addr[16690]= 2128861181;
assign addr[16691]= 2143547897;
assign addr[16692]= 2147361045;
assign addr[16693]= 2140281282;
assign addr[16694]= 2122344521;
assign addr[16695]= 2093641749;
assign addr[16696]= 2054318569;
assign addr[16697]= 2004574453;
assign addr[16698]= 1944661739;
assign addr[16699]= 1874884346;
assign addr[16700]= 1795596234;
assign addr[16701]= 1707199606;
assign addr[16702]= 1610142873;
assign addr[16703]= 1504918373;
assign addr[16704]= 1392059879;
assign addr[16705]= 1272139887;
assign addr[16706]= 1145766716;
assign addr[16707]= 1013581418;
assign addr[16708]= 876254528;
assign addr[16709]= 734482665;
assign addr[16710]= 588984994;
assign addr[16711]= 440499581;
assign addr[16712]= 289779648;
assign addr[16713]= 137589750;
assign addr[16714]= -15298099;
assign addr[16715]= -168108346;
assign addr[16716]= -320065829;
assign addr[16717]= -470399716;
assign addr[16718]= -618347408;
assign addr[16719]= -763158411;
assign addr[16720]= -904098143;
assign addr[16721]= -1040451659;
assign addr[16722]= -1171527280;
assign addr[16723]= -1296660098;
assign addr[16724]= -1415215352;
assign addr[16725]= -1526591649;
assign addr[16726]= -1630224009;
assign addr[16727]= -1725586737;
assign addr[16728]= -1812196087;
assign addr[16729]= -1889612716;
assign addr[16730]= -1957443913;
assign addr[16731]= -2015345591;
assign addr[16732]= -2063024031;
assign addr[16733]= -2100237377;
assign addr[16734]= -2126796855;
assign addr[16735]= -2142567738;
assign addr[16736]= -2147470025;
assign addr[16737]= -2141478848;
assign addr[16738]= -2124624598;
assign addr[16739]= -2096992772;
assign addr[16740]= -2058723538;
assign addr[16741]= -2010011024;
assign addr[16742]= -1951102334;
assign addr[16743]= -1882296293;
assign addr[16744]= -1803941934;
assign addr[16745]= -1716436725;
assign addr[16746]= -1620224553;
assign addr[16747]= -1515793473;
assign addr[16748]= -1403673233;
assign addr[16749]= -1284432584;
assign addr[16750]= -1158676398;
assign addr[16751]= -1027042599;
assign addr[16752]= -890198924;
assign addr[16753]= -748839539;
assign addr[16754]= -603681519;
assign addr[16755]= -455461206;
assign addr[16756]= -304930476;
assign addr[16757]= -152852926;
assign addr[16758]= 0;
assign addr[16759]= 152852926;
assign addr[16760]= 304930476;
assign addr[16761]= 455461206;
assign addr[16762]= 603681519;
assign addr[16763]= 748839539;
assign addr[16764]= 890198924;
assign addr[16765]= 1027042599;
assign addr[16766]= 1158676398;
assign addr[16767]= 1284432584;
assign addr[16768]= 1403673233;
assign addr[16769]= 1515793473;
assign addr[16770]= 1620224553;
assign addr[16771]= 1716436725;
assign addr[16772]= 1803941934;
assign addr[16773]= 1882296293;
assign addr[16774]= 1951102334;
assign addr[16775]= 2010011024;
assign addr[16776]= 2058723538;
assign addr[16777]= 2096992772;
assign addr[16778]= 2124624598;
assign addr[16779]= 2141478848;
assign addr[16780]= 2147470025;
assign addr[16781]= 2142567738;
assign addr[16782]= 2126796855;
assign addr[16783]= 2100237377;
assign addr[16784]= 2063024031;
assign addr[16785]= 2015345591;
assign addr[16786]= 1957443913;
assign addr[16787]= 1889612716;
assign addr[16788]= 1812196087;
assign addr[16789]= 1725586737;
assign addr[16790]= 1630224009;
assign addr[16791]= 1526591649;
assign addr[16792]= 1415215352;
assign addr[16793]= 1296660098;
assign addr[16794]= 1171527280;
assign addr[16795]= 1040451659;
assign addr[16796]= 904098143;
assign addr[16797]= 763158411;
assign addr[16798]= 618347408;
assign addr[16799]= 470399716;
assign addr[16800]= 320065829;
assign addr[16801]= 168108346;
assign addr[16802]= 15298099;
assign addr[16803]= -137589750;
assign addr[16804]= -289779648;
assign addr[16805]= -440499581;
assign addr[16806]= -588984994;
assign addr[16807]= -734482665;
assign addr[16808]= -876254528;
assign addr[16809]= -1013581418;
assign addr[16810]= -1145766716;
assign addr[16811]= -1272139887;
assign addr[16812]= -1392059879;
assign addr[16813]= -1504918373;
assign addr[16814]= -1610142873;
assign addr[16815]= -1707199606;
assign addr[16816]= -1795596234;
assign addr[16817]= -1874884346;
assign addr[16818]= -1944661739;
assign addr[16819]= -2004574453;
assign addr[16820]= -2054318569;
assign addr[16821]= -2093641749;
assign addr[16822]= -2122344521;
assign addr[16823]= -2140281282;
assign addr[16824]= -2147361045;
assign addr[16825]= -2143547897;
assign addr[16826]= -2128861181;
assign addr[16827]= -2103375398;
assign addr[16828]= -2067219829;
assign addr[16829]= -2020577882;
assign addr[16830]= -1963686155;
assign addr[16831]= -1896833245;
assign addr[16832]= -1820358275;
assign addr[16833]= -1734649179;
assign addr[16834]= -1640140734;
assign addr[16835]= -1537312353;
assign addr[16836]= -1426685652;
assign addr[16837]= -1308821808;
assign addr[16838]= -1184318708;
assign addr[16839]= -1053807919;
assign addr[16840]= -917951481;
assign addr[16841]= -777438554;
assign addr[16842]= -632981917;
assign addr[16843]= -485314355;
assign addr[16844]= -335184940;
assign addr[16845]= -183355234;
assign addr[16846]= -30595422;
assign addr[16847]= 122319591;
assign addr[16848]= 274614114;
assign addr[16849]= 425515602;
assign addr[16850]= 574258580;
assign addr[16851]= 720088517;
assign addr[16852]= 862265664;
assign addr[16853]= 1000068799;
assign addr[16854]= 1132798888;
assign addr[16855]= 1259782632;
assign addr[16856]= 1380375881;
assign addr[16857]= 1493966902;
assign addr[16858]= 1599979481;
assign addr[16859]= 1697875851;
assign addr[16860]= 1787159411;
assign addr[16861]= 1867377253;
assign addr[16862]= 1938122457;
assign addr[16863]= 1999036154;
assign addr[16864]= 2049809346;
assign addr[16865]= 2090184478;
assign addr[16866]= 2119956737;
assign addr[16867]= 2138975100;
assign addr[16868]= 2147143090;
assign addr[16869]= 2144419275;
assign addr[16870]= 2130817471;
assign addr[16871]= 2106406677;
assign addr[16872]= 2071310720;
assign addr[16873]= 2025707632;
assign addr[16874]= 1969828744;
assign addr[16875]= 1903957513;
assign addr[16876]= 1828428082;
assign addr[16877]= 1743623590;
assign addr[16878]= 1649974225;
assign addr[16879]= 1547955041;
assign addr[16880]= 1438083551;
assign addr[16881]= 1320917099;
assign addr[16882]= 1197050035;
assign addr[16883]= 1067110699;
assign addr[16884]= 931758235;
assign addr[16885]= 791679244;
assign addr[16886]= 647584304;
assign addr[16887]= 500204365;
assign addr[16888]= 350287041;
assign addr[16889]= 198592817;
assign addr[16890]= 45891193;
assign addr[16891]= -107043224;
assign addr[16892]= -259434643;
assign addr[16893]= -410510029;
assign addr[16894]= -559503022;
assign addr[16895]= -705657826;
assign addr[16896]= -848233042;
assign addr[16897]= -986505429;
assign addr[16898]= -1119773573;
assign addr[16899]= -1247361445;
assign addr[16900]= -1368621831;
assign addr[16901]= -1482939614;
assign addr[16902]= -1589734894;
assign addr[16903]= -1688465931;
assign addr[16904]= -1778631892;
assign addr[16905]= -1859775393;
assign addr[16906]= -1931484818;
assign addr[16907]= -1993396407;
assign addr[16908]= -2045196100;
assign addr[16909]= -2086621133;
assign addr[16910]= -2117461370;
assign addr[16911]= -2137560369;
assign addr[16912]= -2146816171;
assign addr[16913]= -2145181827;
assign addr[16914]= -2132665626;
assign addr[16915]= -2109331059;
assign addr[16916]= -2075296495;
assign addr[16917]= -2030734582;
assign addr[16918]= -1975871368;
assign addr[16919]= -1910985158;
assign addr[16920]= -1836405100;
assign addr[16921]= -1752509516;
assign addr[16922]= -1659723983;
assign addr[16923]= -1558519173;
assign addr[16924]= -1449408469;
assign addr[16925]= -1332945355;
assign addr[16926]= -1209720613;
assign addr[16927]= -1080359326;
assign addr[16928]= -945517704;
assign addr[16929]= -805879757;
assign addr[16930]= -662153826;
assign addr[16931]= -515068990;
assign addr[16932]= -365371365;
assign addr[16933]= -213820322;
assign addr[16934]= -61184634;
assign addr[16935]= 91761426;
assign addr[16936]= 244242007;
assign addr[16937]= 395483624;
assign addr[16938]= 544719071;
assign addr[16939]= 691191324;
assign addr[16940]= 834157373;
assign addr[16941]= 972891995;
assign addr[16942]= 1106691431;
assign addr[16943]= 1234876957;
assign addr[16944]= 1356798326;
assign addr[16945]= 1471837070;
assign addr[16946]= 1579409630;
assign addr[16947]= 1678970324;
assign addr[16948]= 1770014111;
assign addr[16949]= 1852079154;
assign addr[16950]= 1924749160;
assign addr[16951]= 1987655498;
assign addr[16952]= 2040479063;
assign addr[16953]= 2082951896;
assign addr[16954]= 2114858546;
assign addr[16955]= 2136037160;
assign addr[16956]= 2146380306;
assign addr[16957]= 2145835515;
assign addr[16958]= 2134405552;
assign addr[16959]= 2112148396;
assign addr[16960]= 2079176953;
assign addr[16961]= 2035658475;
assign addr[16962]= 1981813720;
assign addr[16963]= 1917915825;
assign addr[16964]= 1844288924;
assign addr[16965]= 1761306505;
assign addr[16966]= 1669389513;
assign addr[16967]= 1569004214;
assign addr[16968]= 1460659832;
assign addr[16969]= 1344905966;
assign addr[16970]= 1222329801;
assign addr[16971]= 1093553126;
assign addr[16972]= 959229189;
assign addr[16973]= 820039373;
assign addr[16974]= 676689746;
assign addr[16975]= 529907477;
assign addr[16976]= 380437148;
assign addr[16977]= 229036977;
assign addr[16978]= 76474970;
assign addr[16979]= -76474970;
assign addr[16980]= -229036977;
assign addr[16981]= -380437148;
assign addr[16982]= -529907477;
assign addr[16983]= -676689746;
assign addr[16984]= -820039373;
assign addr[16985]= -959229189;
assign addr[16986]= -1093553126;
assign addr[16987]= -1222329801;
assign addr[16988]= -1344905966;
assign addr[16989]= -1460659832;
assign addr[16990]= -1569004214;
assign addr[16991]= -1669389513;
assign addr[16992]= -1761306505;
assign addr[16993]= -1844288924;
assign addr[16994]= -1917915825;
assign addr[16995]= -1981813720;
assign addr[16996]= -2035658475;
assign addr[16997]= -2079176953;
assign addr[16998]= -2112148396;
assign addr[16999]= -2134405552;
assign addr[17000]= -2145835515;
assign addr[17001]= -2146380306;
assign addr[17002]= -2136037160;
assign addr[17003]= -2114858546;
assign addr[17004]= -2082951896;
assign addr[17005]= -2040479063;
assign addr[17006]= -1987655498;
assign addr[17007]= -1924749160;
assign addr[17008]= -1852079154;
assign addr[17009]= -1770014111;
assign addr[17010]= -1678970324;
assign addr[17011]= -1579409630;
assign addr[17012]= -1471837070;
assign addr[17013]= -1356798326;
assign addr[17014]= -1234876957;
assign addr[17015]= -1106691431;
assign addr[17016]= -972891995;
assign addr[17017]= -834157373;
assign addr[17018]= -691191324;
assign addr[17019]= -544719071;
assign addr[17020]= -395483624;
assign addr[17021]= -244242007;
assign addr[17022]= -91761426;
assign addr[17023]= 61184634;
assign addr[17024]= 213820322;
assign addr[17025]= 365371365;
assign addr[17026]= 515068990;
assign addr[17027]= 662153826;
assign addr[17028]= 805879757;
assign addr[17029]= 945517704;
assign addr[17030]= 1080359326;
assign addr[17031]= 1209720613;
assign addr[17032]= 1332945355;
assign addr[17033]= 1449408469;
assign addr[17034]= 1558519173;
assign addr[17035]= 1659723983;
assign addr[17036]= 1752509516;
assign addr[17037]= 1836405100;
assign addr[17038]= 1910985158;
assign addr[17039]= 1975871368;
assign addr[17040]= 2030734582;
assign addr[17041]= 2075296495;
assign addr[17042]= 2109331059;
assign addr[17043]= 2132665626;
assign addr[17044]= 2145181827;
assign addr[17045]= 2146816171;
assign addr[17046]= 2137560369;
assign addr[17047]= 2117461370;
assign addr[17048]= 2086621133;
assign addr[17049]= 2045196100;
assign addr[17050]= 1993396407;
assign addr[17051]= 1931484818;
assign addr[17052]= 1859775393;
assign addr[17053]= 1778631892;
assign addr[17054]= 1688465931;
assign addr[17055]= 1589734894;
assign addr[17056]= 1482939614;
assign addr[17057]= 1368621831;
assign addr[17058]= 1247361445;
assign addr[17059]= 1119773573;
assign addr[17060]= 986505429;
assign addr[17061]= 848233042;
assign addr[17062]= 705657826;
assign addr[17063]= 559503022;
assign addr[17064]= 410510029;
assign addr[17065]= 259434643;
assign addr[17066]= 107043224;
assign addr[17067]= -45891193;
assign addr[17068]= -198592817;
assign addr[17069]= -350287041;
assign addr[17070]= -500204365;
assign addr[17071]= -647584304;
assign addr[17072]= -791679244;
assign addr[17073]= -931758235;
assign addr[17074]= -1067110699;
assign addr[17075]= -1197050035;
assign addr[17076]= -1320917099;
assign addr[17077]= -1438083551;
assign addr[17078]= -1547955041;
assign addr[17079]= -1649974225;
assign addr[17080]= -1743623590;
assign addr[17081]= -1828428082;
assign addr[17082]= -1903957513;
assign addr[17083]= -1969828744;
assign addr[17084]= -2025707632;
assign addr[17085]= -2071310720;
assign addr[17086]= -2106406677;
assign addr[17087]= -2130817471;
assign addr[17088]= -2144419275;
assign addr[17089]= -2147143090;
assign addr[17090]= -2138975100;
assign addr[17091]= -2119956737;
assign addr[17092]= -2090184478;
assign addr[17093]= -2049809346;
assign addr[17094]= -1999036154;
assign addr[17095]= -1938122457;
assign addr[17096]= -1867377253;
assign addr[17097]= -1787159411;
assign addr[17098]= -1697875851;
assign addr[17099]= -1599979481;
assign addr[17100]= -1493966902;
assign addr[17101]= -1380375881;
assign addr[17102]= -1259782632;
assign addr[17103]= -1132798888;
assign addr[17104]= -1000068799;
assign addr[17105]= -862265664;
assign addr[17106]= -720088517;
assign addr[17107]= -574258580;
assign addr[17108]= -425515602;
assign addr[17109]= -274614114;
assign addr[17110]= -122319591;
assign addr[17111]= 30595422;
assign addr[17112]= 183355234;
assign addr[17113]= 335184940;
assign addr[17114]= 485314355;
assign addr[17115]= 632981917;
assign addr[17116]= 777438554;
assign addr[17117]= 917951481;
assign addr[17118]= 1053807919;
assign addr[17119]= 1184318708;
assign addr[17120]= 1308821808;
assign addr[17121]= 1426685652;
assign addr[17122]= 1537312353;
assign addr[17123]= 1640140734;
assign addr[17124]= 1734649179;
assign addr[17125]= 1820358275;
assign addr[17126]= 1896833245;
assign addr[17127]= 1963686155;
assign addr[17128]= 2020577882;
assign addr[17129]= 2067219829;
assign addr[17130]= 2103375398;
assign addr[17131]= 2128861181;
assign addr[17132]= 2143547897;
assign addr[17133]= 2147361045;
assign addr[17134]= 2140281282;
assign addr[17135]= 2122344521;
assign addr[17136]= 2093641749;
assign addr[17137]= 2054318569;
assign addr[17138]= 2004574453;
assign addr[17139]= 1944661739;
assign addr[17140]= 1874884346;
assign addr[17141]= 1795596234;
assign addr[17142]= 1707199606;
assign addr[17143]= 1610142873;
assign addr[17144]= 1504918373;
assign addr[17145]= 1392059879;
assign addr[17146]= 1272139887;
assign addr[17147]= 1145766716;
assign addr[17148]= 1013581418;
assign addr[17149]= 876254528;
assign addr[17150]= 734482665;
assign addr[17151]= 588984994;
assign addr[17152]= 440499581;
assign addr[17153]= 289779648;
assign addr[17154]= 137589750;
assign addr[17155]= -15298099;
assign addr[17156]= -168108346;
assign addr[17157]= -320065829;
assign addr[17158]= -470399716;
assign addr[17159]= -618347408;
assign addr[17160]= -763158411;
assign addr[17161]= -904098143;
assign addr[17162]= -1040451659;
assign addr[17163]= -1171527280;
assign addr[17164]= -1296660098;
assign addr[17165]= -1415215352;
assign addr[17166]= -1526591649;
assign addr[17167]= -1630224009;
assign addr[17168]= -1725586737;
assign addr[17169]= -1812196087;
assign addr[17170]= -1889612716;
assign addr[17171]= -1957443913;
assign addr[17172]= -2015345591;
assign addr[17173]= -2063024031;
assign addr[17174]= -2100237377;
assign addr[17175]= -2126796855;
assign addr[17176]= -2142567738;
assign addr[17177]= -2147470025;
assign addr[17178]= -2141478848;
assign addr[17179]= -2124624598;
assign addr[17180]= -2096992772;
assign addr[17181]= -2058723538;
assign addr[17182]= -2010011024;
assign addr[17183]= -1951102334;
assign addr[17184]= -1882296293;
assign addr[17185]= -1803941934;
assign addr[17186]= -1716436725;
assign addr[17187]= -1620224553;
assign addr[17188]= -1515793473;
assign addr[17189]= -1403673233;
assign addr[17190]= -1284432584;
assign addr[17191]= -1158676398;
assign addr[17192]= -1027042599;
assign addr[17193]= -890198924;
assign addr[17194]= -748839539;
assign addr[17195]= -603681519;
assign addr[17196]= -455461206;
assign addr[17197]= -304930476;
assign addr[17198]= -152852926;
assign addr[17199]= 0;
assign addr[17200]= 152852926;
assign addr[17201]= 304930476;
assign addr[17202]= 455461206;
assign addr[17203]= 603681519;
assign addr[17204]= 748839539;
assign addr[17205]= 890198924;
assign addr[17206]= 1027042599;
assign addr[17207]= 1158676398;
assign addr[17208]= 1284432584;
assign addr[17209]= 1403673233;
assign addr[17210]= 1515793473;
assign addr[17211]= 1620224553;
assign addr[17212]= 1716436725;
assign addr[17213]= 1803941934;
assign addr[17214]= 1882296293;
assign addr[17215]= 1951102334;
assign addr[17216]= 2010011024;
assign addr[17217]= 2058723538;
assign addr[17218]= 2096992772;
assign addr[17219]= 2124624598;
assign addr[17220]= 2141478848;
assign addr[17221]= 2147470025;
assign addr[17222]= 2142567738;
assign addr[17223]= 2126796855;
assign addr[17224]= 2100237377;
assign addr[17225]= 2063024031;
assign addr[17226]= 2015345591;
assign addr[17227]= 1957443913;
assign addr[17228]= 1889612716;
assign addr[17229]= 1812196087;
assign addr[17230]= 1725586737;
assign addr[17231]= 1630224009;
assign addr[17232]= 1526591649;
assign addr[17233]= 1415215352;
assign addr[17234]= 1296660098;
assign addr[17235]= 1171527280;
assign addr[17236]= 1040451659;
assign addr[17237]= 904098143;
assign addr[17238]= 763158411;
assign addr[17239]= 618347408;
assign addr[17240]= 470399716;
assign addr[17241]= 320065829;
assign addr[17242]= 168108346;
assign addr[17243]= 15298099;
assign addr[17244]= -137589750;
assign addr[17245]= -289779648;
assign addr[17246]= -440499581;
assign addr[17247]= -588984994;
assign addr[17248]= -734482665;
assign addr[17249]= -876254528;
assign addr[17250]= -1013581418;
assign addr[17251]= -1145766716;
assign addr[17252]= -1272139887;
assign addr[17253]= -1392059879;
assign addr[17254]= -1504918373;
assign addr[17255]= -1610142873;
assign addr[17256]= -1707199606;
assign addr[17257]= -1795596234;
assign addr[17258]= -1874884346;
assign addr[17259]= -1944661739;
assign addr[17260]= -2004574453;
assign addr[17261]= -2054318569;
assign addr[17262]= -2093641749;
assign addr[17263]= -2122344521;
assign addr[17264]= -2140281282;
assign addr[17265]= -2147361045;
assign addr[17266]= -2143547897;
assign addr[17267]= -2128861181;
assign addr[17268]= -2103375398;
assign addr[17269]= -2067219829;
assign addr[17270]= -2020577882;
assign addr[17271]= -1963686155;
assign addr[17272]= -1896833245;
assign addr[17273]= -1820358275;
assign addr[17274]= -1734649179;
assign addr[17275]= -1640140734;
assign addr[17276]= -1537312353;
assign addr[17277]= -1426685652;
assign addr[17278]= -1308821808;
assign addr[17279]= -1184318708;
assign addr[17280]= -1053807919;
assign addr[17281]= -917951481;
assign addr[17282]= -777438554;
assign addr[17283]= -632981917;
assign addr[17284]= -485314355;
assign addr[17285]= -335184940;
assign addr[17286]= -183355234;
assign addr[17287]= -30595422;
assign addr[17288]= 122319591;
assign addr[17289]= 274614114;
assign addr[17290]= 425515602;
assign addr[17291]= 574258580;
assign addr[17292]= 720088517;
assign addr[17293]= 862265664;
assign addr[17294]= 1000068799;
assign addr[17295]= 1132798888;
assign addr[17296]= 1259782632;
assign addr[17297]= 1380375881;
assign addr[17298]= 1493966902;
assign addr[17299]= 1599979481;
assign addr[17300]= 1697875851;
assign addr[17301]= 1787159411;
assign addr[17302]= 1867377253;
assign addr[17303]= 1938122457;
assign addr[17304]= 1999036154;
assign addr[17305]= 2049809346;
assign addr[17306]= 2090184478;
assign addr[17307]= 2119956737;
assign addr[17308]= 2138975100;
assign addr[17309]= 2147143090;
assign addr[17310]= 2144419275;
assign addr[17311]= 2130817471;
assign addr[17312]= 2106406677;
assign addr[17313]= 2071310720;
assign addr[17314]= 2025707632;
assign addr[17315]= 1969828744;
assign addr[17316]= 1903957513;
assign addr[17317]= 1828428082;
assign addr[17318]= 1743623590;
assign addr[17319]= 1649974225;
assign addr[17320]= 1547955041;
assign addr[17321]= 1438083551;
assign addr[17322]= 1320917099;
assign addr[17323]= 1197050035;
assign addr[17324]= 1067110699;
assign addr[17325]= 931758235;
assign addr[17326]= 791679244;
assign addr[17327]= 647584304;
assign addr[17328]= 500204365;
assign addr[17329]= 350287041;
assign addr[17330]= 198592817;
assign addr[17331]= 45891193;
assign addr[17332]= -107043224;
assign addr[17333]= -259434643;
assign addr[17334]= -410510029;
assign addr[17335]= -559503022;
assign addr[17336]= -705657826;
assign addr[17337]= -848233042;
assign addr[17338]= -986505429;
assign addr[17339]= -1119773573;
assign addr[17340]= -1247361445;
assign addr[17341]= -1368621831;
assign addr[17342]= -1482939614;
assign addr[17343]= -1589734894;
assign addr[17344]= -1688465931;
assign addr[17345]= -1778631892;
assign addr[17346]= -1859775393;
assign addr[17347]= -1931484818;
assign addr[17348]= -1993396407;
assign addr[17349]= -2045196100;
assign addr[17350]= -2086621133;
assign addr[17351]= -2117461370;
assign addr[17352]= -2137560369;
assign addr[17353]= -2146816171;
assign addr[17354]= -2145181827;
assign addr[17355]= -2132665626;
assign addr[17356]= -2109331059;
assign addr[17357]= -2075296495;
assign addr[17358]= -2030734582;
assign addr[17359]= -1975871368;
assign addr[17360]= -1910985158;
assign addr[17361]= -1836405100;
assign addr[17362]= -1752509516;
assign addr[17363]= -1659723983;
assign addr[17364]= -1558519173;
assign addr[17365]= -1449408469;
assign addr[17366]= -1332945355;
assign addr[17367]= -1209720613;
assign addr[17368]= -1080359326;
assign addr[17369]= -945517704;
assign addr[17370]= -805879757;
assign addr[17371]= -662153826;
assign addr[17372]= -515068990;
assign addr[17373]= -365371365;
assign addr[17374]= -213820322;
assign addr[17375]= -61184634;
assign addr[17376]= 91761426;
assign addr[17377]= 244242007;
assign addr[17378]= 395483624;
assign addr[17379]= 544719071;
assign addr[17380]= 691191324;
assign addr[17381]= 834157373;
assign addr[17382]= 972891995;
assign addr[17383]= 1106691431;
assign addr[17384]= 1234876957;
assign addr[17385]= 1356798326;
assign addr[17386]= 1471837070;
assign addr[17387]= 1579409630;
assign addr[17388]= 1678970324;
assign addr[17389]= 1770014111;
assign addr[17390]= 1852079154;
assign addr[17391]= 1924749160;
assign addr[17392]= 1987655498;
assign addr[17393]= 2040479063;
assign addr[17394]= 2082951896;
assign addr[17395]= 2114858546;
assign addr[17396]= 2136037160;
assign addr[17397]= 2146380306;
assign addr[17398]= 2145835515;
assign addr[17399]= 2134405552;
assign addr[17400]= 2112148396;
assign addr[17401]= 2079176953;
assign addr[17402]= 2035658475;
assign addr[17403]= 1981813720;
assign addr[17404]= 1917915825;
assign addr[17405]= 1844288924;
assign addr[17406]= 1761306505;
assign addr[17407]= 1669389513;
assign addr[17408]= 1569004214;
assign addr[17409]= 1460659832;
assign addr[17410]= 1344905966;
assign addr[17411]= 1222329801;
assign addr[17412]= 1093553126;
assign addr[17413]= 959229189;
assign addr[17414]= 820039373;
assign addr[17415]= 676689746;
assign addr[17416]= 529907477;
assign addr[17417]= 380437148;
assign addr[17418]= 229036977;
assign addr[17419]= 76474970;
assign addr[17420]= -76474970;
assign addr[17421]= -229036977;
assign addr[17422]= -380437148;
assign addr[17423]= -529907477;
assign addr[17424]= -676689746;
assign addr[17425]= -820039373;
assign addr[17426]= -959229189;
assign addr[17427]= -1093553126;
assign addr[17428]= -1222329801;
assign addr[17429]= -1344905966;
assign addr[17430]= -1460659832;
assign addr[17431]= -1569004214;
assign addr[17432]= -1669389513;
assign addr[17433]= -1761306505;
assign addr[17434]= -1844288924;
assign addr[17435]= -1917915825;
assign addr[17436]= -1981813720;
assign addr[17437]= -2035658475;
assign addr[17438]= -2079176953;
assign addr[17439]= -2112148396;
assign addr[17440]= -2134405552;
assign addr[17441]= -2145835515;
assign addr[17442]= -2146380306;
assign addr[17443]= -2136037160;
assign addr[17444]= -2114858546;
assign addr[17445]= -2082951896;
assign addr[17446]= -2040479063;
assign addr[17447]= -1987655498;
assign addr[17448]= -1924749160;
assign addr[17449]= -1852079154;
assign addr[17450]= -1770014111;
assign addr[17451]= -1678970324;
assign addr[17452]= -1579409630;
assign addr[17453]= -1471837070;
assign addr[17454]= -1356798326;
assign addr[17455]= -1234876957;
assign addr[17456]= -1106691431;
assign addr[17457]= -972891995;
assign addr[17458]= -834157373;
assign addr[17459]= -691191324;
assign addr[17460]= -544719071;
assign addr[17461]= -395483624;
assign addr[17462]= -244242007;
assign addr[17463]= -91761426;
assign addr[17464]= 61184634;
assign addr[17465]= 213820322;
assign addr[17466]= 365371365;
assign addr[17467]= 515068990;
assign addr[17468]= 662153826;
assign addr[17469]= 805879757;
assign addr[17470]= 945517704;
assign addr[17471]= 1080359326;
assign addr[17472]= 1209720613;
assign addr[17473]= 1332945355;
assign addr[17474]= 1449408469;
assign addr[17475]= 1558519173;
assign addr[17476]= 1659723983;
assign addr[17477]= 1752509516;
assign addr[17478]= 1836405100;
assign addr[17479]= 1910985158;
assign addr[17480]= 1975871368;
assign addr[17481]= 2030734582;
assign addr[17482]= 2075296495;
assign addr[17483]= 2109331059;
assign addr[17484]= 2132665626;
assign addr[17485]= 2145181827;
assign addr[17486]= 2146816171;
assign addr[17487]= 2137560369;
assign addr[17488]= 2117461370;
assign addr[17489]= 2086621133;
assign addr[17490]= 2045196100;
assign addr[17491]= 1993396407;
assign addr[17492]= 1931484818;
assign addr[17493]= 1859775393;
assign addr[17494]= 1778631892;
assign addr[17495]= 1688465931;
assign addr[17496]= 1589734894;
assign addr[17497]= 1482939614;
assign addr[17498]= 1368621831;
assign addr[17499]= 1247361445;
assign addr[17500]= 1119773573;
assign addr[17501]= 986505429;
assign addr[17502]= 848233042;
assign addr[17503]= 705657826;
assign addr[17504]= 559503022;
assign addr[17505]= 410510029;
assign addr[17506]= 259434643;
assign addr[17507]= 107043224;
assign addr[17508]= -45891193;
assign addr[17509]= -198592817;
assign addr[17510]= -350287041;
assign addr[17511]= -500204365;
assign addr[17512]= -647584304;
assign addr[17513]= -791679244;
assign addr[17514]= -931758235;
assign addr[17515]= -1067110699;
assign addr[17516]= -1197050035;
assign addr[17517]= -1320917099;
assign addr[17518]= -1438083551;
assign addr[17519]= -1547955041;
assign addr[17520]= -1649974225;
assign addr[17521]= -1743623590;
assign addr[17522]= -1828428082;
assign addr[17523]= -1903957513;
assign addr[17524]= -1969828744;
assign addr[17525]= -2025707632;
assign addr[17526]= -2071310720;
assign addr[17527]= -2106406677;
assign addr[17528]= -2130817471;
assign addr[17529]= -2144419275;
assign addr[17530]= -2147143090;
assign addr[17531]= -2138975100;
assign addr[17532]= -2119956737;
assign addr[17533]= -2090184478;
assign addr[17534]= -2049809346;
assign addr[17535]= -1999036154;
assign addr[17536]= -1938122457;
assign addr[17537]= -1867377253;
assign addr[17538]= -1787159411;
assign addr[17539]= -1697875851;
assign addr[17540]= -1599979481;
assign addr[17541]= -1493966902;
assign addr[17542]= -1380375881;
assign addr[17543]= -1259782632;
assign addr[17544]= -1132798888;
assign addr[17545]= -1000068799;
assign addr[17546]= -862265664;
assign addr[17547]= -720088517;
assign addr[17548]= -574258580;
assign addr[17549]= -425515602;
assign addr[17550]= -274614114;
assign addr[17551]= -122319591;
assign addr[17552]= 30595422;
assign addr[17553]= 183355234;
assign addr[17554]= 335184940;
assign addr[17555]= 485314355;
assign addr[17556]= 632981917;
assign addr[17557]= 777438554;
assign addr[17558]= 917951481;
assign addr[17559]= 1053807919;
assign addr[17560]= 1184318708;
assign addr[17561]= 1308821808;
assign addr[17562]= 1426685652;
assign addr[17563]= 1537312353;
assign addr[17564]= 1640140734;
assign addr[17565]= 1734649179;
assign addr[17566]= 1820358275;
assign addr[17567]= 1896833245;
assign addr[17568]= 1963686155;
assign addr[17569]= 2020577882;
assign addr[17570]= 2067219829;
assign addr[17571]= 2103375398;
assign addr[17572]= 2128861181;
assign addr[17573]= 2143547897;
assign addr[17574]= 2147361045;
assign addr[17575]= 2140281282;
assign addr[17576]= 2122344521;
assign addr[17577]= 2093641749;
assign addr[17578]= 2054318569;
assign addr[17579]= 2004574453;
assign addr[17580]= 1944661739;
assign addr[17581]= 1874884346;
assign addr[17582]= 1795596234;
assign addr[17583]= 1707199606;
assign addr[17584]= 1610142873;
assign addr[17585]= 1504918373;
assign addr[17586]= 1392059879;
assign addr[17587]= 1272139887;
assign addr[17588]= 1145766716;
assign addr[17589]= 1013581418;
assign addr[17590]= 876254528;
assign addr[17591]= 734482665;
assign addr[17592]= 588984994;
assign addr[17593]= 440499581;
assign addr[17594]= 289779648;
assign addr[17595]= 137589750;
assign addr[17596]= -15298099;
assign addr[17597]= -168108346;
assign addr[17598]= -320065829;
assign addr[17599]= -470399716;
assign addr[17600]= -618347408;
assign addr[17601]= -763158411;
assign addr[17602]= -904098143;
assign addr[17603]= -1040451659;
assign addr[17604]= -1171527280;
assign addr[17605]= -1296660098;
assign addr[17606]= -1415215352;
assign addr[17607]= -1526591649;
assign addr[17608]= -1630224009;
assign addr[17609]= -1725586737;
assign addr[17610]= -1812196087;
assign addr[17611]= -1889612716;
assign addr[17612]= -1957443913;
assign addr[17613]= -2015345591;
assign addr[17614]= -2063024031;
assign addr[17615]= -2100237377;
assign addr[17616]= -2126796855;
assign addr[17617]= -2142567738;
assign addr[17618]= -2147470025;
assign addr[17619]= -2141478848;
assign addr[17620]= -2124624598;
assign addr[17621]= -2096992772;
assign addr[17622]= -2058723538;
assign addr[17623]= -2010011024;
assign addr[17624]= -1951102334;
assign addr[17625]= -1882296293;
assign addr[17626]= -1803941934;
assign addr[17627]= -1716436725;
assign addr[17628]= -1620224553;
assign addr[17629]= -1515793473;
assign addr[17630]= -1403673233;
assign addr[17631]= -1284432584;
assign addr[17632]= -1158676398;
assign addr[17633]= -1027042599;
assign addr[17634]= -890198924;
assign addr[17635]= -748839539;
assign addr[17636]= -603681519;
assign addr[17637]= -455461206;
assign addr[17638]= -304930476;
assign addr[17639]= -152852926;
assign addr[17640]= 0;
assign addr[17641]= 152852926;
assign addr[17642]= 304930476;
assign addr[17643]= 455461206;
assign addr[17644]= 603681519;
assign addr[17645]= 748839539;
assign addr[17646]= 890198924;
assign addr[17647]= 1027042599;
assign addr[17648]= 1158676398;
assign addr[17649]= 1284432584;
assign addr[17650]= 1403673233;
assign addr[17651]= 1515793473;
assign addr[17652]= 1620224553;
assign addr[17653]= 1716436725;
assign addr[17654]= 1803941934;
assign addr[17655]= 1882296293;
assign addr[17656]= 1951102334;
assign addr[17657]= 2010011024;
assign addr[17658]= 2058723538;
assign addr[17659]= 2096992772;
assign addr[17660]= 2124624598;
assign addr[17661]= 2141478848;
assign addr[17662]= 2147470025;
assign addr[17663]= 2142567738;
assign addr[17664]= 2126796855;
assign addr[17665]= 2100237377;
assign addr[17666]= 2063024031;
assign addr[17667]= 2015345591;
assign addr[17668]= 1957443913;
assign addr[17669]= 1889612716;
assign addr[17670]= 1812196087;
assign addr[17671]= 1725586737;
assign addr[17672]= 1630224009;
assign addr[17673]= 1526591649;
assign addr[17674]= 1415215352;
assign addr[17675]= 1296660098;
assign addr[17676]= 1171527280;
assign addr[17677]= 1040451659;
assign addr[17678]= 904098143;
assign addr[17679]= 763158411;
assign addr[17680]= 618347408;
assign addr[17681]= 470399716;
assign addr[17682]= 320065829;
assign addr[17683]= 168108346;
assign addr[17684]= 15298099;
assign addr[17685]= -137589750;
assign addr[17686]= -289779648;
assign addr[17687]= -440499581;
assign addr[17688]= -588984994;
assign addr[17689]= -734482665;
assign addr[17690]= -876254528;
assign addr[17691]= -1013581418;
assign addr[17692]= -1145766716;
assign addr[17693]= -1272139887;
assign addr[17694]= -1392059879;
assign addr[17695]= -1504918373;
assign addr[17696]= -1610142873;
assign addr[17697]= -1707199606;
assign addr[17698]= -1795596234;
assign addr[17699]= -1874884346;
assign addr[17700]= -1944661739;
assign addr[17701]= -2004574453;
assign addr[17702]= -2054318569;
assign addr[17703]= -2093641749;
assign addr[17704]= -2122344521;
assign addr[17705]= -2140281282;
assign addr[17706]= -2147361045;
assign addr[17707]= -2143547897;
assign addr[17708]= -2128861181;
assign addr[17709]= -2103375398;
assign addr[17710]= -2067219829;
assign addr[17711]= -2020577882;
assign addr[17712]= -1963686155;
assign addr[17713]= -1896833245;
assign addr[17714]= -1820358275;
assign addr[17715]= -1734649179;
assign addr[17716]= -1640140734;
assign addr[17717]= -1537312353;
assign addr[17718]= -1426685652;
assign addr[17719]= -1308821808;
assign addr[17720]= -1184318708;
assign addr[17721]= -1053807919;
assign addr[17722]= -917951481;
assign addr[17723]= -777438554;
assign addr[17724]= -632981917;
assign addr[17725]= -485314355;
assign addr[17726]= -335184940;
assign addr[17727]= -183355234;
assign addr[17728]= -30595422;
assign addr[17729]= 122319591;
assign addr[17730]= 274614114;
assign addr[17731]= 425515602;
assign addr[17732]= 574258580;
assign addr[17733]= 720088517;
assign addr[17734]= 862265664;
assign addr[17735]= 1000068799;
assign addr[17736]= 1132798888;
assign addr[17737]= 1259782632;
assign addr[17738]= 1380375881;
assign addr[17739]= 1493966902;
assign addr[17740]= 1599979481;
assign addr[17741]= 1697875851;
assign addr[17742]= 1787159411;
assign addr[17743]= 1867377253;
assign addr[17744]= 1938122457;
assign addr[17745]= 1999036154;
assign addr[17746]= 2049809346;
assign addr[17747]= 2090184478;
assign addr[17748]= 2119956737;
assign addr[17749]= 2138975100;
assign addr[17750]= 2147143090;
assign addr[17751]= 2144419275;
assign addr[17752]= 2130817471;
assign addr[17753]= 2106406677;
assign addr[17754]= 2071310720;
assign addr[17755]= 2025707632;
assign addr[17756]= 1969828744;
assign addr[17757]= 1903957513;
assign addr[17758]= 1828428082;
assign addr[17759]= 1743623590;
assign addr[17760]= 1649974225;
assign addr[17761]= 1547955041;
assign addr[17762]= 1438083551;
assign addr[17763]= 1320917099;
assign addr[17764]= 1197050035;
assign addr[17765]= 1067110699;
assign addr[17766]= 931758235;
assign addr[17767]= 791679244;
assign addr[17768]= 647584304;
assign addr[17769]= 500204365;
assign addr[17770]= 350287041;
assign addr[17771]= 198592817;
assign addr[17772]= 45891193;
assign addr[17773]= -107043224;
assign addr[17774]= -259434643;
assign addr[17775]= -410510029;
assign addr[17776]= -559503022;
assign addr[17777]= -705657826;
assign addr[17778]= -848233042;
assign addr[17779]= -986505429;
assign addr[17780]= -1119773573;
assign addr[17781]= -1247361445;
assign addr[17782]= -1368621831;
assign addr[17783]= -1482939614;
assign addr[17784]= -1589734894;
assign addr[17785]= -1688465931;
assign addr[17786]= -1778631892;
assign addr[17787]= -1859775393;
assign addr[17788]= -1931484818;
assign addr[17789]= -1993396407;
assign addr[17790]= -2045196100;
assign addr[17791]= -2086621133;
assign addr[17792]= -2117461370;
assign addr[17793]= -2137560369;
assign addr[17794]= -2146816171;
assign addr[17795]= -2145181827;
assign addr[17796]= -2132665626;
assign addr[17797]= -2109331059;
assign addr[17798]= -2075296495;
assign addr[17799]= -2030734582;
assign addr[17800]= -1975871368;
assign addr[17801]= -1910985158;
assign addr[17802]= -1836405100;
assign addr[17803]= -1752509516;
assign addr[17804]= -1659723983;
assign addr[17805]= -1558519173;
assign addr[17806]= -1449408469;
assign addr[17807]= -1332945355;
assign addr[17808]= -1209720613;
assign addr[17809]= -1080359326;
assign addr[17810]= -945517704;
assign addr[17811]= -805879757;
assign addr[17812]= -662153826;
assign addr[17813]= -515068990;
assign addr[17814]= -365371365;
assign addr[17815]= -213820322;
assign addr[17816]= -61184634;
assign addr[17817]= 91761426;
assign addr[17818]= 244242007;
assign addr[17819]= 395483624;
assign addr[17820]= 544719071;
assign addr[17821]= 691191324;
assign addr[17822]= 834157373;
assign addr[17823]= 972891995;
assign addr[17824]= 1106691431;
assign addr[17825]= 1234876957;
assign addr[17826]= 1356798326;
assign addr[17827]= 1471837070;
assign addr[17828]= 1579409630;
assign addr[17829]= 1678970324;
assign addr[17830]= 1770014111;
assign addr[17831]= 1852079154;
assign addr[17832]= 1924749160;
assign addr[17833]= 1987655498;
assign addr[17834]= 2040479063;
assign addr[17835]= 2082951896;
assign addr[17836]= 2114858546;
assign addr[17837]= 2136037160;
assign addr[17838]= 2146380306;
assign addr[17839]= 2145835515;
assign addr[17840]= 2134405552;
assign addr[17841]= 2112148396;
assign addr[17842]= 2079176953;
assign addr[17843]= 2035658475;
assign addr[17844]= 1981813720;
assign addr[17845]= 1917915825;
assign addr[17846]= 1844288924;
assign addr[17847]= 1761306505;
assign addr[17848]= 1669389513;
assign addr[17849]= 1569004214;
assign addr[17850]= 1460659832;
assign addr[17851]= 1344905966;
assign addr[17852]= 1222329801;
assign addr[17853]= 1093553126;
assign addr[17854]= 959229189;
assign addr[17855]= 820039373;
assign addr[17856]= 676689746;
assign addr[17857]= 529907477;
assign addr[17858]= 380437148;
assign addr[17859]= 229036977;
assign addr[17860]= 76474970;
assign addr[17861]= -76474970;
assign addr[17862]= -229036977;
assign addr[17863]= -380437148;
assign addr[17864]= -529907477;
assign addr[17865]= -676689746;
assign addr[17866]= -820039373;
assign addr[17867]= -959229189;
assign addr[17868]= -1093553126;
assign addr[17869]= -1222329801;
assign addr[17870]= -1344905966;
assign addr[17871]= -1460659832;
assign addr[17872]= -1569004214;
assign addr[17873]= -1669389513;
assign addr[17874]= -1761306505;
assign addr[17875]= -1844288924;
assign addr[17876]= -1917915825;
assign addr[17877]= -1981813720;
assign addr[17878]= -2035658475;
assign addr[17879]= -2079176953;
assign addr[17880]= -2112148396;
assign addr[17881]= -2134405552;
assign addr[17882]= -2145835515;
assign addr[17883]= -2146380306;
assign addr[17884]= -2136037160;
assign addr[17885]= -2114858546;
assign addr[17886]= -2082951896;
assign addr[17887]= -2040479063;
assign addr[17888]= -1987655498;
assign addr[17889]= -1924749160;
assign addr[17890]= -1852079154;
assign addr[17891]= -1770014111;
assign addr[17892]= -1678970324;
assign addr[17893]= -1579409630;
assign addr[17894]= -1471837070;
assign addr[17895]= -1356798326;
assign addr[17896]= -1234876957;
assign addr[17897]= -1106691431;
assign addr[17898]= -972891995;
assign addr[17899]= -834157373;
assign addr[17900]= -691191324;
assign addr[17901]= -544719071;
assign addr[17902]= -395483624;
assign addr[17903]= -244242007;
assign addr[17904]= -91761426;
assign addr[17905]= 61184634;
assign addr[17906]= 213820322;
assign addr[17907]= 365371365;
assign addr[17908]= 515068990;
assign addr[17909]= 662153826;
assign addr[17910]= 805879757;
assign addr[17911]= 945517704;
assign addr[17912]= 1080359326;
assign addr[17913]= 1209720613;
assign addr[17914]= 1332945355;
assign addr[17915]= 1449408469;
assign addr[17916]= 1558519173;
assign addr[17917]= 1659723983;
assign addr[17918]= 1752509516;
assign addr[17919]= 1836405100;
assign addr[17920]= 1910985158;
assign addr[17921]= 1975871368;
assign addr[17922]= 2030734582;
assign addr[17923]= 2075296495;
assign addr[17924]= 2109331059;
assign addr[17925]= 2132665626;
assign addr[17926]= 2145181827;
assign addr[17927]= 2146816171;
assign addr[17928]= 2137560369;
assign addr[17929]= 2117461370;
assign addr[17930]= 2086621133;
assign addr[17931]= 2045196100;
assign addr[17932]= 1993396407;
assign addr[17933]= 1931484818;
assign addr[17934]= 1859775393;
assign addr[17935]= 1778631892;
assign addr[17936]= 1688465931;
assign addr[17937]= 1589734894;
assign addr[17938]= 1482939614;
assign addr[17939]= 1368621831;
assign addr[17940]= 1247361445;
assign addr[17941]= 1119773573;
assign addr[17942]= 986505429;
assign addr[17943]= 848233042;
assign addr[17944]= 705657826;
assign addr[17945]= 559503022;
assign addr[17946]= 410510029;
assign addr[17947]= 259434643;
assign addr[17948]= 107043224;
assign addr[17949]= -45891193;
assign addr[17950]= -198592817;
assign addr[17951]= -350287041;
assign addr[17952]= -500204365;
assign addr[17953]= -647584304;
assign addr[17954]= -791679244;
assign addr[17955]= -931758235;
assign addr[17956]= -1067110699;
assign addr[17957]= -1197050035;
assign addr[17958]= -1320917099;
assign addr[17959]= -1438083551;
assign addr[17960]= -1547955041;
assign addr[17961]= -1649974225;
assign addr[17962]= -1743623590;
assign addr[17963]= -1828428082;
assign addr[17964]= -1903957513;
assign addr[17965]= -1969828744;
assign addr[17966]= -2025707632;
assign addr[17967]= -2071310720;
assign addr[17968]= -2106406677;
assign addr[17969]= -2130817471;
assign addr[17970]= -2144419275;
assign addr[17971]= -2147143090;
assign addr[17972]= -2138975100;
assign addr[17973]= -2119956737;
assign addr[17974]= -2090184478;
assign addr[17975]= -2049809346;
assign addr[17976]= -1999036154;
assign addr[17977]= -1938122457;
assign addr[17978]= -1867377253;
assign addr[17979]= -1787159411;
assign addr[17980]= -1697875851;
assign addr[17981]= -1599979481;
assign addr[17982]= -1493966902;
assign addr[17983]= -1380375881;
assign addr[17984]= -1259782632;
assign addr[17985]= -1132798888;
assign addr[17986]= -1000068799;
assign addr[17987]= -862265664;
assign addr[17988]= -720088517;
assign addr[17989]= -574258580;
assign addr[17990]= -425515602;
assign addr[17991]= -274614114;
assign addr[17992]= -122319591;
assign addr[17993]= 30595422;
assign addr[17994]= 183355234;
assign addr[17995]= 335184940;
assign addr[17996]= 485314355;
assign addr[17997]= 632981917;
assign addr[17998]= 777438554;
assign addr[17999]= 917951481;
assign addr[18000]= 1053807919;
assign addr[18001]= 1184318708;
assign addr[18002]= 1308821808;
assign addr[18003]= 1426685652;
assign addr[18004]= 1537312353;
assign addr[18005]= 1640140734;
assign addr[18006]= 1734649179;
assign addr[18007]= 1820358275;
assign addr[18008]= 1896833245;
assign addr[18009]= 1963686155;
assign addr[18010]= 2020577882;
assign addr[18011]= 2067219829;
assign addr[18012]= 2103375398;
assign addr[18013]= 2128861181;
assign addr[18014]= 2143547897;
assign addr[18015]= 2147361045;
assign addr[18016]= 2140281282;
assign addr[18017]= 2122344521;
assign addr[18018]= 2093641749;
assign addr[18019]= 2054318569;
assign addr[18020]= 2004574453;
assign addr[18021]= 1944661739;
assign addr[18022]= 1874884346;
assign addr[18023]= 1795596234;
assign addr[18024]= 1707199606;
assign addr[18025]= 1610142873;
assign addr[18026]= 1504918373;
assign addr[18027]= 1392059879;
assign addr[18028]= 1272139887;
assign addr[18029]= 1145766716;
assign addr[18030]= 1013581418;
assign addr[18031]= 876254528;
assign addr[18032]= 734482665;
assign addr[18033]= 588984994;
assign addr[18034]= 440499581;
assign addr[18035]= 289779648;
assign addr[18036]= 137589750;
assign addr[18037]= -15298099;
assign addr[18038]= -168108346;
assign addr[18039]= -320065829;
assign addr[18040]= -470399716;
assign addr[18041]= -618347408;
assign addr[18042]= -763158411;
assign addr[18043]= -904098143;
assign addr[18044]= -1040451659;
assign addr[18045]= -1171527280;
assign addr[18046]= -1296660098;
assign addr[18047]= -1415215352;
assign addr[18048]= -1526591649;
assign addr[18049]= -1630224009;
assign addr[18050]= -1725586737;
assign addr[18051]= -1812196087;
assign addr[18052]= -1889612716;
assign addr[18053]= -1957443913;
assign addr[18054]= -2015345591;
assign addr[18055]= -2063024031;
assign addr[18056]= -2100237377;
assign addr[18057]= -2126796855;
assign addr[18058]= -2142567738;
assign addr[18059]= -2147470025;
assign addr[18060]= -2141478848;
assign addr[18061]= -2124624598;
assign addr[18062]= -2096992772;
assign addr[18063]= -2058723538;
assign addr[18064]= -2010011024;
assign addr[18065]= -1951102334;
assign addr[18066]= -1882296293;
assign addr[18067]= -1803941934;
assign addr[18068]= -1716436725;
assign addr[18069]= -1620224553;
assign addr[18070]= -1515793473;
assign addr[18071]= -1403673233;
assign addr[18072]= -1284432584;
assign addr[18073]= -1158676398;
assign addr[18074]= -1027042599;
assign addr[18075]= -890198924;
assign addr[18076]= -748839539;
assign addr[18077]= -603681519;
assign addr[18078]= -455461206;
assign addr[18079]= -304930476;
assign addr[18080]= -152852926;
assign addr[18081]= 0;
assign addr[18082]= 152852926;
assign addr[18083]= 304930476;
assign addr[18084]= 455461206;
assign addr[18085]= 603681519;
assign addr[18086]= 748839539;
assign addr[18087]= 890198924;
assign addr[18088]= 1027042599;
assign addr[18089]= 1158676398;
assign addr[18090]= 1284432584;
assign addr[18091]= 1403673233;
assign addr[18092]= 1515793473;
assign addr[18093]= 1620224553;
assign addr[18094]= 1716436725;
assign addr[18095]= 1803941934;
assign addr[18096]= 1882296293;
assign addr[18097]= 1951102334;
assign addr[18098]= 2010011024;
assign addr[18099]= 2058723538;
assign addr[18100]= 2096992772;
assign addr[18101]= 2124624598;
assign addr[18102]= 2141478848;
assign addr[18103]= 2147470025;
assign addr[18104]= 2142567738;
assign addr[18105]= 2126796855;
assign addr[18106]= 2100237377;
assign addr[18107]= 2063024031;
assign addr[18108]= 2015345591;
assign addr[18109]= 1957443913;
assign addr[18110]= 1889612716;
assign addr[18111]= 1812196087;
assign addr[18112]= 1725586737;
assign addr[18113]= 1630224009;
assign addr[18114]= 1526591649;
assign addr[18115]= 1415215352;
assign addr[18116]= 1296660098;
assign addr[18117]= 1171527280;
assign addr[18118]= 1040451659;
assign addr[18119]= 904098143;
assign addr[18120]= 763158411;
assign addr[18121]= 618347408;
assign addr[18122]= 470399716;
assign addr[18123]= 320065829;
assign addr[18124]= 168108346;
assign addr[18125]= 15298099;
assign addr[18126]= -137589750;
assign addr[18127]= -289779648;
assign addr[18128]= -440499581;
assign addr[18129]= -588984994;
assign addr[18130]= -734482665;
assign addr[18131]= -876254528;
assign addr[18132]= -1013581418;
assign addr[18133]= -1145766716;
assign addr[18134]= -1272139887;
assign addr[18135]= -1392059879;
assign addr[18136]= -1504918373;
assign addr[18137]= -1610142873;
assign addr[18138]= -1707199606;
assign addr[18139]= -1795596234;
assign addr[18140]= -1874884346;
assign addr[18141]= -1944661739;
assign addr[18142]= -2004574453;
assign addr[18143]= -2054318569;
assign addr[18144]= -2093641749;
assign addr[18145]= -2122344521;
assign addr[18146]= -2140281282;
assign addr[18147]= -2147361045;
assign addr[18148]= -2143547897;
assign addr[18149]= -2128861181;
assign addr[18150]= -2103375398;
assign addr[18151]= -2067219829;
assign addr[18152]= -2020577882;
assign addr[18153]= -1963686155;
assign addr[18154]= -1896833245;
assign addr[18155]= -1820358275;
assign addr[18156]= -1734649179;
assign addr[18157]= -1640140734;
assign addr[18158]= -1537312353;
assign addr[18159]= -1426685652;
assign addr[18160]= -1308821808;
assign addr[18161]= -1184318708;
assign addr[18162]= -1053807919;
assign addr[18163]= -917951481;
assign addr[18164]= -777438554;
assign addr[18165]= -632981917;
assign addr[18166]= -485314355;
assign addr[18167]= -335184940;
assign addr[18168]= -183355234;
assign addr[18169]= -30595422;
assign addr[18170]= 122319591;
assign addr[18171]= 274614114;
assign addr[18172]= 425515602;
assign addr[18173]= 574258580;
assign addr[18174]= 720088517;
assign addr[18175]= 862265664;
assign addr[18176]= 1000068799;
assign addr[18177]= 1132798888;
assign addr[18178]= 1259782632;
assign addr[18179]= 1380375881;
assign addr[18180]= 1493966902;
assign addr[18181]= 1599979481;
assign addr[18182]= 1697875851;
assign addr[18183]= 1787159411;
assign addr[18184]= 1867377253;
assign addr[18185]= 1938122457;
assign addr[18186]= 1999036154;
assign addr[18187]= 2049809346;
assign addr[18188]= 2090184478;
assign addr[18189]= 2119956737;
assign addr[18190]= 2138975100;
assign addr[18191]= 2147143090;
assign addr[18192]= 2144419275;
assign addr[18193]= 2130817471;
assign addr[18194]= 2106406677;
assign addr[18195]= 2071310720;
assign addr[18196]= 2025707632;
assign addr[18197]= 1969828744;
assign addr[18198]= 1903957513;
assign addr[18199]= 1828428082;
assign addr[18200]= 1743623590;
assign addr[18201]= 1649974225;
assign addr[18202]= 1547955041;
assign addr[18203]= 1438083551;
assign addr[18204]= 1320917099;
assign addr[18205]= 1197050035;
assign addr[18206]= 1067110699;
assign addr[18207]= 931758235;
assign addr[18208]= 791679244;
assign addr[18209]= 647584304;
assign addr[18210]= 500204365;
assign addr[18211]= 350287041;
assign addr[18212]= 198592817;
assign addr[18213]= 45891193;
assign addr[18214]= -107043224;
assign addr[18215]= -259434643;
assign addr[18216]= -410510029;
assign addr[18217]= -559503022;
assign addr[18218]= -705657826;
assign addr[18219]= -848233042;
assign addr[18220]= -986505429;
assign addr[18221]= -1119773573;
assign addr[18222]= -1247361445;
assign addr[18223]= -1368621831;
assign addr[18224]= -1482939614;
assign addr[18225]= -1589734894;
assign addr[18226]= -1688465931;
assign addr[18227]= -1778631892;
assign addr[18228]= -1859775393;
assign addr[18229]= -1931484818;
assign addr[18230]= -1993396407;
assign addr[18231]= -2045196100;
assign addr[18232]= -2086621133;
assign addr[18233]= -2117461370;
assign addr[18234]= -2137560369;
assign addr[18235]= -2146816171;
assign addr[18236]= -2145181827;
assign addr[18237]= -2132665626;
assign addr[18238]= -2109331059;
assign addr[18239]= -2075296495;
assign addr[18240]= -2030734582;
assign addr[18241]= -1975871368;
assign addr[18242]= -1910985158;
assign addr[18243]= -1836405100;
assign addr[18244]= -1752509516;
assign addr[18245]= -1659723983;
assign addr[18246]= -1558519173;
assign addr[18247]= -1449408469;
assign addr[18248]= -1332945355;
assign addr[18249]= -1209720613;
assign addr[18250]= -1080359326;
assign addr[18251]= -945517704;
assign addr[18252]= -805879757;
assign addr[18253]= -662153826;
assign addr[18254]= -515068990;
assign addr[18255]= -365371365;
assign addr[18256]= -213820322;
assign addr[18257]= -61184634;
assign addr[18258]= 91761426;
assign addr[18259]= 244242007;
assign addr[18260]= 395483624;
assign addr[18261]= 544719071;
assign addr[18262]= 691191324;
assign addr[18263]= 834157373;
assign addr[18264]= 972891995;
assign addr[18265]= 1106691431;
assign addr[18266]= 1234876957;
assign addr[18267]= 1356798326;
assign addr[18268]= 1471837070;
assign addr[18269]= 1579409630;
assign addr[18270]= 1678970324;
assign addr[18271]= 1770014111;
assign addr[18272]= 1852079154;
assign addr[18273]= 1924749160;
assign addr[18274]= 1987655498;
assign addr[18275]= 2040479063;
assign addr[18276]= 2082951896;
assign addr[18277]= 2114858546;
assign addr[18278]= 2136037160;
assign addr[18279]= 2146380306;
assign addr[18280]= 2145835515;
assign addr[18281]= 2134405552;
assign addr[18282]= 2112148396;
assign addr[18283]= 2079176953;
assign addr[18284]= 2035658475;
assign addr[18285]= 1981813720;
assign addr[18286]= 1917915825;
assign addr[18287]= 1844288924;
assign addr[18288]= 1761306505;
assign addr[18289]= 1669389513;
assign addr[18290]= 1569004214;
assign addr[18291]= 1460659832;
assign addr[18292]= 1344905966;
assign addr[18293]= 1222329801;
assign addr[18294]= 1093553126;
assign addr[18295]= 959229189;
assign addr[18296]= 820039373;
assign addr[18297]= 676689746;
assign addr[18298]= 529907477;
assign addr[18299]= 380437148;
assign addr[18300]= 229036977;
assign addr[18301]= 76474970;
assign addr[18302]= -76474970;
assign addr[18303]= -229036977;
assign addr[18304]= -380437148;
assign addr[18305]= -529907477;
assign addr[18306]= -676689746;
assign addr[18307]= -820039373;
assign addr[18308]= -959229189;
assign addr[18309]= -1093553126;
assign addr[18310]= -1222329801;
assign addr[18311]= -1344905966;
assign addr[18312]= -1460659832;
assign addr[18313]= -1569004214;
assign addr[18314]= -1669389513;
assign addr[18315]= -1761306505;
assign addr[18316]= -1844288924;
assign addr[18317]= -1917915825;
assign addr[18318]= -1981813720;
assign addr[18319]= -2035658475;
assign addr[18320]= -2079176953;
assign addr[18321]= -2112148396;
assign addr[18322]= -2134405552;
assign addr[18323]= -2145835515;
assign addr[18324]= -2146380306;
assign addr[18325]= -2136037160;
assign addr[18326]= -2114858546;
assign addr[18327]= -2082951896;
assign addr[18328]= -2040479063;
assign addr[18329]= -1987655498;
assign addr[18330]= -1924749160;
assign addr[18331]= -1852079154;
assign addr[18332]= -1770014111;
assign addr[18333]= -1678970324;
assign addr[18334]= -1579409630;
assign addr[18335]= -1471837070;
assign addr[18336]= -1356798326;
assign addr[18337]= -1234876957;
assign addr[18338]= -1106691431;
assign addr[18339]= -972891995;
assign addr[18340]= -834157373;
assign addr[18341]= -691191324;
assign addr[18342]= -544719071;
assign addr[18343]= -395483624;
assign addr[18344]= -244242007;
assign addr[18345]= -91761426;
assign addr[18346]= 61184634;
assign addr[18347]= 213820322;
assign addr[18348]= 365371365;
assign addr[18349]= 515068990;
assign addr[18350]= 662153826;
assign addr[18351]= 805879757;
assign addr[18352]= 945517704;
assign addr[18353]= 1080359326;
assign addr[18354]= 1209720613;
assign addr[18355]= 1332945355;
assign addr[18356]= 1449408469;
assign addr[18357]= 1558519173;
assign addr[18358]= 1659723983;
assign addr[18359]= 1752509516;
assign addr[18360]= 1836405100;
assign addr[18361]= 1910985158;
assign addr[18362]= 1975871368;
assign addr[18363]= 2030734582;
assign addr[18364]= 2075296495;
assign addr[18365]= 2109331059;
assign addr[18366]= 2132665626;
assign addr[18367]= 2145181827;
assign addr[18368]= 2146816171;
assign addr[18369]= 2137560369;
assign addr[18370]= 2117461370;
assign addr[18371]= 2086621133;
assign addr[18372]= 2045196100;
assign addr[18373]= 1993396407;
assign addr[18374]= 1931484818;
assign addr[18375]= 1859775393;
assign addr[18376]= 1778631892;
assign addr[18377]= 1688465931;
assign addr[18378]= 1589734894;
assign addr[18379]= 1482939614;
assign addr[18380]= 1368621831;
assign addr[18381]= 1247361445;
assign addr[18382]= 1119773573;
assign addr[18383]= 986505429;
assign addr[18384]= 848233042;
assign addr[18385]= 705657826;
assign addr[18386]= 559503022;
assign addr[18387]= 410510029;
assign addr[18388]= 259434643;
assign addr[18389]= 107043224;
assign addr[18390]= -45891193;
assign addr[18391]= -198592817;
assign addr[18392]= -350287041;
assign addr[18393]= -500204365;
assign addr[18394]= -647584304;
assign addr[18395]= -791679244;
assign addr[18396]= -931758235;
assign addr[18397]= -1067110699;
assign addr[18398]= -1197050035;
assign addr[18399]= -1320917099;
assign addr[18400]= -1438083551;
assign addr[18401]= -1547955041;
assign addr[18402]= -1649974225;
assign addr[18403]= -1743623590;
assign addr[18404]= -1828428082;
assign addr[18405]= -1903957513;
assign addr[18406]= -1969828744;
assign addr[18407]= -2025707632;
assign addr[18408]= -2071310720;
assign addr[18409]= -2106406677;
assign addr[18410]= -2130817471;
assign addr[18411]= -2144419275;
assign addr[18412]= -2147143090;
assign addr[18413]= -2138975100;
assign addr[18414]= -2119956737;
assign addr[18415]= -2090184478;
assign addr[18416]= -2049809346;
assign addr[18417]= -1999036154;
assign addr[18418]= -1938122457;
assign addr[18419]= -1867377253;
assign addr[18420]= -1787159411;
assign addr[18421]= -1697875851;
assign addr[18422]= -1599979481;
assign addr[18423]= -1493966902;
assign addr[18424]= -1380375881;
assign addr[18425]= -1259782632;
assign addr[18426]= -1132798888;
assign addr[18427]= -1000068799;
assign addr[18428]= -862265664;
assign addr[18429]= -720088517;
assign addr[18430]= -574258580;
assign addr[18431]= -425515602;
assign addr[18432]= -274614114;
assign addr[18433]= -122319591;
assign addr[18434]= 30595422;
assign addr[18435]= 183355234;
assign addr[18436]= 335184940;
assign addr[18437]= 485314355;
assign addr[18438]= 632981917;
assign addr[18439]= 777438554;
assign addr[18440]= 917951481;
assign addr[18441]= 1053807919;
assign addr[18442]= 1184318708;
assign addr[18443]= 1308821808;
assign addr[18444]= 1426685652;
assign addr[18445]= 1537312353;
assign addr[18446]= 1640140734;
assign addr[18447]= 1734649179;
assign addr[18448]= 1820358275;
assign addr[18449]= 1896833245;
assign addr[18450]= 1963686155;
assign addr[18451]= 2020577882;
assign addr[18452]= 2067219829;
assign addr[18453]= 2103375398;
assign addr[18454]= 2128861181;
assign addr[18455]= 2143547897;
assign addr[18456]= 2147361045;
assign addr[18457]= 2140281282;
assign addr[18458]= 2122344521;
assign addr[18459]= 2093641749;
assign addr[18460]= 2054318569;
assign addr[18461]= 2004574453;
assign addr[18462]= 1944661739;
assign addr[18463]= 1874884346;
assign addr[18464]= 1795596234;
assign addr[18465]= 1707199606;
assign addr[18466]= 1610142873;
assign addr[18467]= 1504918373;
assign addr[18468]= 1392059879;
assign addr[18469]= 1272139887;
assign addr[18470]= 1145766716;
assign addr[18471]= 1013581418;
assign addr[18472]= 876254528;
assign addr[18473]= 734482665;
assign addr[18474]= 588984994;
assign addr[18475]= 440499581;
assign addr[18476]= 289779648;
assign addr[18477]= 137589750;
assign addr[18478]= -15298099;
assign addr[18479]= -168108346;
assign addr[18480]= -320065829;
assign addr[18481]= -470399716;
assign addr[18482]= -618347408;
assign addr[18483]= -763158411;
assign addr[18484]= -904098143;
assign addr[18485]= -1040451659;
assign addr[18486]= -1171527280;
assign addr[18487]= -1296660098;
assign addr[18488]= -1415215352;
assign addr[18489]= -1526591649;
assign addr[18490]= -1630224009;
assign addr[18491]= -1725586737;
assign addr[18492]= -1812196087;
assign addr[18493]= -1889612716;
assign addr[18494]= -1957443913;
assign addr[18495]= -2015345591;
assign addr[18496]= -2063024031;
assign addr[18497]= -2100237377;
assign addr[18498]= -2126796855;
assign addr[18499]= -2142567738;
assign addr[18500]= -2147470025;
assign addr[18501]= -2141478848;
assign addr[18502]= -2124624598;
assign addr[18503]= -2096992772;
assign addr[18504]= -2058723538;
assign addr[18505]= -2010011024;
assign addr[18506]= -1951102334;
assign addr[18507]= -1882296293;
assign addr[18508]= -1803941934;
assign addr[18509]= -1716436725;
assign addr[18510]= -1620224553;
assign addr[18511]= -1515793473;
assign addr[18512]= -1403673233;
assign addr[18513]= -1284432584;
assign addr[18514]= -1158676398;
assign addr[18515]= -1027042599;
assign addr[18516]= -890198924;
assign addr[18517]= -748839539;
assign addr[18518]= -603681519;
assign addr[18519]= -455461206;
assign addr[18520]= -304930476;
assign addr[18521]= -152852926;
assign addr[18522]= 0;
assign addr[18523]= 152852926;
assign addr[18524]= 304930476;
assign addr[18525]= 455461206;
assign addr[18526]= 603681519;
assign addr[18527]= 748839539;
assign addr[18528]= 890198924;
assign addr[18529]= 1027042599;
assign addr[18530]= 1158676398;
assign addr[18531]= 1284432584;
assign addr[18532]= 1403673233;
assign addr[18533]= 1515793473;
assign addr[18534]= 1620224553;
assign addr[18535]= 1716436725;
assign addr[18536]= 1803941934;
assign addr[18537]= 1882296293;
assign addr[18538]= 1951102334;
assign addr[18539]= 2010011024;
assign addr[18540]= 2058723538;
assign addr[18541]= 2096992772;
assign addr[18542]= 2124624598;
assign addr[18543]= 2141478848;
assign addr[18544]= 2147470025;
assign addr[18545]= 2142567738;
assign addr[18546]= 2126796855;
assign addr[18547]= 2100237377;
assign addr[18548]= 2063024031;
assign addr[18549]= 2015345591;
assign addr[18550]= 1957443913;
assign addr[18551]= 1889612716;
assign addr[18552]= 1812196087;
assign addr[18553]= 1725586737;
assign addr[18554]= 1630224009;
assign addr[18555]= 1526591649;
assign addr[18556]= 1415215352;
assign addr[18557]= 1296660098;
assign addr[18558]= 1171527280;
assign addr[18559]= 1040451659;
assign addr[18560]= 904098143;
assign addr[18561]= 763158411;
assign addr[18562]= 618347408;
assign addr[18563]= 470399716;
assign addr[18564]= 320065829;
assign addr[18565]= 168108346;
assign addr[18566]= 15298099;
assign addr[18567]= -137589750;
assign addr[18568]= -289779648;
assign addr[18569]= -440499581;
assign addr[18570]= -588984994;
assign addr[18571]= -734482665;
assign addr[18572]= -876254528;
assign addr[18573]= -1013581418;
assign addr[18574]= -1145766716;
assign addr[18575]= -1272139887;
assign addr[18576]= -1392059879;
assign addr[18577]= -1504918373;
assign addr[18578]= -1610142873;
assign addr[18579]= -1707199606;
assign addr[18580]= -1795596234;
assign addr[18581]= -1874884346;
assign addr[18582]= -1944661739;
assign addr[18583]= -2004574453;
assign addr[18584]= -2054318569;
assign addr[18585]= -2093641749;
assign addr[18586]= -2122344521;
assign addr[18587]= -2140281282;
assign addr[18588]= -2147361045;
assign addr[18589]= -2143547897;
assign addr[18590]= -2128861181;
assign addr[18591]= -2103375398;
assign addr[18592]= -2067219829;
assign addr[18593]= -2020577882;
assign addr[18594]= -1963686155;
assign addr[18595]= -1896833245;
assign addr[18596]= -1820358275;
assign addr[18597]= -1734649179;
assign addr[18598]= -1640140734;
assign addr[18599]= -1537312353;
assign addr[18600]= -1426685652;
assign addr[18601]= -1308821808;
assign addr[18602]= -1184318708;
assign addr[18603]= -1053807919;
assign addr[18604]= -917951481;
assign addr[18605]= -777438554;
assign addr[18606]= -632981917;
assign addr[18607]= -485314355;
assign addr[18608]= -335184940;
assign addr[18609]= -183355234;
assign addr[18610]= -30595422;
assign addr[18611]= 122319591;
assign addr[18612]= 274614114;
assign addr[18613]= 425515602;
assign addr[18614]= 574258580;
assign addr[18615]= 720088517;
assign addr[18616]= 862265664;
assign addr[18617]= 1000068799;
assign addr[18618]= 1132798888;
assign addr[18619]= 1259782632;
assign addr[18620]= 1380375881;
assign addr[18621]= 1493966902;
assign addr[18622]= 1599979481;
assign addr[18623]= 1697875851;
assign addr[18624]= 1787159411;
assign addr[18625]= 1867377253;
assign addr[18626]= 1938122457;
assign addr[18627]= 1999036154;
assign addr[18628]= 2049809346;
assign addr[18629]= 2090184478;
assign addr[18630]= 2119956737;
assign addr[18631]= 2138975100;
assign addr[18632]= 2147143090;
assign addr[18633]= 2144419275;
assign addr[18634]= 2130817471;
assign addr[18635]= 2106406677;
assign addr[18636]= 2071310720;
assign addr[18637]= 2025707632;
assign addr[18638]= 1969828744;
assign addr[18639]= 1903957513;
assign addr[18640]= 1828428082;
assign addr[18641]= 1743623590;
assign addr[18642]= 1649974225;
assign addr[18643]= 1547955041;
assign addr[18644]= 1438083551;
assign addr[18645]= 1320917099;
assign addr[18646]= 1197050035;
assign addr[18647]= 1067110699;
assign addr[18648]= 931758235;
assign addr[18649]= 791679244;
assign addr[18650]= 647584304;
assign addr[18651]= 500204365;
assign addr[18652]= 350287041;
assign addr[18653]= 198592817;
assign addr[18654]= 45891193;
assign addr[18655]= -107043224;
assign addr[18656]= -259434643;
assign addr[18657]= -410510029;
assign addr[18658]= -559503022;
assign addr[18659]= -705657826;
assign addr[18660]= -848233042;
assign addr[18661]= -986505429;
assign addr[18662]= -1119773573;
assign addr[18663]= -1247361445;
assign addr[18664]= -1368621831;
assign addr[18665]= -1482939614;
assign addr[18666]= -1589734894;
assign addr[18667]= -1688465931;
assign addr[18668]= -1778631892;
assign addr[18669]= -1859775393;
assign addr[18670]= -1931484818;
assign addr[18671]= -1993396407;
assign addr[18672]= -2045196100;
assign addr[18673]= -2086621133;
assign addr[18674]= -2117461370;
assign addr[18675]= -2137560369;
assign addr[18676]= -2146816171;
assign addr[18677]= -2145181827;
assign addr[18678]= -2132665626;
assign addr[18679]= -2109331059;
assign addr[18680]= -2075296495;
assign addr[18681]= -2030734582;
assign addr[18682]= -1975871368;
assign addr[18683]= -1910985158;
assign addr[18684]= -1836405100;
assign addr[18685]= -1752509516;
assign addr[18686]= -1659723983;
assign addr[18687]= -1558519173;
assign addr[18688]= -1449408469;
assign addr[18689]= -1332945355;
assign addr[18690]= -1209720613;
assign addr[18691]= -1080359326;
assign addr[18692]= -945517704;
assign addr[18693]= -805879757;
assign addr[18694]= -662153826;
assign addr[18695]= -515068990;
assign addr[18696]= -365371365;
assign addr[18697]= -213820322;
assign addr[18698]= -61184634;
assign addr[18699]= 91761426;
assign addr[18700]= 244242007;
assign addr[18701]= 395483624;
assign addr[18702]= 544719071;
assign addr[18703]= 691191324;
assign addr[18704]= 834157373;
assign addr[18705]= 972891995;
assign addr[18706]= 1106691431;
assign addr[18707]= 1234876957;
assign addr[18708]= 1356798326;
assign addr[18709]= 1471837070;
assign addr[18710]= 1579409630;
assign addr[18711]= 1678970324;
assign addr[18712]= 1770014111;
assign addr[18713]= 1852079154;
assign addr[18714]= 1924749160;
assign addr[18715]= 1987655498;
assign addr[18716]= 2040479063;
assign addr[18717]= 2082951896;
assign addr[18718]= 2114858546;
assign addr[18719]= 2136037160;
assign addr[18720]= 2146380306;
assign addr[18721]= 2145835515;
assign addr[18722]= 2134405552;
assign addr[18723]= 2112148396;
assign addr[18724]= 2079176953;
assign addr[18725]= 2035658475;
assign addr[18726]= 1981813720;
assign addr[18727]= 1917915825;
assign addr[18728]= 1844288924;
assign addr[18729]= 1761306505;
assign addr[18730]= 1669389513;
assign addr[18731]= 1569004214;
assign addr[18732]= 1460659832;
assign addr[18733]= 1344905966;
assign addr[18734]= 1222329801;
assign addr[18735]= 1093553126;
assign addr[18736]= 959229189;
assign addr[18737]= 820039373;
assign addr[18738]= 676689746;
assign addr[18739]= 529907477;
assign addr[18740]= 380437148;
assign addr[18741]= 229036977;
assign addr[18742]= 76474970;
assign addr[18743]= -76474970;
assign addr[18744]= -229036977;
assign addr[18745]= -380437148;
assign addr[18746]= -529907477;
assign addr[18747]= -676689746;
assign addr[18748]= -820039373;
assign addr[18749]= -959229189;
assign addr[18750]= -1093553126;
assign addr[18751]= -1222329801;
assign addr[18752]= -1344905966;
assign addr[18753]= -1460659832;
assign addr[18754]= -1569004214;
assign addr[18755]= -1669389513;
assign addr[18756]= -1761306505;
assign addr[18757]= -1844288924;
assign addr[18758]= -1917915825;
assign addr[18759]= -1981813720;
assign addr[18760]= -2035658475;
assign addr[18761]= -2079176953;
assign addr[18762]= -2112148396;
assign addr[18763]= -2134405552;
assign addr[18764]= -2145835515;
assign addr[18765]= -2146380306;
assign addr[18766]= -2136037160;
assign addr[18767]= -2114858546;
assign addr[18768]= -2082951896;
assign addr[18769]= -2040479063;
assign addr[18770]= -1987655498;
assign addr[18771]= -1924749160;
assign addr[18772]= -1852079154;
assign addr[18773]= -1770014111;
assign addr[18774]= -1678970324;
assign addr[18775]= -1579409630;
assign addr[18776]= -1471837070;
assign addr[18777]= -1356798326;
assign addr[18778]= -1234876957;
assign addr[18779]= -1106691431;
assign addr[18780]= -972891995;
assign addr[18781]= -834157373;
assign addr[18782]= -691191324;
assign addr[18783]= -544719071;
assign addr[18784]= -395483624;
assign addr[18785]= -244242007;
assign addr[18786]= -91761426;
assign addr[18787]= 61184634;
assign addr[18788]= 213820322;
assign addr[18789]= 365371365;
assign addr[18790]= 515068990;
assign addr[18791]= 662153826;
assign addr[18792]= 805879757;
assign addr[18793]= 945517704;
assign addr[18794]= 1080359326;
assign addr[18795]= 1209720613;
assign addr[18796]= 1332945355;
assign addr[18797]= 1449408469;
assign addr[18798]= 1558519173;
assign addr[18799]= 1659723983;
assign addr[18800]= 1752509516;
assign addr[18801]= 1836405100;
assign addr[18802]= 1910985158;
assign addr[18803]= 1975871368;
assign addr[18804]= 2030734582;
assign addr[18805]= 2075296495;
assign addr[18806]= 2109331059;
assign addr[18807]= 2132665626;
assign addr[18808]= 2145181827;
assign addr[18809]= 2146816171;
assign addr[18810]= 2137560369;
assign addr[18811]= 2117461370;
assign addr[18812]= 2086621133;
assign addr[18813]= 2045196100;
assign addr[18814]= 1993396407;
assign addr[18815]= 1931484818;
assign addr[18816]= 1859775393;
assign addr[18817]= 1778631892;
assign addr[18818]= 1688465931;
assign addr[18819]= 1589734894;
assign addr[18820]= 1482939614;
assign addr[18821]= 1368621831;
assign addr[18822]= 1247361445;
assign addr[18823]= 1119773573;
assign addr[18824]= 986505429;
assign addr[18825]= 848233042;
assign addr[18826]= 705657826;
assign addr[18827]= 559503022;
assign addr[18828]= 410510029;
assign addr[18829]= 259434643;
assign addr[18830]= 107043224;
assign addr[18831]= -45891193;
assign addr[18832]= -198592817;
assign addr[18833]= -350287041;
assign addr[18834]= -500204365;
assign addr[18835]= -647584304;
assign addr[18836]= -791679244;
assign addr[18837]= -931758235;
assign addr[18838]= -1067110699;
assign addr[18839]= -1197050035;
assign addr[18840]= -1320917099;
assign addr[18841]= -1438083551;
assign addr[18842]= -1547955041;
assign addr[18843]= -1649974225;
assign addr[18844]= -1743623590;
assign addr[18845]= -1828428082;
assign addr[18846]= -1903957513;
assign addr[18847]= -1969828744;
assign addr[18848]= -2025707632;
assign addr[18849]= -2071310720;
assign addr[18850]= -2106406677;
assign addr[18851]= -2130817471;
assign addr[18852]= -2144419275;
assign addr[18853]= -2147143090;
assign addr[18854]= -2138975100;
assign addr[18855]= -2119956737;
assign addr[18856]= -2090184478;
assign addr[18857]= -2049809346;
assign addr[18858]= -1999036154;
assign addr[18859]= -1938122457;
assign addr[18860]= -1867377253;
assign addr[18861]= -1787159411;
assign addr[18862]= -1697875851;
assign addr[18863]= -1599979481;
assign addr[18864]= -1493966902;
assign addr[18865]= -1380375881;
assign addr[18866]= -1259782632;
assign addr[18867]= -1132798888;
assign addr[18868]= -1000068799;
assign addr[18869]= -862265664;
assign addr[18870]= -720088517;
assign addr[18871]= -574258580;
assign addr[18872]= -425515602;
assign addr[18873]= -274614114;
assign addr[18874]= -122319591;
assign addr[18875]= 30595422;
assign addr[18876]= 183355234;
assign addr[18877]= 335184940;
assign addr[18878]= 485314355;
assign addr[18879]= 632981917;
assign addr[18880]= 777438554;
assign addr[18881]= 917951481;
assign addr[18882]= 1053807919;
assign addr[18883]= 1184318708;
assign addr[18884]= 1308821808;
assign addr[18885]= 1426685652;
assign addr[18886]= 1537312353;
assign addr[18887]= 1640140734;
assign addr[18888]= 1734649179;
assign addr[18889]= 1820358275;
assign addr[18890]= 1896833245;
assign addr[18891]= 1963686155;
assign addr[18892]= 2020577882;
assign addr[18893]= 2067219829;
assign addr[18894]= 2103375398;
assign addr[18895]= 2128861181;
assign addr[18896]= 2143547897;
assign addr[18897]= 2147361045;
assign addr[18898]= 2140281282;
assign addr[18899]= 2122344521;
assign addr[18900]= 2093641749;
assign addr[18901]= 2054318569;
assign addr[18902]= 2004574453;
assign addr[18903]= 1944661739;
assign addr[18904]= 1874884346;
assign addr[18905]= 1795596234;
assign addr[18906]= 1707199606;
assign addr[18907]= 1610142873;
assign addr[18908]= 1504918373;
assign addr[18909]= 1392059879;
assign addr[18910]= 1272139887;
assign addr[18911]= 1145766716;
assign addr[18912]= 1013581418;
assign addr[18913]= 876254528;
assign addr[18914]= 734482665;
assign addr[18915]= 588984994;
assign addr[18916]= 440499581;
assign addr[18917]= 289779648;
assign addr[18918]= 137589750;
assign addr[18919]= -15298099;
assign addr[18920]= -168108346;
assign addr[18921]= -320065829;
assign addr[18922]= -470399716;
assign addr[18923]= -618347408;
assign addr[18924]= -763158411;
assign addr[18925]= -904098143;
assign addr[18926]= -1040451659;
assign addr[18927]= -1171527280;
assign addr[18928]= -1296660098;
assign addr[18929]= -1415215352;
assign addr[18930]= -1526591649;
assign addr[18931]= -1630224009;
assign addr[18932]= -1725586737;
assign addr[18933]= -1812196087;
assign addr[18934]= -1889612716;
assign addr[18935]= -1957443913;
assign addr[18936]= -2015345591;
assign addr[18937]= -2063024031;
assign addr[18938]= -2100237377;
assign addr[18939]= -2126796855;
assign addr[18940]= -2142567738;
assign addr[18941]= -2147470025;
assign addr[18942]= -2141478848;
assign addr[18943]= -2124624598;
assign addr[18944]= -2096992772;
assign addr[18945]= -2058723538;
assign addr[18946]= -2010011024;
assign addr[18947]= -1951102334;
assign addr[18948]= -1882296293;
assign addr[18949]= -1803941934;
assign addr[18950]= -1716436725;
assign addr[18951]= -1620224553;
assign addr[18952]= -1515793473;
assign addr[18953]= -1403673233;
assign addr[18954]= -1284432584;
assign addr[18955]= -1158676398;
assign addr[18956]= -1027042599;
assign addr[18957]= -890198924;
assign addr[18958]= -748839539;
assign addr[18959]= -603681519;
assign addr[18960]= -455461206;
assign addr[18961]= -304930476;
assign addr[18962]= -152852926;
assign addr[18963]= 0;
assign addr[18964]= 152852926;
assign addr[18965]= 304930476;
assign addr[18966]= 455461206;
assign addr[18967]= 603681519;
assign addr[18968]= 748839539;
assign addr[18969]= 890198924;
assign addr[18970]= 1027042599;
assign addr[18971]= 1158676398;
assign addr[18972]= 1284432584;
assign addr[18973]= 1403673233;
assign addr[18974]= 1515793473;
assign addr[18975]= 1620224553;
assign addr[18976]= 1716436725;
assign addr[18977]= 1803941934;
assign addr[18978]= 1882296293;
assign addr[18979]= 1951102334;
assign addr[18980]= 2010011024;
assign addr[18981]= 2058723538;
assign addr[18982]= 2096992772;
assign addr[18983]= 2124624598;
assign addr[18984]= 2141478848;
assign addr[18985]= 2147470025;
assign addr[18986]= 2142567738;
assign addr[18987]= 2126796855;
assign addr[18988]= 2100237377;
assign addr[18989]= 2063024031;
assign addr[18990]= 2015345591;
assign addr[18991]= 1957443913;
assign addr[18992]= 1889612716;
assign addr[18993]= 1812196087;
assign addr[18994]= 1725586737;
assign addr[18995]= 1630224009;
assign addr[18996]= 1526591649;
assign addr[18997]= 1415215352;
assign addr[18998]= 1296660098;
assign addr[18999]= 1171527280;
assign addr[19000]= 1040451659;
assign addr[19001]= 904098143;
assign addr[19002]= 763158411;
assign addr[19003]= 618347408;
assign addr[19004]= 470399716;
assign addr[19005]= 320065829;
assign addr[19006]= 168108346;
assign addr[19007]= 15298099;
assign addr[19008]= -137589750;
assign addr[19009]= -289779648;
assign addr[19010]= -440499581;
assign addr[19011]= -588984994;
assign addr[19012]= -734482665;
assign addr[19013]= -876254528;
assign addr[19014]= -1013581418;
assign addr[19015]= -1145766716;
assign addr[19016]= -1272139887;
assign addr[19017]= -1392059879;
assign addr[19018]= -1504918373;
assign addr[19019]= -1610142873;
assign addr[19020]= -1707199606;
assign addr[19021]= -1795596234;
assign addr[19022]= -1874884346;
assign addr[19023]= -1944661739;
assign addr[19024]= -2004574453;
assign addr[19025]= -2054318569;
assign addr[19026]= -2093641749;
assign addr[19027]= -2122344521;
assign addr[19028]= -2140281282;
assign addr[19029]= -2147361045;
assign addr[19030]= -2143547897;
assign addr[19031]= -2128861181;
assign addr[19032]= -2103375398;
assign addr[19033]= -2067219829;
assign addr[19034]= -2020577882;
assign addr[19035]= -1963686155;
assign addr[19036]= -1896833245;
assign addr[19037]= -1820358275;
assign addr[19038]= -1734649179;
assign addr[19039]= -1640140734;
assign addr[19040]= -1537312353;
assign addr[19041]= -1426685652;
assign addr[19042]= -1308821808;
assign addr[19043]= -1184318708;
assign addr[19044]= -1053807919;
assign addr[19045]= -917951481;
assign addr[19046]= -777438554;
assign addr[19047]= -632981917;
assign addr[19048]= -485314355;
assign addr[19049]= -335184940;
assign addr[19050]= -183355234;
assign addr[19051]= -30595422;
assign addr[19052]= 122319591;
assign addr[19053]= 274614114;
assign addr[19054]= 425515602;
assign addr[19055]= 574258580;
assign addr[19056]= 720088517;
assign addr[19057]= 862265664;
assign addr[19058]= 1000068799;
assign addr[19059]= 1132798888;
assign addr[19060]= 1259782632;
assign addr[19061]= 1380375881;
assign addr[19062]= 1493966902;
assign addr[19063]= 1599979481;
assign addr[19064]= 1697875851;
assign addr[19065]= 1787159411;
assign addr[19066]= 1867377253;
assign addr[19067]= 1938122457;
assign addr[19068]= 1999036154;
assign addr[19069]= 2049809346;
assign addr[19070]= 2090184478;
assign addr[19071]= 2119956737;
assign addr[19072]= 2138975100;
assign addr[19073]= 2147143090;
assign addr[19074]= 2144419275;
assign addr[19075]= 2130817471;
assign addr[19076]= 2106406677;
assign addr[19077]= 2071310720;
assign addr[19078]= 2025707632;
assign addr[19079]= 1969828744;
assign addr[19080]= 1903957513;
assign addr[19081]= 1828428082;
assign addr[19082]= 1743623590;
assign addr[19083]= 1649974225;
assign addr[19084]= 1547955041;
assign addr[19085]= 1438083551;
assign addr[19086]= 1320917099;
assign addr[19087]= 1197050035;
assign addr[19088]= 1067110699;
assign addr[19089]= 931758235;
assign addr[19090]= 791679244;
assign addr[19091]= 647584304;
assign addr[19092]= 500204365;
assign addr[19093]= 350287041;
assign addr[19094]= 198592817;
assign addr[19095]= 45891193;
assign addr[19096]= -107043224;
assign addr[19097]= -259434643;
assign addr[19098]= -410510029;
assign addr[19099]= -559503022;
assign addr[19100]= -705657826;
assign addr[19101]= -848233042;
assign addr[19102]= -986505429;
assign addr[19103]= -1119773573;
assign addr[19104]= -1247361445;
assign addr[19105]= -1368621831;
assign addr[19106]= -1482939614;
assign addr[19107]= -1589734894;
assign addr[19108]= -1688465931;
assign addr[19109]= -1778631892;
assign addr[19110]= -1859775393;
assign addr[19111]= -1931484818;
assign addr[19112]= -1993396407;
assign addr[19113]= -2045196100;
assign addr[19114]= -2086621133;
assign addr[19115]= -2117461370;
assign addr[19116]= -2137560369;
assign addr[19117]= -2146816171;
assign addr[19118]= -2145181827;
assign addr[19119]= -2132665626;
assign addr[19120]= -2109331059;
assign addr[19121]= -2075296495;
assign addr[19122]= -2030734582;
assign addr[19123]= -1975871368;
assign addr[19124]= -1910985158;
assign addr[19125]= -1836405100;
assign addr[19126]= -1752509516;
assign addr[19127]= -1659723983;
assign addr[19128]= -1558519173;
assign addr[19129]= -1449408469;
assign addr[19130]= -1332945355;
assign addr[19131]= -1209720613;
assign addr[19132]= -1080359326;
assign addr[19133]= -945517704;
assign addr[19134]= -805879757;
assign addr[19135]= -662153826;
assign addr[19136]= -515068990;
assign addr[19137]= -365371365;
assign addr[19138]= -213820322;
assign addr[19139]= -61184634;
assign addr[19140]= 91761426;
assign addr[19141]= 244242007;
assign addr[19142]= 395483624;
assign addr[19143]= 544719071;
assign addr[19144]= 691191324;
assign addr[19145]= 834157373;
assign addr[19146]= 972891995;
assign addr[19147]= 1106691431;
assign addr[19148]= 1234876957;
assign addr[19149]= 1356798326;
assign addr[19150]= 1471837070;
assign addr[19151]= 1579409630;
assign addr[19152]= 1678970324;
assign addr[19153]= 1770014111;
assign addr[19154]= 1852079154;
assign addr[19155]= 1924749160;
assign addr[19156]= 1987655498;
assign addr[19157]= 2040479063;
assign addr[19158]= 2082951896;
assign addr[19159]= 2114858546;
assign addr[19160]= 2136037160;
assign addr[19161]= 2146380306;
assign addr[19162]= 2145835515;
assign addr[19163]= 2134405552;
assign addr[19164]= 2112148396;
assign addr[19165]= 2079176953;
assign addr[19166]= 2035658475;
assign addr[19167]= 1981813720;
assign addr[19168]= 1917915825;
assign addr[19169]= 1844288924;
assign addr[19170]= 1761306505;
assign addr[19171]= 1669389513;
assign addr[19172]= 1569004214;
assign addr[19173]= 1460659832;
assign addr[19174]= 1344905966;
assign addr[19175]= 1222329801;
assign addr[19176]= 1093553126;
assign addr[19177]= 959229189;
assign addr[19178]= 820039373;
assign addr[19179]= 676689746;
assign addr[19180]= 529907477;
assign addr[19181]= 380437148;
assign addr[19182]= 229036977;
assign addr[19183]= 76474970;
assign addr[19184]= -76474970;
assign addr[19185]= -229036977;
assign addr[19186]= -380437148;
assign addr[19187]= -529907477;
assign addr[19188]= -676689746;
assign addr[19189]= -820039373;
assign addr[19190]= -959229189;
assign addr[19191]= -1093553126;
assign addr[19192]= -1222329801;
assign addr[19193]= -1344905966;
assign addr[19194]= -1460659832;
assign addr[19195]= -1569004214;
assign addr[19196]= -1669389513;
assign addr[19197]= -1761306505;
assign addr[19198]= -1844288924;
assign addr[19199]= -1917915825;
assign addr[19200]= -1981813720;
assign addr[19201]= -2035658475;
assign addr[19202]= -2079176953;
assign addr[19203]= -2112148396;
assign addr[19204]= -2134405552;
assign addr[19205]= -2145835515;
assign addr[19206]= -2146380306;
assign addr[19207]= -2136037160;
assign addr[19208]= -2114858546;
assign addr[19209]= -2082951896;
assign addr[19210]= -2040479063;
assign addr[19211]= -1987655498;
assign addr[19212]= -1924749160;
assign addr[19213]= -1852079154;
assign addr[19214]= -1770014111;
assign addr[19215]= -1678970324;
assign addr[19216]= -1579409630;
assign addr[19217]= -1471837070;
assign addr[19218]= -1356798326;
assign addr[19219]= -1234876957;
assign addr[19220]= -1106691431;
assign addr[19221]= -972891995;
assign addr[19222]= -834157373;
assign addr[19223]= -691191324;
assign addr[19224]= -544719071;
assign addr[19225]= -395483624;
assign addr[19226]= -244242007;
assign addr[19227]= -91761426;
assign addr[19228]= 61184634;
assign addr[19229]= 213820322;
assign addr[19230]= 365371365;
assign addr[19231]= 515068990;
assign addr[19232]= 662153826;
assign addr[19233]= 805879757;
assign addr[19234]= 945517704;
assign addr[19235]= 1080359326;
assign addr[19236]= 1209720613;
assign addr[19237]= 1332945355;
assign addr[19238]= 1449408469;
assign addr[19239]= 1558519173;
assign addr[19240]= 1659723983;
assign addr[19241]= 1752509516;
assign addr[19242]= 1836405100;
assign addr[19243]= 1910985158;
assign addr[19244]= 1975871368;
assign addr[19245]= 2030734582;
assign addr[19246]= 2075296495;
assign addr[19247]= 2109331059;
assign addr[19248]= 2132665626;
assign addr[19249]= 2145181827;
assign addr[19250]= 2146816171;
assign addr[19251]= 2137560369;
assign addr[19252]= 2117461370;
assign addr[19253]= 2086621133;
assign addr[19254]= 2045196100;
assign addr[19255]= 1993396407;
assign addr[19256]= 1931484818;
assign addr[19257]= 1859775393;
assign addr[19258]= 1778631892;
assign addr[19259]= 1688465931;
assign addr[19260]= 1589734894;
assign addr[19261]= 1482939614;
assign addr[19262]= 1368621831;
assign addr[19263]= 1247361445;
assign addr[19264]= 1119773573;
assign addr[19265]= 986505429;
assign addr[19266]= 848233042;
assign addr[19267]= 705657826;
assign addr[19268]= 559503022;
assign addr[19269]= 410510029;
assign addr[19270]= 259434643;
assign addr[19271]= 107043224;
assign addr[19272]= -45891193;
assign addr[19273]= -198592817;
assign addr[19274]= -350287041;
assign addr[19275]= -500204365;
assign addr[19276]= -647584304;
assign addr[19277]= -791679244;
assign addr[19278]= -931758235;
assign addr[19279]= -1067110699;
assign addr[19280]= -1197050035;
assign addr[19281]= -1320917099;
assign addr[19282]= -1438083551;
assign addr[19283]= -1547955041;
assign addr[19284]= -1649974225;
assign addr[19285]= -1743623590;
assign addr[19286]= -1828428082;
assign addr[19287]= -1903957513;
assign addr[19288]= -1969828744;
assign addr[19289]= -2025707632;
assign addr[19290]= -2071310720;
assign addr[19291]= -2106406677;
assign addr[19292]= -2130817471;
assign addr[19293]= -2144419275;
assign addr[19294]= -2147143090;
assign addr[19295]= -2138975100;
assign addr[19296]= -2119956737;
assign addr[19297]= -2090184478;
assign addr[19298]= -2049809346;
assign addr[19299]= -1999036154;
assign addr[19300]= -1938122457;
assign addr[19301]= -1867377253;
assign addr[19302]= -1787159411;
assign addr[19303]= -1697875851;
assign addr[19304]= -1599979481;
assign addr[19305]= -1493966902;
assign addr[19306]= -1380375881;
assign addr[19307]= -1259782632;
assign addr[19308]= -1132798888;
assign addr[19309]= -1000068799;
assign addr[19310]= -862265664;
assign addr[19311]= -720088517;
assign addr[19312]= -574258580;
assign addr[19313]= -425515602;
assign addr[19314]= -274614114;
assign addr[19315]= -122319591;
assign addr[19316]= 30595422;
assign addr[19317]= 183355234;
assign addr[19318]= 335184940;
assign addr[19319]= 485314355;
assign addr[19320]= 632981917;
assign addr[19321]= 777438554;
assign addr[19322]= 917951481;
assign addr[19323]= 1053807919;
assign addr[19324]= 1184318708;
assign addr[19325]= 1308821808;
assign addr[19326]= 1426685652;
assign addr[19327]= 1537312353;
assign addr[19328]= 1640140734;
assign addr[19329]= 1734649179;
assign addr[19330]= 1820358275;
assign addr[19331]= 1896833245;
assign addr[19332]= 1963686155;
assign addr[19333]= 2020577882;
assign addr[19334]= 2067219829;
assign addr[19335]= 2103375398;
assign addr[19336]= 2128861181;
assign addr[19337]= 2143547897;
assign addr[19338]= 2147361045;
assign addr[19339]= 2140281282;
assign addr[19340]= 2122344521;
assign addr[19341]= 2093641749;
assign addr[19342]= 2054318569;
assign addr[19343]= 2004574453;
assign addr[19344]= 1944661739;
assign addr[19345]= 1874884346;
assign addr[19346]= 1795596234;
assign addr[19347]= 1707199606;
assign addr[19348]= 1610142873;
assign addr[19349]= 1504918373;
assign addr[19350]= 1392059879;
assign addr[19351]= 1272139887;
assign addr[19352]= 1145766716;
assign addr[19353]= 1013581418;
assign addr[19354]= 876254528;
assign addr[19355]= 734482665;
assign addr[19356]= 588984994;
assign addr[19357]= 440499581;
assign addr[19358]= 289779648;
assign addr[19359]= 137589750;
assign addr[19360]= -15298099;
assign addr[19361]= -168108346;
assign addr[19362]= -320065829;
assign addr[19363]= -470399716;
assign addr[19364]= -618347408;
assign addr[19365]= -763158411;
assign addr[19366]= -904098143;
assign addr[19367]= -1040451659;
assign addr[19368]= -1171527280;
assign addr[19369]= -1296660098;
assign addr[19370]= -1415215352;
assign addr[19371]= -1526591649;
assign addr[19372]= -1630224009;
assign addr[19373]= -1725586737;
assign addr[19374]= -1812196087;
assign addr[19375]= -1889612716;
assign addr[19376]= -1957443913;
assign addr[19377]= -2015345591;
assign addr[19378]= -2063024031;
assign addr[19379]= -2100237377;
assign addr[19380]= -2126796855;
assign addr[19381]= -2142567738;
assign addr[19382]= -2147470025;
assign addr[19383]= -2141478848;
assign addr[19384]= -2124624598;
assign addr[19385]= -2096992772;
assign addr[19386]= -2058723538;
assign addr[19387]= -2010011024;
assign addr[19388]= -1951102334;
assign addr[19389]= -1882296293;
assign addr[19390]= -1803941934;
assign addr[19391]= -1716436725;
assign addr[19392]= -1620224553;
assign addr[19393]= -1515793473;
assign addr[19394]= -1403673233;
assign addr[19395]= -1284432584;
assign addr[19396]= -1158676398;
assign addr[19397]= -1027042599;
assign addr[19398]= -890198924;
assign addr[19399]= -748839539;
assign addr[19400]= -603681519;
assign addr[19401]= -455461206;
assign addr[19402]= -304930476;
assign addr[19403]= -152852926;
assign addr[19404]= 0;
assign addr[19405]= 152852926;
assign addr[19406]= 304930476;
assign addr[19407]= 455461206;
assign addr[19408]= 603681519;
assign addr[19409]= 748839539;
assign addr[19410]= 890198924;
assign addr[19411]= 1027042599;
assign addr[19412]= 1158676398;
assign addr[19413]= 1284432584;
assign addr[19414]= 1403673233;
assign addr[19415]= 1515793473;
assign addr[19416]= 1620224553;
assign addr[19417]= 1716436725;
assign addr[19418]= 1803941934;
assign addr[19419]= 1882296293;
assign addr[19420]= 1951102334;
assign addr[19421]= 2010011024;
assign addr[19422]= 2058723538;
assign addr[19423]= 2096992772;
assign addr[19424]= 2124624598;
assign addr[19425]= 2141478848;
assign addr[19426]= 2147470025;
assign addr[19427]= 2142567738;
assign addr[19428]= 2126796855;
assign addr[19429]= 2100237377;
assign addr[19430]= 2063024031;
assign addr[19431]= 2015345591;
assign addr[19432]= 1957443913;
assign addr[19433]= 1889612716;
assign addr[19434]= 1812196087;
assign addr[19435]= 1725586737;
assign addr[19436]= 1630224009;
assign addr[19437]= 1526591649;
assign addr[19438]= 1415215352;
assign addr[19439]= 1296660098;
assign addr[19440]= 1171527280;
assign addr[19441]= 1040451659;
assign addr[19442]= 904098143;
assign addr[19443]= 763158411;
assign addr[19444]= 618347408;
assign addr[19445]= 470399716;
assign addr[19446]= 320065829;
assign addr[19447]= 168108346;
assign addr[19448]= 15298099;
assign addr[19449]= -137589750;
assign addr[19450]= -289779648;
assign addr[19451]= -440499581;
assign addr[19452]= -588984994;
assign addr[19453]= -734482665;
assign addr[19454]= -876254528;
assign addr[19455]= -1013581418;
assign addr[19456]= -1145766716;
assign addr[19457]= -1272139887;
assign addr[19458]= -1392059879;
assign addr[19459]= -1504918373;
assign addr[19460]= -1610142873;
assign addr[19461]= -1707199606;
assign addr[19462]= -1795596234;
assign addr[19463]= -1874884346;
assign addr[19464]= -1944661739;
assign addr[19465]= -2004574453;
assign addr[19466]= -2054318569;
assign addr[19467]= -2093641749;
assign addr[19468]= -2122344521;
assign addr[19469]= -2140281282;
assign addr[19470]= -2147361045;
assign addr[19471]= -2143547897;
assign addr[19472]= -2128861181;
assign addr[19473]= -2103375398;
assign addr[19474]= -2067219829;
assign addr[19475]= -2020577882;
assign addr[19476]= -1963686155;
assign addr[19477]= -1896833245;
assign addr[19478]= -1820358275;
assign addr[19479]= -1734649179;
assign addr[19480]= -1640140734;
assign addr[19481]= -1537312353;
assign addr[19482]= -1426685652;
assign addr[19483]= -1308821808;
assign addr[19484]= -1184318708;
assign addr[19485]= -1053807919;
assign addr[19486]= -917951481;
assign addr[19487]= -777438554;
assign addr[19488]= -632981917;
assign addr[19489]= -485314355;
assign addr[19490]= -335184940;
assign addr[19491]= -183355234;
assign addr[19492]= -30595422;
assign addr[19493]= 122319591;
assign addr[19494]= 274614114;
assign addr[19495]= 425515602;
assign addr[19496]= 574258580;
assign addr[19497]= 720088517;
assign addr[19498]= 862265664;
assign addr[19499]= 1000068799;
assign addr[19500]= 1132798888;
assign addr[19501]= 1259782632;
assign addr[19502]= 1380375881;
assign addr[19503]= 1493966902;
assign addr[19504]= 1599979481;
assign addr[19505]= 1697875851;
assign addr[19506]= 1787159411;
assign addr[19507]= 1867377253;
assign addr[19508]= 1938122457;
assign addr[19509]= 1999036154;
assign addr[19510]= 2049809346;
assign addr[19511]= 2090184478;
assign addr[19512]= 2119956737;
assign addr[19513]= 2138975100;
assign addr[19514]= 2147143090;
assign addr[19515]= 2144419275;
assign addr[19516]= 2130817471;
assign addr[19517]= 2106406677;
assign addr[19518]= 2071310720;
assign addr[19519]= 2025707632;
assign addr[19520]= 1969828744;
assign addr[19521]= 1903957513;
assign addr[19522]= 1828428082;
assign addr[19523]= 1743623590;
assign addr[19524]= 1649974225;
assign addr[19525]= 1547955041;
assign addr[19526]= 1438083551;
assign addr[19527]= 1320917099;
assign addr[19528]= 1197050035;
assign addr[19529]= 1067110699;
assign addr[19530]= 931758235;
assign addr[19531]= 791679244;
assign addr[19532]= 647584304;
assign addr[19533]= 500204365;
assign addr[19534]= 350287041;
assign addr[19535]= 198592817;
assign addr[19536]= 45891193;
assign addr[19537]= -107043224;
assign addr[19538]= -259434643;
assign addr[19539]= -410510029;
assign addr[19540]= -559503022;
assign addr[19541]= -705657826;
assign addr[19542]= -848233042;
assign addr[19543]= -986505429;
assign addr[19544]= -1119773573;
assign addr[19545]= -1247361445;
assign addr[19546]= -1368621831;
assign addr[19547]= -1482939614;
assign addr[19548]= -1589734894;
assign addr[19549]= -1688465931;
assign addr[19550]= -1778631892;
assign addr[19551]= -1859775393;
assign addr[19552]= -1931484818;
assign addr[19553]= -1993396407;
assign addr[19554]= -2045196100;
assign addr[19555]= -2086621133;
assign addr[19556]= -2117461370;
assign addr[19557]= -2137560369;
assign addr[19558]= -2146816171;
assign addr[19559]= -2145181827;
assign addr[19560]= -2132665626;
assign addr[19561]= -2109331059;
assign addr[19562]= -2075296495;
assign addr[19563]= -2030734582;
assign addr[19564]= -1975871368;
assign addr[19565]= -1910985158;
assign addr[19566]= -1836405100;
assign addr[19567]= -1752509516;
assign addr[19568]= -1659723983;
assign addr[19569]= -1558519173;
assign addr[19570]= -1449408469;
assign addr[19571]= -1332945355;
assign addr[19572]= -1209720613;
assign addr[19573]= -1080359326;
assign addr[19574]= -945517704;
assign addr[19575]= -805879757;
assign addr[19576]= -662153826;
assign addr[19577]= -515068990;
assign addr[19578]= -365371365;
assign addr[19579]= -213820322;
assign addr[19580]= -61184634;
assign addr[19581]= 91761426;
assign addr[19582]= 244242007;
assign addr[19583]= 395483624;
assign addr[19584]= 544719071;
assign addr[19585]= 691191324;
assign addr[19586]= 834157373;
assign addr[19587]= 972891995;
assign addr[19588]= 1106691431;
assign addr[19589]= 1234876957;
assign addr[19590]= 1356798326;
assign addr[19591]= 1471837070;
assign addr[19592]= 1579409630;
assign addr[19593]= 1678970324;
assign addr[19594]= 1770014111;
assign addr[19595]= 1852079154;
assign addr[19596]= 1924749160;
assign addr[19597]= 1987655498;
assign addr[19598]= 2040479063;
assign addr[19599]= 2082951896;
assign addr[19600]= 2114858546;
assign addr[19601]= 2136037160;
assign addr[19602]= 2146380306;
assign addr[19603]= 2145835515;
assign addr[19604]= 2134405552;
assign addr[19605]= 2112148396;
assign addr[19606]= 2079176953;
assign addr[19607]= 2035658475;
assign addr[19608]= 1981813720;
assign addr[19609]= 1917915825;
assign addr[19610]= 1844288924;
assign addr[19611]= 1761306505;
assign addr[19612]= 1669389513;
assign addr[19613]= 1569004214;
assign addr[19614]= 1460659832;
assign addr[19615]= 1344905966;
assign addr[19616]= 1222329801;
assign addr[19617]= 1093553126;
assign addr[19618]= 959229189;
assign addr[19619]= 820039373;
assign addr[19620]= 676689746;
assign addr[19621]= 529907477;
assign addr[19622]= 380437148;
assign addr[19623]= 229036977;
assign addr[19624]= 76474970;
assign addr[19625]= -76474970;
assign addr[19626]= -229036977;
assign addr[19627]= -380437148;
assign addr[19628]= -529907477;
assign addr[19629]= -676689746;
assign addr[19630]= -820039373;
assign addr[19631]= -959229189;
assign addr[19632]= -1093553126;
assign addr[19633]= -1222329801;
assign addr[19634]= -1344905966;
assign addr[19635]= -1460659832;
assign addr[19636]= -1569004214;
assign addr[19637]= -1669389513;
assign addr[19638]= -1761306505;
assign addr[19639]= -1844288924;
assign addr[19640]= -1917915825;
assign addr[19641]= -1981813720;
assign addr[19642]= -2035658475;
assign addr[19643]= -2079176953;
assign addr[19644]= -2112148396;
assign addr[19645]= -2134405552;
assign addr[19646]= -2145835515;
assign addr[19647]= -2146380306;
assign addr[19648]= -2136037160;
assign addr[19649]= -2114858546;
assign addr[19650]= -2082951896;
assign addr[19651]= -2040479063;
assign addr[19652]= -1987655498;
assign addr[19653]= -1924749160;
assign addr[19654]= -1852079154;
assign addr[19655]= -1770014111;
assign addr[19656]= -1678970324;
assign addr[19657]= -1579409630;
assign addr[19658]= -1471837070;
assign addr[19659]= -1356798326;
assign addr[19660]= -1234876957;
assign addr[19661]= -1106691431;
assign addr[19662]= -972891995;
assign addr[19663]= -834157373;
assign addr[19664]= -691191324;
assign addr[19665]= -544719071;
assign addr[19666]= -395483624;
assign addr[19667]= -244242007;
assign addr[19668]= -91761426;
assign addr[19669]= 61184634;
assign addr[19670]= 213820322;
assign addr[19671]= 365371365;
assign addr[19672]= 515068990;
assign addr[19673]= 662153826;
assign addr[19674]= 805879757;
assign addr[19675]= 945517704;
assign addr[19676]= 1080359326;
assign addr[19677]= 1209720613;
assign addr[19678]= 1332945355;
assign addr[19679]= 1449408469;
assign addr[19680]= 1558519173;
assign addr[19681]= 1659723983;
assign addr[19682]= 1752509516;
assign addr[19683]= 1836405100;
assign addr[19684]= 1910985158;
assign addr[19685]= 1975871368;
assign addr[19686]= 2030734582;
assign addr[19687]= 2075296495;
assign addr[19688]= 2109331059;
assign addr[19689]= 2132665626;
assign addr[19690]= 2145181827;
assign addr[19691]= 2146816171;
assign addr[19692]= 2137560369;
assign addr[19693]= 2117461370;
assign addr[19694]= 2086621133;
assign addr[19695]= 2045196100;
assign addr[19696]= 1993396407;
assign addr[19697]= 1931484818;
assign addr[19698]= 1859775393;
assign addr[19699]= 1778631892;
assign addr[19700]= 1688465931;
assign addr[19701]= 1589734894;
assign addr[19702]= 1482939614;
assign addr[19703]= 1368621831;
assign addr[19704]= 1247361445;
assign addr[19705]= 1119773573;
assign addr[19706]= 986505429;
assign addr[19707]= 848233042;
assign addr[19708]= 705657826;
assign addr[19709]= 559503022;
assign addr[19710]= 410510029;
assign addr[19711]= 259434643;
assign addr[19712]= 107043224;
assign addr[19713]= -45891193;
assign addr[19714]= -198592817;
assign addr[19715]= -350287041;
assign addr[19716]= -500204365;
assign addr[19717]= -647584304;
assign addr[19718]= -791679244;
assign addr[19719]= -931758235;
assign addr[19720]= -1067110699;
assign addr[19721]= -1197050035;
assign addr[19722]= -1320917099;
assign addr[19723]= -1438083551;
assign addr[19724]= -1547955041;
assign addr[19725]= -1649974225;
assign addr[19726]= -1743623590;
assign addr[19727]= -1828428082;
assign addr[19728]= -1903957513;
assign addr[19729]= -1969828744;
assign addr[19730]= -2025707632;
assign addr[19731]= -2071310720;
assign addr[19732]= -2106406677;
assign addr[19733]= -2130817471;
assign addr[19734]= -2144419275;
assign addr[19735]= -2147143090;
assign addr[19736]= -2138975100;
assign addr[19737]= -2119956737;
assign addr[19738]= -2090184478;
assign addr[19739]= -2049809346;
assign addr[19740]= -1999036154;
assign addr[19741]= -1938122457;
assign addr[19742]= -1867377253;
assign addr[19743]= -1787159411;
assign addr[19744]= -1697875851;
assign addr[19745]= -1599979481;
assign addr[19746]= -1493966902;
assign addr[19747]= -1380375881;
assign addr[19748]= -1259782632;
assign addr[19749]= -1132798888;
assign addr[19750]= -1000068799;
assign addr[19751]= -862265664;
assign addr[19752]= -720088517;
assign addr[19753]= -574258580;
assign addr[19754]= -425515602;
assign addr[19755]= -274614114;
assign addr[19756]= -122319591;
assign addr[19757]= 30595422;
assign addr[19758]= 183355234;
assign addr[19759]= 335184940;
assign addr[19760]= 485314355;
assign addr[19761]= 632981917;
assign addr[19762]= 777438554;
assign addr[19763]= 917951481;
assign addr[19764]= 1053807919;
assign addr[19765]= 1184318708;
assign addr[19766]= 1308821808;
assign addr[19767]= 1426685652;
assign addr[19768]= 1537312353;
assign addr[19769]= 1640140734;
assign addr[19770]= 1734649179;
assign addr[19771]= 1820358275;
assign addr[19772]= 1896833245;
assign addr[19773]= 1963686155;
assign addr[19774]= 2020577882;
assign addr[19775]= 2067219829;
assign addr[19776]= 2103375398;
assign addr[19777]= 2128861181;
assign addr[19778]= 2143547897;
assign addr[19779]= 2147361045;
assign addr[19780]= 2140281282;
assign addr[19781]= 2122344521;
assign addr[19782]= 2093641749;
assign addr[19783]= 2054318569;
assign addr[19784]= 2004574453;
assign addr[19785]= 1944661739;
assign addr[19786]= 1874884346;
assign addr[19787]= 1795596234;
assign addr[19788]= 1707199606;
assign addr[19789]= 1610142873;
assign addr[19790]= 1504918373;
assign addr[19791]= 1392059879;
assign addr[19792]= 1272139887;
assign addr[19793]= 1145766716;
assign addr[19794]= 1013581418;
assign addr[19795]= 876254528;
assign addr[19796]= 734482665;
assign addr[19797]= 588984994;
assign addr[19798]= 440499581;
assign addr[19799]= 289779648;
assign addr[19800]= 137589750;
assign addr[19801]= -15298099;
assign addr[19802]= -168108346;
assign addr[19803]= -320065829;
assign addr[19804]= -470399716;
assign addr[19805]= -618347408;
assign addr[19806]= -763158411;
assign addr[19807]= -904098143;
assign addr[19808]= -1040451659;
assign addr[19809]= -1171527280;
assign addr[19810]= -1296660098;
assign addr[19811]= -1415215352;
assign addr[19812]= -1526591649;
assign addr[19813]= -1630224009;
assign addr[19814]= -1725586737;
assign addr[19815]= -1812196087;
assign addr[19816]= -1889612716;
assign addr[19817]= -1957443913;
assign addr[19818]= -2015345591;
assign addr[19819]= -2063024031;
assign addr[19820]= -2100237377;
assign addr[19821]= -2126796855;
assign addr[19822]= -2142567738;
assign addr[19823]= -2147470025;
assign addr[19824]= -2141478848;
assign addr[19825]= -2124624598;
assign addr[19826]= -2096992772;
assign addr[19827]= -2058723538;
assign addr[19828]= -2010011024;
assign addr[19829]= -1951102334;
assign addr[19830]= -1882296293;
assign addr[19831]= -1803941934;
assign addr[19832]= -1716436725;
assign addr[19833]= -1620224553;
assign addr[19834]= -1515793473;
assign addr[19835]= -1403673233;
assign addr[19836]= -1284432584;
assign addr[19837]= -1158676398;
assign addr[19838]= -1027042599;
assign addr[19839]= -890198924;
assign addr[19840]= -748839539;
assign addr[19841]= -603681519;
assign addr[19842]= -455461206;
assign addr[19843]= -304930476;
assign addr[19844]= -152852926;
assign addr[19845]= 0;
assign addr[19846]= 152852926;
assign addr[19847]= 304930476;
assign addr[19848]= 455461206;
assign addr[19849]= 603681519;
assign addr[19850]= 748839539;
assign addr[19851]= 890198924;
assign addr[19852]= 1027042599;
assign addr[19853]= 1158676398;
assign addr[19854]= 1284432584;
assign addr[19855]= 1403673233;
assign addr[19856]= 1515793473;
assign addr[19857]= 1620224553;
assign addr[19858]= 1716436725;
assign addr[19859]= 1803941934;
assign addr[19860]= 1882296293;
assign addr[19861]= 1951102334;
assign addr[19862]= 2010011024;
assign addr[19863]= 2058723538;
assign addr[19864]= 2096992772;
assign addr[19865]= 2124624598;
assign addr[19866]= 2141478848;
assign addr[19867]= 2147470025;
assign addr[19868]= 2142567738;
assign addr[19869]= 2126796855;
assign addr[19870]= 2100237377;
assign addr[19871]= 2063024031;
assign addr[19872]= 2015345591;
assign addr[19873]= 1957443913;
assign addr[19874]= 1889612716;
assign addr[19875]= 1812196087;
assign addr[19876]= 1725586737;
assign addr[19877]= 1630224009;
assign addr[19878]= 1526591649;
assign addr[19879]= 1415215352;
assign addr[19880]= 1296660098;
assign addr[19881]= 1171527280;
assign addr[19882]= 1040451659;
assign addr[19883]= 904098143;
assign addr[19884]= 763158411;
assign addr[19885]= 618347408;
assign addr[19886]= 470399716;
assign addr[19887]= 320065829;
assign addr[19888]= 168108346;
assign addr[19889]= 15298099;
assign addr[19890]= -137589750;
assign addr[19891]= -289779648;
assign addr[19892]= -440499581;
assign addr[19893]= -588984994;
assign addr[19894]= -734482665;
assign addr[19895]= -876254528;
assign addr[19896]= -1013581418;
assign addr[19897]= -1145766716;
assign addr[19898]= -1272139887;
assign addr[19899]= -1392059879;
assign addr[19900]= -1504918373;
assign addr[19901]= -1610142873;
assign addr[19902]= -1707199606;
assign addr[19903]= -1795596234;
assign addr[19904]= -1874884346;
assign addr[19905]= -1944661739;
assign addr[19906]= -2004574453;
assign addr[19907]= -2054318569;
assign addr[19908]= -2093641749;
assign addr[19909]= -2122344521;
assign addr[19910]= -2140281282;
assign addr[19911]= -2147361045;
assign addr[19912]= -2143547897;
assign addr[19913]= -2128861181;
assign addr[19914]= -2103375398;
assign addr[19915]= -2067219829;
assign addr[19916]= -2020577882;
assign addr[19917]= -1963686155;
assign addr[19918]= -1896833245;
assign addr[19919]= -1820358275;
assign addr[19920]= -1734649179;
assign addr[19921]= -1640140734;
assign addr[19922]= -1537312353;
assign addr[19923]= -1426685652;
assign addr[19924]= -1308821808;
assign addr[19925]= -1184318708;
assign addr[19926]= -1053807919;
assign addr[19927]= -917951481;
assign addr[19928]= -777438554;
assign addr[19929]= -632981917;
assign addr[19930]= -485314355;
assign addr[19931]= -335184940;
assign addr[19932]= -183355234;
assign addr[19933]= -30595422;
assign addr[19934]= 122319591;
assign addr[19935]= 274614114;
assign addr[19936]= 425515602;
assign addr[19937]= 574258580;
assign addr[19938]= 720088517;
assign addr[19939]= 862265664;
assign addr[19940]= 1000068799;
assign addr[19941]= 1132798888;
assign addr[19942]= 1259782632;
assign addr[19943]= 1380375881;
assign addr[19944]= 1493966902;
assign addr[19945]= 1599979481;
assign addr[19946]= 1697875851;
assign addr[19947]= 1787159411;
assign addr[19948]= 1867377253;
assign addr[19949]= 1938122457;
assign addr[19950]= 1999036154;
assign addr[19951]= 2049809346;
assign addr[19952]= 2090184478;
assign addr[19953]= 2119956737;
assign addr[19954]= 2138975100;
assign addr[19955]= 2147143090;
assign addr[19956]= 2144419275;
assign addr[19957]= 2130817471;
assign addr[19958]= 2106406677;
assign addr[19959]= 2071310720;
assign addr[19960]= 2025707632;
assign addr[19961]= 1969828744;
assign addr[19962]= 1903957513;
assign addr[19963]= 1828428082;
assign addr[19964]= 1743623590;
assign addr[19965]= 1649974225;
assign addr[19966]= 1547955041;
assign addr[19967]= 1438083551;
assign addr[19968]= 1320917099;
assign addr[19969]= 1197050035;
assign addr[19970]= 1067110699;
assign addr[19971]= 931758235;
assign addr[19972]= 791679244;
assign addr[19973]= 647584304;
assign addr[19974]= 500204365;
assign addr[19975]= 350287041;
assign addr[19976]= 198592817;
assign addr[19977]= 45891193;
assign addr[19978]= -107043224;
assign addr[19979]= -259434643;
assign addr[19980]= -410510029;
assign addr[19981]= -559503022;
assign addr[19982]= -705657826;
assign addr[19983]= -848233042;
assign addr[19984]= -986505429;
assign addr[19985]= -1119773573;
assign addr[19986]= -1247361445;
assign addr[19987]= -1368621831;
assign addr[19988]= -1482939614;
assign addr[19989]= -1589734894;
assign addr[19990]= -1688465931;
assign addr[19991]= -1778631892;
assign addr[19992]= -1859775393;
assign addr[19993]= -1931484818;
assign addr[19994]= -1993396407;
assign addr[19995]= -2045196100;
assign addr[19996]= -2086621133;
assign addr[19997]= -2117461370;
assign addr[19998]= -2137560369;
assign addr[19999]= -2146816171;
assign addr[20000]= -2145181827;
assign addr[20001]= -2132665626;
assign addr[20002]= -2109331059;
assign addr[20003]= -2075296495;
assign addr[20004]= -2030734582;
assign addr[20005]= -1975871368;
assign addr[20006]= -1910985158;
assign addr[20007]= -1836405100;
assign addr[20008]= -1752509516;
assign addr[20009]= -1659723983;
assign addr[20010]= -1558519173;
assign addr[20011]= -1449408469;
assign addr[20012]= -1332945355;
assign addr[20013]= -1209720613;
assign addr[20014]= -1080359326;
assign addr[20015]= -945517704;
assign addr[20016]= -805879757;
assign addr[20017]= -662153826;
assign addr[20018]= -515068990;
assign addr[20019]= -365371365;
assign addr[20020]= -213820322;
assign addr[20021]= -61184634;
assign addr[20022]= 91761426;
assign addr[20023]= 244242007;
assign addr[20024]= 395483624;
assign addr[20025]= 544719071;
assign addr[20026]= 691191324;
assign addr[20027]= 834157373;
assign addr[20028]= 972891995;
assign addr[20029]= 1106691431;
assign addr[20030]= 1234876957;
assign addr[20031]= 1356798326;
assign addr[20032]= 1471837070;
assign addr[20033]= 1579409630;
assign addr[20034]= 1678970324;
assign addr[20035]= 1770014111;
assign addr[20036]= 1852079154;
assign addr[20037]= 1924749160;
assign addr[20038]= 1987655498;
assign addr[20039]= 2040479063;
assign addr[20040]= 2082951896;
assign addr[20041]= 2114858546;
assign addr[20042]= 2136037160;
assign addr[20043]= 2146380306;
assign addr[20044]= 2145835515;
assign addr[20045]= 2134405552;
assign addr[20046]= 2112148396;
assign addr[20047]= 2079176953;
assign addr[20048]= 2035658475;
assign addr[20049]= 1981813720;
assign addr[20050]= 1917915825;
assign addr[20051]= 1844288924;
assign addr[20052]= 1761306505;
assign addr[20053]= 1669389513;
assign addr[20054]= 1569004214;
assign addr[20055]= 1460659832;
assign addr[20056]= 1344905966;
assign addr[20057]= 1222329801;
assign addr[20058]= 1093553126;
assign addr[20059]= 959229189;
assign addr[20060]= 820039373;
assign addr[20061]= 676689746;
assign addr[20062]= 529907477;
assign addr[20063]= 380437148;
assign addr[20064]= 229036977;
assign addr[20065]= 76474970;
assign addr[20066]= -76474970;
assign addr[20067]= -229036977;
assign addr[20068]= -380437148;
assign addr[20069]= -529907477;
assign addr[20070]= -676689746;
assign addr[20071]= -820039373;
assign addr[20072]= -959229189;
assign addr[20073]= -1093553126;
assign addr[20074]= -1222329801;
assign addr[20075]= -1344905966;
assign addr[20076]= -1460659832;
assign addr[20077]= -1569004214;
assign addr[20078]= -1669389513;
assign addr[20079]= -1761306505;
assign addr[20080]= -1844288924;
assign addr[20081]= -1917915825;
assign addr[20082]= -1981813720;
assign addr[20083]= -2035658475;
assign addr[20084]= -2079176953;
assign addr[20085]= -2112148396;
assign addr[20086]= -2134405552;
assign addr[20087]= -2145835515;
assign addr[20088]= -2146380306;
assign addr[20089]= -2136037160;
assign addr[20090]= -2114858546;
assign addr[20091]= -2082951896;
assign addr[20092]= -2040479063;
assign addr[20093]= -1987655498;
assign addr[20094]= -1924749160;
assign addr[20095]= -1852079154;
assign addr[20096]= -1770014111;
assign addr[20097]= -1678970324;
assign addr[20098]= -1579409630;
assign addr[20099]= -1471837070;
assign addr[20100]= -1356798326;
assign addr[20101]= -1234876957;
assign addr[20102]= -1106691431;
assign addr[20103]= -972891995;
assign addr[20104]= -834157373;
assign addr[20105]= -691191324;
assign addr[20106]= -544719071;
assign addr[20107]= -395483624;
assign addr[20108]= -244242007;
assign addr[20109]= -91761426;
assign addr[20110]= 61184634;
assign addr[20111]= 213820322;
assign addr[20112]= 365371365;
assign addr[20113]= 515068990;
assign addr[20114]= 662153826;
assign addr[20115]= 805879757;
assign addr[20116]= 945517704;
assign addr[20117]= 1080359326;
assign addr[20118]= 1209720613;
assign addr[20119]= 1332945355;
assign addr[20120]= 1449408469;
assign addr[20121]= 1558519173;
assign addr[20122]= 1659723983;
assign addr[20123]= 1752509516;
assign addr[20124]= 1836405100;
assign addr[20125]= 1910985158;
assign addr[20126]= 1975871368;
assign addr[20127]= 2030734582;
assign addr[20128]= 2075296495;
assign addr[20129]= 2109331059;
assign addr[20130]= 2132665626;
assign addr[20131]= 2145181827;
assign addr[20132]= 2146816171;
assign addr[20133]= 2137560369;
assign addr[20134]= 2117461370;
assign addr[20135]= 2086621133;
assign addr[20136]= 2045196100;
assign addr[20137]= 1993396407;
assign addr[20138]= 1931484818;
assign addr[20139]= 1859775393;
assign addr[20140]= 1778631892;
assign addr[20141]= 1688465931;
assign addr[20142]= 1589734894;
assign addr[20143]= 1482939614;
assign addr[20144]= 1368621831;
assign addr[20145]= 1247361445;
assign addr[20146]= 1119773573;
assign addr[20147]= 986505429;
assign addr[20148]= 848233042;
assign addr[20149]= 705657826;
assign addr[20150]= 559503022;
assign addr[20151]= 410510029;
assign addr[20152]= 259434643;
assign addr[20153]= 107043224;
assign addr[20154]= -45891193;
assign addr[20155]= -198592817;
assign addr[20156]= -350287041;
assign addr[20157]= -500204365;
assign addr[20158]= -647584304;
assign addr[20159]= -791679244;
assign addr[20160]= -931758235;
assign addr[20161]= -1067110699;
assign addr[20162]= -1197050035;
assign addr[20163]= -1320917099;
assign addr[20164]= -1438083551;
assign addr[20165]= -1547955041;
assign addr[20166]= -1649974225;
assign addr[20167]= -1743623590;
assign addr[20168]= -1828428082;
assign addr[20169]= -1903957513;
assign addr[20170]= -1969828744;
assign addr[20171]= -2025707632;
assign addr[20172]= -2071310720;
assign addr[20173]= -2106406677;
assign addr[20174]= -2130817471;
assign addr[20175]= -2144419275;
assign addr[20176]= -2147143090;
assign addr[20177]= -2138975100;
assign addr[20178]= -2119956737;
assign addr[20179]= -2090184478;
assign addr[20180]= -2049809346;
assign addr[20181]= -1999036154;
assign addr[20182]= -1938122457;
assign addr[20183]= -1867377253;
assign addr[20184]= -1787159411;
assign addr[20185]= -1697875851;
assign addr[20186]= -1599979481;
assign addr[20187]= -1493966902;
assign addr[20188]= -1380375881;
assign addr[20189]= -1259782632;
assign addr[20190]= -1132798888;
assign addr[20191]= -1000068799;
assign addr[20192]= -862265664;
assign addr[20193]= -720088517;
assign addr[20194]= -574258580;
assign addr[20195]= -425515602;
assign addr[20196]= -274614114;
assign addr[20197]= -122319591;
assign addr[20198]= 30595422;
assign addr[20199]= 183355234;
assign addr[20200]= 335184940;
assign addr[20201]= 485314355;
assign addr[20202]= 632981917;
assign addr[20203]= 777438554;
assign addr[20204]= 917951481;
assign addr[20205]= 1053807919;
assign addr[20206]= 1184318708;
assign addr[20207]= 1308821808;
assign addr[20208]= 1426685652;
assign addr[20209]= 1537312353;
assign addr[20210]= 1640140734;
assign addr[20211]= 1734649179;
assign addr[20212]= 1820358275;
assign addr[20213]= 1896833245;
assign addr[20214]= 1963686155;
assign addr[20215]= 2020577882;
assign addr[20216]= 2067219829;
assign addr[20217]= 2103375398;
assign addr[20218]= 2128861181;
assign addr[20219]= 2143547897;
assign addr[20220]= 2147361045;
assign addr[20221]= 2140281282;
assign addr[20222]= 2122344521;
assign addr[20223]= 2093641749;
assign addr[20224]= 2054318569;
assign addr[20225]= 2004574453;
assign addr[20226]= 1944661739;
assign addr[20227]= 1874884346;
assign addr[20228]= 1795596234;
assign addr[20229]= 1707199606;
assign addr[20230]= 1610142873;
assign addr[20231]= 1504918373;
assign addr[20232]= 1392059879;
assign addr[20233]= 1272139887;
assign addr[20234]= 1145766716;
assign addr[20235]= 1013581418;
assign addr[20236]= 876254528;
assign addr[20237]= 734482665;
assign addr[20238]= 588984994;
assign addr[20239]= 440499581;
assign addr[20240]= 289779648;
assign addr[20241]= 137589750;
assign addr[20242]= -15298099;
assign addr[20243]= -168108346;
assign addr[20244]= -320065829;
assign addr[20245]= -470399716;
assign addr[20246]= -618347408;
assign addr[20247]= -763158411;
assign addr[20248]= -904098143;
assign addr[20249]= -1040451659;
assign addr[20250]= -1171527280;
assign addr[20251]= -1296660098;
assign addr[20252]= -1415215352;
assign addr[20253]= -1526591649;
assign addr[20254]= -1630224009;
assign addr[20255]= -1725586737;
assign addr[20256]= -1812196087;
assign addr[20257]= -1889612716;
assign addr[20258]= -1957443913;
assign addr[20259]= -2015345591;
assign addr[20260]= -2063024031;
assign addr[20261]= -2100237377;
assign addr[20262]= -2126796855;
assign addr[20263]= -2142567738;
assign addr[20264]= -2147470025;
assign addr[20265]= -2141478848;
assign addr[20266]= -2124624598;
assign addr[20267]= -2096992772;
assign addr[20268]= -2058723538;
assign addr[20269]= -2010011024;
assign addr[20270]= -1951102334;
assign addr[20271]= -1882296293;
assign addr[20272]= -1803941934;
assign addr[20273]= -1716436725;
assign addr[20274]= -1620224553;
assign addr[20275]= -1515793473;
assign addr[20276]= -1403673233;
assign addr[20277]= -1284432584;
assign addr[20278]= -1158676398;
assign addr[20279]= -1027042599;
assign addr[20280]= -890198924;
assign addr[20281]= -748839539;
assign addr[20282]= -603681519;
assign addr[20283]= -455461206;
assign addr[20284]= -304930476;
assign addr[20285]= -152852926;
assign addr[20286]= 0;
assign addr[20287]= 152852926;
assign addr[20288]= 304930476;
assign addr[20289]= 455461206;
assign addr[20290]= 603681519;
assign addr[20291]= 748839539;
assign addr[20292]= 890198924;
assign addr[20293]= 1027042599;
assign addr[20294]= 1158676398;
assign addr[20295]= 1284432584;
assign addr[20296]= 1403673233;
assign addr[20297]= 1515793473;
assign addr[20298]= 1620224553;
assign addr[20299]= 1716436725;
assign addr[20300]= 1803941934;
assign addr[20301]= 1882296293;
assign addr[20302]= 1951102334;
assign addr[20303]= 2010011024;
assign addr[20304]= 2058723538;
assign addr[20305]= 2096992772;
assign addr[20306]= 2124624598;
assign addr[20307]= 2141478848;
assign addr[20308]= 2147470025;
assign addr[20309]= 2142567738;
assign addr[20310]= 2126796855;
assign addr[20311]= 2100237377;
assign addr[20312]= 2063024031;
assign addr[20313]= 2015345591;
assign addr[20314]= 1957443913;
assign addr[20315]= 1889612716;
assign addr[20316]= 1812196087;
assign addr[20317]= 1725586737;
assign addr[20318]= 1630224009;
assign addr[20319]= 1526591649;
assign addr[20320]= 1415215352;
assign addr[20321]= 1296660098;
assign addr[20322]= 1171527280;
assign addr[20323]= 1040451659;
assign addr[20324]= 904098143;
assign addr[20325]= 763158411;
assign addr[20326]= 618347408;
assign addr[20327]= 470399716;
assign addr[20328]= 320065829;
assign addr[20329]= 168108346;
assign addr[20330]= 15298099;
assign addr[20331]= -137589750;
assign addr[20332]= -289779648;
assign addr[20333]= -440499581;
assign addr[20334]= -588984994;
assign addr[20335]= -734482665;
assign addr[20336]= -876254528;
assign addr[20337]= -1013581418;
assign addr[20338]= -1145766716;
assign addr[20339]= -1272139887;
assign addr[20340]= -1392059879;
assign addr[20341]= -1504918373;
assign addr[20342]= -1610142873;
assign addr[20343]= -1707199606;
assign addr[20344]= -1795596234;
assign addr[20345]= -1874884346;
assign addr[20346]= -1944661739;
assign addr[20347]= -2004574453;
assign addr[20348]= -2054318569;
assign addr[20349]= -2093641749;
assign addr[20350]= -2122344521;
assign addr[20351]= -2140281282;
assign addr[20352]= -2147361045;
assign addr[20353]= -2143547897;
assign addr[20354]= -2128861181;
assign addr[20355]= -2103375398;
assign addr[20356]= -2067219829;
assign addr[20357]= -2020577882;
assign addr[20358]= -1963686155;
assign addr[20359]= -1896833245;
assign addr[20360]= -1820358275;
assign addr[20361]= -1734649179;
assign addr[20362]= -1640140734;
assign addr[20363]= -1537312353;
assign addr[20364]= -1426685652;
assign addr[20365]= -1308821808;
assign addr[20366]= -1184318708;
assign addr[20367]= -1053807919;
assign addr[20368]= -917951481;
assign addr[20369]= -777438554;
assign addr[20370]= -632981917;
assign addr[20371]= -485314355;
assign addr[20372]= -335184940;
assign addr[20373]= -183355234;
assign addr[20374]= -30595422;
assign addr[20375]= 122319591;
assign addr[20376]= 274614114;
assign addr[20377]= 425515602;
assign addr[20378]= 574258580;
assign addr[20379]= 720088517;
assign addr[20380]= 862265664;
assign addr[20381]= 1000068799;
assign addr[20382]= 1132798888;
assign addr[20383]= 1259782632;
assign addr[20384]= 1380375881;
assign addr[20385]= 1493966902;
assign addr[20386]= 1599979481;
assign addr[20387]= 1697875851;
assign addr[20388]= 1787159411;
assign addr[20389]= 1867377253;
assign addr[20390]= 1938122457;
assign addr[20391]= 1999036154;
assign addr[20392]= 2049809346;
assign addr[20393]= 2090184478;
assign addr[20394]= 2119956737;
assign addr[20395]= 2138975100;
assign addr[20396]= 2147143090;
assign addr[20397]= 2144419275;
assign addr[20398]= 2130817471;
assign addr[20399]= 2106406677;
assign addr[20400]= 2071310720;
assign addr[20401]= 2025707632;
assign addr[20402]= 1969828744;
assign addr[20403]= 1903957513;
assign addr[20404]= 1828428082;
assign addr[20405]= 1743623590;
assign addr[20406]= 1649974225;
assign addr[20407]= 1547955041;
assign addr[20408]= 1438083551;
assign addr[20409]= 1320917099;
assign addr[20410]= 1197050035;
assign addr[20411]= 1067110699;
assign addr[20412]= 931758235;
assign addr[20413]= 791679244;
assign addr[20414]= 647584304;
assign addr[20415]= 500204365;
assign addr[20416]= 350287041;
assign addr[20417]= 198592817;
assign addr[20418]= 45891193;
assign addr[20419]= -107043224;
assign addr[20420]= -259434643;
assign addr[20421]= -410510029;
assign addr[20422]= -559503022;
assign addr[20423]= -705657826;
assign addr[20424]= -848233042;
assign addr[20425]= -986505429;
assign addr[20426]= -1119773573;
assign addr[20427]= -1247361445;
assign addr[20428]= -1368621831;
assign addr[20429]= -1482939614;
assign addr[20430]= -1589734894;
assign addr[20431]= -1688465931;
assign addr[20432]= -1778631892;
assign addr[20433]= -1859775393;
assign addr[20434]= -1931484818;
assign addr[20435]= -1993396407;
assign addr[20436]= -2045196100;
assign addr[20437]= -2086621133;
assign addr[20438]= -2117461370;
assign addr[20439]= -2137560369;
assign addr[20440]= -2146816171;
assign addr[20441]= -2145181827;
assign addr[20442]= -2132665626;
assign addr[20443]= -2109331059;
assign addr[20444]= -2075296495;
assign addr[20445]= -2030734582;
assign addr[20446]= -1975871368;
assign addr[20447]= -1910985158;
assign addr[20448]= -1836405100;
assign addr[20449]= -1752509516;
assign addr[20450]= -1659723983;
assign addr[20451]= -1558519173;
assign addr[20452]= -1449408469;
assign addr[20453]= -1332945355;
assign addr[20454]= -1209720613;
assign addr[20455]= -1080359326;
assign addr[20456]= -945517704;
assign addr[20457]= -805879757;
assign addr[20458]= -662153826;
assign addr[20459]= -515068990;
assign addr[20460]= -365371365;
assign addr[20461]= -213820322;
assign addr[20462]= -61184634;
assign addr[20463]= 91761426;
assign addr[20464]= 244242007;
assign addr[20465]= 395483624;
assign addr[20466]= 544719071;
assign addr[20467]= 691191324;
assign addr[20468]= 834157373;
assign addr[20469]= 972891995;
assign addr[20470]= 1106691431;
assign addr[20471]= 1234876957;
assign addr[20472]= 1356798326;
assign addr[20473]= 1471837070;
assign addr[20474]= 1579409630;
assign addr[20475]= 1678970324;
assign addr[20476]= 1770014111;
assign addr[20477]= 1852079154;
assign addr[20478]= 1924749160;
assign addr[20479]= 1987655498;
assign addr[20480]= 2040479063;
assign addr[20481]= 2082951896;
assign addr[20482]= 2114858546;
assign addr[20483]= 2136037160;
assign addr[20484]= 2146380306;
assign addr[20485]= 2145835515;
assign addr[20486]= 2134405552;
assign addr[20487]= 2112148396;
assign addr[20488]= 2079176953;
assign addr[20489]= 2035658475;
assign addr[20490]= 1981813720;
assign addr[20491]= 1917915825;
assign addr[20492]= 1844288924;
assign addr[20493]= 1761306505;
assign addr[20494]= 1669389513;
assign addr[20495]= 1569004214;
assign addr[20496]= 1460659832;
assign addr[20497]= 1344905966;
assign addr[20498]= 1222329801;
assign addr[20499]= 1093553126;
assign addr[20500]= 959229189;
assign addr[20501]= 820039373;
assign addr[20502]= 676689746;
assign addr[20503]= 529907477;
assign addr[20504]= 380437148;
assign addr[20505]= 229036977;
assign addr[20506]= 76474970;
assign addr[20507]= -76474970;
assign addr[20508]= -229036977;
assign addr[20509]= -380437148;
assign addr[20510]= -529907477;
assign addr[20511]= -676689746;
assign addr[20512]= -820039373;
assign addr[20513]= -959229189;
assign addr[20514]= -1093553126;
assign addr[20515]= -1222329801;
assign addr[20516]= -1344905966;
assign addr[20517]= -1460659832;
assign addr[20518]= -1569004214;
assign addr[20519]= -1669389513;
assign addr[20520]= -1761306505;
assign addr[20521]= -1844288924;
assign addr[20522]= -1917915825;
assign addr[20523]= -1981813720;
assign addr[20524]= -2035658475;
assign addr[20525]= -2079176953;
assign addr[20526]= -2112148396;
assign addr[20527]= -2134405552;
assign addr[20528]= -2145835515;
assign addr[20529]= -2146380306;
assign addr[20530]= -2136037160;
assign addr[20531]= -2114858546;
assign addr[20532]= -2082951896;
assign addr[20533]= -2040479063;
assign addr[20534]= -1987655498;
assign addr[20535]= -1924749160;
assign addr[20536]= -1852079154;
assign addr[20537]= -1770014111;
assign addr[20538]= -1678970324;
assign addr[20539]= -1579409630;
assign addr[20540]= -1471837070;
assign addr[20541]= -1356798326;
assign addr[20542]= -1234876957;
assign addr[20543]= -1106691431;
assign addr[20544]= -972891995;
assign addr[20545]= -834157373;
assign addr[20546]= -691191324;
assign addr[20547]= -544719071;
assign addr[20548]= -395483624;
assign addr[20549]= -244242007;
assign addr[20550]= -91761426;
assign addr[20551]= 61184634;
assign addr[20552]= 213820322;
assign addr[20553]= 365371365;
assign addr[20554]= 515068990;
assign addr[20555]= 662153826;
assign addr[20556]= 805879757;
assign addr[20557]= 945517704;
assign addr[20558]= 1080359326;
assign addr[20559]= 1209720613;
assign addr[20560]= 1332945355;
assign addr[20561]= 1449408469;
assign addr[20562]= 1558519173;
assign addr[20563]= 1659723983;
assign addr[20564]= 1752509516;
assign addr[20565]= 1836405100;
assign addr[20566]= 1910985158;
assign addr[20567]= 1975871368;
assign addr[20568]= 2030734582;
assign addr[20569]= 2075296495;
assign addr[20570]= 2109331059;
assign addr[20571]= 2132665626;
assign addr[20572]= 2145181827;
assign addr[20573]= 2146816171;
assign addr[20574]= 2137560369;
assign addr[20575]= 2117461370;
assign addr[20576]= 2086621133;
assign addr[20577]= 2045196100;
assign addr[20578]= 1993396407;
assign addr[20579]= 1931484818;
assign addr[20580]= 1859775393;
assign addr[20581]= 1778631892;
assign addr[20582]= 1688465931;
assign addr[20583]= 1589734894;
assign addr[20584]= 1482939614;
assign addr[20585]= 1368621831;
assign addr[20586]= 1247361445;
assign addr[20587]= 1119773573;
assign addr[20588]= 986505429;
assign addr[20589]= 848233042;
assign addr[20590]= 705657826;
assign addr[20591]= 559503022;
assign addr[20592]= 410510029;
assign addr[20593]= 259434643;
assign addr[20594]= 107043224;
assign addr[20595]= -45891193;
assign addr[20596]= -198592817;
assign addr[20597]= -350287041;
assign addr[20598]= -500204365;
assign addr[20599]= -647584304;
assign addr[20600]= -791679244;
assign addr[20601]= -931758235;
assign addr[20602]= -1067110699;
assign addr[20603]= -1197050035;
assign addr[20604]= -1320917099;
assign addr[20605]= -1438083551;
assign addr[20606]= -1547955041;
assign addr[20607]= -1649974225;
assign addr[20608]= -1743623590;
assign addr[20609]= -1828428082;
assign addr[20610]= -1903957513;
assign addr[20611]= -1969828744;
assign addr[20612]= -2025707632;
assign addr[20613]= -2071310720;
assign addr[20614]= -2106406677;
assign addr[20615]= -2130817471;
assign addr[20616]= -2144419275;
assign addr[20617]= -2147143090;
assign addr[20618]= -2138975100;
assign addr[20619]= -2119956737;
assign addr[20620]= -2090184478;
assign addr[20621]= -2049809346;
assign addr[20622]= -1999036154;
assign addr[20623]= -1938122457;
assign addr[20624]= -1867377253;
assign addr[20625]= -1787159411;
assign addr[20626]= -1697875851;
assign addr[20627]= -1599979481;
assign addr[20628]= -1493966902;
assign addr[20629]= -1380375881;
assign addr[20630]= -1259782632;
assign addr[20631]= -1132798888;
assign addr[20632]= -1000068799;
assign addr[20633]= -862265664;
assign addr[20634]= -720088517;
assign addr[20635]= -574258580;
assign addr[20636]= -425515602;
assign addr[20637]= -274614114;
assign addr[20638]= -122319591;
assign addr[20639]= 30595422;
assign addr[20640]= 183355234;
assign addr[20641]= 335184940;
assign addr[20642]= 485314355;
assign addr[20643]= 632981917;
assign addr[20644]= 777438554;
assign addr[20645]= 917951481;
assign addr[20646]= 1053807919;
assign addr[20647]= 1184318708;
assign addr[20648]= 1308821808;
assign addr[20649]= 1426685652;
assign addr[20650]= 1537312353;
assign addr[20651]= 1640140734;
assign addr[20652]= 1734649179;
assign addr[20653]= 1820358275;
assign addr[20654]= 1896833245;
assign addr[20655]= 1963686155;
assign addr[20656]= 2020577882;
assign addr[20657]= 2067219829;
assign addr[20658]= 2103375398;
assign addr[20659]= 2128861181;
assign addr[20660]= 2143547897;
assign addr[20661]= 2147361045;
assign addr[20662]= 2140281282;
assign addr[20663]= 2122344521;
assign addr[20664]= 2093641749;
assign addr[20665]= 2054318569;
assign addr[20666]= 2004574453;
assign addr[20667]= 1944661739;
assign addr[20668]= 1874884346;
assign addr[20669]= 1795596234;
assign addr[20670]= 1707199606;
assign addr[20671]= 1610142873;
assign addr[20672]= 1504918373;
assign addr[20673]= 1392059879;
assign addr[20674]= 1272139887;
assign addr[20675]= 1145766716;
assign addr[20676]= 1013581418;
assign addr[20677]= 876254528;
assign addr[20678]= 734482665;
assign addr[20679]= 588984994;
assign addr[20680]= 440499581;
assign addr[20681]= 289779648;
assign addr[20682]= 137589750;
assign addr[20683]= -15298099;
assign addr[20684]= -168108346;
assign addr[20685]= -320065829;
assign addr[20686]= -470399716;
assign addr[20687]= -618347408;
assign addr[20688]= -763158411;
assign addr[20689]= -904098143;
assign addr[20690]= -1040451659;
assign addr[20691]= -1171527280;
assign addr[20692]= -1296660098;
assign addr[20693]= -1415215352;
assign addr[20694]= -1526591649;
assign addr[20695]= -1630224009;
assign addr[20696]= -1725586737;
assign addr[20697]= -1812196087;
assign addr[20698]= -1889612716;
assign addr[20699]= -1957443913;
assign addr[20700]= -2015345591;
assign addr[20701]= -2063024031;
assign addr[20702]= -2100237377;
assign addr[20703]= -2126796855;
assign addr[20704]= -2142567738;
assign addr[20705]= -2147470025;
assign addr[20706]= -2141478848;
assign addr[20707]= -2124624598;
assign addr[20708]= -2096992772;
assign addr[20709]= -2058723538;
assign addr[20710]= -2010011024;
assign addr[20711]= -1951102334;
assign addr[20712]= -1882296293;
assign addr[20713]= -1803941934;
assign addr[20714]= -1716436725;
assign addr[20715]= -1620224553;
assign addr[20716]= -1515793473;
assign addr[20717]= -1403673233;
assign addr[20718]= -1284432584;
assign addr[20719]= -1158676398;
assign addr[20720]= -1027042599;
assign addr[20721]= -890198924;
assign addr[20722]= -748839539;
assign addr[20723]= -603681519;
assign addr[20724]= -455461206;
assign addr[20725]= -304930476;
assign addr[20726]= -152852926;
assign addr[20727]= 0;
assign addr[20728]= 152852926;
assign addr[20729]= 304930476;
assign addr[20730]= 455461206;
assign addr[20731]= 603681519;
assign addr[20732]= 748839539;
assign addr[20733]= 890198924;
assign addr[20734]= 1027042599;
assign addr[20735]= 1158676398;
assign addr[20736]= 1284432584;
assign addr[20737]= 1403673233;
assign addr[20738]= 1515793473;
assign addr[20739]= 1620224553;
assign addr[20740]= 1716436725;
assign addr[20741]= 1803941934;
assign addr[20742]= 1882296293;
assign addr[20743]= 1951102334;
assign addr[20744]= 2010011024;
assign addr[20745]= 2058723538;
assign addr[20746]= 2096992772;
assign addr[20747]= 2124624598;
assign addr[20748]= 2141478848;
assign addr[20749]= 2147470025;
assign addr[20750]= 2142567738;
assign addr[20751]= 2126796855;
assign addr[20752]= 2100237377;
assign addr[20753]= 2063024031;
assign addr[20754]= 2015345591;
assign addr[20755]= 1957443913;
assign addr[20756]= 1889612716;
assign addr[20757]= 1812196087;
assign addr[20758]= 1725586737;
assign addr[20759]= 1630224009;
assign addr[20760]= 1526591649;
assign addr[20761]= 1415215352;
assign addr[20762]= 1296660098;
assign addr[20763]= 1171527280;
assign addr[20764]= 1040451659;
assign addr[20765]= 904098143;
assign addr[20766]= 763158411;
assign addr[20767]= 618347408;
assign addr[20768]= 470399716;
assign addr[20769]= 320065829;
assign addr[20770]= 168108346;
assign addr[20771]= 15298099;
assign addr[20772]= -137589750;
assign addr[20773]= -289779648;
assign addr[20774]= -440499581;
assign addr[20775]= -588984994;
assign addr[20776]= -734482665;
assign addr[20777]= -876254528;
assign addr[20778]= -1013581418;
assign addr[20779]= -1145766716;
assign addr[20780]= -1272139887;
assign addr[20781]= -1392059879;
assign addr[20782]= -1504918373;
assign addr[20783]= -1610142873;
assign addr[20784]= -1707199606;
assign addr[20785]= -1795596234;
assign addr[20786]= -1874884346;
assign addr[20787]= -1944661739;
assign addr[20788]= -2004574453;
assign addr[20789]= -2054318569;
assign addr[20790]= -2093641749;
assign addr[20791]= -2122344521;
assign addr[20792]= -2140281282;
assign addr[20793]= -2147361045;
assign addr[20794]= -2143547897;
assign addr[20795]= -2128861181;
assign addr[20796]= -2103375398;
assign addr[20797]= -2067219829;
assign addr[20798]= -2020577882;
assign addr[20799]= -1963686155;
assign addr[20800]= -1896833245;
assign addr[20801]= -1820358275;
assign addr[20802]= -1734649179;
assign addr[20803]= -1640140734;
assign addr[20804]= -1537312353;
assign addr[20805]= -1426685652;
assign addr[20806]= -1308821808;
assign addr[20807]= -1184318708;
assign addr[20808]= -1053807919;
assign addr[20809]= -917951481;
assign addr[20810]= -777438554;
assign addr[20811]= -632981917;
assign addr[20812]= -485314355;
assign addr[20813]= -335184940;
assign addr[20814]= -183355234;
assign addr[20815]= -30595422;
assign addr[20816]= 122319591;
assign addr[20817]= 274614114;
assign addr[20818]= 425515602;
assign addr[20819]= 574258580;
assign addr[20820]= 720088517;
assign addr[20821]= 862265664;
assign addr[20822]= 1000068799;
assign addr[20823]= 1132798888;
assign addr[20824]= 1259782632;
assign addr[20825]= 1380375881;
assign addr[20826]= 1493966902;
assign addr[20827]= 1599979481;
assign addr[20828]= 1697875851;
assign addr[20829]= 1787159411;
assign addr[20830]= 1867377253;
assign addr[20831]= 1938122457;
assign addr[20832]= 1999036154;
assign addr[20833]= 2049809346;
assign addr[20834]= 2090184478;
assign addr[20835]= 2119956737;
assign addr[20836]= 2138975100;
assign addr[20837]= 2147143090;
assign addr[20838]= 2144419275;
assign addr[20839]= 2130817471;
assign addr[20840]= 2106406677;
assign addr[20841]= 2071310720;
assign addr[20842]= 2025707632;
assign addr[20843]= 1969828744;
assign addr[20844]= 1903957513;
assign addr[20845]= 1828428082;
assign addr[20846]= 1743623590;
assign addr[20847]= 1649974225;
assign addr[20848]= 1547955041;
assign addr[20849]= 1438083551;
assign addr[20850]= 1320917099;
assign addr[20851]= 1197050035;
assign addr[20852]= 1067110699;
assign addr[20853]= 931758235;
assign addr[20854]= 791679244;
assign addr[20855]= 647584304;
assign addr[20856]= 500204365;
assign addr[20857]= 350287041;
assign addr[20858]= 198592817;
assign addr[20859]= 45891193;
assign addr[20860]= -107043224;
assign addr[20861]= -259434643;
assign addr[20862]= -410510029;
assign addr[20863]= -559503022;
assign addr[20864]= -705657826;
assign addr[20865]= -848233042;
assign addr[20866]= -986505429;
assign addr[20867]= -1119773573;
assign addr[20868]= -1247361445;
assign addr[20869]= -1368621831;
assign addr[20870]= -1482939614;
assign addr[20871]= -1589734894;
assign addr[20872]= -1688465931;
assign addr[20873]= -1778631892;
assign addr[20874]= -1859775393;
assign addr[20875]= -1931484818;
assign addr[20876]= -1993396407;
assign addr[20877]= -2045196100;
assign addr[20878]= -2086621133;
assign addr[20879]= -2117461370;
assign addr[20880]= -2137560369;
assign addr[20881]= -2146816171;
assign addr[20882]= -2145181827;
assign addr[20883]= -2132665626;
assign addr[20884]= -2109331059;
assign addr[20885]= -2075296495;
assign addr[20886]= -2030734582;
assign addr[20887]= -1975871368;
assign addr[20888]= -1910985158;
assign addr[20889]= -1836405100;
assign addr[20890]= -1752509516;
assign addr[20891]= -1659723983;
assign addr[20892]= -1558519173;
assign addr[20893]= -1449408469;
assign addr[20894]= -1332945355;
assign addr[20895]= -1209720613;
assign addr[20896]= -1080359326;
assign addr[20897]= -945517704;
assign addr[20898]= -805879757;
assign addr[20899]= -662153826;
assign addr[20900]= -515068990;
assign addr[20901]= -365371365;
assign addr[20902]= -213820322;
assign addr[20903]= -61184634;
assign addr[20904]= 91761426;
assign addr[20905]= 244242007;
assign addr[20906]= 395483624;
assign addr[20907]= 544719071;
assign addr[20908]= 691191324;
assign addr[20909]= 834157373;
assign addr[20910]= 972891995;
assign addr[20911]= 1106691431;
assign addr[20912]= 1234876957;
assign addr[20913]= 1356798326;
assign addr[20914]= 1471837070;
assign addr[20915]= 1579409630;
assign addr[20916]= 1678970324;
assign addr[20917]= 1770014111;
assign addr[20918]= 1852079154;
assign addr[20919]= 1924749160;
assign addr[20920]= 1987655498;
assign addr[20921]= 2040479063;
assign addr[20922]= 2082951896;
assign addr[20923]= 2114858546;
assign addr[20924]= 2136037160;
assign addr[20925]= 2146380306;
assign addr[20926]= 2145835515;
assign addr[20927]= 2134405552;
assign addr[20928]= 2112148396;
assign addr[20929]= 2079176953;
assign addr[20930]= 2035658475;
assign addr[20931]= 1981813720;
assign addr[20932]= 1917915825;
assign addr[20933]= 1844288924;
assign addr[20934]= 1761306505;
assign addr[20935]= 1669389513;
assign addr[20936]= 1569004214;
assign addr[20937]= 1460659832;
assign addr[20938]= 1344905966;
assign addr[20939]= 1222329801;
assign addr[20940]= 1093553126;
assign addr[20941]= 959229189;
assign addr[20942]= 820039373;
assign addr[20943]= 676689746;
assign addr[20944]= 529907477;
assign addr[20945]= 380437148;
assign addr[20946]= 229036977;
assign addr[20947]= 76474970;
assign addr[20948]= -76474970;
assign addr[20949]= -229036977;
assign addr[20950]= -380437148;
assign addr[20951]= -529907477;
assign addr[20952]= -676689746;
assign addr[20953]= -820039373;
assign addr[20954]= -959229189;
assign addr[20955]= -1093553126;
assign addr[20956]= -1222329801;
assign addr[20957]= -1344905966;
assign addr[20958]= -1460659832;
assign addr[20959]= -1569004214;
assign addr[20960]= -1669389513;
assign addr[20961]= -1761306505;
assign addr[20962]= -1844288924;
assign addr[20963]= -1917915825;
assign addr[20964]= -1981813720;
assign addr[20965]= -2035658475;
assign addr[20966]= -2079176953;
assign addr[20967]= -2112148396;
assign addr[20968]= -2134405552;
assign addr[20969]= -2145835515;
assign addr[20970]= -2146380306;
assign addr[20971]= -2136037160;
assign addr[20972]= -2114858546;
assign addr[20973]= -2082951896;
assign addr[20974]= -2040479063;
assign addr[20975]= -1987655498;
assign addr[20976]= -1924749160;
assign addr[20977]= -1852079154;
assign addr[20978]= -1770014111;
assign addr[20979]= -1678970324;
assign addr[20980]= -1579409630;
assign addr[20981]= -1471837070;
assign addr[20982]= -1356798326;
assign addr[20983]= -1234876957;
assign addr[20984]= -1106691431;
assign addr[20985]= -972891995;
assign addr[20986]= -834157373;
assign addr[20987]= -691191324;
assign addr[20988]= -544719071;
assign addr[20989]= -395483624;
assign addr[20990]= -244242007;
assign addr[20991]= -91761426;
assign addr[20992]= 61184634;
assign addr[20993]= 213820322;
assign addr[20994]= 365371365;
assign addr[20995]= 515068990;
assign addr[20996]= 662153826;
assign addr[20997]= 805879757;
assign addr[20998]= 945517704;
assign addr[20999]= 1080359326;
assign addr[21000]= 1209720613;
assign addr[21001]= 1332945355;
assign addr[21002]= 1449408469;
assign addr[21003]= 1558519173;
assign addr[21004]= 1659723983;
assign addr[21005]= 1752509516;
assign addr[21006]= 1836405100;
assign addr[21007]= 1910985158;
assign addr[21008]= 1975871368;
assign addr[21009]= 2030734582;
assign addr[21010]= 2075296495;
assign addr[21011]= 2109331059;
assign addr[21012]= 2132665626;
assign addr[21013]= 2145181827;
assign addr[21014]= 2146816171;
assign addr[21015]= 2137560369;
assign addr[21016]= 2117461370;
assign addr[21017]= 2086621133;
assign addr[21018]= 2045196100;
assign addr[21019]= 1993396407;
assign addr[21020]= 1931484818;
assign addr[21021]= 1859775393;
assign addr[21022]= 1778631892;
assign addr[21023]= 1688465931;
assign addr[21024]= 1589734894;
assign addr[21025]= 1482939614;
assign addr[21026]= 1368621831;
assign addr[21027]= 1247361445;
assign addr[21028]= 1119773573;
assign addr[21029]= 986505429;
assign addr[21030]= 848233042;
assign addr[21031]= 705657826;
assign addr[21032]= 559503022;
assign addr[21033]= 410510029;
assign addr[21034]= 259434643;
assign addr[21035]= 107043224;
assign addr[21036]= -45891193;
assign addr[21037]= -198592817;
assign addr[21038]= -350287041;
assign addr[21039]= -500204365;
assign addr[21040]= -647584304;
assign addr[21041]= -791679244;
assign addr[21042]= -931758235;
assign addr[21043]= -1067110699;
assign addr[21044]= -1197050035;
assign addr[21045]= -1320917099;
assign addr[21046]= -1438083551;
assign addr[21047]= -1547955041;
assign addr[21048]= -1649974225;
assign addr[21049]= -1743623590;
assign addr[21050]= -1828428082;
assign addr[21051]= -1903957513;
assign addr[21052]= -1969828744;
assign addr[21053]= -2025707632;
assign addr[21054]= -2071310720;
assign addr[21055]= -2106406677;
assign addr[21056]= -2130817471;
assign addr[21057]= -2144419275;
assign addr[21058]= -2147143090;
assign addr[21059]= -2138975100;
assign addr[21060]= -2119956737;
assign addr[21061]= -2090184478;
assign addr[21062]= -2049809346;
assign addr[21063]= -1999036154;
assign addr[21064]= -1938122457;
assign addr[21065]= -1867377253;
assign addr[21066]= -1787159411;
assign addr[21067]= -1697875851;
assign addr[21068]= -1599979481;
assign addr[21069]= -1493966902;
assign addr[21070]= -1380375881;
assign addr[21071]= -1259782632;
assign addr[21072]= -1132798888;
assign addr[21073]= -1000068799;
assign addr[21074]= -862265664;
assign addr[21075]= -720088517;
assign addr[21076]= -574258580;
assign addr[21077]= -425515602;
assign addr[21078]= -274614114;
assign addr[21079]= -122319591;
assign addr[21080]= 30595422;
assign addr[21081]= 183355234;
assign addr[21082]= 335184940;
assign addr[21083]= 485314355;
assign addr[21084]= 632981917;
assign addr[21085]= 777438554;
assign addr[21086]= 917951481;
assign addr[21087]= 1053807919;
assign addr[21088]= 1184318708;
assign addr[21089]= 1308821808;
assign addr[21090]= 1426685652;
assign addr[21091]= 1537312353;
assign addr[21092]= 1640140734;
assign addr[21093]= 1734649179;
assign addr[21094]= 1820358275;
assign addr[21095]= 1896833245;
assign addr[21096]= 1963686155;
assign addr[21097]= 2020577882;
assign addr[21098]= 2067219829;
assign addr[21099]= 2103375398;
assign addr[21100]= 2128861181;
assign addr[21101]= 2143547897;
assign addr[21102]= 2147361045;
assign addr[21103]= 2140281282;
assign addr[21104]= 2122344521;
assign addr[21105]= 2093641749;
assign addr[21106]= 2054318569;
assign addr[21107]= 2004574453;
assign addr[21108]= 1944661739;
assign addr[21109]= 1874884346;
assign addr[21110]= 1795596234;
assign addr[21111]= 1707199606;
assign addr[21112]= 1610142873;
assign addr[21113]= 1504918373;
assign addr[21114]= 1392059879;
assign addr[21115]= 1272139887;
assign addr[21116]= 1145766716;
assign addr[21117]= 1013581418;
assign addr[21118]= 876254528;
assign addr[21119]= 734482665;
assign addr[21120]= 588984994;
assign addr[21121]= 440499581;
assign addr[21122]= 289779648;
assign addr[21123]= 137589750;
assign addr[21124]= -15298099;
assign addr[21125]= -168108346;
assign addr[21126]= -320065829;
assign addr[21127]= -470399716;
assign addr[21128]= -618347408;
assign addr[21129]= -763158411;
assign addr[21130]= -904098143;
assign addr[21131]= -1040451659;
assign addr[21132]= -1171527280;
assign addr[21133]= -1296660098;
assign addr[21134]= -1415215352;
assign addr[21135]= -1526591649;
assign addr[21136]= -1630224009;
assign addr[21137]= -1725586737;
assign addr[21138]= -1812196087;
assign addr[21139]= -1889612716;
assign addr[21140]= -1957443913;
assign addr[21141]= -2015345591;
assign addr[21142]= -2063024031;
assign addr[21143]= -2100237377;
assign addr[21144]= -2126796855;
assign addr[21145]= -2142567738;
assign addr[21146]= -2147470025;
assign addr[21147]= -2141478848;
assign addr[21148]= -2124624598;
assign addr[21149]= -2096992772;
assign addr[21150]= -2058723538;
assign addr[21151]= -2010011024;
assign addr[21152]= -1951102334;
assign addr[21153]= -1882296293;
assign addr[21154]= -1803941934;
assign addr[21155]= -1716436725;
assign addr[21156]= -1620224553;
assign addr[21157]= -1515793473;
assign addr[21158]= -1403673233;
assign addr[21159]= -1284432584;
assign addr[21160]= -1158676398;
assign addr[21161]= -1027042599;
assign addr[21162]= -890198924;
assign addr[21163]= -748839539;
assign addr[21164]= -603681519;
assign addr[21165]= -455461206;
assign addr[21166]= -304930476;
assign addr[21167]= -152852926;
assign addr[21168]= 0;
assign addr[21169]= 152852926;
assign addr[21170]= 304930476;
assign addr[21171]= 455461206;
assign addr[21172]= 603681519;
assign addr[21173]= 748839539;
assign addr[21174]= 890198924;
assign addr[21175]= 1027042599;
assign addr[21176]= 1158676398;
assign addr[21177]= 1284432584;
assign addr[21178]= 1403673233;
assign addr[21179]= 1515793473;
assign addr[21180]= 1620224553;
assign addr[21181]= 1716436725;
assign addr[21182]= 1803941934;
assign addr[21183]= 1882296293;
assign addr[21184]= 1951102334;
assign addr[21185]= 2010011024;
assign addr[21186]= 2058723538;
assign addr[21187]= 2096992772;
assign addr[21188]= 2124624598;
assign addr[21189]= 2141478848;
assign addr[21190]= 2147470025;
assign addr[21191]= 2142567738;
assign addr[21192]= 2126796855;
assign addr[21193]= 2100237377;
assign addr[21194]= 2063024031;
assign addr[21195]= 2015345591;
assign addr[21196]= 1957443913;
assign addr[21197]= 1889612716;
assign addr[21198]= 1812196087;
assign addr[21199]= 1725586737;
assign addr[21200]= 1630224009;
assign addr[21201]= 1526591649;
assign addr[21202]= 1415215352;
assign addr[21203]= 1296660098;
assign addr[21204]= 1171527280;
assign addr[21205]= 1040451659;
assign addr[21206]= 904098143;
assign addr[21207]= 763158411;
assign addr[21208]= 618347408;
assign addr[21209]= 470399716;
assign addr[21210]= 320065829;
assign addr[21211]= 168108346;
assign addr[21212]= 15298099;
assign addr[21213]= -137589750;
assign addr[21214]= -289779648;
assign addr[21215]= -440499581;
assign addr[21216]= -588984994;
assign addr[21217]= -734482665;
assign addr[21218]= -876254528;
assign addr[21219]= -1013581418;
assign addr[21220]= -1145766716;
assign addr[21221]= -1272139887;
assign addr[21222]= -1392059879;
assign addr[21223]= -1504918373;
assign addr[21224]= -1610142873;
assign addr[21225]= -1707199606;
assign addr[21226]= -1795596234;
assign addr[21227]= -1874884346;
assign addr[21228]= -1944661739;
assign addr[21229]= -2004574453;
assign addr[21230]= -2054318569;
assign addr[21231]= -2093641749;
assign addr[21232]= -2122344521;
assign addr[21233]= -2140281282;
assign addr[21234]= -2147361045;
assign addr[21235]= -2143547897;
assign addr[21236]= -2128861181;
assign addr[21237]= -2103375398;
assign addr[21238]= -2067219829;
assign addr[21239]= -2020577882;
assign addr[21240]= -1963686155;
assign addr[21241]= -1896833245;
assign addr[21242]= -1820358275;
assign addr[21243]= -1734649179;
assign addr[21244]= -1640140734;
assign addr[21245]= -1537312353;
assign addr[21246]= -1426685652;
assign addr[21247]= -1308821808;
assign addr[21248]= -1184318708;
assign addr[21249]= -1053807919;
assign addr[21250]= -917951481;
assign addr[21251]= -777438554;
assign addr[21252]= -632981917;
assign addr[21253]= -485314355;
assign addr[21254]= -335184940;
assign addr[21255]= -183355234;
assign addr[21256]= -30595422;
assign addr[21257]= 122319591;
assign addr[21258]= 274614114;
assign addr[21259]= 425515602;
assign addr[21260]= 574258580;
assign addr[21261]= 720088517;
assign addr[21262]= 862265664;
assign addr[21263]= 1000068799;
assign addr[21264]= 1132798888;
assign addr[21265]= 1259782632;
assign addr[21266]= 1380375881;
assign addr[21267]= 1493966902;
assign addr[21268]= 1599979481;
assign addr[21269]= 1697875851;
assign addr[21270]= 1787159411;
assign addr[21271]= 1867377253;
assign addr[21272]= 1938122457;
assign addr[21273]= 1999036154;
assign addr[21274]= 2049809346;
assign addr[21275]= 2090184478;
assign addr[21276]= 2119956737;
assign addr[21277]= 2138975100;
assign addr[21278]= 2147143090;
assign addr[21279]= 2144419275;
assign addr[21280]= 2130817471;
assign addr[21281]= 2106406677;
assign addr[21282]= 2071310720;
assign addr[21283]= 2025707632;
assign addr[21284]= 1969828744;
assign addr[21285]= 1903957513;
assign addr[21286]= 1828428082;
assign addr[21287]= 1743623590;
assign addr[21288]= 1649974225;
assign addr[21289]= 1547955041;
assign addr[21290]= 1438083551;
assign addr[21291]= 1320917099;
assign addr[21292]= 1197050035;
assign addr[21293]= 1067110699;
assign addr[21294]= 931758235;
assign addr[21295]= 791679244;
assign addr[21296]= 647584304;
assign addr[21297]= 500204365;
assign addr[21298]= 350287041;
assign addr[21299]= 198592817;
assign addr[21300]= 45891193;
assign addr[21301]= -107043224;
assign addr[21302]= -259434643;
assign addr[21303]= -410510029;
assign addr[21304]= -559503022;
assign addr[21305]= -705657826;
assign addr[21306]= -848233042;
assign addr[21307]= -986505429;
assign addr[21308]= -1119773573;
assign addr[21309]= -1247361445;
assign addr[21310]= -1368621831;
assign addr[21311]= -1482939614;
assign addr[21312]= -1589734894;
assign addr[21313]= -1688465931;
assign addr[21314]= -1778631892;
assign addr[21315]= -1859775393;
assign addr[21316]= -1931484818;
assign addr[21317]= -1993396407;
assign addr[21318]= -2045196100;
assign addr[21319]= -2086621133;
assign addr[21320]= -2117461370;
assign addr[21321]= -2137560369;
assign addr[21322]= -2146816171;
assign addr[21323]= -2145181827;
assign addr[21324]= -2132665626;
assign addr[21325]= -2109331059;
assign addr[21326]= -2075296495;
assign addr[21327]= -2030734582;
assign addr[21328]= -1975871368;
assign addr[21329]= -1910985158;
assign addr[21330]= -1836405100;
assign addr[21331]= -1752509516;
assign addr[21332]= -1659723983;
assign addr[21333]= -1558519173;
assign addr[21334]= -1449408469;
assign addr[21335]= -1332945355;
assign addr[21336]= -1209720613;
assign addr[21337]= -1080359326;
assign addr[21338]= -945517704;
assign addr[21339]= -805879757;
assign addr[21340]= -662153826;
assign addr[21341]= -515068990;
assign addr[21342]= -365371365;
assign addr[21343]= -213820322;
assign addr[21344]= -61184634;
assign addr[21345]= 91761426;
assign addr[21346]= 244242007;
assign addr[21347]= 395483624;
assign addr[21348]= 544719071;
assign addr[21349]= 691191324;
assign addr[21350]= 834157373;
assign addr[21351]= 972891995;
assign addr[21352]= 1106691431;
assign addr[21353]= 1234876957;
assign addr[21354]= 1356798326;
assign addr[21355]= 1471837070;
assign addr[21356]= 1579409630;
assign addr[21357]= 1678970324;
assign addr[21358]= 1770014111;
assign addr[21359]= 1852079154;
assign addr[21360]= 1924749160;
assign addr[21361]= 1987655498;
assign addr[21362]= 2040479063;
assign addr[21363]= 2082951896;
assign addr[21364]= 2114858546;
assign addr[21365]= 2136037160;
assign addr[21366]= 2146380306;
assign addr[21367]= 2145835515;
assign addr[21368]= 2134405552;
assign addr[21369]= 2112148396;
assign addr[21370]= 2079176953;
assign addr[21371]= 2035658475;
assign addr[21372]= 1981813720;
assign addr[21373]= 1917915825;
assign addr[21374]= 1844288924;
assign addr[21375]= 1761306505;
assign addr[21376]= 1669389513;
assign addr[21377]= 1569004214;
assign addr[21378]= 1460659832;
assign addr[21379]= 1344905966;
assign addr[21380]= 1222329801;
assign addr[21381]= 1093553126;
assign addr[21382]= 959229189;
assign addr[21383]= 820039373;
assign addr[21384]= 676689746;
assign addr[21385]= 529907477;
assign addr[21386]= 380437148;
assign addr[21387]= 229036977;
assign addr[21388]= 76474970;
assign addr[21389]= -76474970;
assign addr[21390]= -229036977;
assign addr[21391]= -380437148;
assign addr[21392]= -529907477;
assign addr[21393]= -676689746;
assign addr[21394]= -820039373;
assign addr[21395]= -959229189;
assign addr[21396]= -1093553126;
assign addr[21397]= -1222329801;
assign addr[21398]= -1344905966;
assign addr[21399]= -1460659832;
assign addr[21400]= -1569004214;
assign addr[21401]= -1669389513;
assign addr[21402]= -1761306505;
assign addr[21403]= -1844288924;
assign addr[21404]= -1917915825;
assign addr[21405]= -1981813720;
assign addr[21406]= -2035658475;
assign addr[21407]= -2079176953;
assign addr[21408]= -2112148396;
assign addr[21409]= -2134405552;
assign addr[21410]= -2145835515;
assign addr[21411]= -2146380306;
assign addr[21412]= -2136037160;
assign addr[21413]= -2114858546;
assign addr[21414]= -2082951896;
assign addr[21415]= -2040479063;
assign addr[21416]= -1987655498;
assign addr[21417]= -1924749160;
assign addr[21418]= -1852079154;
assign addr[21419]= -1770014111;
assign addr[21420]= -1678970324;
assign addr[21421]= -1579409630;
assign addr[21422]= -1471837070;
assign addr[21423]= -1356798326;
assign addr[21424]= -1234876957;
assign addr[21425]= -1106691431;
assign addr[21426]= -972891995;
assign addr[21427]= -834157373;
assign addr[21428]= -691191324;
assign addr[21429]= -544719071;
assign addr[21430]= -395483624;
assign addr[21431]= -244242007;
assign addr[21432]= -91761426;
assign addr[21433]= 61184634;
assign addr[21434]= 213820322;
assign addr[21435]= 365371365;
assign addr[21436]= 515068990;
assign addr[21437]= 662153826;
assign addr[21438]= 805879757;
assign addr[21439]= 945517704;
assign addr[21440]= 1080359326;
assign addr[21441]= 1209720613;
assign addr[21442]= 1332945355;
assign addr[21443]= 1449408469;
assign addr[21444]= 1558519173;
assign addr[21445]= 1659723983;
assign addr[21446]= 1752509516;
assign addr[21447]= 1836405100;
assign addr[21448]= 1910985158;
assign addr[21449]= 1975871368;
assign addr[21450]= 2030734582;
assign addr[21451]= 2075296495;
assign addr[21452]= 2109331059;
assign addr[21453]= 2132665626;
assign addr[21454]= 2145181827;
assign addr[21455]= 2146816171;
assign addr[21456]= 2137560369;
assign addr[21457]= 2117461370;
assign addr[21458]= 2086621133;
assign addr[21459]= 2045196100;
assign addr[21460]= 1993396407;
assign addr[21461]= 1931484818;
assign addr[21462]= 1859775393;
assign addr[21463]= 1778631892;
assign addr[21464]= 1688465931;
assign addr[21465]= 1589734894;
assign addr[21466]= 1482939614;
assign addr[21467]= 1368621831;
assign addr[21468]= 1247361445;
assign addr[21469]= 1119773573;
assign addr[21470]= 986505429;
assign addr[21471]= 848233042;
assign addr[21472]= 705657826;
assign addr[21473]= 559503022;
assign addr[21474]= 410510029;
assign addr[21475]= 259434643;
assign addr[21476]= 107043224;
assign addr[21477]= -45891193;
assign addr[21478]= -198592817;
assign addr[21479]= -350287041;
assign addr[21480]= -500204365;
assign addr[21481]= -647584304;
assign addr[21482]= -791679244;
assign addr[21483]= -931758235;
assign addr[21484]= -1067110699;
assign addr[21485]= -1197050035;
assign addr[21486]= -1320917099;
assign addr[21487]= -1438083551;
assign addr[21488]= -1547955041;
assign addr[21489]= -1649974225;
assign addr[21490]= -1743623590;
assign addr[21491]= -1828428082;
assign addr[21492]= -1903957513;
assign addr[21493]= -1969828744;
assign addr[21494]= -2025707632;
assign addr[21495]= -2071310720;
assign addr[21496]= -2106406677;
assign addr[21497]= -2130817471;
assign addr[21498]= -2144419275;
assign addr[21499]= -2147143090;
assign addr[21500]= -2138975100;
assign addr[21501]= -2119956737;
assign addr[21502]= -2090184478;
assign addr[21503]= -2049809346;
assign addr[21504]= -1999036154;
assign addr[21505]= -1938122457;
assign addr[21506]= -1867377253;
assign addr[21507]= -1787159411;
assign addr[21508]= -1697875851;
assign addr[21509]= -1599979481;
assign addr[21510]= -1493966902;
assign addr[21511]= -1380375881;
assign addr[21512]= -1259782632;
assign addr[21513]= -1132798888;
assign addr[21514]= -1000068799;
assign addr[21515]= -862265664;
assign addr[21516]= -720088517;
assign addr[21517]= -574258580;
assign addr[21518]= -425515602;
assign addr[21519]= -274614114;
assign addr[21520]= -122319591;
assign addr[21521]= 30595422;
assign addr[21522]= 183355234;
assign addr[21523]= 335184940;
assign addr[21524]= 485314355;
assign addr[21525]= 632981917;
assign addr[21526]= 777438554;
assign addr[21527]= 917951481;
assign addr[21528]= 1053807919;
assign addr[21529]= 1184318708;
assign addr[21530]= 1308821808;
assign addr[21531]= 1426685652;
assign addr[21532]= 1537312353;
assign addr[21533]= 1640140734;
assign addr[21534]= 1734649179;
assign addr[21535]= 1820358275;
assign addr[21536]= 1896833245;
assign addr[21537]= 1963686155;
assign addr[21538]= 2020577882;
assign addr[21539]= 2067219829;
assign addr[21540]= 2103375398;
assign addr[21541]= 2128861181;
assign addr[21542]= 2143547897;
assign addr[21543]= 2147361045;
assign addr[21544]= 2140281282;
assign addr[21545]= 2122344521;
assign addr[21546]= 2093641749;
assign addr[21547]= 2054318569;
assign addr[21548]= 2004574453;
assign addr[21549]= 1944661739;
assign addr[21550]= 1874884346;
assign addr[21551]= 1795596234;
assign addr[21552]= 1707199606;
assign addr[21553]= 1610142873;
assign addr[21554]= 1504918373;
assign addr[21555]= 1392059879;
assign addr[21556]= 1272139887;
assign addr[21557]= 1145766716;
assign addr[21558]= 1013581418;
assign addr[21559]= 876254528;
assign addr[21560]= 734482665;
assign addr[21561]= 588984994;
assign addr[21562]= 440499581;
assign addr[21563]= 289779648;
assign addr[21564]= 137589750;
assign addr[21565]= -15298099;
assign addr[21566]= -168108346;
assign addr[21567]= -320065829;
assign addr[21568]= -470399716;
assign addr[21569]= -618347408;
assign addr[21570]= -763158411;
assign addr[21571]= -904098143;
assign addr[21572]= -1040451659;
assign addr[21573]= -1171527280;
assign addr[21574]= -1296660098;
assign addr[21575]= -1415215352;
assign addr[21576]= -1526591649;
assign addr[21577]= -1630224009;
assign addr[21578]= -1725586737;
assign addr[21579]= -1812196087;
assign addr[21580]= -1889612716;
assign addr[21581]= -1957443913;
assign addr[21582]= -2015345591;
assign addr[21583]= -2063024031;
assign addr[21584]= -2100237377;
assign addr[21585]= -2126796855;
assign addr[21586]= -2142567738;
assign addr[21587]= -2147470025;
assign addr[21588]= -2141478848;
assign addr[21589]= -2124624598;
assign addr[21590]= -2096992772;
assign addr[21591]= -2058723538;
assign addr[21592]= -2010011024;
assign addr[21593]= -1951102334;
assign addr[21594]= -1882296293;
assign addr[21595]= -1803941934;
assign addr[21596]= -1716436725;
assign addr[21597]= -1620224553;
assign addr[21598]= -1515793473;
assign addr[21599]= -1403673233;
assign addr[21600]= -1284432584;
assign addr[21601]= -1158676398;
assign addr[21602]= -1027042599;
assign addr[21603]= -890198924;
assign addr[21604]= -748839539;
assign addr[21605]= -603681519;
assign addr[21606]= -455461206;
assign addr[21607]= -304930476;
assign addr[21608]= -152852926;
assign addr[21609]= 0;
assign addr[21610]= 152852926;
assign addr[21611]= 304930476;
assign addr[21612]= 455461206;
assign addr[21613]= 603681519;
assign addr[21614]= 748839539;
assign addr[21615]= 890198924;
assign addr[21616]= 1027042599;
assign addr[21617]= 1158676398;
assign addr[21618]= 1284432584;
assign addr[21619]= 1403673233;
assign addr[21620]= 1515793473;
assign addr[21621]= 1620224553;
assign addr[21622]= 1716436725;
assign addr[21623]= 1803941934;
assign addr[21624]= 1882296293;
assign addr[21625]= 1951102334;
assign addr[21626]= 2010011024;
assign addr[21627]= 2058723538;
assign addr[21628]= 2096992772;
assign addr[21629]= 2124624598;
assign addr[21630]= 2141478848;
assign addr[21631]= 2147470025;
assign addr[21632]= 2142567738;
assign addr[21633]= 2126796855;
assign addr[21634]= 2100237377;
assign addr[21635]= 2063024031;
assign addr[21636]= 2015345591;
assign addr[21637]= 1957443913;
assign addr[21638]= 1889612716;
assign addr[21639]= 1812196087;
assign addr[21640]= 1725586737;
assign addr[21641]= 1630224009;
assign addr[21642]= 1526591649;
assign addr[21643]= 1415215352;
assign addr[21644]= 1296660098;
assign addr[21645]= 1171527280;
assign addr[21646]= 1040451659;
assign addr[21647]= 904098143;
assign addr[21648]= 763158411;
assign addr[21649]= 618347408;
assign addr[21650]= 470399716;
assign addr[21651]= 320065829;
assign addr[21652]= 168108346;
assign addr[21653]= 15298099;
assign addr[21654]= -137589750;
assign addr[21655]= -289779648;
assign addr[21656]= -440499581;
assign addr[21657]= -588984994;
assign addr[21658]= -734482665;
assign addr[21659]= -876254528;
assign addr[21660]= -1013581418;
assign addr[21661]= -1145766716;
assign addr[21662]= -1272139887;
assign addr[21663]= -1392059879;
assign addr[21664]= -1504918373;
assign addr[21665]= -1610142873;
assign addr[21666]= -1707199606;
assign addr[21667]= -1795596234;
assign addr[21668]= -1874884346;
assign addr[21669]= -1944661739;
assign addr[21670]= -2004574453;
assign addr[21671]= -2054318569;
assign addr[21672]= -2093641749;
assign addr[21673]= -2122344521;
assign addr[21674]= -2140281282;
assign addr[21675]= -2147361045;
assign addr[21676]= -2143547897;
assign addr[21677]= -2128861181;
assign addr[21678]= -2103375398;
assign addr[21679]= -2067219829;
assign addr[21680]= -2020577882;
assign addr[21681]= -1963686155;
assign addr[21682]= -1896833245;
assign addr[21683]= -1820358275;
assign addr[21684]= -1734649179;
assign addr[21685]= -1640140734;
assign addr[21686]= -1537312353;
assign addr[21687]= -1426685652;
assign addr[21688]= -1308821808;
assign addr[21689]= -1184318708;
assign addr[21690]= -1053807919;
assign addr[21691]= -917951481;
assign addr[21692]= -777438554;
assign addr[21693]= -632981917;
assign addr[21694]= -485314355;
assign addr[21695]= -335184940;
assign addr[21696]= -183355234;
assign addr[21697]= -30595422;
assign addr[21698]= 122319591;
assign addr[21699]= 274614114;
assign addr[21700]= 425515602;
assign addr[21701]= 574258580;
assign addr[21702]= 720088517;
assign addr[21703]= 862265664;
assign addr[21704]= 1000068799;
assign addr[21705]= 1132798888;
assign addr[21706]= 1259782632;
assign addr[21707]= 1380375881;
assign addr[21708]= 1493966902;
assign addr[21709]= 1599979481;
assign addr[21710]= 1697875851;
assign addr[21711]= 1787159411;
assign addr[21712]= 1867377253;
assign addr[21713]= 1938122457;
assign addr[21714]= 1999036154;
assign addr[21715]= 2049809346;
assign addr[21716]= 2090184478;
assign addr[21717]= 2119956737;
assign addr[21718]= 2138975100;
assign addr[21719]= 2147143090;
assign addr[21720]= 2144419275;
assign addr[21721]= 2130817471;
assign addr[21722]= 2106406677;
assign addr[21723]= 2071310720;
assign addr[21724]= 2025707632;
assign addr[21725]= 1969828744;
assign addr[21726]= 1903957513;
assign addr[21727]= 1828428082;
assign addr[21728]= 1743623590;
assign addr[21729]= 1649974225;
assign addr[21730]= 1547955041;
assign addr[21731]= 1438083551;
assign addr[21732]= 1320917099;
assign addr[21733]= 1197050035;
assign addr[21734]= 1067110699;
assign addr[21735]= 931758235;
assign addr[21736]= 791679244;
assign addr[21737]= 647584304;
assign addr[21738]= 500204365;
assign addr[21739]= 350287041;
assign addr[21740]= 198592817;
assign addr[21741]= 45891193;
assign addr[21742]= -107043224;
assign addr[21743]= -259434643;
assign addr[21744]= -410510029;
assign addr[21745]= -559503022;
assign addr[21746]= -705657826;
assign addr[21747]= -848233042;
assign addr[21748]= -986505429;
assign addr[21749]= -1119773573;
assign addr[21750]= -1247361445;
assign addr[21751]= -1368621831;
assign addr[21752]= -1482939614;
assign addr[21753]= -1589734894;
assign addr[21754]= -1688465931;
assign addr[21755]= -1778631892;
assign addr[21756]= -1859775393;
assign addr[21757]= -1931484818;
assign addr[21758]= -1993396407;
assign addr[21759]= -2045196100;
assign addr[21760]= -2086621133;
assign addr[21761]= -2117461370;
assign addr[21762]= -2137560369;
assign addr[21763]= -2146816171;
assign addr[21764]= -2145181827;
assign addr[21765]= -2132665626;
assign addr[21766]= -2109331059;
assign addr[21767]= -2075296495;
assign addr[21768]= -2030734582;
assign addr[21769]= -1975871368;
assign addr[21770]= -1910985158;
assign addr[21771]= -1836405100;
assign addr[21772]= -1752509516;
assign addr[21773]= -1659723983;
assign addr[21774]= -1558519173;
assign addr[21775]= -1449408469;
assign addr[21776]= -1332945355;
assign addr[21777]= -1209720613;
assign addr[21778]= -1080359326;
assign addr[21779]= -945517704;
assign addr[21780]= -805879757;
assign addr[21781]= -662153826;
assign addr[21782]= -515068990;
assign addr[21783]= -365371365;
assign addr[21784]= -213820322;
assign addr[21785]= -61184634;
assign addr[21786]= 91761426;
assign addr[21787]= 244242007;
assign addr[21788]= 395483624;
assign addr[21789]= 544719071;
assign addr[21790]= 691191324;
assign addr[21791]= 834157373;
assign addr[21792]= 972891995;
assign addr[21793]= 1106691431;
assign addr[21794]= 1234876957;
assign addr[21795]= 1356798326;
assign addr[21796]= 1471837070;
assign addr[21797]= 1579409630;
assign addr[21798]= 1678970324;
assign addr[21799]= 1770014111;
assign addr[21800]= 1852079154;
assign addr[21801]= 1924749160;
assign addr[21802]= 1987655498;
assign addr[21803]= 2040479063;
assign addr[21804]= 2082951896;
assign addr[21805]= 2114858546;
assign addr[21806]= 2136037160;
assign addr[21807]= 2146380306;
assign addr[21808]= 2145835515;
assign addr[21809]= 2134405552;
assign addr[21810]= 2112148396;
assign addr[21811]= 2079176953;
assign addr[21812]= 2035658475;
assign addr[21813]= 1981813720;
assign addr[21814]= 1917915825;
assign addr[21815]= 1844288924;
assign addr[21816]= 1761306505;
assign addr[21817]= 1669389513;
assign addr[21818]= 1569004214;
assign addr[21819]= 1460659832;
assign addr[21820]= 1344905966;
assign addr[21821]= 1222329801;
assign addr[21822]= 1093553126;
assign addr[21823]= 959229189;
assign addr[21824]= 820039373;
assign addr[21825]= 676689746;
assign addr[21826]= 529907477;
assign addr[21827]= 380437148;
assign addr[21828]= 229036977;
assign addr[21829]= 76474970;
assign addr[21830]= -76474970;
assign addr[21831]= -229036977;
assign addr[21832]= -380437148;
assign addr[21833]= -529907477;
assign addr[21834]= -676689746;
assign addr[21835]= -820039373;
assign addr[21836]= -959229189;
assign addr[21837]= -1093553126;
assign addr[21838]= -1222329801;
assign addr[21839]= -1344905966;
assign addr[21840]= -1460659832;
assign addr[21841]= -1569004214;
assign addr[21842]= -1669389513;
assign addr[21843]= -1761306505;
assign addr[21844]= -1844288924;
assign addr[21845]= -1917915825;
assign addr[21846]= -1981813720;
assign addr[21847]= -2035658475;
assign addr[21848]= -2079176953;
assign addr[21849]= -2112148396;
assign addr[21850]= -2134405552;
assign addr[21851]= -2145835515;
assign addr[21852]= -2146380306;
assign addr[21853]= -2136037160;
assign addr[21854]= -2114858546;
assign addr[21855]= -2082951896;
assign addr[21856]= -2040479063;
assign addr[21857]= -1987655498;
assign addr[21858]= -1924749160;
assign addr[21859]= -1852079154;
assign addr[21860]= -1770014111;
assign addr[21861]= -1678970324;
assign addr[21862]= -1579409630;
assign addr[21863]= -1471837070;
assign addr[21864]= -1356798326;
assign addr[21865]= -1234876957;
assign addr[21866]= -1106691431;
assign addr[21867]= -972891995;
assign addr[21868]= -834157373;
assign addr[21869]= -691191324;
assign addr[21870]= -544719071;
assign addr[21871]= -395483624;
assign addr[21872]= -244242007;
assign addr[21873]= -91761426;
assign addr[21874]= 61184634;
assign addr[21875]= 213820322;
assign addr[21876]= 365371365;
assign addr[21877]= 515068990;
assign addr[21878]= 662153826;
assign addr[21879]= 805879757;
assign addr[21880]= 945517704;
assign addr[21881]= 1080359326;
assign addr[21882]= 1209720613;
assign addr[21883]= 1332945355;
assign addr[21884]= 1449408469;
assign addr[21885]= 1558519173;
assign addr[21886]= 1659723983;
assign addr[21887]= 1752509516;
assign addr[21888]= 1836405100;
assign addr[21889]= 1910985158;
assign addr[21890]= 1975871368;
assign addr[21891]= 2030734582;
assign addr[21892]= 2075296495;
assign addr[21893]= 2109331059;
assign addr[21894]= 2132665626;
assign addr[21895]= 2145181827;
assign addr[21896]= 2146816171;
assign addr[21897]= 2137560369;
assign addr[21898]= 2117461370;
assign addr[21899]= 2086621133;
assign addr[21900]= 2045196100;
assign addr[21901]= 1993396407;
assign addr[21902]= 1931484818;
assign addr[21903]= 1859775393;
assign addr[21904]= 1778631892;
assign addr[21905]= 1688465931;
assign addr[21906]= 1589734894;
assign addr[21907]= 1482939614;
assign addr[21908]= 1368621831;
assign addr[21909]= 1247361445;
assign addr[21910]= 1119773573;
assign addr[21911]= 986505429;
assign addr[21912]= 848233042;
assign addr[21913]= 705657826;
assign addr[21914]= 559503022;
assign addr[21915]= 410510029;
assign addr[21916]= 259434643;
assign addr[21917]= 107043224;
assign addr[21918]= -45891193;
assign addr[21919]= -198592817;
assign addr[21920]= -350287041;
assign addr[21921]= -500204365;
assign addr[21922]= -647584304;
assign addr[21923]= -791679244;
assign addr[21924]= -931758235;
assign addr[21925]= -1067110699;
assign addr[21926]= -1197050035;
assign addr[21927]= -1320917099;
assign addr[21928]= -1438083551;
assign addr[21929]= -1547955041;
assign addr[21930]= -1649974225;
assign addr[21931]= -1743623590;
assign addr[21932]= -1828428082;
assign addr[21933]= -1903957513;
assign addr[21934]= -1969828744;
assign addr[21935]= -2025707632;
assign addr[21936]= -2071310720;
assign addr[21937]= -2106406677;
assign addr[21938]= -2130817471;
assign addr[21939]= -2144419275;
assign addr[21940]= -2147143090;
assign addr[21941]= -2138975100;
assign addr[21942]= -2119956737;
assign addr[21943]= -2090184478;
assign addr[21944]= -2049809346;
assign addr[21945]= -1999036154;
assign addr[21946]= -1938122457;
assign addr[21947]= -1867377253;
assign addr[21948]= -1787159411;
assign addr[21949]= -1697875851;
assign addr[21950]= -1599979481;
assign addr[21951]= -1493966902;
assign addr[21952]= -1380375881;
assign addr[21953]= -1259782632;
assign addr[21954]= -1132798888;
assign addr[21955]= -1000068799;
assign addr[21956]= -862265664;
assign addr[21957]= -720088517;
assign addr[21958]= -574258580;
assign addr[21959]= -425515602;
assign addr[21960]= -274614114;
assign addr[21961]= -122319591;
assign addr[21962]= 30595422;
assign addr[21963]= 183355234;
assign addr[21964]= 335184940;
assign addr[21965]= 485314355;
assign addr[21966]= 632981917;
assign addr[21967]= 777438554;
assign addr[21968]= 917951481;
assign addr[21969]= 1053807919;
assign addr[21970]= 1184318708;
assign addr[21971]= 1308821808;
assign addr[21972]= 1426685652;
assign addr[21973]= 1537312353;
assign addr[21974]= 1640140734;
assign addr[21975]= 1734649179;
assign addr[21976]= 1820358275;
assign addr[21977]= 1896833245;
assign addr[21978]= 1963686155;
assign addr[21979]= 2020577882;
assign addr[21980]= 2067219829;
assign addr[21981]= 2103375398;
assign addr[21982]= 2128861181;
assign addr[21983]= 2143547897;
assign addr[21984]= 2147361045;
assign addr[21985]= 2140281282;
assign addr[21986]= 2122344521;
assign addr[21987]= 2093641749;
assign addr[21988]= 2054318569;
assign addr[21989]= 2004574453;
assign addr[21990]= 1944661739;
assign addr[21991]= 1874884346;
assign addr[21992]= 1795596234;
assign addr[21993]= 1707199606;
assign addr[21994]= 1610142873;
assign addr[21995]= 1504918373;
assign addr[21996]= 1392059879;
assign addr[21997]= 1272139887;
assign addr[21998]= 1145766716;
assign addr[21999]= 1013581418;
assign addr[22000]= 876254528;
assign addr[22001]= 734482665;
assign addr[22002]= 588984994;
assign addr[22003]= 440499581;
assign addr[22004]= 289779648;
assign addr[22005]= 137589750;
assign addr[22006]= -15298099;
assign addr[22007]= -168108346;
assign addr[22008]= -320065829;
assign addr[22009]= -470399716;
assign addr[22010]= -618347408;
assign addr[22011]= -763158411;
assign addr[22012]= -904098143;
assign addr[22013]= -1040451659;
assign addr[22014]= -1171527280;
assign addr[22015]= -1296660098;
assign addr[22016]= -1415215352;
assign addr[22017]= -1526591649;
assign addr[22018]= -1630224009;
assign addr[22019]= -1725586737;
assign addr[22020]= -1812196087;
assign addr[22021]= -1889612716;
assign addr[22022]= -1957443913;
assign addr[22023]= -2015345591;
assign addr[22024]= -2063024031;
assign addr[22025]= -2100237377;
assign addr[22026]= -2126796855;
assign addr[22027]= -2142567738;
assign addr[22028]= -2147470025;
assign addr[22029]= -2141478848;
assign addr[22030]= -2124624598;
assign addr[22031]= -2096992772;
assign addr[22032]= -2058723538;
assign addr[22033]= -2010011024;
assign addr[22034]= -1951102334;
assign addr[22035]= -1882296293;
assign addr[22036]= -1803941934;
assign addr[22037]= -1716436725;
assign addr[22038]= -1620224553;
assign addr[22039]= -1515793473;
assign addr[22040]= -1403673233;
assign addr[22041]= -1284432584;
assign addr[22042]= -1158676398;
assign addr[22043]= -1027042599;
assign addr[22044]= -890198924;
assign addr[22045]= -748839539;
assign addr[22046]= -603681519;
assign addr[22047]= -455461206;
assign addr[22048]= -304930476;
assign addr[22049]= -152852926;
assign addr[22050]= 0;
assign addr[22051]= 152852926;
assign addr[22052]= 304930476;
assign addr[22053]= 455461206;
assign addr[22054]= 603681519;
assign addr[22055]= 748839539;
assign addr[22056]= 890198924;
assign addr[22057]= 1027042599;
assign addr[22058]= 1158676398;
assign addr[22059]= 1284432584;
assign addr[22060]= 1403673233;
assign addr[22061]= 1515793473;
assign addr[22062]= 1620224553;
assign addr[22063]= 1716436725;
assign addr[22064]= 1803941934;
assign addr[22065]= 1882296293;
assign addr[22066]= 1951102334;
assign addr[22067]= 2010011024;
assign addr[22068]= 2058723538;
assign addr[22069]= 2096992772;
assign addr[22070]= 2124624598;
assign addr[22071]= 2141478848;
assign addr[22072]= 2147470025;
assign addr[22073]= 2142567738;
assign addr[22074]= 2126796855;
assign addr[22075]= 2100237377;
assign addr[22076]= 2063024031;
assign addr[22077]= 2015345591;
assign addr[22078]= 1957443913;
assign addr[22079]= 1889612716;
assign addr[22080]= 1812196087;
assign addr[22081]= 1725586737;
assign addr[22082]= 1630224009;
assign addr[22083]= 1526591649;
assign addr[22084]= 1415215352;
assign addr[22085]= 1296660098;
assign addr[22086]= 1171527280;
assign addr[22087]= 1040451659;
assign addr[22088]= 904098143;
assign addr[22089]= 763158411;
assign addr[22090]= 618347408;
assign addr[22091]= 470399716;
assign addr[22092]= 320065829;
assign addr[22093]= 168108346;
assign addr[22094]= 15298099;
assign addr[22095]= -137589750;
assign addr[22096]= -289779648;
assign addr[22097]= -440499581;
assign addr[22098]= -588984994;
assign addr[22099]= -734482665;
assign addr[22100]= -876254528;
assign addr[22101]= -1013581418;
assign addr[22102]= -1145766716;
assign addr[22103]= -1272139887;
assign addr[22104]= -1392059879;
assign addr[22105]= -1504918373;
assign addr[22106]= -1610142873;
assign addr[22107]= -1707199606;
assign addr[22108]= -1795596234;
assign addr[22109]= -1874884346;
assign addr[22110]= -1944661739;
assign addr[22111]= -2004574453;
assign addr[22112]= -2054318569;
assign addr[22113]= -2093641749;
assign addr[22114]= -2122344521;
assign addr[22115]= -2140281282;
assign addr[22116]= -2147361045;
assign addr[22117]= -2143547897;
assign addr[22118]= -2128861181;
assign addr[22119]= -2103375398;
assign addr[22120]= -2067219829;
assign addr[22121]= -2020577882;
assign addr[22122]= -1963686155;
assign addr[22123]= -1896833245;
assign addr[22124]= -1820358275;
assign addr[22125]= -1734649179;
assign addr[22126]= -1640140734;
assign addr[22127]= -1537312353;
assign addr[22128]= -1426685652;
assign addr[22129]= -1308821808;
assign addr[22130]= -1184318708;
assign addr[22131]= -1053807919;
assign addr[22132]= -917951481;
assign addr[22133]= -777438554;
assign addr[22134]= -632981917;
assign addr[22135]= -485314355;
assign addr[22136]= -335184940;
assign addr[22137]= -183355234;
assign addr[22138]= -30595422;
assign addr[22139]= 122319591;
assign addr[22140]= 274614114;
assign addr[22141]= 425515602;
assign addr[22142]= 574258580;
assign addr[22143]= 720088517;
assign addr[22144]= 862265664;
assign addr[22145]= 1000068799;
assign addr[22146]= 1132798888;
assign addr[22147]= 1259782632;
assign addr[22148]= 1380375881;
assign addr[22149]= 1493966902;
assign addr[22150]= 1599979481;
assign addr[22151]= 1697875851;
assign addr[22152]= 1787159411;
assign addr[22153]= 1867377253;
assign addr[22154]= 1938122457;
assign addr[22155]= 1999036154;
assign addr[22156]= 2049809346;
assign addr[22157]= 2090184478;
assign addr[22158]= 2119956737;
assign addr[22159]= 2138975100;
assign addr[22160]= 2147143090;
assign addr[22161]= 2144419275;
assign addr[22162]= 2130817471;
assign addr[22163]= 2106406677;
assign addr[22164]= 2071310720;
assign addr[22165]= 2025707632;
assign addr[22166]= 1969828744;
assign addr[22167]= 1903957513;
assign addr[22168]= 1828428082;
assign addr[22169]= 1743623590;
assign addr[22170]= 1649974225;
assign addr[22171]= 1547955041;
assign addr[22172]= 1438083551;
assign addr[22173]= 1320917099;
assign addr[22174]= 1197050035;
assign addr[22175]= 1067110699;
assign addr[22176]= 931758235;
assign addr[22177]= 791679244;
assign addr[22178]= 647584304;
assign addr[22179]= 500204365;
assign addr[22180]= 350287041;
assign addr[22181]= 198592817;
assign addr[22182]= 45891193;
assign addr[22183]= -107043224;
assign addr[22184]= -259434643;
assign addr[22185]= -410510029;
assign addr[22186]= -559503022;
assign addr[22187]= -705657826;
assign addr[22188]= -848233042;
assign addr[22189]= -986505429;
assign addr[22190]= -1119773573;
assign addr[22191]= -1247361445;
assign addr[22192]= -1368621831;
assign addr[22193]= -1482939614;
assign addr[22194]= -1589734894;
assign addr[22195]= -1688465931;
assign addr[22196]= -1778631892;
assign addr[22197]= -1859775393;
assign addr[22198]= -1931484818;
assign addr[22199]= -1993396407;
assign addr[22200]= -2045196100;
assign addr[22201]= -2086621133;
assign addr[22202]= -2117461370;
assign addr[22203]= -2137560369;
assign addr[22204]= -2146816171;
assign addr[22205]= -2145181827;
assign addr[22206]= -2132665626;
assign addr[22207]= -2109331059;
assign addr[22208]= -2075296495;
assign addr[22209]= -2030734582;
assign addr[22210]= -1975871368;
assign addr[22211]= -1910985158;
assign addr[22212]= -1836405100;
assign addr[22213]= -1752509516;
assign addr[22214]= -1659723983;
assign addr[22215]= -1558519173;
assign addr[22216]= -1449408469;
assign addr[22217]= -1332945355;
assign addr[22218]= -1209720613;
assign addr[22219]= -1080359326;
assign addr[22220]= -945517704;
assign addr[22221]= -805879757;
assign addr[22222]= -662153826;
assign addr[22223]= -515068990;
assign addr[22224]= -365371365;
assign addr[22225]= -213820322;
assign addr[22226]= -61184634;
assign addr[22227]= 91761426;
assign addr[22228]= 244242007;
assign addr[22229]= 395483624;
assign addr[22230]= 544719071;
assign addr[22231]= 691191324;
assign addr[22232]= 834157373;
assign addr[22233]= 972891995;
assign addr[22234]= 1106691431;
assign addr[22235]= 1234876957;
assign addr[22236]= 1356798326;
assign addr[22237]= 1471837070;
assign addr[22238]= 1579409630;
assign addr[22239]= 1678970324;
assign addr[22240]= 1770014111;
assign addr[22241]= 1852079154;
assign addr[22242]= 1924749160;
assign addr[22243]= 1987655498;
assign addr[22244]= 2040479063;
assign addr[22245]= 2082951896;
assign addr[22246]= 2114858546;
assign addr[22247]= 2136037160;
assign addr[22248]= 2146380306;
assign addr[22249]= 2145835515;
assign addr[22250]= 2134405552;
assign addr[22251]= 2112148396;
assign addr[22252]= 2079176953;
assign addr[22253]= 2035658475;
assign addr[22254]= 1981813720;
assign addr[22255]= 1917915825;
assign addr[22256]= 1844288924;
assign addr[22257]= 1761306505;
assign addr[22258]= 1669389513;
assign addr[22259]= 1569004214;
assign addr[22260]= 1460659832;
assign addr[22261]= 1344905966;
assign addr[22262]= 1222329801;
assign addr[22263]= 1093553126;
assign addr[22264]= 959229189;
assign addr[22265]= 820039373;
assign addr[22266]= 676689746;
assign addr[22267]= 529907477;
assign addr[22268]= 380437148;
assign addr[22269]= 229036977;
assign addr[22270]= 76474970;
assign addr[22271]= -76474970;
assign addr[22272]= -229036977;
assign addr[22273]= -380437148;
assign addr[22274]= -529907477;
assign addr[22275]= -676689746;
assign addr[22276]= -820039373;
assign addr[22277]= -959229189;
assign addr[22278]= -1093553126;
assign addr[22279]= -1222329801;
assign addr[22280]= -1344905966;
assign addr[22281]= -1460659832;
assign addr[22282]= -1569004214;
assign addr[22283]= -1669389513;
assign addr[22284]= -1761306505;
assign addr[22285]= -1844288924;
assign addr[22286]= -1917915825;
assign addr[22287]= -1981813720;
assign addr[22288]= -2035658475;
assign addr[22289]= -2079176953;
assign addr[22290]= -2112148396;
assign addr[22291]= -2134405552;
assign addr[22292]= -2145835515;
assign addr[22293]= -2146380306;
assign addr[22294]= -2136037160;
assign addr[22295]= -2114858546;
assign addr[22296]= -2082951896;
assign addr[22297]= -2040479063;
assign addr[22298]= -1987655498;
assign addr[22299]= -1924749160;
assign addr[22300]= -1852079154;
assign addr[22301]= -1770014111;
assign addr[22302]= -1678970324;
assign addr[22303]= -1579409630;
assign addr[22304]= -1471837070;
assign addr[22305]= -1356798326;
assign addr[22306]= -1234876957;
assign addr[22307]= -1106691431;
assign addr[22308]= -972891995;
assign addr[22309]= -834157373;
assign addr[22310]= -691191324;
assign addr[22311]= -544719071;
assign addr[22312]= -395483624;
assign addr[22313]= -244242007;
assign addr[22314]= -91761426;
assign addr[22315]= 61184634;
assign addr[22316]= 213820322;
assign addr[22317]= 365371365;
assign addr[22318]= 515068990;
assign addr[22319]= 662153826;
assign addr[22320]= 805879757;
assign addr[22321]= 945517704;
assign addr[22322]= 1080359326;
assign addr[22323]= 1209720613;
assign addr[22324]= 1332945355;
assign addr[22325]= 1449408469;
assign addr[22326]= 1558519173;
assign addr[22327]= 1659723983;
assign addr[22328]= 1752509516;
assign addr[22329]= 1836405100;
assign addr[22330]= 1910985158;
assign addr[22331]= 1975871368;
assign addr[22332]= 2030734582;
assign addr[22333]= 2075296495;
assign addr[22334]= 2109331059;
assign addr[22335]= 2132665626;
assign addr[22336]= 2145181827;
assign addr[22337]= 2146816171;
assign addr[22338]= 2137560369;
assign addr[22339]= 2117461370;
assign addr[22340]= 2086621133;
assign addr[22341]= 2045196100;
assign addr[22342]= 1993396407;
assign addr[22343]= 1931484818;
assign addr[22344]= 1859775393;
assign addr[22345]= 1778631892;
assign addr[22346]= 1688465931;
assign addr[22347]= 1589734894;
assign addr[22348]= 1482939614;
assign addr[22349]= 1368621831;
assign addr[22350]= 1247361445;
assign addr[22351]= 1119773573;
assign addr[22352]= 986505429;
assign addr[22353]= 848233042;
assign addr[22354]= 705657826;
assign addr[22355]= 559503022;
assign addr[22356]= 410510029;
assign addr[22357]= 259434643;
assign addr[22358]= 107043224;
assign addr[22359]= -45891193;
assign addr[22360]= -198592817;
assign addr[22361]= -350287041;
assign addr[22362]= -500204365;
assign addr[22363]= -647584304;
assign addr[22364]= -791679244;
assign addr[22365]= -931758235;
assign addr[22366]= -1067110699;
assign addr[22367]= -1197050035;
assign addr[22368]= -1320917099;
assign addr[22369]= -1438083551;
assign addr[22370]= -1547955041;
assign addr[22371]= -1649974225;
assign addr[22372]= -1743623590;
assign addr[22373]= -1828428082;
assign addr[22374]= -1903957513;
assign addr[22375]= -1969828744;
assign addr[22376]= -2025707632;
assign addr[22377]= -2071310720;
assign addr[22378]= -2106406677;
assign addr[22379]= -2130817471;
assign addr[22380]= -2144419275;
assign addr[22381]= -2147143090;
assign addr[22382]= -2138975100;
assign addr[22383]= -2119956737;
assign addr[22384]= -2090184478;
assign addr[22385]= -2049809346;
assign addr[22386]= -1999036154;
assign addr[22387]= -1938122457;
assign addr[22388]= -1867377253;
assign addr[22389]= -1787159411;
assign addr[22390]= -1697875851;
assign addr[22391]= -1599979481;
assign addr[22392]= -1493966902;
assign addr[22393]= -1380375881;
assign addr[22394]= -1259782632;
assign addr[22395]= -1132798888;
assign addr[22396]= -1000068799;
assign addr[22397]= -862265664;
assign addr[22398]= -720088517;
assign addr[22399]= -574258580;
assign addr[22400]= -425515602;
assign addr[22401]= -274614114;
assign addr[22402]= -122319591;
assign addr[22403]= 30595422;
assign addr[22404]= 183355234;
assign addr[22405]= 335184940;
assign addr[22406]= 485314355;
assign addr[22407]= 632981917;
assign addr[22408]= 777438554;
assign addr[22409]= 917951481;
assign addr[22410]= 1053807919;
assign addr[22411]= 1184318708;
assign addr[22412]= 1308821808;
assign addr[22413]= 1426685652;
assign addr[22414]= 1537312353;
assign addr[22415]= 1640140734;
assign addr[22416]= 1734649179;
assign addr[22417]= 1820358275;
assign addr[22418]= 1896833245;
assign addr[22419]= 1963686155;
assign addr[22420]= 2020577882;
assign addr[22421]= 2067219829;
assign addr[22422]= 2103375398;
assign addr[22423]= 2128861181;
assign addr[22424]= 2143547897;
assign addr[22425]= 2147361045;
assign addr[22426]= 2140281282;
assign addr[22427]= 2122344521;
assign addr[22428]= 2093641749;
assign addr[22429]= 2054318569;
assign addr[22430]= 2004574453;
assign addr[22431]= 1944661739;
assign addr[22432]= 1874884346;
assign addr[22433]= 1795596234;
assign addr[22434]= 1707199606;
assign addr[22435]= 1610142873;
assign addr[22436]= 1504918373;
assign addr[22437]= 1392059879;
assign addr[22438]= 1272139887;
assign addr[22439]= 1145766716;
assign addr[22440]= 1013581418;
assign addr[22441]= 876254528;
assign addr[22442]= 734482665;
assign addr[22443]= 588984994;
assign addr[22444]= 440499581;
assign addr[22445]= 289779648;
assign addr[22446]= 137589750;
assign addr[22447]= -15298099;
assign addr[22448]= -168108346;
assign addr[22449]= -320065829;
assign addr[22450]= -470399716;
assign addr[22451]= -618347408;
assign addr[22452]= -763158411;
assign addr[22453]= -904098143;
assign addr[22454]= -1040451659;
assign addr[22455]= -1171527280;
assign addr[22456]= -1296660098;
assign addr[22457]= -1415215352;
assign addr[22458]= -1526591649;
assign addr[22459]= -1630224009;
assign addr[22460]= -1725586737;
assign addr[22461]= -1812196087;
assign addr[22462]= -1889612716;
assign addr[22463]= -1957443913;
assign addr[22464]= -2015345591;
assign addr[22465]= -2063024031;
assign addr[22466]= -2100237377;
assign addr[22467]= -2126796855;
assign addr[22468]= -2142567738;
assign addr[22469]= -2147470025;
assign addr[22470]= -2141478848;
assign addr[22471]= -2124624598;
assign addr[22472]= -2096992772;
assign addr[22473]= -2058723538;
assign addr[22474]= -2010011024;
assign addr[22475]= -1951102334;
assign addr[22476]= -1882296293;
assign addr[22477]= -1803941934;
assign addr[22478]= -1716436725;
assign addr[22479]= -1620224553;
assign addr[22480]= -1515793473;
assign addr[22481]= -1403673233;
assign addr[22482]= -1284432584;
assign addr[22483]= -1158676398;
assign addr[22484]= -1027042599;
assign addr[22485]= -890198924;
assign addr[22486]= -748839539;
assign addr[22487]= -603681519;
assign addr[22488]= -455461206;
assign addr[22489]= -304930476;
assign addr[22490]= -152852926;
assign addr[22491]= 0;
assign addr[22492]= 152852926;
assign addr[22493]= 304930476;
assign addr[22494]= 455461206;
assign addr[22495]= 603681519;
assign addr[22496]= 748839539;
assign addr[22497]= 890198924;
assign addr[22498]= 1027042599;
assign addr[22499]= 1158676398;
assign addr[22500]= 1284432584;
assign addr[22501]= 1403673233;
assign addr[22502]= 1515793473;
assign addr[22503]= 1620224553;
assign addr[22504]= 1716436725;
assign addr[22505]= 1803941934;
assign addr[22506]= 1882296293;
assign addr[22507]= 1951102334;
assign addr[22508]= 2010011024;
assign addr[22509]= 2058723538;
assign addr[22510]= 2096992772;
assign addr[22511]= 2124624598;
assign addr[22512]= 2141478848;
assign addr[22513]= 2147470025;
assign addr[22514]= 2142567738;
assign addr[22515]= 2126796855;
assign addr[22516]= 2100237377;
assign addr[22517]= 2063024031;
assign addr[22518]= 2015345591;
assign addr[22519]= 1957443913;
assign addr[22520]= 1889612716;
assign addr[22521]= 1812196087;
assign addr[22522]= 1725586737;
assign addr[22523]= 1630224009;
assign addr[22524]= 1526591649;
assign addr[22525]= 1415215352;
assign addr[22526]= 1296660098;
assign addr[22527]= 1171527280;
assign addr[22528]= 1040451659;
assign addr[22529]= 904098143;
assign addr[22530]= 763158411;
assign addr[22531]= 618347408;
assign addr[22532]= 470399716;
assign addr[22533]= 320065829;
assign addr[22534]= 168108346;
assign addr[22535]= 15298099;
assign addr[22536]= -137589750;
assign addr[22537]= -289779648;
assign addr[22538]= -440499581;
assign addr[22539]= -588984994;
assign addr[22540]= -734482665;
assign addr[22541]= -876254528;
assign addr[22542]= -1013581418;
assign addr[22543]= -1145766716;
assign addr[22544]= -1272139887;
assign addr[22545]= -1392059879;
assign addr[22546]= -1504918373;
assign addr[22547]= -1610142873;
assign addr[22548]= -1707199606;
assign addr[22549]= -1795596234;
assign addr[22550]= -1874884346;
assign addr[22551]= -1944661739;
assign addr[22552]= -2004574453;
assign addr[22553]= -2054318569;
assign addr[22554]= -2093641749;
assign addr[22555]= -2122344521;
assign addr[22556]= -2140281282;
assign addr[22557]= -2147361045;
assign addr[22558]= -2143547897;
assign addr[22559]= -2128861181;
assign addr[22560]= -2103375398;
assign addr[22561]= -2067219829;
assign addr[22562]= -2020577882;
assign addr[22563]= -1963686155;
assign addr[22564]= -1896833245;
assign addr[22565]= -1820358275;
assign addr[22566]= -1734649179;
assign addr[22567]= -1640140734;
assign addr[22568]= -1537312353;
assign addr[22569]= -1426685652;
assign addr[22570]= -1308821808;
assign addr[22571]= -1184318708;
assign addr[22572]= -1053807919;
assign addr[22573]= -917951481;
assign addr[22574]= -777438554;
assign addr[22575]= -632981917;
assign addr[22576]= -485314355;
assign addr[22577]= -335184940;
assign addr[22578]= -183355234;
assign addr[22579]= -30595422;
assign addr[22580]= 122319591;
assign addr[22581]= 274614114;
assign addr[22582]= 425515602;
assign addr[22583]= 574258580;
assign addr[22584]= 720088517;
assign addr[22585]= 862265664;
assign addr[22586]= 1000068799;
assign addr[22587]= 1132798888;
assign addr[22588]= 1259782632;
assign addr[22589]= 1380375881;
assign addr[22590]= 1493966902;
assign addr[22591]= 1599979481;
assign addr[22592]= 1697875851;
assign addr[22593]= 1787159411;
assign addr[22594]= 1867377253;
assign addr[22595]= 1938122457;
assign addr[22596]= 1999036154;
assign addr[22597]= 2049809346;
assign addr[22598]= 2090184478;
assign addr[22599]= 2119956737;
assign addr[22600]= 2138975100;
assign addr[22601]= 2147143090;
assign addr[22602]= 2144419275;
assign addr[22603]= 2130817471;
assign addr[22604]= 2106406677;
assign addr[22605]= 2071310720;
assign addr[22606]= 2025707632;
assign addr[22607]= 1969828744;
assign addr[22608]= 1903957513;
assign addr[22609]= 1828428082;
assign addr[22610]= 1743623590;
assign addr[22611]= 1649974225;
assign addr[22612]= 1547955041;
assign addr[22613]= 1438083551;
assign addr[22614]= 1320917099;
assign addr[22615]= 1197050035;
assign addr[22616]= 1067110699;
assign addr[22617]= 931758235;
assign addr[22618]= 791679244;
assign addr[22619]= 647584304;
assign addr[22620]= 500204365;
assign addr[22621]= 350287041;
assign addr[22622]= 198592817;
assign addr[22623]= 45891193;
assign addr[22624]= -107043224;
assign addr[22625]= -259434643;
assign addr[22626]= -410510029;
assign addr[22627]= -559503022;
assign addr[22628]= -705657826;
assign addr[22629]= -848233042;
assign addr[22630]= -986505429;
assign addr[22631]= -1119773573;
assign addr[22632]= -1247361445;
assign addr[22633]= -1368621831;
assign addr[22634]= -1482939614;
assign addr[22635]= -1589734894;
assign addr[22636]= -1688465931;
assign addr[22637]= -1778631892;
assign addr[22638]= -1859775393;
assign addr[22639]= -1931484818;
assign addr[22640]= -1993396407;
assign addr[22641]= -2045196100;
assign addr[22642]= -2086621133;
assign addr[22643]= -2117461370;
assign addr[22644]= -2137560369;
assign addr[22645]= -2146816171;
assign addr[22646]= -2145181827;
assign addr[22647]= -2132665626;
assign addr[22648]= -2109331059;
assign addr[22649]= -2075296495;
assign addr[22650]= -2030734582;
assign addr[22651]= -1975871368;
assign addr[22652]= -1910985158;
assign addr[22653]= -1836405100;
assign addr[22654]= -1752509516;
assign addr[22655]= -1659723983;
assign addr[22656]= -1558519173;
assign addr[22657]= -1449408469;
assign addr[22658]= -1332945355;
assign addr[22659]= -1209720613;
assign addr[22660]= -1080359326;
assign addr[22661]= -945517704;
assign addr[22662]= -805879757;
assign addr[22663]= -662153826;
assign addr[22664]= -515068990;
assign addr[22665]= -365371365;
assign addr[22666]= -213820322;
assign addr[22667]= -61184634;
assign addr[22668]= 91761426;
assign addr[22669]= 244242007;
assign addr[22670]= 395483624;
assign addr[22671]= 544719071;
assign addr[22672]= 691191324;
assign addr[22673]= 834157373;
assign addr[22674]= 972891995;
assign addr[22675]= 1106691431;
assign addr[22676]= 1234876957;
assign addr[22677]= 1356798326;
assign addr[22678]= 1471837070;
assign addr[22679]= 1579409630;
assign addr[22680]= 1678970324;
assign addr[22681]= 1770014111;
assign addr[22682]= 1852079154;
assign addr[22683]= 1924749160;
assign addr[22684]= 1987655498;
assign addr[22685]= 2040479063;
assign addr[22686]= 2082951896;
assign addr[22687]= 2114858546;
assign addr[22688]= 2136037160;
assign addr[22689]= 2146380306;
assign addr[22690]= 2145835515;
assign addr[22691]= 2134405552;
assign addr[22692]= 2112148396;
assign addr[22693]= 2079176953;
assign addr[22694]= 2035658475;
assign addr[22695]= 1981813720;
assign addr[22696]= 1917915825;
assign addr[22697]= 1844288924;
assign addr[22698]= 1761306505;
assign addr[22699]= 1669389513;
assign addr[22700]= 1569004214;
assign addr[22701]= 1460659832;
assign addr[22702]= 1344905966;
assign addr[22703]= 1222329801;
assign addr[22704]= 1093553126;
assign addr[22705]= 959229189;
assign addr[22706]= 820039373;
assign addr[22707]= 676689746;
assign addr[22708]= 529907477;
assign addr[22709]= 380437148;
assign addr[22710]= 229036977;
assign addr[22711]= 76474970;
assign addr[22712]= -76474970;
assign addr[22713]= -229036977;
assign addr[22714]= -380437148;
assign addr[22715]= -529907477;
assign addr[22716]= -676689746;
assign addr[22717]= -820039373;
assign addr[22718]= -959229189;
assign addr[22719]= -1093553126;
assign addr[22720]= -1222329801;
assign addr[22721]= -1344905966;
assign addr[22722]= -1460659832;
assign addr[22723]= -1569004214;
assign addr[22724]= -1669389513;
assign addr[22725]= -1761306505;
assign addr[22726]= -1844288924;
assign addr[22727]= -1917915825;
assign addr[22728]= -1981813720;
assign addr[22729]= -2035658475;
assign addr[22730]= -2079176953;
assign addr[22731]= -2112148396;
assign addr[22732]= -2134405552;
assign addr[22733]= -2145835515;
assign addr[22734]= -2146380306;
assign addr[22735]= -2136037160;
assign addr[22736]= -2114858546;
assign addr[22737]= -2082951896;
assign addr[22738]= -2040479063;
assign addr[22739]= -1987655498;
assign addr[22740]= -1924749160;
assign addr[22741]= -1852079154;
assign addr[22742]= -1770014111;
assign addr[22743]= -1678970324;
assign addr[22744]= -1579409630;
assign addr[22745]= -1471837070;
assign addr[22746]= -1356798326;
assign addr[22747]= -1234876957;
assign addr[22748]= -1106691431;
assign addr[22749]= -972891995;
assign addr[22750]= -834157373;
assign addr[22751]= -691191324;
assign addr[22752]= -544719071;
assign addr[22753]= -395483624;
assign addr[22754]= -244242007;
assign addr[22755]= -91761426;
assign addr[22756]= 61184634;
assign addr[22757]= 213820322;
assign addr[22758]= 365371365;
assign addr[22759]= 515068990;
assign addr[22760]= 662153826;
assign addr[22761]= 805879757;
assign addr[22762]= 945517704;
assign addr[22763]= 1080359326;
assign addr[22764]= 1209720613;
assign addr[22765]= 1332945355;
assign addr[22766]= 1449408469;
assign addr[22767]= 1558519173;
assign addr[22768]= 1659723983;
assign addr[22769]= 1752509516;
assign addr[22770]= 1836405100;
assign addr[22771]= 1910985158;
assign addr[22772]= 1975871368;
assign addr[22773]= 2030734582;
assign addr[22774]= 2075296495;
assign addr[22775]= 2109331059;
assign addr[22776]= 2132665626;
assign addr[22777]= 2145181827;
assign addr[22778]= 2146816171;
assign addr[22779]= 2137560369;
assign addr[22780]= 2117461370;
assign addr[22781]= 2086621133;
assign addr[22782]= 2045196100;
assign addr[22783]= 1993396407;
assign addr[22784]= 1931484818;
assign addr[22785]= 1859775393;
assign addr[22786]= 1778631892;
assign addr[22787]= 1688465931;
assign addr[22788]= 1589734894;
assign addr[22789]= 1482939614;
assign addr[22790]= 1368621831;
assign addr[22791]= 1247361445;
assign addr[22792]= 1119773573;
assign addr[22793]= 986505429;
assign addr[22794]= 848233042;
assign addr[22795]= 705657826;
assign addr[22796]= 559503022;
assign addr[22797]= 410510029;
assign addr[22798]= 259434643;
assign addr[22799]= 107043224;
assign addr[22800]= -45891193;
assign addr[22801]= -198592817;
assign addr[22802]= -350287041;
assign addr[22803]= -500204365;
assign addr[22804]= -647584304;
assign addr[22805]= -791679244;
assign addr[22806]= -931758235;
assign addr[22807]= -1067110699;
assign addr[22808]= -1197050035;
assign addr[22809]= -1320917099;
assign addr[22810]= -1438083551;
assign addr[22811]= -1547955041;
assign addr[22812]= -1649974225;
assign addr[22813]= -1743623590;
assign addr[22814]= -1828428082;
assign addr[22815]= -1903957513;
assign addr[22816]= -1969828744;
assign addr[22817]= -2025707632;
assign addr[22818]= -2071310720;
assign addr[22819]= -2106406677;
assign addr[22820]= -2130817471;
assign addr[22821]= -2144419275;
assign addr[22822]= -2147143090;
assign addr[22823]= -2138975100;
assign addr[22824]= -2119956737;
assign addr[22825]= -2090184478;
assign addr[22826]= -2049809346;
assign addr[22827]= -1999036154;
assign addr[22828]= -1938122457;
assign addr[22829]= -1867377253;
assign addr[22830]= -1787159411;
assign addr[22831]= -1697875851;
assign addr[22832]= -1599979481;
assign addr[22833]= -1493966902;
assign addr[22834]= -1380375881;
assign addr[22835]= -1259782632;
assign addr[22836]= -1132798888;
assign addr[22837]= -1000068799;
assign addr[22838]= -862265664;
assign addr[22839]= -720088517;
assign addr[22840]= -574258580;
assign addr[22841]= -425515602;
assign addr[22842]= -274614114;
assign addr[22843]= -122319591;
assign addr[22844]= 30595422;
assign addr[22845]= 183355234;
assign addr[22846]= 335184940;
assign addr[22847]= 485314355;
assign addr[22848]= 632981917;
assign addr[22849]= 777438554;
assign addr[22850]= 917951481;
assign addr[22851]= 1053807919;
assign addr[22852]= 1184318708;
assign addr[22853]= 1308821808;
assign addr[22854]= 1426685652;
assign addr[22855]= 1537312353;
assign addr[22856]= 1640140734;
assign addr[22857]= 1734649179;
assign addr[22858]= 1820358275;
assign addr[22859]= 1896833245;
assign addr[22860]= 1963686155;
assign addr[22861]= 2020577882;
assign addr[22862]= 2067219829;
assign addr[22863]= 2103375398;
assign addr[22864]= 2128861181;
assign addr[22865]= 2143547897;
assign addr[22866]= 2147361045;
assign addr[22867]= 2140281282;
assign addr[22868]= 2122344521;
assign addr[22869]= 2093641749;
assign addr[22870]= 2054318569;
assign addr[22871]= 2004574453;
assign addr[22872]= 1944661739;
assign addr[22873]= 1874884346;
assign addr[22874]= 1795596234;
assign addr[22875]= 1707199606;
assign addr[22876]= 1610142873;
assign addr[22877]= 1504918373;
assign addr[22878]= 1392059879;
assign addr[22879]= 1272139887;
assign addr[22880]= 1145766716;
assign addr[22881]= 1013581418;
assign addr[22882]= 876254528;
assign addr[22883]= 734482665;
assign addr[22884]= 588984994;
assign addr[22885]= 440499581;
assign addr[22886]= 289779648;
assign addr[22887]= 137589750;
assign addr[22888]= -15298099;
assign addr[22889]= -168108346;
assign addr[22890]= -320065829;
assign addr[22891]= -470399716;
assign addr[22892]= -618347408;
assign addr[22893]= -763158411;
assign addr[22894]= -904098143;
assign addr[22895]= -1040451659;
assign addr[22896]= -1171527280;
assign addr[22897]= -1296660098;
assign addr[22898]= -1415215352;
assign addr[22899]= -1526591649;
assign addr[22900]= -1630224009;
assign addr[22901]= -1725586737;
assign addr[22902]= -1812196087;
assign addr[22903]= -1889612716;
assign addr[22904]= -1957443913;
assign addr[22905]= -2015345591;
assign addr[22906]= -2063024031;
assign addr[22907]= -2100237377;
assign addr[22908]= -2126796855;
assign addr[22909]= -2142567738;
assign addr[22910]= -2147470025;
assign addr[22911]= -2141478848;
assign addr[22912]= -2124624598;
assign addr[22913]= -2096992772;
assign addr[22914]= -2058723538;
assign addr[22915]= -2010011024;
assign addr[22916]= -1951102334;
assign addr[22917]= -1882296293;
assign addr[22918]= -1803941934;
assign addr[22919]= -1716436725;
assign addr[22920]= -1620224553;
assign addr[22921]= -1515793473;
assign addr[22922]= -1403673233;
assign addr[22923]= -1284432584;
assign addr[22924]= -1158676398;
assign addr[22925]= -1027042599;
assign addr[22926]= -890198924;
assign addr[22927]= -748839539;
assign addr[22928]= -603681519;
assign addr[22929]= -455461206;
assign addr[22930]= -304930476;
assign addr[22931]= -152852926;
assign addr[22932]= 0;
assign addr[22933]= 152852926;
assign addr[22934]= 304930476;
assign addr[22935]= 455461206;
assign addr[22936]= 603681519;
assign addr[22937]= 748839539;
assign addr[22938]= 890198924;
assign addr[22939]= 1027042599;
assign addr[22940]= 1158676398;
assign addr[22941]= 1284432584;
assign addr[22942]= 1403673233;
assign addr[22943]= 1515793473;
assign addr[22944]= 1620224553;
assign addr[22945]= 1716436725;
assign addr[22946]= 1803941934;
assign addr[22947]= 1882296293;
assign addr[22948]= 1951102334;
assign addr[22949]= 2010011024;
assign addr[22950]= 2058723538;
assign addr[22951]= 2096992772;
assign addr[22952]= 2124624598;
assign addr[22953]= 2141478848;
assign addr[22954]= 2147470025;
assign addr[22955]= 2142567738;
assign addr[22956]= 2126796855;
assign addr[22957]= 2100237377;
assign addr[22958]= 2063024031;
assign addr[22959]= 2015345591;
assign addr[22960]= 1957443913;
assign addr[22961]= 1889612716;
assign addr[22962]= 1812196087;
assign addr[22963]= 1725586737;
assign addr[22964]= 1630224009;
assign addr[22965]= 1526591649;
assign addr[22966]= 1415215352;
assign addr[22967]= 1296660098;
assign addr[22968]= 1171527280;
assign addr[22969]= 1040451659;
assign addr[22970]= 904098143;
assign addr[22971]= 763158411;
assign addr[22972]= 618347408;
assign addr[22973]= 470399716;
assign addr[22974]= 320065829;
assign addr[22975]= 168108346;
assign addr[22976]= 15298099;
assign addr[22977]= -137589750;
assign addr[22978]= -289779648;
assign addr[22979]= -440499581;
assign addr[22980]= -588984994;
assign addr[22981]= -734482665;
assign addr[22982]= -876254528;
assign addr[22983]= -1013581418;
assign addr[22984]= -1145766716;
assign addr[22985]= -1272139887;
assign addr[22986]= -1392059879;
assign addr[22987]= -1504918373;
assign addr[22988]= -1610142873;
assign addr[22989]= -1707199606;
assign addr[22990]= -1795596234;
assign addr[22991]= -1874884346;
assign addr[22992]= -1944661739;
assign addr[22993]= -2004574453;
assign addr[22994]= -2054318569;
assign addr[22995]= -2093641749;
assign addr[22996]= -2122344521;
assign addr[22997]= -2140281282;
assign addr[22998]= -2147361045;
assign addr[22999]= -2143547897;
assign addr[23000]= -2128861181;
assign addr[23001]= -2103375398;
assign addr[23002]= -2067219829;
assign addr[23003]= -2020577882;
assign addr[23004]= -1963686155;
assign addr[23005]= -1896833245;
assign addr[23006]= -1820358275;
assign addr[23007]= -1734649179;
assign addr[23008]= -1640140734;
assign addr[23009]= -1537312353;
assign addr[23010]= -1426685652;
assign addr[23011]= -1308821808;
assign addr[23012]= -1184318708;
assign addr[23013]= -1053807919;
assign addr[23014]= -917951481;
assign addr[23015]= -777438554;
assign addr[23016]= -632981917;
assign addr[23017]= -485314355;
assign addr[23018]= -335184940;
assign addr[23019]= -183355234;
assign addr[23020]= -30595422;
assign addr[23021]= 122319591;
assign addr[23022]= 274614114;
assign addr[23023]= 425515602;
assign addr[23024]= 574258580;
assign addr[23025]= 720088517;
assign addr[23026]= 862265664;
assign addr[23027]= 1000068799;
assign addr[23028]= 1132798888;
assign addr[23029]= 1259782632;
assign addr[23030]= 1380375881;
assign addr[23031]= 1493966902;
assign addr[23032]= 1599979481;
assign addr[23033]= 1697875851;
assign addr[23034]= 1787159411;
assign addr[23035]= 1867377253;
assign addr[23036]= 1938122457;
assign addr[23037]= 1999036154;
assign addr[23038]= 2049809346;
assign addr[23039]= 2090184478;
assign addr[23040]= 2119956737;
assign addr[23041]= 2138975100;
assign addr[23042]= 2147143090;
assign addr[23043]= 2144419275;
assign addr[23044]= 2130817471;
assign addr[23045]= 2106406677;
assign addr[23046]= 2071310720;
assign addr[23047]= 2025707632;
assign addr[23048]= 1969828744;
assign addr[23049]= 1903957513;
assign addr[23050]= 1828428082;
assign addr[23051]= 1743623590;
assign addr[23052]= 1649974225;
assign addr[23053]= 1547955041;
assign addr[23054]= 1438083551;
assign addr[23055]= 1320917099;
assign addr[23056]= 1197050035;
assign addr[23057]= 1067110699;
assign addr[23058]= 931758235;
assign addr[23059]= 791679244;
assign addr[23060]= 647584304;
assign addr[23061]= 500204365;
assign addr[23062]= 350287041;
assign addr[23063]= 198592817;
assign addr[23064]= 45891193;
assign addr[23065]= -107043224;
assign addr[23066]= -259434643;
assign addr[23067]= -410510029;
assign addr[23068]= -559503022;
assign addr[23069]= -705657826;
assign addr[23070]= -848233042;
assign addr[23071]= -986505429;
assign addr[23072]= -1119773573;
assign addr[23073]= -1247361445;
assign addr[23074]= -1368621831;
assign addr[23075]= -1482939614;
assign addr[23076]= -1589734894;
assign addr[23077]= -1688465931;
assign addr[23078]= -1778631892;
assign addr[23079]= -1859775393;
assign addr[23080]= -1931484818;
assign addr[23081]= -1993396407;
assign addr[23082]= -2045196100;
assign addr[23083]= -2086621133;
assign addr[23084]= -2117461370;
assign addr[23085]= -2137560369;
assign addr[23086]= -2146816171;
assign addr[23087]= -2145181827;
assign addr[23088]= -2132665626;
assign addr[23089]= -2109331059;
assign addr[23090]= -2075296495;
assign addr[23091]= -2030734582;
assign addr[23092]= -1975871368;
assign addr[23093]= -1910985158;
assign addr[23094]= -1836405100;
assign addr[23095]= -1752509516;
assign addr[23096]= -1659723983;
assign addr[23097]= -1558519173;
assign addr[23098]= -1449408469;
assign addr[23099]= -1332945355;
assign addr[23100]= -1209720613;
assign addr[23101]= -1080359326;
assign addr[23102]= -945517704;
assign addr[23103]= -805879757;
assign addr[23104]= -662153826;
assign addr[23105]= -515068990;
assign addr[23106]= -365371365;
assign addr[23107]= -213820322;
assign addr[23108]= -61184634;
assign addr[23109]= 91761426;
assign addr[23110]= 244242007;
assign addr[23111]= 395483624;
assign addr[23112]= 544719071;
assign addr[23113]= 691191324;
assign addr[23114]= 834157373;
assign addr[23115]= 972891995;
assign addr[23116]= 1106691431;
assign addr[23117]= 1234876957;
assign addr[23118]= 1356798326;
assign addr[23119]= 1471837070;
assign addr[23120]= 1579409630;
assign addr[23121]= 1678970324;
assign addr[23122]= 1770014111;
assign addr[23123]= 1852079154;
assign addr[23124]= 1924749160;
assign addr[23125]= 1987655498;
assign addr[23126]= 2040479063;
assign addr[23127]= 2082951896;
assign addr[23128]= 2114858546;
assign addr[23129]= 2136037160;
assign addr[23130]= 2146380306;
assign addr[23131]= 2145835515;
assign addr[23132]= 2134405552;
assign addr[23133]= 2112148396;
assign addr[23134]= 2079176953;
assign addr[23135]= 2035658475;
assign addr[23136]= 1981813720;
assign addr[23137]= 1917915825;
assign addr[23138]= 1844288924;
assign addr[23139]= 1761306505;
assign addr[23140]= 1669389513;
assign addr[23141]= 1569004214;
assign addr[23142]= 1460659832;
assign addr[23143]= 1344905966;
assign addr[23144]= 1222329801;
assign addr[23145]= 1093553126;
assign addr[23146]= 959229189;
assign addr[23147]= 820039373;
assign addr[23148]= 676689746;
assign addr[23149]= 529907477;
assign addr[23150]= 380437148;
assign addr[23151]= 229036977;
assign addr[23152]= 76474970;
assign addr[23153]= -76474970;
assign addr[23154]= -229036977;
assign addr[23155]= -380437148;
assign addr[23156]= -529907477;
assign addr[23157]= -676689746;
assign addr[23158]= -820039373;
assign addr[23159]= -959229189;
assign addr[23160]= -1093553126;
assign addr[23161]= -1222329801;
assign addr[23162]= -1344905966;
assign addr[23163]= -1460659832;
assign addr[23164]= -1569004214;
assign addr[23165]= -1669389513;
assign addr[23166]= -1761306505;
assign addr[23167]= -1844288924;
assign addr[23168]= -1917915825;
assign addr[23169]= -1981813720;
assign addr[23170]= -2035658475;
assign addr[23171]= -2079176953;
assign addr[23172]= -2112148396;
assign addr[23173]= -2134405552;
assign addr[23174]= -2145835515;
assign addr[23175]= -2146380306;
assign addr[23176]= -2136037160;
assign addr[23177]= -2114858546;
assign addr[23178]= -2082951896;
assign addr[23179]= -2040479063;
assign addr[23180]= -1987655498;
assign addr[23181]= -1924749160;
assign addr[23182]= -1852079154;
assign addr[23183]= -1770014111;
assign addr[23184]= -1678970324;
assign addr[23185]= -1579409630;
assign addr[23186]= -1471837070;
assign addr[23187]= -1356798326;
assign addr[23188]= -1234876957;
assign addr[23189]= -1106691431;
assign addr[23190]= -972891995;
assign addr[23191]= -834157373;
assign addr[23192]= -691191324;
assign addr[23193]= -544719071;
assign addr[23194]= -395483624;
assign addr[23195]= -244242007;
assign addr[23196]= -91761426;
assign addr[23197]= 61184634;
assign addr[23198]= 213820322;
assign addr[23199]= 365371365;
assign addr[23200]= 515068990;
assign addr[23201]= 662153826;
assign addr[23202]= 805879757;
assign addr[23203]= 945517704;
assign addr[23204]= 1080359326;
assign addr[23205]= 1209720613;
assign addr[23206]= 1332945355;
assign addr[23207]= 1449408469;
assign addr[23208]= 1558519173;
assign addr[23209]= 1659723983;
assign addr[23210]= 1752509516;
assign addr[23211]= 1836405100;
assign addr[23212]= 1910985158;
assign addr[23213]= 1975871368;
assign addr[23214]= 2030734582;
assign addr[23215]= 2075296495;
assign addr[23216]= 2109331059;
assign addr[23217]= 2132665626;
assign addr[23218]= 2145181827;
assign addr[23219]= 2146816171;
assign addr[23220]= 2137560369;
assign addr[23221]= 2117461370;
assign addr[23222]= 2086621133;
assign addr[23223]= 2045196100;
assign addr[23224]= 1993396407;
assign addr[23225]= 1931484818;
assign addr[23226]= 1859775393;
assign addr[23227]= 1778631892;
assign addr[23228]= 1688465931;
assign addr[23229]= 1589734894;
assign addr[23230]= 1482939614;
assign addr[23231]= 1368621831;
assign addr[23232]= 1247361445;
assign addr[23233]= 1119773573;
assign addr[23234]= 986505429;
assign addr[23235]= 848233042;
assign addr[23236]= 705657826;
assign addr[23237]= 559503022;
assign addr[23238]= 410510029;
assign addr[23239]= 259434643;
assign addr[23240]= 107043224;
assign addr[23241]= -45891193;
assign addr[23242]= -198592817;
assign addr[23243]= -350287041;
assign addr[23244]= -500204365;
assign addr[23245]= -647584304;
assign addr[23246]= -791679244;
assign addr[23247]= -931758235;
assign addr[23248]= -1067110699;
assign addr[23249]= -1197050035;
assign addr[23250]= -1320917099;
assign addr[23251]= -1438083551;
assign addr[23252]= -1547955041;
assign addr[23253]= -1649974225;
assign addr[23254]= -1743623590;
assign addr[23255]= -1828428082;
assign addr[23256]= -1903957513;
assign addr[23257]= -1969828744;
assign addr[23258]= -2025707632;
assign addr[23259]= -2071310720;
assign addr[23260]= -2106406677;
assign addr[23261]= -2130817471;
assign addr[23262]= -2144419275;
assign addr[23263]= -2147143090;
assign addr[23264]= -2138975100;
assign addr[23265]= -2119956737;
assign addr[23266]= -2090184478;
assign addr[23267]= -2049809346;
assign addr[23268]= -1999036154;
assign addr[23269]= -1938122457;
assign addr[23270]= -1867377253;
assign addr[23271]= -1787159411;
assign addr[23272]= -1697875851;
assign addr[23273]= -1599979481;
assign addr[23274]= -1493966902;
assign addr[23275]= -1380375881;
assign addr[23276]= -1259782632;
assign addr[23277]= -1132798888;
assign addr[23278]= -1000068799;
assign addr[23279]= -862265664;
assign addr[23280]= -720088517;
assign addr[23281]= -574258580;
assign addr[23282]= -425515602;
assign addr[23283]= -274614114;
assign addr[23284]= -122319591;
assign addr[23285]= 30595422;
assign addr[23286]= 183355234;
assign addr[23287]= 335184940;
assign addr[23288]= 485314355;
assign addr[23289]= 632981917;
assign addr[23290]= 777438554;
assign addr[23291]= 917951481;
assign addr[23292]= 1053807919;
assign addr[23293]= 1184318708;
assign addr[23294]= 1308821808;
assign addr[23295]= 1426685652;
assign addr[23296]= 1537312353;
assign addr[23297]= 1640140734;
assign addr[23298]= 1734649179;
assign addr[23299]= 1820358275;
assign addr[23300]= 1896833245;
assign addr[23301]= 1963686155;
assign addr[23302]= 2020577882;
assign addr[23303]= 2067219829;
assign addr[23304]= 2103375398;
assign addr[23305]= 2128861181;
assign addr[23306]= 2143547897;
assign addr[23307]= 2147361045;
assign addr[23308]= 2140281282;
assign addr[23309]= 2122344521;
assign addr[23310]= 2093641749;
assign addr[23311]= 2054318569;
assign addr[23312]= 2004574453;
assign addr[23313]= 1944661739;
assign addr[23314]= 1874884346;
assign addr[23315]= 1795596234;
assign addr[23316]= 1707199606;
assign addr[23317]= 1610142873;
assign addr[23318]= 1504918373;
assign addr[23319]= 1392059879;
assign addr[23320]= 1272139887;
assign addr[23321]= 1145766716;
assign addr[23322]= 1013581418;
assign addr[23323]= 876254528;
assign addr[23324]= 734482665;
assign addr[23325]= 588984994;
assign addr[23326]= 440499581;
assign addr[23327]= 289779648;
assign addr[23328]= 137589750;
assign addr[23329]= -15298099;
assign addr[23330]= -168108346;
assign addr[23331]= -320065829;
assign addr[23332]= -470399716;
assign addr[23333]= -618347408;
assign addr[23334]= -763158411;
assign addr[23335]= -904098143;
assign addr[23336]= -1040451659;
assign addr[23337]= -1171527280;
assign addr[23338]= -1296660098;
assign addr[23339]= -1415215352;
assign addr[23340]= -1526591649;
assign addr[23341]= -1630224009;
assign addr[23342]= -1725586737;
assign addr[23343]= -1812196087;
assign addr[23344]= -1889612716;
assign addr[23345]= -1957443913;
assign addr[23346]= -2015345591;
assign addr[23347]= -2063024031;
assign addr[23348]= -2100237377;
assign addr[23349]= -2126796855;
assign addr[23350]= -2142567738;
assign addr[23351]= -2147470025;
assign addr[23352]= -2141478848;
assign addr[23353]= -2124624598;
assign addr[23354]= -2096992772;
assign addr[23355]= -2058723538;
assign addr[23356]= -2010011024;
assign addr[23357]= -1951102334;
assign addr[23358]= -1882296293;
assign addr[23359]= -1803941934;
assign addr[23360]= -1716436725;
assign addr[23361]= -1620224553;
assign addr[23362]= -1515793473;
assign addr[23363]= -1403673233;
assign addr[23364]= -1284432584;
assign addr[23365]= -1158676398;
assign addr[23366]= -1027042599;
assign addr[23367]= -890198924;
assign addr[23368]= -748839539;
assign addr[23369]= -603681519;
assign addr[23370]= -455461206;
assign addr[23371]= -304930476;
assign addr[23372]= -152852926;
assign addr[23373]= 0;
assign addr[23374]= 152852926;
assign addr[23375]= 304930476;
assign addr[23376]= 455461206;
assign addr[23377]= 603681519;
assign addr[23378]= 748839539;
assign addr[23379]= 890198924;
assign addr[23380]= 1027042599;
assign addr[23381]= 1158676398;
assign addr[23382]= 1284432584;
assign addr[23383]= 1403673233;
assign addr[23384]= 1515793473;
assign addr[23385]= 1620224553;
assign addr[23386]= 1716436725;
assign addr[23387]= 1803941934;
assign addr[23388]= 1882296293;
assign addr[23389]= 1951102334;
assign addr[23390]= 2010011024;
assign addr[23391]= 2058723538;
assign addr[23392]= 2096992772;
assign addr[23393]= 2124624598;
assign addr[23394]= 2141478848;
assign addr[23395]= 2147470025;
assign addr[23396]= 2142567738;
assign addr[23397]= 2126796855;
assign addr[23398]= 2100237377;
assign addr[23399]= 2063024031;
assign addr[23400]= 2015345591;
assign addr[23401]= 1957443913;
assign addr[23402]= 1889612716;
assign addr[23403]= 1812196087;
assign addr[23404]= 1725586737;
assign addr[23405]= 1630224009;
assign addr[23406]= 1526591649;
assign addr[23407]= 1415215352;
assign addr[23408]= 1296660098;
assign addr[23409]= 1171527280;
assign addr[23410]= 1040451659;
assign addr[23411]= 904098143;
assign addr[23412]= 763158411;
assign addr[23413]= 618347408;
assign addr[23414]= 470399716;
assign addr[23415]= 320065829;
assign addr[23416]= 168108346;
assign addr[23417]= 15298099;
assign addr[23418]= -137589750;
assign addr[23419]= -289779648;
assign addr[23420]= -440499581;
assign addr[23421]= -588984994;
assign addr[23422]= -734482665;
assign addr[23423]= -876254528;
assign addr[23424]= -1013581418;
assign addr[23425]= -1145766716;
assign addr[23426]= -1272139887;
assign addr[23427]= -1392059879;
assign addr[23428]= -1504918373;
assign addr[23429]= -1610142873;
assign addr[23430]= -1707199606;
assign addr[23431]= -1795596234;
assign addr[23432]= -1874884346;
assign addr[23433]= -1944661739;
assign addr[23434]= -2004574453;
assign addr[23435]= -2054318569;
assign addr[23436]= -2093641749;
assign addr[23437]= -2122344521;
assign addr[23438]= -2140281282;
assign addr[23439]= -2147361045;
assign addr[23440]= -2143547897;
assign addr[23441]= -2128861181;
assign addr[23442]= -2103375398;
assign addr[23443]= -2067219829;
assign addr[23444]= -2020577882;
assign addr[23445]= -1963686155;
assign addr[23446]= -1896833245;
assign addr[23447]= -1820358275;
assign addr[23448]= -1734649179;
assign addr[23449]= -1640140734;
assign addr[23450]= -1537312353;
assign addr[23451]= -1426685652;
assign addr[23452]= -1308821808;
assign addr[23453]= -1184318708;
assign addr[23454]= -1053807919;
assign addr[23455]= -917951481;
assign addr[23456]= -777438554;
assign addr[23457]= -632981917;
assign addr[23458]= -485314355;
assign addr[23459]= -335184940;
assign addr[23460]= -183355234;
assign addr[23461]= -30595422;
assign addr[23462]= 122319591;
assign addr[23463]= 274614114;
assign addr[23464]= 425515602;
assign addr[23465]= 574258580;
assign addr[23466]= 720088517;
assign addr[23467]= 862265664;
assign addr[23468]= 1000068799;
assign addr[23469]= 1132798888;
assign addr[23470]= 1259782632;
assign addr[23471]= 1380375881;
assign addr[23472]= 1493966902;
assign addr[23473]= 1599979481;
assign addr[23474]= 1697875851;
assign addr[23475]= 1787159411;
assign addr[23476]= 1867377253;
assign addr[23477]= 1938122457;
assign addr[23478]= 1999036154;
assign addr[23479]= 2049809346;
assign addr[23480]= 2090184478;
assign addr[23481]= 2119956737;
assign addr[23482]= 2138975100;
assign addr[23483]= 2147143090;
assign addr[23484]= 2144419275;
assign addr[23485]= 2130817471;
assign addr[23486]= 2106406677;
assign addr[23487]= 2071310720;
assign addr[23488]= 2025707632;
assign addr[23489]= 1969828744;
assign addr[23490]= 1903957513;
assign addr[23491]= 1828428082;
assign addr[23492]= 1743623590;
assign addr[23493]= 1649974225;
assign addr[23494]= 1547955041;
assign addr[23495]= 1438083551;
assign addr[23496]= 1320917099;
assign addr[23497]= 1197050035;
assign addr[23498]= 1067110699;
assign addr[23499]= 931758235;
assign addr[23500]= 791679244;
assign addr[23501]= 647584304;
assign addr[23502]= 500204365;
assign addr[23503]= 350287041;
assign addr[23504]= 198592817;
assign addr[23505]= 45891193;
assign addr[23506]= -107043224;
assign addr[23507]= -259434643;
assign addr[23508]= -410510029;
assign addr[23509]= -559503022;
assign addr[23510]= -705657826;
assign addr[23511]= -848233042;
assign addr[23512]= -986505429;
assign addr[23513]= -1119773573;
assign addr[23514]= -1247361445;
assign addr[23515]= -1368621831;
assign addr[23516]= -1482939614;
assign addr[23517]= -1589734894;
assign addr[23518]= -1688465931;
assign addr[23519]= -1778631892;
assign addr[23520]= -1859775393;
assign addr[23521]= -1931484818;
assign addr[23522]= -1993396407;
assign addr[23523]= -2045196100;
assign addr[23524]= -2086621133;
assign addr[23525]= -2117461370;
assign addr[23526]= -2137560369;
assign addr[23527]= -2146816171;
assign addr[23528]= -2145181827;
assign addr[23529]= -2132665626;
assign addr[23530]= -2109331059;
assign addr[23531]= -2075296495;
assign addr[23532]= -2030734582;
assign addr[23533]= -1975871368;
assign addr[23534]= -1910985158;
assign addr[23535]= -1836405100;
assign addr[23536]= -1752509516;
assign addr[23537]= -1659723983;
assign addr[23538]= -1558519173;
assign addr[23539]= -1449408469;
assign addr[23540]= -1332945355;
assign addr[23541]= -1209720613;
assign addr[23542]= -1080359326;
assign addr[23543]= -945517704;
assign addr[23544]= -805879757;
assign addr[23545]= -662153826;
assign addr[23546]= -515068990;
assign addr[23547]= -365371365;
assign addr[23548]= -213820322;
assign addr[23549]= -61184634;
assign addr[23550]= 91761426;
assign addr[23551]= 244242007;
assign addr[23552]= 395483624;
assign addr[23553]= 544719071;
assign addr[23554]= 691191324;
assign addr[23555]= 834157373;
assign addr[23556]= 972891995;
assign addr[23557]= 1106691431;
assign addr[23558]= 1234876957;
assign addr[23559]= 1356798326;
assign addr[23560]= 1471837070;
assign addr[23561]= 1579409630;
assign addr[23562]= 1678970324;
assign addr[23563]= 1770014111;
assign addr[23564]= 1852079154;
assign addr[23565]= 1924749160;
assign addr[23566]= 1987655498;
assign addr[23567]= 2040479063;
assign addr[23568]= 2082951896;
assign addr[23569]= 2114858546;
assign addr[23570]= 2136037160;
assign addr[23571]= 2146380306;
assign addr[23572]= 2145835515;
assign addr[23573]= 2134405552;
assign addr[23574]= 2112148396;
assign addr[23575]= 2079176953;
assign addr[23576]= 2035658475;
assign addr[23577]= 1981813720;
assign addr[23578]= 1917915825;
assign addr[23579]= 1844288924;
assign addr[23580]= 1761306505;
assign addr[23581]= 1669389513;
assign addr[23582]= 1569004214;
assign addr[23583]= 1460659832;
assign addr[23584]= 1344905966;
assign addr[23585]= 1222329801;
assign addr[23586]= 1093553126;
assign addr[23587]= 959229189;
assign addr[23588]= 820039373;
assign addr[23589]= 676689746;
assign addr[23590]= 529907477;
assign addr[23591]= 380437148;
assign addr[23592]= 229036977;
assign addr[23593]= 76474970;
assign addr[23594]= -76474970;
assign addr[23595]= -229036977;
assign addr[23596]= -380437148;
assign addr[23597]= -529907477;
assign addr[23598]= -676689746;
assign addr[23599]= -820039373;
assign addr[23600]= -959229189;
assign addr[23601]= -1093553126;
assign addr[23602]= -1222329801;
assign addr[23603]= -1344905966;
assign addr[23604]= -1460659832;
assign addr[23605]= -1569004214;
assign addr[23606]= -1669389513;
assign addr[23607]= -1761306505;
assign addr[23608]= -1844288924;
assign addr[23609]= -1917915825;
assign addr[23610]= -1981813720;
assign addr[23611]= -2035658475;
assign addr[23612]= -2079176953;
assign addr[23613]= -2112148396;
assign addr[23614]= -2134405552;
assign addr[23615]= -2145835515;
assign addr[23616]= -2146380306;
assign addr[23617]= -2136037160;
assign addr[23618]= -2114858546;
assign addr[23619]= -2082951896;
assign addr[23620]= -2040479063;
assign addr[23621]= -1987655498;
assign addr[23622]= -1924749160;
assign addr[23623]= -1852079154;
assign addr[23624]= -1770014111;
assign addr[23625]= -1678970324;
assign addr[23626]= -1579409630;
assign addr[23627]= -1471837070;
assign addr[23628]= -1356798326;
assign addr[23629]= -1234876957;
assign addr[23630]= -1106691431;
assign addr[23631]= -972891995;
assign addr[23632]= -834157373;
assign addr[23633]= -691191324;
assign addr[23634]= -544719071;
assign addr[23635]= -395483624;
assign addr[23636]= -244242007;
assign addr[23637]= -91761426;
assign addr[23638]= 61184634;
assign addr[23639]= 213820322;
assign addr[23640]= 365371365;
assign addr[23641]= 515068990;
assign addr[23642]= 662153826;
assign addr[23643]= 805879757;
assign addr[23644]= 945517704;
assign addr[23645]= 1080359326;
assign addr[23646]= 1209720613;
assign addr[23647]= 1332945355;
assign addr[23648]= 1449408469;
assign addr[23649]= 1558519173;
assign addr[23650]= 1659723983;
assign addr[23651]= 1752509516;
assign addr[23652]= 1836405100;
assign addr[23653]= 1910985158;
assign addr[23654]= 1975871368;
assign addr[23655]= 2030734582;
assign addr[23656]= 2075296495;
assign addr[23657]= 2109331059;
assign addr[23658]= 2132665626;
assign addr[23659]= 2145181827;
assign addr[23660]= 2146816171;
assign addr[23661]= 2137560369;
assign addr[23662]= 2117461370;
assign addr[23663]= 2086621133;
assign addr[23664]= 2045196100;
assign addr[23665]= 1993396407;
assign addr[23666]= 1931484818;
assign addr[23667]= 1859775393;
assign addr[23668]= 1778631892;
assign addr[23669]= 1688465931;
assign addr[23670]= 1589734894;
assign addr[23671]= 1482939614;
assign addr[23672]= 1368621831;
assign addr[23673]= 1247361445;
assign addr[23674]= 1119773573;
assign addr[23675]= 986505429;
assign addr[23676]= 848233042;
assign addr[23677]= 705657826;
assign addr[23678]= 559503022;
assign addr[23679]= 410510029;
assign addr[23680]= 259434643;
assign addr[23681]= 107043224;
assign addr[23682]= -45891193;
assign addr[23683]= -198592817;
assign addr[23684]= -350287041;
assign addr[23685]= -500204365;
assign addr[23686]= -647584304;
assign addr[23687]= -791679244;
assign addr[23688]= -931758235;
assign addr[23689]= -1067110699;
assign addr[23690]= -1197050035;
assign addr[23691]= -1320917099;
assign addr[23692]= -1438083551;
assign addr[23693]= -1547955041;
assign addr[23694]= -1649974225;
assign addr[23695]= -1743623590;
assign addr[23696]= -1828428082;
assign addr[23697]= -1903957513;
assign addr[23698]= -1969828744;
assign addr[23699]= -2025707632;
assign addr[23700]= -2071310720;
assign addr[23701]= -2106406677;
assign addr[23702]= -2130817471;
assign addr[23703]= -2144419275;
assign addr[23704]= -2147143090;
assign addr[23705]= -2138975100;
assign addr[23706]= -2119956737;
assign addr[23707]= -2090184478;
assign addr[23708]= -2049809346;
assign addr[23709]= -1999036154;
assign addr[23710]= -1938122457;
assign addr[23711]= -1867377253;
assign addr[23712]= -1787159411;
assign addr[23713]= -1697875851;
assign addr[23714]= -1599979481;
assign addr[23715]= -1493966902;
assign addr[23716]= -1380375881;
assign addr[23717]= -1259782632;
assign addr[23718]= -1132798888;
assign addr[23719]= -1000068799;
assign addr[23720]= -862265664;
assign addr[23721]= -720088517;
assign addr[23722]= -574258580;
assign addr[23723]= -425515602;
assign addr[23724]= -274614114;
assign addr[23725]= -122319591;
assign addr[23726]= 30595422;
assign addr[23727]= 183355234;
assign addr[23728]= 335184940;
assign addr[23729]= 485314355;
assign addr[23730]= 632981917;
assign addr[23731]= 777438554;
assign addr[23732]= 917951481;
assign addr[23733]= 1053807919;
assign addr[23734]= 1184318708;
assign addr[23735]= 1308821808;
assign addr[23736]= 1426685652;
assign addr[23737]= 1537312353;
assign addr[23738]= 1640140734;
assign addr[23739]= 1734649179;
assign addr[23740]= 1820358275;
assign addr[23741]= 1896833245;
assign addr[23742]= 1963686155;
assign addr[23743]= 2020577882;
assign addr[23744]= 2067219829;
assign addr[23745]= 2103375398;
assign addr[23746]= 2128861181;
assign addr[23747]= 2143547897;
assign addr[23748]= 2147361045;
assign addr[23749]= 2140281282;
assign addr[23750]= 2122344521;
assign addr[23751]= 2093641749;
assign addr[23752]= 2054318569;
assign addr[23753]= 2004574453;
assign addr[23754]= 1944661739;
assign addr[23755]= 1874884346;
assign addr[23756]= 1795596234;
assign addr[23757]= 1707199606;
assign addr[23758]= 1610142873;
assign addr[23759]= 1504918373;
assign addr[23760]= 1392059879;
assign addr[23761]= 1272139887;
assign addr[23762]= 1145766716;
assign addr[23763]= 1013581418;
assign addr[23764]= 876254528;
assign addr[23765]= 734482665;
assign addr[23766]= 588984994;
assign addr[23767]= 440499581;
assign addr[23768]= 289779648;
assign addr[23769]= 137589750;
assign addr[23770]= -15298099;
assign addr[23771]= -168108346;
assign addr[23772]= -320065829;
assign addr[23773]= -470399716;
assign addr[23774]= -618347408;
assign addr[23775]= -763158411;
assign addr[23776]= -904098143;
assign addr[23777]= -1040451659;
assign addr[23778]= -1171527280;
assign addr[23779]= -1296660098;
assign addr[23780]= -1415215352;
assign addr[23781]= -1526591649;
assign addr[23782]= -1630224009;
assign addr[23783]= -1725586737;
assign addr[23784]= -1812196087;
assign addr[23785]= -1889612716;
assign addr[23786]= -1957443913;
assign addr[23787]= -2015345591;
assign addr[23788]= -2063024031;
assign addr[23789]= -2100237377;
assign addr[23790]= -2126796855;
assign addr[23791]= -2142567738;
assign addr[23792]= -2147470025;
assign addr[23793]= -2141478848;
assign addr[23794]= -2124624598;
assign addr[23795]= -2096992772;
assign addr[23796]= -2058723538;
assign addr[23797]= -2010011024;
assign addr[23798]= -1951102334;
assign addr[23799]= -1882296293;
assign addr[23800]= -1803941934;
assign addr[23801]= -1716436725;
assign addr[23802]= -1620224553;
assign addr[23803]= -1515793473;
assign addr[23804]= -1403673233;
assign addr[23805]= -1284432584;
assign addr[23806]= -1158676398;
assign addr[23807]= -1027042599;
assign addr[23808]= -890198924;
assign addr[23809]= -748839539;
assign addr[23810]= -603681519;
assign addr[23811]= -455461206;
assign addr[23812]= -304930476;
assign addr[23813]= -152852926;
assign addr[23814]= 0;
assign addr[23815]= 152852926;
assign addr[23816]= 304930476;
assign addr[23817]= 455461206;
assign addr[23818]= 603681519;
assign addr[23819]= 748839539;
assign addr[23820]= 890198924;
assign addr[23821]= 1027042599;
assign addr[23822]= 1158676398;
assign addr[23823]= 1284432584;
assign addr[23824]= 1403673233;
assign addr[23825]= 1515793473;
assign addr[23826]= 1620224553;
assign addr[23827]= 1716436725;
assign addr[23828]= 1803941934;
assign addr[23829]= 1882296293;
assign addr[23830]= 1951102334;
assign addr[23831]= 2010011024;
assign addr[23832]= 2058723538;
assign addr[23833]= 2096992772;
assign addr[23834]= 2124624598;
assign addr[23835]= 2141478848;
assign addr[23836]= 2147470025;
assign addr[23837]= 2142567738;
assign addr[23838]= 2126796855;
assign addr[23839]= 2100237377;
assign addr[23840]= 2063024031;
assign addr[23841]= 2015345591;
assign addr[23842]= 1957443913;
assign addr[23843]= 1889612716;
assign addr[23844]= 1812196087;
assign addr[23845]= 1725586737;
assign addr[23846]= 1630224009;
assign addr[23847]= 1526591649;
assign addr[23848]= 1415215352;
assign addr[23849]= 1296660098;
assign addr[23850]= 1171527280;
assign addr[23851]= 1040451659;
assign addr[23852]= 904098143;
assign addr[23853]= 763158411;
assign addr[23854]= 618347408;
assign addr[23855]= 470399716;
assign addr[23856]= 320065829;
assign addr[23857]= 168108346;
assign addr[23858]= 15298099;
assign addr[23859]= -137589750;
assign addr[23860]= -289779648;
assign addr[23861]= -440499581;
assign addr[23862]= -588984994;
assign addr[23863]= -734482665;
assign addr[23864]= -876254528;
assign addr[23865]= -1013581418;
assign addr[23866]= -1145766716;
assign addr[23867]= -1272139887;
assign addr[23868]= -1392059879;
assign addr[23869]= -1504918373;
assign addr[23870]= -1610142873;
assign addr[23871]= -1707199606;
assign addr[23872]= -1795596234;
assign addr[23873]= -1874884346;
assign addr[23874]= -1944661739;
assign addr[23875]= -2004574453;
assign addr[23876]= -2054318569;
assign addr[23877]= -2093641749;
assign addr[23878]= -2122344521;
assign addr[23879]= -2140281282;
assign addr[23880]= -2147361045;
assign addr[23881]= -2143547897;
assign addr[23882]= -2128861181;
assign addr[23883]= -2103375398;
assign addr[23884]= -2067219829;
assign addr[23885]= -2020577882;
assign addr[23886]= -1963686155;
assign addr[23887]= -1896833245;
assign addr[23888]= -1820358275;
assign addr[23889]= -1734649179;
assign addr[23890]= -1640140734;
assign addr[23891]= -1537312353;
assign addr[23892]= -1426685652;
assign addr[23893]= -1308821808;
assign addr[23894]= -1184318708;
assign addr[23895]= -1053807919;
assign addr[23896]= -917951481;
assign addr[23897]= -777438554;
assign addr[23898]= -632981917;
assign addr[23899]= -485314355;
assign addr[23900]= -335184940;
assign addr[23901]= -183355234;
assign addr[23902]= -30595422;
assign addr[23903]= 122319591;
assign addr[23904]= 274614114;
assign addr[23905]= 425515602;
assign addr[23906]= 574258580;
assign addr[23907]= 720088517;
assign addr[23908]= 862265664;
assign addr[23909]= 1000068799;
assign addr[23910]= 1132798888;
assign addr[23911]= 1259782632;
assign addr[23912]= 1380375881;
assign addr[23913]= 1493966902;
assign addr[23914]= 1599979481;
assign addr[23915]= 1697875851;
assign addr[23916]= 1787159411;
assign addr[23917]= 1867377253;
assign addr[23918]= 1938122457;
assign addr[23919]= 1999036154;
assign addr[23920]= 2049809346;
assign addr[23921]= 2090184478;
assign addr[23922]= 2119956737;
assign addr[23923]= 2138975100;
assign addr[23924]= 2147143090;
assign addr[23925]= 2144419275;
assign addr[23926]= 2130817471;
assign addr[23927]= 2106406677;
assign addr[23928]= 2071310720;
assign addr[23929]= 2025707632;
assign addr[23930]= 1969828744;
assign addr[23931]= 1903957513;
assign addr[23932]= 1828428082;
assign addr[23933]= 1743623590;
assign addr[23934]= 1649974225;
assign addr[23935]= 1547955041;
assign addr[23936]= 1438083551;
assign addr[23937]= 1320917099;
assign addr[23938]= 1197050035;
assign addr[23939]= 1067110699;
assign addr[23940]= 931758235;
assign addr[23941]= 791679244;
assign addr[23942]= 647584304;
assign addr[23943]= 500204365;
assign addr[23944]= 350287041;
assign addr[23945]= 198592817;
assign addr[23946]= 45891193;
assign addr[23947]= -107043224;
assign addr[23948]= -259434643;
assign addr[23949]= -410510029;
assign addr[23950]= -559503022;
assign addr[23951]= -705657826;
assign addr[23952]= -848233042;
assign addr[23953]= -986505429;
assign addr[23954]= -1119773573;
assign addr[23955]= -1247361445;
assign addr[23956]= -1368621831;
assign addr[23957]= -1482939614;
assign addr[23958]= -1589734894;
assign addr[23959]= -1688465931;
assign addr[23960]= -1778631892;
assign addr[23961]= -1859775393;
assign addr[23962]= -1931484818;
assign addr[23963]= -1993396407;
assign addr[23964]= -2045196100;
assign addr[23965]= -2086621133;
assign addr[23966]= -2117461370;
assign addr[23967]= -2137560369;
assign addr[23968]= -2146816171;
assign addr[23969]= -2145181827;
assign addr[23970]= -2132665626;
assign addr[23971]= -2109331059;
assign addr[23972]= -2075296495;
assign addr[23973]= -2030734582;
assign addr[23974]= -1975871368;
assign addr[23975]= -1910985158;
assign addr[23976]= -1836405100;
assign addr[23977]= -1752509516;
assign addr[23978]= -1659723983;
assign addr[23979]= -1558519173;
assign addr[23980]= -1449408469;
assign addr[23981]= -1332945355;
assign addr[23982]= -1209720613;
assign addr[23983]= -1080359326;
assign addr[23984]= -945517704;
assign addr[23985]= -805879757;
assign addr[23986]= -662153826;
assign addr[23987]= -515068990;
assign addr[23988]= -365371365;
assign addr[23989]= -213820322;
assign addr[23990]= -61184634;
assign addr[23991]= 91761426;
assign addr[23992]= 244242007;
assign addr[23993]= 395483624;
assign addr[23994]= 544719071;
assign addr[23995]= 691191324;
assign addr[23996]= 834157373;
assign addr[23997]= 972891995;
assign addr[23998]= 1106691431;
assign addr[23999]= 1234876957;
assign addr[24000]= 1356798326;
assign addr[24001]= 1471837070;
assign addr[24002]= 1579409630;
assign addr[24003]= 1678970324;
assign addr[24004]= 1770014111;
assign addr[24005]= 1852079154;
assign addr[24006]= 1924749160;
assign addr[24007]= 1987655498;
assign addr[24008]= 2040479063;
assign addr[24009]= 2082951896;
assign addr[24010]= 2114858546;
assign addr[24011]= 2136037160;
assign addr[24012]= 2146380306;
assign addr[24013]= 2145835515;
assign addr[24014]= 2134405552;
assign addr[24015]= 2112148396;
assign addr[24016]= 2079176953;
assign addr[24017]= 2035658475;
assign addr[24018]= 1981813720;
assign addr[24019]= 1917915825;
assign addr[24020]= 1844288924;
assign addr[24021]= 1761306505;
assign addr[24022]= 1669389513;
assign addr[24023]= 1569004214;
assign addr[24024]= 1460659832;
assign addr[24025]= 1344905966;
assign addr[24026]= 1222329801;
assign addr[24027]= 1093553126;
assign addr[24028]= 959229189;
assign addr[24029]= 820039373;
assign addr[24030]= 676689746;
assign addr[24031]= 529907477;
assign addr[24032]= 380437148;
assign addr[24033]= 229036977;
assign addr[24034]= 76474970;
assign addr[24035]= -76474970;
assign addr[24036]= -229036977;
assign addr[24037]= -380437148;
assign addr[24038]= -529907477;
assign addr[24039]= -676689746;
assign addr[24040]= -820039373;
assign addr[24041]= -959229189;
assign addr[24042]= -1093553126;
assign addr[24043]= -1222329801;
assign addr[24044]= -1344905966;
assign addr[24045]= -1460659832;
assign addr[24046]= -1569004214;
assign addr[24047]= -1669389513;
assign addr[24048]= -1761306505;
assign addr[24049]= -1844288924;
assign addr[24050]= -1917915825;
assign addr[24051]= -1981813720;
assign addr[24052]= -2035658475;
assign addr[24053]= -2079176953;
assign addr[24054]= -2112148396;
assign addr[24055]= -2134405552;
assign addr[24056]= -2145835515;
assign addr[24057]= -2146380306;
assign addr[24058]= -2136037160;
assign addr[24059]= -2114858546;
assign addr[24060]= -2082951896;
assign addr[24061]= -2040479063;
assign addr[24062]= -1987655498;
assign addr[24063]= -1924749160;
assign addr[24064]= -1852079154;
assign addr[24065]= -1770014111;
assign addr[24066]= -1678970324;
assign addr[24067]= -1579409630;
assign addr[24068]= -1471837070;
assign addr[24069]= -1356798326;
assign addr[24070]= -1234876957;
assign addr[24071]= -1106691431;
assign addr[24072]= -972891995;
assign addr[24073]= -834157373;
assign addr[24074]= -691191324;
assign addr[24075]= -544719071;
assign addr[24076]= -395483624;
assign addr[24077]= -244242007;
assign addr[24078]= -91761426;
assign addr[24079]= 61184634;
assign addr[24080]= 213820322;
assign addr[24081]= 365371365;
assign addr[24082]= 515068990;
assign addr[24083]= 662153826;
assign addr[24084]= 805879757;
assign addr[24085]= 945517704;
assign addr[24086]= 1080359326;
assign addr[24087]= 1209720613;
assign addr[24088]= 1332945355;
assign addr[24089]= 1449408469;
assign addr[24090]= 1558519173;
assign addr[24091]= 1659723983;
assign addr[24092]= 1752509516;
assign addr[24093]= 1836405100;
assign addr[24094]= 1910985158;
assign addr[24095]= 1975871368;
assign addr[24096]= 2030734582;
assign addr[24097]= 2075296495;
assign addr[24098]= 2109331059;
assign addr[24099]= 2132665626;
assign addr[24100]= 2145181827;
assign addr[24101]= 2146816171;
assign addr[24102]= 2137560369;
assign addr[24103]= 2117461370;
assign addr[24104]= 2086621133;
assign addr[24105]= 2045196100;
assign addr[24106]= 1993396407;
assign addr[24107]= 1931484818;
assign addr[24108]= 1859775393;
assign addr[24109]= 1778631892;
assign addr[24110]= 1688465931;
assign addr[24111]= 1589734894;
assign addr[24112]= 1482939614;
assign addr[24113]= 1368621831;
assign addr[24114]= 1247361445;
assign addr[24115]= 1119773573;
assign addr[24116]= 986505429;
assign addr[24117]= 848233042;
assign addr[24118]= 705657826;
assign addr[24119]= 559503022;
assign addr[24120]= 410510029;
assign addr[24121]= 259434643;
assign addr[24122]= 107043224;
assign addr[24123]= -45891193;
assign addr[24124]= -198592817;
assign addr[24125]= -350287041;
assign addr[24126]= -500204365;
assign addr[24127]= -647584304;
assign addr[24128]= -791679244;
assign addr[24129]= -931758235;
assign addr[24130]= -1067110699;
assign addr[24131]= -1197050035;
assign addr[24132]= -1320917099;
assign addr[24133]= -1438083551;
assign addr[24134]= -1547955041;
assign addr[24135]= -1649974225;
assign addr[24136]= -1743623590;
assign addr[24137]= -1828428082;
assign addr[24138]= -1903957513;
assign addr[24139]= -1969828744;
assign addr[24140]= -2025707632;
assign addr[24141]= -2071310720;
assign addr[24142]= -2106406677;
assign addr[24143]= -2130817471;
assign addr[24144]= -2144419275;
assign addr[24145]= -2147143090;
assign addr[24146]= -2138975100;
assign addr[24147]= -2119956737;
assign addr[24148]= -2090184478;
assign addr[24149]= -2049809346;
assign addr[24150]= -1999036154;
assign addr[24151]= -1938122457;
assign addr[24152]= -1867377253;
assign addr[24153]= -1787159411;
assign addr[24154]= -1697875851;
assign addr[24155]= -1599979481;
assign addr[24156]= -1493966902;
assign addr[24157]= -1380375881;
assign addr[24158]= -1259782632;
assign addr[24159]= -1132798888;
assign addr[24160]= -1000068799;
assign addr[24161]= -862265664;
assign addr[24162]= -720088517;
assign addr[24163]= -574258580;
assign addr[24164]= -425515602;
assign addr[24165]= -274614114;
assign addr[24166]= -122319591;
assign addr[24167]= 30595422;
assign addr[24168]= 183355234;
assign addr[24169]= 335184940;
assign addr[24170]= 485314355;
assign addr[24171]= 632981917;
assign addr[24172]= 777438554;
assign addr[24173]= 917951481;
assign addr[24174]= 1053807919;
assign addr[24175]= 1184318708;
assign addr[24176]= 1308821808;
assign addr[24177]= 1426685652;
assign addr[24178]= 1537312353;
assign addr[24179]= 1640140734;
assign addr[24180]= 1734649179;
assign addr[24181]= 1820358275;
assign addr[24182]= 1896833245;
assign addr[24183]= 1963686155;
assign addr[24184]= 2020577882;
assign addr[24185]= 2067219829;
assign addr[24186]= 2103375398;
assign addr[24187]= 2128861181;
assign addr[24188]= 2143547897;
assign addr[24189]= 2147361045;
assign addr[24190]= 2140281282;
assign addr[24191]= 2122344521;
assign addr[24192]= 2093641749;
assign addr[24193]= 2054318569;
assign addr[24194]= 2004574453;
assign addr[24195]= 1944661739;
assign addr[24196]= 1874884346;
assign addr[24197]= 1795596234;
assign addr[24198]= 1707199606;
assign addr[24199]= 1610142873;
assign addr[24200]= 1504918373;
assign addr[24201]= 1392059879;
assign addr[24202]= 1272139887;
assign addr[24203]= 1145766716;
assign addr[24204]= 1013581418;
assign addr[24205]= 876254528;
assign addr[24206]= 734482665;
assign addr[24207]= 588984994;
assign addr[24208]= 440499581;
assign addr[24209]= 289779648;
assign addr[24210]= 137589750;
assign addr[24211]= -15298099;
assign addr[24212]= -168108346;
assign addr[24213]= -320065829;
assign addr[24214]= -470399716;
assign addr[24215]= -618347408;
assign addr[24216]= -763158411;
assign addr[24217]= -904098143;
assign addr[24218]= -1040451659;
assign addr[24219]= -1171527280;
assign addr[24220]= -1296660098;
assign addr[24221]= -1415215352;
assign addr[24222]= -1526591649;
assign addr[24223]= -1630224009;
assign addr[24224]= -1725586737;
assign addr[24225]= -1812196087;
assign addr[24226]= -1889612716;
assign addr[24227]= -1957443913;
assign addr[24228]= -2015345591;
assign addr[24229]= -2063024031;
assign addr[24230]= -2100237377;
assign addr[24231]= -2126796855;
assign addr[24232]= -2142567738;
assign addr[24233]= -2147470025;
assign addr[24234]= -2141478848;
assign addr[24235]= -2124624598;
assign addr[24236]= -2096992772;
assign addr[24237]= -2058723538;
assign addr[24238]= -2010011024;
assign addr[24239]= -1951102334;
assign addr[24240]= -1882296293;
assign addr[24241]= -1803941934;
assign addr[24242]= -1716436725;
assign addr[24243]= -1620224553;
assign addr[24244]= -1515793473;
assign addr[24245]= -1403673233;
assign addr[24246]= -1284432584;
assign addr[24247]= -1158676398;
assign addr[24248]= -1027042599;
assign addr[24249]= -890198924;
assign addr[24250]= -748839539;
assign addr[24251]= -603681519;
assign addr[24252]= -455461206;
assign addr[24253]= -304930476;
assign addr[24254]= -152852926;
assign addr[24255]= 0;
assign addr[24256]= 152852926;
assign addr[24257]= 304930476;
assign addr[24258]= 455461206;
assign addr[24259]= 603681519;
assign addr[24260]= 748839539;
assign addr[24261]= 890198924;
assign addr[24262]= 1027042599;
assign addr[24263]= 1158676398;
assign addr[24264]= 1284432584;
assign addr[24265]= 1403673233;
assign addr[24266]= 1515793473;
assign addr[24267]= 1620224553;
assign addr[24268]= 1716436725;
assign addr[24269]= 1803941934;
assign addr[24270]= 1882296293;
assign addr[24271]= 1951102334;
assign addr[24272]= 2010011024;
assign addr[24273]= 2058723538;
assign addr[24274]= 2096992772;
assign addr[24275]= 2124624598;
assign addr[24276]= 2141478848;
assign addr[24277]= 2147470025;
assign addr[24278]= 2142567738;
assign addr[24279]= 2126796855;
assign addr[24280]= 2100237377;
assign addr[24281]= 2063024031;
assign addr[24282]= 2015345591;
assign addr[24283]= 1957443913;
assign addr[24284]= 1889612716;
assign addr[24285]= 1812196087;
assign addr[24286]= 1725586737;
assign addr[24287]= 1630224009;
assign addr[24288]= 1526591649;
assign addr[24289]= 1415215352;
assign addr[24290]= 1296660098;
assign addr[24291]= 1171527280;
assign addr[24292]= 1040451659;
assign addr[24293]= 904098143;
assign addr[24294]= 763158411;
assign addr[24295]= 618347408;
assign addr[24296]= 470399716;
assign addr[24297]= 320065829;
assign addr[24298]= 168108346;
assign addr[24299]= 15298099;
assign addr[24300]= -137589750;
assign addr[24301]= -289779648;
assign addr[24302]= -440499581;
assign addr[24303]= -588984994;
assign addr[24304]= -734482665;
assign addr[24305]= -876254528;
assign addr[24306]= -1013581418;
assign addr[24307]= -1145766716;
assign addr[24308]= -1272139887;
assign addr[24309]= -1392059879;
assign addr[24310]= -1504918373;
assign addr[24311]= -1610142873;
assign addr[24312]= -1707199606;
assign addr[24313]= -1795596234;
assign addr[24314]= -1874884346;
assign addr[24315]= -1944661739;
assign addr[24316]= -2004574453;
assign addr[24317]= -2054318569;
assign addr[24318]= -2093641749;
assign addr[24319]= -2122344521;
assign addr[24320]= -2140281282;
assign addr[24321]= -2147361045;
assign addr[24322]= -2143547897;
assign addr[24323]= -2128861181;
assign addr[24324]= -2103375398;
assign addr[24325]= -2067219829;
assign addr[24326]= -2020577882;
assign addr[24327]= -1963686155;
assign addr[24328]= -1896833245;
assign addr[24329]= -1820358275;
assign addr[24330]= -1734649179;
assign addr[24331]= -1640140734;
assign addr[24332]= -1537312353;
assign addr[24333]= -1426685652;
assign addr[24334]= -1308821808;
assign addr[24335]= -1184318708;
assign addr[24336]= -1053807919;
assign addr[24337]= -917951481;
assign addr[24338]= -777438554;
assign addr[24339]= -632981917;
assign addr[24340]= -485314355;
assign addr[24341]= -335184940;
assign addr[24342]= -183355234;
assign addr[24343]= -30595422;
assign addr[24344]= 122319591;
assign addr[24345]= 274614114;
assign addr[24346]= 425515602;
assign addr[24347]= 574258580;
assign addr[24348]= 720088517;
assign addr[24349]= 862265664;
assign addr[24350]= 1000068799;
assign addr[24351]= 1132798888;
assign addr[24352]= 1259782632;
assign addr[24353]= 1380375881;
assign addr[24354]= 1493966902;
assign addr[24355]= 1599979481;
assign addr[24356]= 1697875851;
assign addr[24357]= 1787159411;
assign addr[24358]= 1867377253;
assign addr[24359]= 1938122457;
assign addr[24360]= 1999036154;
assign addr[24361]= 2049809346;
assign addr[24362]= 2090184478;
assign addr[24363]= 2119956737;
assign addr[24364]= 2138975100;
assign addr[24365]= 2147143090;
assign addr[24366]= 2144419275;
assign addr[24367]= 2130817471;
assign addr[24368]= 2106406677;
assign addr[24369]= 2071310720;
assign addr[24370]= 2025707632;
assign addr[24371]= 1969828744;
assign addr[24372]= 1903957513;
assign addr[24373]= 1828428082;
assign addr[24374]= 1743623590;
assign addr[24375]= 1649974225;
assign addr[24376]= 1547955041;
assign addr[24377]= 1438083551;
assign addr[24378]= 1320917099;
assign addr[24379]= 1197050035;
assign addr[24380]= 1067110699;
assign addr[24381]= 931758235;
assign addr[24382]= 791679244;
assign addr[24383]= 647584304;
assign addr[24384]= 500204365;
assign addr[24385]= 350287041;
assign addr[24386]= 198592817;
assign addr[24387]= 45891193;
assign addr[24388]= -107043224;
assign addr[24389]= -259434643;
assign addr[24390]= -410510029;
assign addr[24391]= -559503022;
assign addr[24392]= -705657826;
assign addr[24393]= -848233042;
assign addr[24394]= -986505429;
assign addr[24395]= -1119773573;
assign addr[24396]= -1247361445;
assign addr[24397]= -1368621831;
assign addr[24398]= -1482939614;
assign addr[24399]= -1589734894;
assign addr[24400]= -1688465931;
assign addr[24401]= -1778631892;
assign addr[24402]= -1859775393;
assign addr[24403]= -1931484818;
assign addr[24404]= -1993396407;
assign addr[24405]= -2045196100;
assign addr[24406]= -2086621133;
assign addr[24407]= -2117461370;
assign addr[24408]= -2137560369;
assign addr[24409]= -2146816171;
assign addr[24410]= -2145181827;
assign addr[24411]= -2132665626;
assign addr[24412]= -2109331059;
assign addr[24413]= -2075296495;
assign addr[24414]= -2030734582;
assign addr[24415]= -1975871368;
assign addr[24416]= -1910985158;
assign addr[24417]= -1836405100;
assign addr[24418]= -1752509516;
assign addr[24419]= -1659723983;
assign addr[24420]= -1558519173;
assign addr[24421]= -1449408469;
assign addr[24422]= -1332945355;
assign addr[24423]= -1209720613;
assign addr[24424]= -1080359326;
assign addr[24425]= -945517704;
assign addr[24426]= -805879757;
assign addr[24427]= -662153826;
assign addr[24428]= -515068990;
assign addr[24429]= -365371365;
assign addr[24430]= -213820322;
assign addr[24431]= -61184634;
assign addr[24432]= 91761426;
assign addr[24433]= 244242007;
assign addr[24434]= 395483624;
assign addr[24435]= 544719071;
assign addr[24436]= 691191324;
assign addr[24437]= 834157373;
assign addr[24438]= 972891995;
assign addr[24439]= 1106691431;
assign addr[24440]= 1234876957;
assign addr[24441]= 1356798326;
assign addr[24442]= 1471837070;
assign addr[24443]= 1579409630;
assign addr[24444]= 1678970324;
assign addr[24445]= 1770014111;
assign addr[24446]= 1852079154;
assign addr[24447]= 1924749160;
assign addr[24448]= 1987655498;
assign addr[24449]= 2040479063;
assign addr[24450]= 2082951896;
assign addr[24451]= 2114858546;
assign addr[24452]= 2136037160;
assign addr[24453]= 2146380306;
assign addr[24454]= 2145835515;
assign addr[24455]= 2134405552;
assign addr[24456]= 2112148396;
assign addr[24457]= 2079176953;
assign addr[24458]= 2035658475;
assign addr[24459]= 1981813720;
assign addr[24460]= 1917915825;
assign addr[24461]= 1844288924;
assign addr[24462]= 1761306505;
assign addr[24463]= 1669389513;
assign addr[24464]= 1569004214;
assign addr[24465]= 1460659832;
assign addr[24466]= 1344905966;
assign addr[24467]= 1222329801;
assign addr[24468]= 1093553126;
assign addr[24469]= 959229189;
assign addr[24470]= 820039373;
assign addr[24471]= 676689746;
assign addr[24472]= 529907477;
assign addr[24473]= 380437148;
assign addr[24474]= 229036977;
assign addr[24475]= 76474970;
assign addr[24476]= -76474970;
assign addr[24477]= -229036977;
assign addr[24478]= -380437148;
assign addr[24479]= -529907477;
assign addr[24480]= -676689746;
assign addr[24481]= -820039373;
assign addr[24482]= -959229189;
assign addr[24483]= -1093553126;
assign addr[24484]= -1222329801;
assign addr[24485]= -1344905966;
assign addr[24486]= -1460659832;
assign addr[24487]= -1569004214;
assign addr[24488]= -1669389513;
assign addr[24489]= -1761306505;
assign addr[24490]= -1844288924;
assign addr[24491]= -1917915825;
assign addr[24492]= -1981813720;
assign addr[24493]= -2035658475;
assign addr[24494]= -2079176953;
assign addr[24495]= -2112148396;
assign addr[24496]= -2134405552;
assign addr[24497]= -2145835515;
assign addr[24498]= -2146380306;
assign addr[24499]= -2136037160;
assign addr[24500]= -2114858546;
assign addr[24501]= -2082951896;
assign addr[24502]= -2040479063;
assign addr[24503]= -1987655498;
assign addr[24504]= -1924749160;
assign addr[24505]= -1852079154;
assign addr[24506]= -1770014111;
assign addr[24507]= -1678970324;
assign addr[24508]= -1579409630;
assign addr[24509]= -1471837070;
assign addr[24510]= -1356798326;
assign addr[24511]= -1234876957;
assign addr[24512]= -1106691431;
assign addr[24513]= -972891995;
assign addr[24514]= -834157373;
assign addr[24515]= -691191324;
assign addr[24516]= -544719071;
assign addr[24517]= -395483624;
assign addr[24518]= -244242007;
assign addr[24519]= -91761426;
assign addr[24520]= 61184634;
assign addr[24521]= 213820322;
assign addr[24522]= 365371365;
assign addr[24523]= 515068990;
assign addr[24524]= 662153826;
assign addr[24525]= 805879757;
assign addr[24526]= 945517704;
assign addr[24527]= 1080359326;
assign addr[24528]= 1209720613;
assign addr[24529]= 1332945355;
assign addr[24530]= 1449408469;
assign addr[24531]= 1558519173;
assign addr[24532]= 1659723983;
assign addr[24533]= 1752509516;
assign addr[24534]= 1836405100;
assign addr[24535]= 1910985158;
assign addr[24536]= 1975871368;
assign addr[24537]= 2030734582;
assign addr[24538]= 2075296495;
assign addr[24539]= 2109331059;
assign addr[24540]= 2132665626;
assign addr[24541]= 2145181827;
assign addr[24542]= 2146816171;
assign addr[24543]= 2137560369;
assign addr[24544]= 2117461370;
assign addr[24545]= 2086621133;
assign addr[24546]= 2045196100;
assign addr[24547]= 1993396407;
assign addr[24548]= 1931484818;
assign addr[24549]= 1859775393;
assign addr[24550]= 1778631892;
assign addr[24551]= 1688465931;
assign addr[24552]= 1589734894;
assign addr[24553]= 1482939614;
assign addr[24554]= 1368621831;
assign addr[24555]= 1247361445;
assign addr[24556]= 1119773573;
assign addr[24557]= 986505429;
assign addr[24558]= 848233042;
assign addr[24559]= 705657826;
assign addr[24560]= 559503022;
assign addr[24561]= 410510029;
assign addr[24562]= 259434643;
assign addr[24563]= 107043224;
assign addr[24564]= -45891193;
assign addr[24565]= -198592817;
assign addr[24566]= -350287041;
assign addr[24567]= -500204365;
assign addr[24568]= -647584304;
assign addr[24569]= -791679244;
assign addr[24570]= -931758235;
assign addr[24571]= -1067110699;
assign addr[24572]= -1197050035;
assign addr[24573]= -1320917099;
assign addr[24574]= -1438083551;
assign addr[24575]= -1547955041;
assign addr[24576]= -1649974225;
assign addr[24577]= -1743623590;
assign addr[24578]= -1828428082;
assign addr[24579]= -1903957513;
assign addr[24580]= -1969828744;
assign addr[24581]= -2025707632;
assign addr[24582]= -2071310720;
assign addr[24583]= -2106406677;
assign addr[24584]= -2130817471;
assign addr[24585]= -2144419275;
assign addr[24586]= -2147143090;
assign addr[24587]= -2138975100;
assign addr[24588]= -2119956737;
assign addr[24589]= -2090184478;
assign addr[24590]= -2049809346;
assign addr[24591]= -1999036154;
assign addr[24592]= -1938122457;
assign addr[24593]= -1867377253;
assign addr[24594]= -1787159411;
assign addr[24595]= -1697875851;
assign addr[24596]= -1599979481;
assign addr[24597]= -1493966902;
assign addr[24598]= -1380375881;
assign addr[24599]= -1259782632;
assign addr[24600]= -1132798888;
assign addr[24601]= -1000068799;
assign addr[24602]= -862265664;
assign addr[24603]= -720088517;
assign addr[24604]= -574258580;
assign addr[24605]= -425515602;
assign addr[24606]= -274614114;
assign addr[24607]= -122319591;
assign addr[24608]= 30595422;
assign addr[24609]= 183355234;
assign addr[24610]= 335184940;
assign addr[24611]= 485314355;
assign addr[24612]= 632981917;
assign addr[24613]= 777438554;
assign addr[24614]= 917951481;
assign addr[24615]= 1053807919;
assign addr[24616]= 1184318708;
assign addr[24617]= 1308821808;
assign addr[24618]= 1426685652;
assign addr[24619]= 1537312353;
assign addr[24620]= 1640140734;
assign addr[24621]= 1734649179;
assign addr[24622]= 1820358275;
assign addr[24623]= 1896833245;
assign addr[24624]= 1963686155;
assign addr[24625]= 2020577882;
assign addr[24626]= 2067219829;
assign addr[24627]= 2103375398;
assign addr[24628]= 2128861181;
assign addr[24629]= 2143547897;
assign addr[24630]= 2147361045;
assign addr[24631]= 2140281282;
assign addr[24632]= 2122344521;
assign addr[24633]= 2093641749;
assign addr[24634]= 2054318569;
assign addr[24635]= 2004574453;
assign addr[24636]= 1944661739;
assign addr[24637]= 1874884346;
assign addr[24638]= 1795596234;
assign addr[24639]= 1707199606;
assign addr[24640]= 1610142873;
assign addr[24641]= 1504918373;
assign addr[24642]= 1392059879;
assign addr[24643]= 1272139887;
assign addr[24644]= 1145766716;
assign addr[24645]= 1013581418;
assign addr[24646]= 876254528;
assign addr[24647]= 734482665;
assign addr[24648]= 588984994;
assign addr[24649]= 440499581;
assign addr[24650]= 289779648;
assign addr[24651]= 137589750;
assign addr[24652]= -15298099;
assign addr[24653]= -168108346;
assign addr[24654]= -320065829;
assign addr[24655]= -470399716;
assign addr[24656]= -618347408;
assign addr[24657]= -763158411;
assign addr[24658]= -904098143;
assign addr[24659]= -1040451659;
assign addr[24660]= -1171527280;
assign addr[24661]= -1296660098;
assign addr[24662]= -1415215352;
assign addr[24663]= -1526591649;
assign addr[24664]= -1630224009;
assign addr[24665]= -1725586737;
assign addr[24666]= -1812196087;
assign addr[24667]= -1889612716;
assign addr[24668]= -1957443913;
assign addr[24669]= -2015345591;
assign addr[24670]= -2063024031;
assign addr[24671]= -2100237377;
assign addr[24672]= -2126796855;
assign addr[24673]= -2142567738;
assign addr[24674]= -2147470025;
assign addr[24675]= -2141478848;
assign addr[24676]= -2124624598;
assign addr[24677]= -2096992772;
assign addr[24678]= -2058723538;
assign addr[24679]= -2010011024;
assign addr[24680]= -1951102334;
assign addr[24681]= -1882296293;
assign addr[24682]= -1803941934;
assign addr[24683]= -1716436725;
assign addr[24684]= -1620224553;
assign addr[24685]= -1515793473;
assign addr[24686]= -1403673233;
assign addr[24687]= -1284432584;
assign addr[24688]= -1158676398;
assign addr[24689]= -1027042599;
assign addr[24690]= -890198924;
assign addr[24691]= -748839539;
assign addr[24692]= -603681519;
assign addr[24693]= -455461206;
assign addr[24694]= -304930476;
assign addr[24695]= -152852926;
assign addr[24696]= 0;
assign addr[24697]= 152852926;
assign addr[24698]= 304930476;
assign addr[24699]= 455461206;
assign addr[24700]= 603681519;
assign addr[24701]= 748839539;
assign addr[24702]= 890198924;
assign addr[24703]= 1027042599;
assign addr[24704]= 1158676398;
assign addr[24705]= 1284432584;
assign addr[24706]= 1403673233;
assign addr[24707]= 1515793473;
assign addr[24708]= 1620224553;
assign addr[24709]= 1716436725;
assign addr[24710]= 1803941934;
assign addr[24711]= 1882296293;
assign addr[24712]= 1951102334;
assign addr[24713]= 2010011024;
assign addr[24714]= 2058723538;
assign addr[24715]= 2096992772;
assign addr[24716]= 2124624598;
assign addr[24717]= 2141478848;
assign addr[24718]= 2147470025;
assign addr[24719]= 2142567738;
assign addr[24720]= 2126796855;
assign addr[24721]= 2100237377;
assign addr[24722]= 2063024031;
assign addr[24723]= 2015345591;
assign addr[24724]= 1957443913;
assign addr[24725]= 1889612716;
assign addr[24726]= 1812196087;
assign addr[24727]= 1725586737;
assign addr[24728]= 1630224009;
assign addr[24729]= 1526591649;
assign addr[24730]= 1415215352;
assign addr[24731]= 1296660098;
assign addr[24732]= 1171527280;
assign addr[24733]= 1040451659;
assign addr[24734]= 904098143;
assign addr[24735]= 763158411;
assign addr[24736]= 618347408;
assign addr[24737]= 470399716;
assign addr[24738]= 320065829;
assign addr[24739]= 168108346;
assign addr[24740]= 15298099;
assign addr[24741]= -137589750;
assign addr[24742]= -289779648;
assign addr[24743]= -440499581;
assign addr[24744]= -588984994;
assign addr[24745]= -734482665;
assign addr[24746]= -876254528;
assign addr[24747]= -1013581418;
assign addr[24748]= -1145766716;
assign addr[24749]= -1272139887;
assign addr[24750]= -1392059879;
assign addr[24751]= -1504918373;
assign addr[24752]= -1610142873;
assign addr[24753]= -1707199606;
assign addr[24754]= -1795596234;
assign addr[24755]= -1874884346;
assign addr[24756]= -1944661739;
assign addr[24757]= -2004574453;
assign addr[24758]= -2054318569;
assign addr[24759]= -2093641749;
assign addr[24760]= -2122344521;
assign addr[24761]= -2140281282;
assign addr[24762]= -2147361045;
assign addr[24763]= -2143547897;
assign addr[24764]= -2128861181;
assign addr[24765]= -2103375398;
assign addr[24766]= -2067219829;
assign addr[24767]= -2020577882;
assign addr[24768]= -1963686155;
assign addr[24769]= -1896833245;
assign addr[24770]= -1820358275;
assign addr[24771]= -1734649179;
assign addr[24772]= -1640140734;
assign addr[24773]= -1537312353;
assign addr[24774]= -1426685652;
assign addr[24775]= -1308821808;
assign addr[24776]= -1184318708;
assign addr[24777]= -1053807919;
assign addr[24778]= -917951481;
assign addr[24779]= -777438554;
assign addr[24780]= -632981917;
assign addr[24781]= -485314355;
assign addr[24782]= -335184940;
assign addr[24783]= -183355234;
assign addr[24784]= -30595422;
assign addr[24785]= 122319591;
assign addr[24786]= 274614114;
assign addr[24787]= 425515602;
assign addr[24788]= 574258580;
assign addr[24789]= 720088517;
assign addr[24790]= 862265664;
assign addr[24791]= 1000068799;
assign addr[24792]= 1132798888;
assign addr[24793]= 1259782632;
assign addr[24794]= 1380375881;
assign addr[24795]= 1493966902;
assign addr[24796]= 1599979481;
assign addr[24797]= 1697875851;
assign addr[24798]= 1787159411;
assign addr[24799]= 1867377253;
assign addr[24800]= 1938122457;
assign addr[24801]= 1999036154;
assign addr[24802]= 2049809346;
assign addr[24803]= 2090184478;
assign addr[24804]= 2119956737;
assign addr[24805]= 2138975100;
assign addr[24806]= 2147143090;
assign addr[24807]= 2144419275;
assign addr[24808]= 2130817471;
assign addr[24809]= 2106406677;
assign addr[24810]= 2071310720;
assign addr[24811]= 2025707632;
assign addr[24812]= 1969828744;
assign addr[24813]= 1903957513;
assign addr[24814]= 1828428082;
assign addr[24815]= 1743623590;
assign addr[24816]= 1649974225;
assign addr[24817]= 1547955041;
assign addr[24818]= 1438083551;
assign addr[24819]= 1320917099;
assign addr[24820]= 1197050035;
assign addr[24821]= 1067110699;
assign addr[24822]= 931758235;
assign addr[24823]= 791679244;
assign addr[24824]= 647584304;
assign addr[24825]= 500204365;
assign addr[24826]= 350287041;
assign addr[24827]= 198592817;
assign addr[24828]= 45891193;
assign addr[24829]= -107043224;
assign addr[24830]= -259434643;
assign addr[24831]= -410510029;
assign addr[24832]= -559503022;
assign addr[24833]= -705657826;
assign addr[24834]= -848233042;
assign addr[24835]= -986505429;
assign addr[24836]= -1119773573;
assign addr[24837]= -1247361445;
assign addr[24838]= -1368621831;
assign addr[24839]= -1482939614;
assign addr[24840]= -1589734894;
assign addr[24841]= -1688465931;
assign addr[24842]= -1778631892;
assign addr[24843]= -1859775393;
assign addr[24844]= -1931484818;
assign addr[24845]= -1993396407;
assign addr[24846]= -2045196100;
assign addr[24847]= -2086621133;
assign addr[24848]= -2117461370;
assign addr[24849]= -2137560369;
assign addr[24850]= -2146816171;
assign addr[24851]= -2145181827;
assign addr[24852]= -2132665626;
assign addr[24853]= -2109331059;
assign addr[24854]= -2075296495;
assign addr[24855]= -2030734582;
assign addr[24856]= -1975871368;
assign addr[24857]= -1910985158;
assign addr[24858]= -1836405100;
assign addr[24859]= -1752509516;
assign addr[24860]= -1659723983;
assign addr[24861]= -1558519173;
assign addr[24862]= -1449408469;
assign addr[24863]= -1332945355;
assign addr[24864]= -1209720613;
assign addr[24865]= -1080359326;
assign addr[24866]= -945517704;
assign addr[24867]= -805879757;
assign addr[24868]= -662153826;
assign addr[24869]= -515068990;
assign addr[24870]= -365371365;
assign addr[24871]= -213820322;
assign addr[24872]= -61184634;
assign addr[24873]= 91761426;
assign addr[24874]= 244242007;
assign addr[24875]= 395483624;
assign addr[24876]= 544719071;
assign addr[24877]= 691191324;
assign addr[24878]= 834157373;
assign addr[24879]= 972891995;
assign addr[24880]= 1106691431;
assign addr[24881]= 1234876957;
assign addr[24882]= 1356798326;
assign addr[24883]= 1471837070;
assign addr[24884]= 1579409630;
assign addr[24885]= 1678970324;
assign addr[24886]= 1770014111;
assign addr[24887]= 1852079154;
assign addr[24888]= 1924749160;
assign addr[24889]= 1987655498;
assign addr[24890]= 2040479063;
assign addr[24891]= 2082951896;
assign addr[24892]= 2114858546;
assign addr[24893]= 2136037160;
assign addr[24894]= 2146380306;
assign addr[24895]= 2145835515;
assign addr[24896]= 2134405552;
assign addr[24897]= 2112148396;
assign addr[24898]= 2079176953;
assign addr[24899]= 2035658475;
assign addr[24900]= 1981813720;
assign addr[24901]= 1917915825;
assign addr[24902]= 1844288924;
assign addr[24903]= 1761306505;
assign addr[24904]= 1669389513;
assign addr[24905]= 1569004214;
assign addr[24906]= 1460659832;
assign addr[24907]= 1344905966;
assign addr[24908]= 1222329801;
assign addr[24909]= 1093553126;
assign addr[24910]= 959229189;
assign addr[24911]= 820039373;
assign addr[24912]= 676689746;
assign addr[24913]= 529907477;
assign addr[24914]= 380437148;
assign addr[24915]= 229036977;
assign addr[24916]= 76474970;
assign addr[24917]= -76474970;
assign addr[24918]= -229036977;
assign addr[24919]= -380437148;
assign addr[24920]= -529907477;
assign addr[24921]= -676689746;
assign addr[24922]= -820039373;
assign addr[24923]= -959229189;
assign addr[24924]= -1093553126;
assign addr[24925]= -1222329801;
assign addr[24926]= -1344905966;
assign addr[24927]= -1460659832;
assign addr[24928]= -1569004214;
assign addr[24929]= -1669389513;
assign addr[24930]= -1761306505;
assign addr[24931]= -1844288924;
assign addr[24932]= -1917915825;
assign addr[24933]= -1981813720;
assign addr[24934]= -2035658475;
assign addr[24935]= -2079176953;
assign addr[24936]= -2112148396;
assign addr[24937]= -2134405552;
assign addr[24938]= -2145835515;
assign addr[24939]= -2146380306;
assign addr[24940]= -2136037160;
assign addr[24941]= -2114858546;
assign addr[24942]= -2082951896;
assign addr[24943]= -2040479063;
assign addr[24944]= -1987655498;
assign addr[24945]= -1924749160;
assign addr[24946]= -1852079154;
assign addr[24947]= -1770014111;
assign addr[24948]= -1678970324;
assign addr[24949]= -1579409630;
assign addr[24950]= -1471837070;
assign addr[24951]= -1356798326;
assign addr[24952]= -1234876957;
assign addr[24953]= -1106691431;
assign addr[24954]= -972891995;
assign addr[24955]= -834157373;
assign addr[24956]= -691191324;
assign addr[24957]= -544719071;
assign addr[24958]= -395483624;
assign addr[24959]= -244242007;
assign addr[24960]= -91761426;
assign addr[24961]= 61184634;
assign addr[24962]= 213820322;
assign addr[24963]= 365371365;
assign addr[24964]= 515068990;
assign addr[24965]= 662153826;
assign addr[24966]= 805879757;
assign addr[24967]= 945517704;
assign addr[24968]= 1080359326;
assign addr[24969]= 1209720613;
assign addr[24970]= 1332945355;
assign addr[24971]= 1449408469;
assign addr[24972]= 1558519173;
assign addr[24973]= 1659723983;
assign addr[24974]= 1752509516;
assign addr[24975]= 1836405100;
assign addr[24976]= 1910985158;
assign addr[24977]= 1975871368;
assign addr[24978]= 2030734582;
assign addr[24979]= 2075296495;
assign addr[24980]= 2109331059;
assign addr[24981]= 2132665626;
assign addr[24982]= 2145181827;
assign addr[24983]= 2146816171;
assign addr[24984]= 2137560369;
assign addr[24985]= 2117461370;
assign addr[24986]= 2086621133;
assign addr[24987]= 2045196100;
assign addr[24988]= 1993396407;
assign addr[24989]= 1931484818;
assign addr[24990]= 1859775393;
assign addr[24991]= 1778631892;
assign addr[24992]= 1688465931;
assign addr[24993]= 1589734894;
assign addr[24994]= 1482939614;
assign addr[24995]= 1368621831;
assign addr[24996]= 1247361445;
assign addr[24997]= 1119773573;
assign addr[24998]= 986505429;
assign addr[24999]= 848233042;
assign addr[25000]= 705657826;
assign addr[25001]= 559503022;
assign addr[25002]= 410510029;
assign addr[25003]= 259434643;
assign addr[25004]= 107043224;
assign addr[25005]= -45891193;
assign addr[25006]= -198592817;
assign addr[25007]= -350287041;
assign addr[25008]= -500204365;
assign addr[25009]= -647584304;
assign addr[25010]= -791679244;
assign addr[25011]= -931758235;
assign addr[25012]= -1067110699;
assign addr[25013]= -1197050035;
assign addr[25014]= -1320917099;
assign addr[25015]= -1438083551;
assign addr[25016]= -1547955041;
assign addr[25017]= -1649974225;
assign addr[25018]= -1743623590;
assign addr[25019]= -1828428082;
assign addr[25020]= -1903957513;
assign addr[25021]= -1969828744;
assign addr[25022]= -2025707632;
assign addr[25023]= -2071310720;
assign addr[25024]= -2106406677;
assign addr[25025]= -2130817471;
assign addr[25026]= -2144419275;
assign addr[25027]= -2147143090;
assign addr[25028]= -2138975100;
assign addr[25029]= -2119956737;
assign addr[25030]= -2090184478;
assign addr[25031]= -2049809346;
assign addr[25032]= -1999036154;
assign addr[25033]= -1938122457;
assign addr[25034]= -1867377253;
assign addr[25035]= -1787159411;
assign addr[25036]= -1697875851;
assign addr[25037]= -1599979481;
assign addr[25038]= -1493966902;
assign addr[25039]= -1380375881;
assign addr[25040]= -1259782632;
assign addr[25041]= -1132798888;
assign addr[25042]= -1000068799;
assign addr[25043]= -862265664;
assign addr[25044]= -720088517;
assign addr[25045]= -574258580;
assign addr[25046]= -425515602;
assign addr[25047]= -274614114;
assign addr[25048]= -122319591;
assign addr[25049]= 30595422;
assign addr[25050]= 183355234;
assign addr[25051]= 335184940;
assign addr[25052]= 485314355;
assign addr[25053]= 632981917;
assign addr[25054]= 777438554;
assign addr[25055]= 917951481;
assign addr[25056]= 1053807919;
assign addr[25057]= 1184318708;
assign addr[25058]= 1308821808;
assign addr[25059]= 1426685652;
assign addr[25060]= 1537312353;
assign addr[25061]= 1640140734;
assign addr[25062]= 1734649179;
assign addr[25063]= 1820358275;
assign addr[25064]= 1896833245;
assign addr[25065]= 1963686155;
assign addr[25066]= 2020577882;
assign addr[25067]= 2067219829;
assign addr[25068]= 2103375398;
assign addr[25069]= 2128861181;
assign addr[25070]= 2143547897;
assign addr[25071]= 2147361045;
assign addr[25072]= 2140281282;
assign addr[25073]= 2122344521;
assign addr[25074]= 2093641749;
assign addr[25075]= 2054318569;
assign addr[25076]= 2004574453;
assign addr[25077]= 1944661739;
assign addr[25078]= 1874884346;
assign addr[25079]= 1795596234;
assign addr[25080]= 1707199606;
assign addr[25081]= 1610142873;
assign addr[25082]= 1504918373;
assign addr[25083]= 1392059879;
assign addr[25084]= 1272139887;
assign addr[25085]= 1145766716;
assign addr[25086]= 1013581418;
assign addr[25087]= 876254528;
assign addr[25088]= 734482665;
assign addr[25089]= 588984994;
assign addr[25090]= 440499581;
assign addr[25091]= 289779648;
assign addr[25092]= 137589750;
assign addr[25093]= -15298099;
assign addr[25094]= -168108346;
assign addr[25095]= -320065829;
assign addr[25096]= -470399716;
assign addr[25097]= -618347408;
assign addr[25098]= -763158411;
assign addr[25099]= -904098143;
assign addr[25100]= -1040451659;
assign addr[25101]= -1171527280;
assign addr[25102]= -1296660098;
assign addr[25103]= -1415215352;
assign addr[25104]= -1526591649;
assign addr[25105]= -1630224009;
assign addr[25106]= -1725586737;
assign addr[25107]= -1812196087;
assign addr[25108]= -1889612716;
assign addr[25109]= -1957443913;
assign addr[25110]= -2015345591;
assign addr[25111]= -2063024031;
assign addr[25112]= -2100237377;
assign addr[25113]= -2126796855;
assign addr[25114]= -2142567738;
assign addr[25115]= -2147470025;
assign addr[25116]= -2141478848;
assign addr[25117]= -2124624598;
assign addr[25118]= -2096992772;
assign addr[25119]= -2058723538;
assign addr[25120]= -2010011024;
assign addr[25121]= -1951102334;
assign addr[25122]= -1882296293;
assign addr[25123]= -1803941934;
assign addr[25124]= -1716436725;
assign addr[25125]= -1620224553;
assign addr[25126]= -1515793473;
assign addr[25127]= -1403673233;
assign addr[25128]= -1284432584;
assign addr[25129]= -1158676398;
assign addr[25130]= -1027042599;
assign addr[25131]= -890198924;
assign addr[25132]= -748839539;
assign addr[25133]= -603681519;
assign addr[25134]= -455461206;
assign addr[25135]= -304930476;
assign addr[25136]= -152852926;
assign addr[25137]= 0;
assign addr[25138]= 152852926;
assign addr[25139]= 304930476;
assign addr[25140]= 455461206;
assign addr[25141]= 603681519;
assign addr[25142]= 748839539;
assign addr[25143]= 890198924;
assign addr[25144]= 1027042599;
assign addr[25145]= 1158676398;
assign addr[25146]= 1284432584;
assign addr[25147]= 1403673233;
assign addr[25148]= 1515793473;
assign addr[25149]= 1620224553;
assign addr[25150]= 1716436725;
assign addr[25151]= 1803941934;
assign addr[25152]= 1882296293;
assign addr[25153]= 1951102334;
assign addr[25154]= 2010011024;
assign addr[25155]= 2058723538;
assign addr[25156]= 2096992772;
assign addr[25157]= 2124624598;
assign addr[25158]= 2141478848;
assign addr[25159]= 2147470025;
assign addr[25160]= 2142567738;
assign addr[25161]= 2126796855;
assign addr[25162]= 2100237377;
assign addr[25163]= 2063024031;
assign addr[25164]= 2015345591;
assign addr[25165]= 1957443913;
assign addr[25166]= 1889612716;
assign addr[25167]= 1812196087;
assign addr[25168]= 1725586737;
assign addr[25169]= 1630224009;
assign addr[25170]= 1526591649;
assign addr[25171]= 1415215352;
assign addr[25172]= 1296660098;
assign addr[25173]= 1171527280;
assign addr[25174]= 1040451659;
assign addr[25175]= 904098143;
assign addr[25176]= 763158411;
assign addr[25177]= 618347408;
assign addr[25178]= 470399716;
assign addr[25179]= 320065829;
assign addr[25180]= 168108346;
assign addr[25181]= 15298099;
assign addr[25182]= -137589750;
assign addr[25183]= -289779648;
assign addr[25184]= -440499581;
assign addr[25185]= -588984994;
assign addr[25186]= -734482665;
assign addr[25187]= -876254528;
assign addr[25188]= -1013581418;
assign addr[25189]= -1145766716;
assign addr[25190]= -1272139887;
assign addr[25191]= -1392059879;
assign addr[25192]= -1504918373;
assign addr[25193]= -1610142873;
assign addr[25194]= -1707199606;
assign addr[25195]= -1795596234;
assign addr[25196]= -1874884346;
assign addr[25197]= -1944661739;
assign addr[25198]= -2004574453;
assign addr[25199]= -2054318569;
assign addr[25200]= -2093641749;
assign addr[25201]= -2122344521;
assign addr[25202]= -2140281282;
assign addr[25203]= -2147361045;
assign addr[25204]= -2143547897;
assign addr[25205]= -2128861181;
assign addr[25206]= -2103375398;
assign addr[25207]= -2067219829;
assign addr[25208]= -2020577882;
assign addr[25209]= -1963686155;
assign addr[25210]= -1896833245;
assign addr[25211]= -1820358275;
assign addr[25212]= -1734649179;
assign addr[25213]= -1640140734;
assign addr[25214]= -1537312353;
assign addr[25215]= -1426685652;
assign addr[25216]= -1308821808;
assign addr[25217]= -1184318708;
assign addr[25218]= -1053807919;
assign addr[25219]= -917951481;
assign addr[25220]= -777438554;
assign addr[25221]= -632981917;
assign addr[25222]= -485314355;
assign addr[25223]= -335184940;
assign addr[25224]= -183355234;
assign addr[25225]= -30595422;
assign addr[25226]= 122319591;
assign addr[25227]= 274614114;
assign addr[25228]= 425515602;
assign addr[25229]= 574258580;
assign addr[25230]= 720088517;
assign addr[25231]= 862265664;
assign addr[25232]= 1000068799;
assign addr[25233]= 1132798888;
assign addr[25234]= 1259782632;
assign addr[25235]= 1380375881;
assign addr[25236]= 1493966902;
assign addr[25237]= 1599979481;
assign addr[25238]= 1697875851;
assign addr[25239]= 1787159411;
assign addr[25240]= 1867377253;
assign addr[25241]= 1938122457;
assign addr[25242]= 1999036154;
assign addr[25243]= 2049809346;
assign addr[25244]= 2090184478;
assign addr[25245]= 2119956737;
assign addr[25246]= 2138975100;
assign addr[25247]= 2147143090;
assign addr[25248]= 2144419275;
assign addr[25249]= 2130817471;
assign addr[25250]= 2106406677;
assign addr[25251]= 2071310720;
assign addr[25252]= 2025707632;
assign addr[25253]= 1969828744;
assign addr[25254]= 1903957513;
assign addr[25255]= 1828428082;
assign addr[25256]= 1743623590;
assign addr[25257]= 1649974225;
assign addr[25258]= 1547955041;
assign addr[25259]= 1438083551;
assign addr[25260]= 1320917099;
assign addr[25261]= 1197050035;
assign addr[25262]= 1067110699;
assign addr[25263]= 931758235;
assign addr[25264]= 791679244;
assign addr[25265]= 647584304;
assign addr[25266]= 500204365;
assign addr[25267]= 350287041;
assign addr[25268]= 198592817;
assign addr[25269]= 45891193;
assign addr[25270]= -107043224;
assign addr[25271]= -259434643;
assign addr[25272]= -410510029;
assign addr[25273]= -559503022;
assign addr[25274]= -705657826;
assign addr[25275]= -848233042;
assign addr[25276]= -986505429;
assign addr[25277]= -1119773573;
assign addr[25278]= -1247361445;
assign addr[25279]= -1368621831;
assign addr[25280]= -1482939614;
assign addr[25281]= -1589734894;
assign addr[25282]= -1688465931;
assign addr[25283]= -1778631892;
assign addr[25284]= -1859775393;
assign addr[25285]= -1931484818;
assign addr[25286]= -1993396407;
assign addr[25287]= -2045196100;
assign addr[25288]= -2086621133;
assign addr[25289]= -2117461370;
assign addr[25290]= -2137560369;
assign addr[25291]= -2146816171;
assign addr[25292]= -2145181827;
assign addr[25293]= -2132665626;
assign addr[25294]= -2109331059;
assign addr[25295]= -2075296495;
assign addr[25296]= -2030734582;
assign addr[25297]= -1975871368;
assign addr[25298]= -1910985158;
assign addr[25299]= -1836405100;
assign addr[25300]= -1752509516;
assign addr[25301]= -1659723983;
assign addr[25302]= -1558519173;
assign addr[25303]= -1449408469;
assign addr[25304]= -1332945355;
assign addr[25305]= -1209720613;
assign addr[25306]= -1080359326;
assign addr[25307]= -945517704;
assign addr[25308]= -805879757;
assign addr[25309]= -662153826;
assign addr[25310]= -515068990;
assign addr[25311]= -365371365;
assign addr[25312]= -213820322;
assign addr[25313]= -61184634;
assign addr[25314]= 91761426;
assign addr[25315]= 244242007;
assign addr[25316]= 395483624;
assign addr[25317]= 544719071;
assign addr[25318]= 691191324;
assign addr[25319]= 834157373;
assign addr[25320]= 972891995;
assign addr[25321]= 1106691431;
assign addr[25322]= 1234876957;
assign addr[25323]= 1356798326;
assign addr[25324]= 1471837070;
assign addr[25325]= 1579409630;
assign addr[25326]= 1678970324;
assign addr[25327]= 1770014111;
assign addr[25328]= 1852079154;
assign addr[25329]= 1924749160;
assign addr[25330]= 1987655498;
assign addr[25331]= 2040479063;
assign addr[25332]= 2082951896;
assign addr[25333]= 2114858546;
assign addr[25334]= 2136037160;
assign addr[25335]= 2146380306;
assign addr[25336]= 2145835515;
assign addr[25337]= 2134405552;
assign addr[25338]= 2112148396;
assign addr[25339]= 2079176953;
assign addr[25340]= 2035658475;
assign addr[25341]= 1981813720;
assign addr[25342]= 1917915825;
assign addr[25343]= 1844288924;
assign addr[25344]= 1761306505;
assign addr[25345]= 1669389513;
assign addr[25346]= 1569004214;
assign addr[25347]= 1460659832;
assign addr[25348]= 1344905966;
assign addr[25349]= 1222329801;
assign addr[25350]= 1093553126;
assign addr[25351]= 959229189;
assign addr[25352]= 820039373;
assign addr[25353]= 676689746;
assign addr[25354]= 529907477;
assign addr[25355]= 380437148;
assign addr[25356]= 229036977;
assign addr[25357]= 76474970;
assign addr[25358]= -76474970;
assign addr[25359]= -229036977;
assign addr[25360]= -380437148;
assign addr[25361]= -529907477;
assign addr[25362]= -676689746;
assign addr[25363]= -820039373;
assign addr[25364]= -959229189;
assign addr[25365]= -1093553126;
assign addr[25366]= -1222329801;
assign addr[25367]= -1344905966;
assign addr[25368]= -1460659832;
assign addr[25369]= -1569004214;
assign addr[25370]= -1669389513;
assign addr[25371]= -1761306505;
assign addr[25372]= -1844288924;
assign addr[25373]= -1917915825;
assign addr[25374]= -1981813720;
assign addr[25375]= -2035658475;
assign addr[25376]= -2079176953;
assign addr[25377]= -2112148396;
assign addr[25378]= -2134405552;
assign addr[25379]= -2145835515;
assign addr[25380]= -2146380306;
assign addr[25381]= -2136037160;
assign addr[25382]= -2114858546;
assign addr[25383]= -2082951896;
assign addr[25384]= -2040479063;
assign addr[25385]= -1987655498;
assign addr[25386]= -1924749160;
assign addr[25387]= -1852079154;
assign addr[25388]= -1770014111;
assign addr[25389]= -1678970324;
assign addr[25390]= -1579409630;
assign addr[25391]= -1471837070;
assign addr[25392]= -1356798326;
assign addr[25393]= -1234876957;
assign addr[25394]= -1106691431;
assign addr[25395]= -972891995;
assign addr[25396]= -834157373;
assign addr[25397]= -691191324;
assign addr[25398]= -544719071;
assign addr[25399]= -395483624;
assign addr[25400]= -244242007;
assign addr[25401]= -91761426;
assign addr[25402]= 61184634;
assign addr[25403]= 213820322;
assign addr[25404]= 365371365;
assign addr[25405]= 515068990;
assign addr[25406]= 662153826;
assign addr[25407]= 805879757;
assign addr[25408]= 945517704;
assign addr[25409]= 1080359326;
assign addr[25410]= 1209720613;
assign addr[25411]= 1332945355;
assign addr[25412]= 1449408469;
assign addr[25413]= 1558519173;
assign addr[25414]= 1659723983;
assign addr[25415]= 1752509516;
assign addr[25416]= 1836405100;
assign addr[25417]= 1910985158;
assign addr[25418]= 1975871368;
assign addr[25419]= 2030734582;
assign addr[25420]= 2075296495;
assign addr[25421]= 2109331059;
assign addr[25422]= 2132665626;
assign addr[25423]= 2145181827;
assign addr[25424]= 2146816171;
assign addr[25425]= 2137560369;
assign addr[25426]= 2117461370;
assign addr[25427]= 2086621133;
assign addr[25428]= 2045196100;
assign addr[25429]= 1993396407;
assign addr[25430]= 1931484818;
assign addr[25431]= 1859775393;
assign addr[25432]= 1778631892;
assign addr[25433]= 1688465931;
assign addr[25434]= 1589734894;
assign addr[25435]= 1482939614;
assign addr[25436]= 1368621831;
assign addr[25437]= 1247361445;
assign addr[25438]= 1119773573;
assign addr[25439]= 986505429;
assign addr[25440]= 848233042;
assign addr[25441]= 705657826;
assign addr[25442]= 559503022;
assign addr[25443]= 410510029;
assign addr[25444]= 259434643;
assign addr[25445]= 107043224;
assign addr[25446]= -45891193;
assign addr[25447]= -198592817;
assign addr[25448]= -350287041;
assign addr[25449]= -500204365;
assign addr[25450]= -647584304;
assign addr[25451]= -791679244;
assign addr[25452]= -931758235;
assign addr[25453]= -1067110699;
assign addr[25454]= -1197050035;
assign addr[25455]= -1320917099;
assign addr[25456]= -1438083551;
assign addr[25457]= -1547955041;
assign addr[25458]= -1649974225;
assign addr[25459]= -1743623590;
assign addr[25460]= -1828428082;
assign addr[25461]= -1903957513;
assign addr[25462]= -1969828744;
assign addr[25463]= -2025707632;
assign addr[25464]= -2071310720;
assign addr[25465]= -2106406677;
assign addr[25466]= -2130817471;
assign addr[25467]= -2144419275;
assign addr[25468]= -2147143090;
assign addr[25469]= -2138975100;
assign addr[25470]= -2119956737;
assign addr[25471]= -2090184478;
assign addr[25472]= -2049809346;
assign addr[25473]= -1999036154;
assign addr[25474]= -1938122457;
assign addr[25475]= -1867377253;
assign addr[25476]= -1787159411;
assign addr[25477]= -1697875851;
assign addr[25478]= -1599979481;
assign addr[25479]= -1493966902;
assign addr[25480]= -1380375881;
assign addr[25481]= -1259782632;
assign addr[25482]= -1132798888;
assign addr[25483]= -1000068799;
assign addr[25484]= -862265664;
assign addr[25485]= -720088517;
assign addr[25486]= -574258580;
assign addr[25487]= -425515602;
assign addr[25488]= -274614114;
assign addr[25489]= -122319591;
assign addr[25490]= 30595422;
assign addr[25491]= 183355234;
assign addr[25492]= 335184940;
assign addr[25493]= 485314355;
assign addr[25494]= 632981917;
assign addr[25495]= 777438554;
assign addr[25496]= 917951481;
assign addr[25497]= 1053807919;
assign addr[25498]= 1184318708;
assign addr[25499]= 1308821808;
assign addr[25500]= 1426685652;
assign addr[25501]= 1537312353;
assign addr[25502]= 1640140734;
assign addr[25503]= 1734649179;
assign addr[25504]= 1820358275;
assign addr[25505]= 1896833245;
assign addr[25506]= 1963686155;
assign addr[25507]= 2020577882;
assign addr[25508]= 2067219829;
assign addr[25509]= 2103375398;
assign addr[25510]= 2128861181;
assign addr[25511]= 2143547897;
assign addr[25512]= 2147361045;
assign addr[25513]= 2140281282;
assign addr[25514]= 2122344521;
assign addr[25515]= 2093641749;
assign addr[25516]= 2054318569;
assign addr[25517]= 2004574453;
assign addr[25518]= 1944661739;
assign addr[25519]= 1874884346;
assign addr[25520]= 1795596234;
assign addr[25521]= 1707199606;
assign addr[25522]= 1610142873;
assign addr[25523]= 1504918373;
assign addr[25524]= 1392059879;
assign addr[25525]= 1272139887;
assign addr[25526]= 1145766716;
assign addr[25527]= 1013581418;
assign addr[25528]= 876254528;
assign addr[25529]= 734482665;
assign addr[25530]= 588984994;
assign addr[25531]= 440499581;
assign addr[25532]= 289779648;
assign addr[25533]= 137589750;
assign addr[25534]= -15298099;
assign addr[25535]= -168108346;
assign addr[25536]= -320065829;
assign addr[25537]= -470399716;
assign addr[25538]= -618347408;
assign addr[25539]= -763158411;
assign addr[25540]= -904098143;
assign addr[25541]= -1040451659;
assign addr[25542]= -1171527280;
assign addr[25543]= -1296660098;
assign addr[25544]= -1415215352;
assign addr[25545]= -1526591649;
assign addr[25546]= -1630224009;
assign addr[25547]= -1725586737;
assign addr[25548]= -1812196087;
assign addr[25549]= -1889612716;
assign addr[25550]= -1957443913;
assign addr[25551]= -2015345591;
assign addr[25552]= -2063024031;
assign addr[25553]= -2100237377;
assign addr[25554]= -2126796855;
assign addr[25555]= -2142567738;
assign addr[25556]= -2147470025;
assign addr[25557]= -2141478848;
assign addr[25558]= -2124624598;
assign addr[25559]= -2096992772;
assign addr[25560]= -2058723538;
assign addr[25561]= -2010011024;
assign addr[25562]= -1951102334;
assign addr[25563]= -1882296293;
assign addr[25564]= -1803941934;
assign addr[25565]= -1716436725;
assign addr[25566]= -1620224553;
assign addr[25567]= -1515793473;
assign addr[25568]= -1403673233;
assign addr[25569]= -1284432584;
assign addr[25570]= -1158676398;
assign addr[25571]= -1027042599;
assign addr[25572]= -890198924;
assign addr[25573]= -748839539;
assign addr[25574]= -603681519;
assign addr[25575]= -455461206;
assign addr[25576]= -304930476;
assign addr[25577]= -152852926;
assign addr[25578]= 0;
assign addr[25579]= 152852926;
assign addr[25580]= 304930476;
assign addr[25581]= 455461206;
assign addr[25582]= 603681519;
assign addr[25583]= 748839539;
assign addr[25584]= 890198924;
assign addr[25585]= 1027042599;
assign addr[25586]= 1158676398;
assign addr[25587]= 1284432584;
assign addr[25588]= 1403673233;
assign addr[25589]= 1515793473;
assign addr[25590]= 1620224553;
assign addr[25591]= 1716436725;
assign addr[25592]= 1803941934;
assign addr[25593]= 1882296293;
assign addr[25594]= 1951102334;
assign addr[25595]= 2010011024;
assign addr[25596]= 2058723538;
assign addr[25597]= 2096992772;
assign addr[25598]= 2124624598;
assign addr[25599]= 2141478848;
assign addr[25600]= 2147470025;
assign addr[25601]= 2142567738;
assign addr[25602]= 2126796855;
assign addr[25603]= 2100237377;
assign addr[25604]= 2063024031;
assign addr[25605]= 2015345591;
assign addr[25606]= 1957443913;
assign addr[25607]= 1889612716;
assign addr[25608]= 1812196087;
assign addr[25609]= 1725586737;
assign addr[25610]= 1630224009;
assign addr[25611]= 1526591649;
assign addr[25612]= 1415215352;
assign addr[25613]= 1296660098;
assign addr[25614]= 1171527280;
assign addr[25615]= 1040451659;
assign addr[25616]= 904098143;
assign addr[25617]= 763158411;
assign addr[25618]= 618347408;
assign addr[25619]= 470399716;
assign addr[25620]= 320065829;
assign addr[25621]= 168108346;
assign addr[25622]= 15298099;
assign addr[25623]= -137589750;
assign addr[25624]= -289779648;
assign addr[25625]= -440499581;
assign addr[25626]= -588984994;
assign addr[25627]= -734482665;
assign addr[25628]= -876254528;
assign addr[25629]= -1013581418;
assign addr[25630]= -1145766716;
assign addr[25631]= -1272139887;
assign addr[25632]= -1392059879;
assign addr[25633]= -1504918373;
assign addr[25634]= -1610142873;
assign addr[25635]= -1707199606;
assign addr[25636]= -1795596234;
assign addr[25637]= -1874884346;
assign addr[25638]= -1944661739;
assign addr[25639]= -2004574453;
assign addr[25640]= -2054318569;
assign addr[25641]= -2093641749;
assign addr[25642]= -2122344521;
assign addr[25643]= -2140281282;
assign addr[25644]= -2147361045;
assign addr[25645]= -2143547897;
assign addr[25646]= -2128861181;
assign addr[25647]= -2103375398;
assign addr[25648]= -2067219829;
assign addr[25649]= -2020577882;
assign addr[25650]= -1963686155;
assign addr[25651]= -1896833245;
assign addr[25652]= -1820358275;
assign addr[25653]= -1734649179;
assign addr[25654]= -1640140734;
assign addr[25655]= -1537312353;
assign addr[25656]= -1426685652;
assign addr[25657]= -1308821808;
assign addr[25658]= -1184318708;
assign addr[25659]= -1053807919;
assign addr[25660]= -917951481;
assign addr[25661]= -777438554;
assign addr[25662]= -632981917;
assign addr[25663]= -485314355;
assign addr[25664]= -335184940;
assign addr[25665]= -183355234;
assign addr[25666]= -30595422;
assign addr[25667]= 122319591;
assign addr[25668]= 274614114;
assign addr[25669]= 425515602;
assign addr[25670]= 574258580;
assign addr[25671]= 720088517;
assign addr[25672]= 862265664;
assign addr[25673]= 1000068799;
assign addr[25674]= 1132798888;
assign addr[25675]= 1259782632;
assign addr[25676]= 1380375881;
assign addr[25677]= 1493966902;
assign addr[25678]= 1599979481;
assign addr[25679]= 1697875851;
assign addr[25680]= 1787159411;
assign addr[25681]= 1867377253;
assign addr[25682]= 1938122457;
assign addr[25683]= 1999036154;
assign addr[25684]= 2049809346;
assign addr[25685]= 2090184478;
assign addr[25686]= 2119956737;
assign addr[25687]= 2138975100;
assign addr[25688]= 2147143090;
assign addr[25689]= 2144419275;
assign addr[25690]= 2130817471;
assign addr[25691]= 2106406677;
assign addr[25692]= 2071310720;
assign addr[25693]= 2025707632;
assign addr[25694]= 1969828744;
assign addr[25695]= 1903957513;
assign addr[25696]= 1828428082;
assign addr[25697]= 1743623590;
assign addr[25698]= 1649974225;
assign addr[25699]= 1547955041;
assign addr[25700]= 1438083551;
assign addr[25701]= 1320917099;
assign addr[25702]= 1197050035;
assign addr[25703]= 1067110699;
assign addr[25704]= 931758235;
assign addr[25705]= 791679244;
assign addr[25706]= 647584304;
assign addr[25707]= 500204365;
assign addr[25708]= 350287041;
assign addr[25709]= 198592817;
assign addr[25710]= 45891193;
assign addr[25711]= -107043224;
assign addr[25712]= -259434643;
assign addr[25713]= -410510029;
assign addr[25714]= -559503022;
assign addr[25715]= -705657826;
assign addr[25716]= -848233042;
assign addr[25717]= -986505429;
assign addr[25718]= -1119773573;
assign addr[25719]= -1247361445;
assign addr[25720]= -1368621831;
assign addr[25721]= -1482939614;
assign addr[25722]= -1589734894;
assign addr[25723]= -1688465931;
assign addr[25724]= -1778631892;
assign addr[25725]= -1859775393;
assign addr[25726]= -1931484818;
assign addr[25727]= -1993396407;
assign addr[25728]= -2045196100;
assign addr[25729]= -2086621133;
assign addr[25730]= -2117461370;
assign addr[25731]= -2137560369;
assign addr[25732]= -2146816171;
assign addr[25733]= -2145181827;
assign addr[25734]= -2132665626;
assign addr[25735]= -2109331059;
assign addr[25736]= -2075296495;
assign addr[25737]= -2030734582;
assign addr[25738]= -1975871368;
assign addr[25739]= -1910985158;
assign addr[25740]= -1836405100;
assign addr[25741]= -1752509516;
assign addr[25742]= -1659723983;
assign addr[25743]= -1558519173;
assign addr[25744]= -1449408469;
assign addr[25745]= -1332945355;
assign addr[25746]= -1209720613;
assign addr[25747]= -1080359326;
assign addr[25748]= -945517704;
assign addr[25749]= -805879757;
assign addr[25750]= -662153826;
assign addr[25751]= -515068990;
assign addr[25752]= -365371365;
assign addr[25753]= -213820322;
assign addr[25754]= -61184634;
assign addr[25755]= 91761426;
assign addr[25756]= 244242007;
assign addr[25757]= 395483624;
assign addr[25758]= 544719071;
assign addr[25759]= 691191324;
assign addr[25760]= 834157373;
assign addr[25761]= 972891995;
assign addr[25762]= 1106691431;
assign addr[25763]= 1234876957;
assign addr[25764]= 1356798326;
assign addr[25765]= 1471837070;
assign addr[25766]= 1579409630;
assign addr[25767]= 1678970324;
assign addr[25768]= 1770014111;
assign addr[25769]= 1852079154;
assign addr[25770]= 1924749160;
assign addr[25771]= 1987655498;
assign addr[25772]= 2040479063;
assign addr[25773]= 2082951896;
assign addr[25774]= 2114858546;
assign addr[25775]= 2136037160;
assign addr[25776]= 2146380306;
assign addr[25777]= 2145835515;
assign addr[25778]= 2134405552;
assign addr[25779]= 2112148396;
assign addr[25780]= 2079176953;
assign addr[25781]= 2035658475;
assign addr[25782]= 1981813720;
assign addr[25783]= 1917915825;
assign addr[25784]= 1844288924;
assign addr[25785]= 1761306505;
assign addr[25786]= 1669389513;
assign addr[25787]= 1569004214;
assign addr[25788]= 1460659832;
assign addr[25789]= 1344905966;
assign addr[25790]= 1222329801;
assign addr[25791]= 1093553126;
assign addr[25792]= 959229189;
assign addr[25793]= 820039373;
assign addr[25794]= 676689746;
assign addr[25795]= 529907477;
assign addr[25796]= 380437148;
assign addr[25797]= 229036977;
assign addr[25798]= 76474970;
assign addr[25799]= -76474970;
assign addr[25800]= -229036977;
assign addr[25801]= -380437148;
assign addr[25802]= -529907477;
assign addr[25803]= -676689746;
assign addr[25804]= -820039373;
assign addr[25805]= -959229189;
assign addr[25806]= -1093553126;
assign addr[25807]= -1222329801;
assign addr[25808]= -1344905966;
assign addr[25809]= -1460659832;
assign addr[25810]= -1569004214;
assign addr[25811]= -1669389513;
assign addr[25812]= -1761306505;
assign addr[25813]= -1844288924;
assign addr[25814]= -1917915825;
assign addr[25815]= -1981813720;
assign addr[25816]= -2035658475;
assign addr[25817]= -2079176953;
assign addr[25818]= -2112148396;
assign addr[25819]= -2134405552;
assign addr[25820]= -2145835515;
assign addr[25821]= -2146380306;
assign addr[25822]= -2136037160;
assign addr[25823]= -2114858546;
assign addr[25824]= -2082951896;
assign addr[25825]= -2040479063;
assign addr[25826]= -1987655498;
assign addr[25827]= -1924749160;
assign addr[25828]= -1852079154;
assign addr[25829]= -1770014111;
assign addr[25830]= -1678970324;
assign addr[25831]= -1579409630;
assign addr[25832]= -1471837070;
assign addr[25833]= -1356798326;
assign addr[25834]= -1234876957;
assign addr[25835]= -1106691431;
assign addr[25836]= -972891995;
assign addr[25837]= -834157373;
assign addr[25838]= -691191324;
assign addr[25839]= -544719071;
assign addr[25840]= -395483624;
assign addr[25841]= -244242007;
assign addr[25842]= -91761426;
assign addr[25843]= 61184634;
assign addr[25844]= 213820322;
assign addr[25845]= 365371365;
assign addr[25846]= 515068990;
assign addr[25847]= 662153826;
assign addr[25848]= 805879757;
assign addr[25849]= 945517704;
assign addr[25850]= 1080359326;
assign addr[25851]= 1209720613;
assign addr[25852]= 1332945355;
assign addr[25853]= 1449408469;
assign addr[25854]= 1558519173;
assign addr[25855]= 1659723983;
assign addr[25856]= 1752509516;
assign addr[25857]= 1836405100;
assign addr[25858]= 1910985158;
assign addr[25859]= 1975871368;
assign addr[25860]= 2030734582;
assign addr[25861]= 2075296495;
assign addr[25862]= 2109331059;
assign addr[25863]= 2132665626;
assign addr[25864]= 2145181827;
assign addr[25865]= 2146816171;
assign addr[25866]= 2137560369;
assign addr[25867]= 2117461370;
assign addr[25868]= 2086621133;
assign addr[25869]= 2045196100;
assign addr[25870]= 1993396407;
assign addr[25871]= 1931484818;
assign addr[25872]= 1859775393;
assign addr[25873]= 1778631892;
assign addr[25874]= 1688465931;
assign addr[25875]= 1589734894;
assign addr[25876]= 1482939614;
assign addr[25877]= 1368621831;
assign addr[25878]= 1247361445;
assign addr[25879]= 1119773573;
assign addr[25880]= 986505429;
assign addr[25881]= 848233042;
assign addr[25882]= 705657826;
assign addr[25883]= 559503022;
assign addr[25884]= 410510029;
assign addr[25885]= 259434643;
assign addr[25886]= 107043224;
assign addr[25887]= -45891193;
assign addr[25888]= -198592817;
assign addr[25889]= -350287041;
assign addr[25890]= -500204365;
assign addr[25891]= -647584304;
assign addr[25892]= -791679244;
assign addr[25893]= -931758235;
assign addr[25894]= -1067110699;
assign addr[25895]= -1197050035;
assign addr[25896]= -1320917099;
assign addr[25897]= -1438083551;
assign addr[25898]= -1547955041;
assign addr[25899]= -1649974225;
assign addr[25900]= -1743623590;
assign addr[25901]= -1828428082;
assign addr[25902]= -1903957513;
assign addr[25903]= -1969828744;
assign addr[25904]= -2025707632;
assign addr[25905]= -2071310720;
assign addr[25906]= -2106406677;
assign addr[25907]= -2130817471;
assign addr[25908]= -2144419275;
assign addr[25909]= -2147143090;
assign addr[25910]= -2138975100;
assign addr[25911]= -2119956737;
assign addr[25912]= -2090184478;
assign addr[25913]= -2049809346;
assign addr[25914]= -1999036154;
assign addr[25915]= -1938122457;
assign addr[25916]= -1867377253;
assign addr[25917]= -1787159411;
assign addr[25918]= -1697875851;
assign addr[25919]= -1599979481;
assign addr[25920]= -1493966902;
assign addr[25921]= -1380375881;
assign addr[25922]= -1259782632;
assign addr[25923]= -1132798888;
assign addr[25924]= -1000068799;
assign addr[25925]= -862265664;
assign addr[25926]= -720088517;
assign addr[25927]= -574258580;
assign addr[25928]= -425515602;
assign addr[25929]= -274614114;
assign addr[25930]= -122319591;
assign addr[25931]= 30595422;
assign addr[25932]= 183355234;
assign addr[25933]= 335184940;
assign addr[25934]= 485314355;
assign addr[25935]= 632981917;
assign addr[25936]= 777438554;
assign addr[25937]= 917951481;
assign addr[25938]= 1053807919;
assign addr[25939]= 1184318708;
assign addr[25940]= 1308821808;
assign addr[25941]= 1426685652;
assign addr[25942]= 1537312353;
assign addr[25943]= 1640140734;
assign addr[25944]= 1734649179;
assign addr[25945]= 1820358275;
assign addr[25946]= 1896833245;
assign addr[25947]= 1963686155;
assign addr[25948]= 2020577882;
assign addr[25949]= 2067219829;
assign addr[25950]= 2103375398;
assign addr[25951]= 2128861181;
assign addr[25952]= 2143547897;
assign addr[25953]= 2147361045;
assign addr[25954]= 2140281282;
assign addr[25955]= 2122344521;
assign addr[25956]= 2093641749;
assign addr[25957]= 2054318569;
assign addr[25958]= 2004574453;
assign addr[25959]= 1944661739;
assign addr[25960]= 1874884346;
assign addr[25961]= 1795596234;
assign addr[25962]= 1707199606;
assign addr[25963]= 1610142873;
assign addr[25964]= 1504918373;
assign addr[25965]= 1392059879;
assign addr[25966]= 1272139887;
assign addr[25967]= 1145766716;
assign addr[25968]= 1013581418;
assign addr[25969]= 876254528;
assign addr[25970]= 734482665;
assign addr[25971]= 588984994;
assign addr[25972]= 440499581;
assign addr[25973]= 289779648;
assign addr[25974]= 137589750;
assign addr[25975]= -15298099;
assign addr[25976]= -168108346;
assign addr[25977]= -320065829;
assign addr[25978]= -470399716;
assign addr[25979]= -618347408;
assign addr[25980]= -763158411;
assign addr[25981]= -904098143;
assign addr[25982]= -1040451659;
assign addr[25983]= -1171527280;
assign addr[25984]= -1296660098;
assign addr[25985]= -1415215352;
assign addr[25986]= -1526591649;
assign addr[25987]= -1630224009;
assign addr[25988]= -1725586737;
assign addr[25989]= -1812196087;
assign addr[25990]= -1889612716;
assign addr[25991]= -1957443913;
assign addr[25992]= -2015345591;
assign addr[25993]= -2063024031;
assign addr[25994]= -2100237377;
assign addr[25995]= -2126796855;
assign addr[25996]= -2142567738;
assign addr[25997]= -2147470025;
assign addr[25998]= -2141478848;
assign addr[25999]= -2124624598;
assign addr[26000]= -2096992772;
assign addr[26001]= -2058723538;
assign addr[26002]= -2010011024;
assign addr[26003]= -1951102334;
assign addr[26004]= -1882296293;
assign addr[26005]= -1803941934;
assign addr[26006]= -1716436725;
assign addr[26007]= -1620224553;
assign addr[26008]= -1515793473;
assign addr[26009]= -1403673233;
assign addr[26010]= -1284432584;
assign addr[26011]= -1158676398;
assign addr[26012]= -1027042599;
assign addr[26013]= -890198924;
assign addr[26014]= -748839539;
assign addr[26015]= -603681519;
assign addr[26016]= -455461206;
assign addr[26017]= -304930476;
assign addr[26018]= -152852926;
assign addr[26019]= 0;
assign addr[26020]= 152852926;
assign addr[26021]= 304930476;
assign addr[26022]= 455461206;
assign addr[26023]= 603681519;
assign addr[26024]= 748839539;
assign addr[26025]= 890198924;
assign addr[26026]= 1027042599;
assign addr[26027]= 1158676398;
assign addr[26028]= 1284432584;
assign addr[26029]= 1403673233;
assign addr[26030]= 1515793473;
assign addr[26031]= 1620224553;
assign addr[26032]= 1716436725;
assign addr[26033]= 1803941934;
assign addr[26034]= 1882296293;
assign addr[26035]= 1951102334;
assign addr[26036]= 2010011024;
assign addr[26037]= 2058723538;
assign addr[26038]= 2096992772;
assign addr[26039]= 2124624598;
assign addr[26040]= 2141478848;
assign addr[26041]= 2147470025;
assign addr[26042]= 2142567738;
assign addr[26043]= 2126796855;
assign addr[26044]= 2100237377;
assign addr[26045]= 2063024031;
assign addr[26046]= 2015345591;
assign addr[26047]= 1957443913;
assign addr[26048]= 1889612716;
assign addr[26049]= 1812196087;
assign addr[26050]= 1725586737;
assign addr[26051]= 1630224009;
assign addr[26052]= 1526591649;
assign addr[26053]= 1415215352;
assign addr[26054]= 1296660098;
assign addr[26055]= 1171527280;
assign addr[26056]= 1040451659;
assign addr[26057]= 904098143;
assign addr[26058]= 763158411;
assign addr[26059]= 618347408;
assign addr[26060]= 470399716;
assign addr[26061]= 320065829;
assign addr[26062]= 168108346;
assign addr[26063]= 15298099;
assign addr[26064]= -137589750;
assign addr[26065]= -289779648;
assign addr[26066]= -440499581;
assign addr[26067]= -588984994;
assign addr[26068]= -734482665;
assign addr[26069]= -876254528;
assign addr[26070]= -1013581418;
assign addr[26071]= -1145766716;
assign addr[26072]= -1272139887;
assign addr[26073]= -1392059879;
assign addr[26074]= -1504918373;
assign addr[26075]= -1610142873;
assign addr[26076]= -1707199606;
assign addr[26077]= -1795596234;
assign addr[26078]= -1874884346;
assign addr[26079]= -1944661739;
assign addr[26080]= -2004574453;
assign addr[26081]= -2054318569;
assign addr[26082]= -2093641749;
assign addr[26083]= -2122344521;
assign addr[26084]= -2140281282;
assign addr[26085]= -2147361045;
assign addr[26086]= -2143547897;
assign addr[26087]= -2128861181;
assign addr[26088]= -2103375398;
assign addr[26089]= -2067219829;
assign addr[26090]= -2020577882;
assign addr[26091]= -1963686155;
assign addr[26092]= -1896833245;
assign addr[26093]= -1820358275;
assign addr[26094]= -1734649179;
assign addr[26095]= -1640140734;
assign addr[26096]= -1537312353;
assign addr[26097]= -1426685652;
assign addr[26098]= -1308821808;
assign addr[26099]= -1184318708;
assign addr[26100]= -1053807919;
assign addr[26101]= -917951481;
assign addr[26102]= -777438554;
assign addr[26103]= -632981917;
assign addr[26104]= -485314355;
assign addr[26105]= -335184940;
assign addr[26106]= -183355234;
assign addr[26107]= -30595422;
assign addr[26108]= 122319591;
assign addr[26109]= 274614114;
assign addr[26110]= 425515602;
assign addr[26111]= 574258580;
assign addr[26112]= 720088517;
assign addr[26113]= 862265664;
assign addr[26114]= 1000068799;
assign addr[26115]= 1132798888;
assign addr[26116]= 1259782632;
assign addr[26117]= 1380375881;
assign addr[26118]= 1493966902;
assign addr[26119]= 1599979481;
assign addr[26120]= 1697875851;
assign addr[26121]= 1787159411;
assign addr[26122]= 1867377253;
assign addr[26123]= 1938122457;
assign addr[26124]= 1999036154;
assign addr[26125]= 2049809346;
assign addr[26126]= 2090184478;
assign addr[26127]= 2119956737;
assign addr[26128]= 2138975100;
assign addr[26129]= 2147143090;
assign addr[26130]= 2144419275;
assign addr[26131]= 2130817471;
assign addr[26132]= 2106406677;
assign addr[26133]= 2071310720;
assign addr[26134]= 2025707632;
assign addr[26135]= 1969828744;
assign addr[26136]= 1903957513;
assign addr[26137]= 1828428082;
assign addr[26138]= 1743623590;
assign addr[26139]= 1649974225;
assign addr[26140]= 1547955041;
assign addr[26141]= 1438083551;
assign addr[26142]= 1320917099;
assign addr[26143]= 1197050035;
assign addr[26144]= 1067110699;
assign addr[26145]= 931758235;
assign addr[26146]= 791679244;
assign addr[26147]= 647584304;
assign addr[26148]= 500204365;
assign addr[26149]= 350287041;
assign addr[26150]= 198592817;
assign addr[26151]= 45891193;
assign addr[26152]= -107043224;
assign addr[26153]= -259434643;
assign addr[26154]= -410510029;
assign addr[26155]= -559503022;
assign addr[26156]= -705657826;
assign addr[26157]= -848233042;
assign addr[26158]= -986505429;
assign addr[26159]= -1119773573;
assign addr[26160]= -1247361445;
assign addr[26161]= -1368621831;
assign addr[26162]= -1482939614;
assign addr[26163]= -1589734894;
assign addr[26164]= -1688465931;
assign addr[26165]= -1778631892;
assign addr[26166]= -1859775393;
assign addr[26167]= -1931484818;
assign addr[26168]= -1993396407;
assign addr[26169]= -2045196100;
assign addr[26170]= -2086621133;
assign addr[26171]= -2117461370;
assign addr[26172]= -2137560369;
assign addr[26173]= -2146816171;
assign addr[26174]= -2145181827;
assign addr[26175]= -2132665626;
assign addr[26176]= -2109331059;
assign addr[26177]= -2075296495;
assign addr[26178]= -2030734582;
assign addr[26179]= -1975871368;
assign addr[26180]= -1910985158;
assign addr[26181]= -1836405100;
assign addr[26182]= -1752509516;
assign addr[26183]= -1659723983;
assign addr[26184]= -1558519173;
assign addr[26185]= -1449408469;
assign addr[26186]= -1332945355;
assign addr[26187]= -1209720613;
assign addr[26188]= -1080359326;
assign addr[26189]= -945517704;
assign addr[26190]= -805879757;
assign addr[26191]= -662153826;
assign addr[26192]= -515068990;
assign addr[26193]= -365371365;
assign addr[26194]= -213820322;
assign addr[26195]= -61184634;
assign addr[26196]= 91761426;
assign addr[26197]= 244242007;
assign addr[26198]= 395483624;
assign addr[26199]= 544719071;
assign addr[26200]= 691191324;
assign addr[26201]= 834157373;
assign addr[26202]= 972891995;
assign addr[26203]= 1106691431;
assign addr[26204]= 1234876957;
assign addr[26205]= 1356798326;
assign addr[26206]= 1471837070;
assign addr[26207]= 1579409630;
assign addr[26208]= 1678970324;
assign addr[26209]= 1770014111;
assign addr[26210]= 1852079154;
assign addr[26211]= 1924749160;
assign addr[26212]= 1987655498;
assign addr[26213]= 2040479063;
assign addr[26214]= 2082951896;
assign addr[26215]= 2114858546;
assign addr[26216]= 2136037160;
assign addr[26217]= 2146380306;
assign addr[26218]= 2145835515;
assign addr[26219]= 2134405552;
assign addr[26220]= 2112148396;
assign addr[26221]= 2079176953;
assign addr[26222]= 2035658475;
assign addr[26223]= 1981813720;
assign addr[26224]= 1917915825;
assign addr[26225]= 1844288924;
assign addr[26226]= 1761306505;
assign addr[26227]= 1669389513;
assign addr[26228]= 1569004214;
assign addr[26229]= 1460659832;
assign addr[26230]= 1344905966;
assign addr[26231]= 1222329801;
assign addr[26232]= 1093553126;
assign addr[26233]= 959229189;
assign addr[26234]= 820039373;
assign addr[26235]= 676689746;
assign addr[26236]= 529907477;
assign addr[26237]= 380437148;
assign addr[26238]= 229036977;
assign addr[26239]= 76474970;
assign addr[26240]= -76474970;
assign addr[26241]= -229036977;
assign addr[26242]= -380437148;
assign addr[26243]= -529907477;
assign addr[26244]= -676689746;
assign addr[26245]= -820039373;
assign addr[26246]= -959229189;
assign addr[26247]= -1093553126;
assign addr[26248]= -1222329801;
assign addr[26249]= -1344905966;
assign addr[26250]= -1460659832;
assign addr[26251]= -1569004214;
assign addr[26252]= -1669389513;
assign addr[26253]= -1761306505;
assign addr[26254]= -1844288924;
assign addr[26255]= -1917915825;
assign addr[26256]= -1981813720;
assign addr[26257]= -2035658475;
assign addr[26258]= -2079176953;
assign addr[26259]= -2112148396;
assign addr[26260]= -2134405552;
assign addr[26261]= -2145835515;
assign addr[26262]= -2146380306;
assign addr[26263]= -2136037160;
assign addr[26264]= -2114858546;
assign addr[26265]= -2082951896;
assign addr[26266]= -2040479063;
assign addr[26267]= -1987655498;
assign addr[26268]= -1924749160;
assign addr[26269]= -1852079154;
assign addr[26270]= -1770014111;
assign addr[26271]= -1678970324;
assign addr[26272]= -1579409630;
assign addr[26273]= -1471837070;
assign addr[26274]= -1356798326;
assign addr[26275]= -1234876957;
assign addr[26276]= -1106691431;
assign addr[26277]= -972891995;
assign addr[26278]= -834157373;
assign addr[26279]= -691191324;
assign addr[26280]= -544719071;
assign addr[26281]= -395483624;
assign addr[26282]= -244242007;
assign addr[26283]= -91761426;
assign addr[26284]= 61184634;
assign addr[26285]= 213820322;
assign addr[26286]= 365371365;
assign addr[26287]= 515068990;
assign addr[26288]= 662153826;
assign addr[26289]= 805879757;
assign addr[26290]= 945517704;
assign addr[26291]= 1080359326;
assign addr[26292]= 1209720613;
assign addr[26293]= 1332945355;
assign addr[26294]= 1449408469;
assign addr[26295]= 1558519173;
assign addr[26296]= 1659723983;
assign addr[26297]= 1752509516;
assign addr[26298]= 1836405100;
assign addr[26299]= 1910985158;
assign addr[26300]= 1975871368;
assign addr[26301]= 2030734582;
assign addr[26302]= 2075296495;
assign addr[26303]= 2109331059;
assign addr[26304]= 2132665626;
assign addr[26305]= 2145181827;
assign addr[26306]= 2146816171;
assign addr[26307]= 2137560369;
assign addr[26308]= 2117461370;
assign addr[26309]= 2086621133;
assign addr[26310]= 2045196100;
assign addr[26311]= 1993396407;
assign addr[26312]= 1931484818;
assign addr[26313]= 1859775393;
assign addr[26314]= 1778631892;
assign addr[26315]= 1688465931;
assign addr[26316]= 1589734894;
assign addr[26317]= 1482939614;
assign addr[26318]= 1368621831;
assign addr[26319]= 1247361445;
assign addr[26320]= 1119773573;
assign addr[26321]= 986505429;
assign addr[26322]= 848233042;
assign addr[26323]= 705657826;
assign addr[26324]= 559503022;
assign addr[26325]= 410510029;
assign addr[26326]= 259434643;
assign addr[26327]= 107043224;
assign addr[26328]= -45891193;
assign addr[26329]= -198592817;
assign addr[26330]= -350287041;
assign addr[26331]= -500204365;
assign addr[26332]= -647584304;
assign addr[26333]= -791679244;
assign addr[26334]= -931758235;
assign addr[26335]= -1067110699;
assign addr[26336]= -1197050035;
assign addr[26337]= -1320917099;
assign addr[26338]= -1438083551;
assign addr[26339]= -1547955041;
assign addr[26340]= -1649974225;
assign addr[26341]= -1743623590;
assign addr[26342]= -1828428082;
assign addr[26343]= -1903957513;
assign addr[26344]= -1969828744;
assign addr[26345]= -2025707632;
assign addr[26346]= -2071310720;
assign addr[26347]= -2106406677;
assign addr[26348]= -2130817471;
assign addr[26349]= -2144419275;
assign addr[26350]= -2147143090;
assign addr[26351]= -2138975100;
assign addr[26352]= -2119956737;
assign addr[26353]= -2090184478;
assign addr[26354]= -2049809346;
assign addr[26355]= -1999036154;
assign addr[26356]= -1938122457;
assign addr[26357]= -1867377253;
assign addr[26358]= -1787159411;
assign addr[26359]= -1697875851;
assign addr[26360]= -1599979481;
assign addr[26361]= -1493966902;
assign addr[26362]= -1380375881;
assign addr[26363]= -1259782632;
assign addr[26364]= -1132798888;
assign addr[26365]= -1000068799;
assign addr[26366]= -862265664;
assign addr[26367]= -720088517;
assign addr[26368]= -574258580;
assign addr[26369]= -425515602;
assign addr[26370]= -274614114;
assign addr[26371]= -122319591;
assign addr[26372]= 30595422;
assign addr[26373]= 183355234;
assign addr[26374]= 335184940;
assign addr[26375]= 485314355;
assign addr[26376]= 632981917;
assign addr[26377]= 777438554;
assign addr[26378]= 917951481;
assign addr[26379]= 1053807919;
assign addr[26380]= 1184318708;
assign addr[26381]= 1308821808;
assign addr[26382]= 1426685652;
assign addr[26383]= 1537312353;
assign addr[26384]= 1640140734;
assign addr[26385]= 1734649179;
assign addr[26386]= 1820358275;
assign addr[26387]= 1896833245;
assign addr[26388]= 1963686155;
assign addr[26389]= 2020577882;
assign addr[26390]= 2067219829;
assign addr[26391]= 2103375398;
assign addr[26392]= 2128861181;
assign addr[26393]= 2143547897;
assign addr[26394]= 2147361045;
assign addr[26395]= 2140281282;
assign addr[26396]= 2122344521;
assign addr[26397]= 2093641749;
assign addr[26398]= 2054318569;
assign addr[26399]= 2004574453;
assign addr[26400]= 1944661739;
assign addr[26401]= 1874884346;
assign addr[26402]= 1795596234;
assign addr[26403]= 1707199606;
assign addr[26404]= 1610142873;
assign addr[26405]= 1504918373;
assign addr[26406]= 1392059879;
assign addr[26407]= 1272139887;
assign addr[26408]= 1145766716;
assign addr[26409]= 1013581418;
assign addr[26410]= 876254528;
assign addr[26411]= 734482665;
assign addr[26412]= 588984994;
assign addr[26413]= 440499581;
assign addr[26414]= 289779648;
assign addr[26415]= 137589750;
assign addr[26416]= -15298099;
assign addr[26417]= -168108346;
assign addr[26418]= -320065829;
assign addr[26419]= -470399716;
assign addr[26420]= -618347408;
assign addr[26421]= -763158411;
assign addr[26422]= -904098143;
assign addr[26423]= -1040451659;
assign addr[26424]= -1171527280;
assign addr[26425]= -1296660098;
assign addr[26426]= -1415215352;
assign addr[26427]= -1526591649;
assign addr[26428]= -1630224009;
assign addr[26429]= -1725586737;
assign addr[26430]= -1812196087;
assign addr[26431]= -1889612716;
assign addr[26432]= -1957443913;
assign addr[26433]= -2015345591;
assign addr[26434]= -2063024031;
assign addr[26435]= -2100237377;
assign addr[26436]= -2126796855;
assign addr[26437]= -2142567738;
assign addr[26438]= -2147470025;
assign addr[26439]= -2141478848;
assign addr[26440]= -2124624598;
assign addr[26441]= -2096992772;
assign addr[26442]= -2058723538;
assign addr[26443]= -2010011024;
assign addr[26444]= -1951102334;
assign addr[26445]= -1882296293;
assign addr[26446]= -1803941934;
assign addr[26447]= -1716436725;
assign addr[26448]= -1620224553;
assign addr[26449]= -1515793473;
assign addr[26450]= -1403673233;
assign addr[26451]= -1284432584;
assign addr[26452]= -1158676398;
assign addr[26453]= -1027042599;
assign addr[26454]= -890198924;
assign addr[26455]= -748839539;
assign addr[26456]= -603681519;
assign addr[26457]= -455461206;
assign addr[26458]= -304930476;
assign addr[26459]= -152852926;
assign addr[26460]= 0;
assign addr[26461]= 152852926;
assign addr[26462]= 304930476;
assign addr[26463]= 455461206;
assign addr[26464]= 603681519;
assign addr[26465]= 748839539;
assign addr[26466]= 890198924;
assign addr[26467]= 1027042599;
assign addr[26468]= 1158676398;
assign addr[26469]= 1284432584;
assign addr[26470]= 1403673233;
assign addr[26471]= 1515793473;
assign addr[26472]= 1620224553;
assign addr[26473]= 1716436725;
assign addr[26474]= 1803941934;
assign addr[26475]= 1882296293;
assign addr[26476]= 1951102334;
assign addr[26477]= 2010011024;
assign addr[26478]= 2058723538;
assign addr[26479]= 2096992772;
assign addr[26480]= 2124624598;
assign addr[26481]= 2141478848;
assign addr[26482]= 2147470025;
assign addr[26483]= 2142567738;
assign addr[26484]= 2126796855;
assign addr[26485]= 2100237377;
assign addr[26486]= 2063024031;
assign addr[26487]= 2015345591;
assign addr[26488]= 1957443913;
assign addr[26489]= 1889612716;
assign addr[26490]= 1812196087;
assign addr[26491]= 1725586737;
assign addr[26492]= 1630224009;
assign addr[26493]= 1526591649;
assign addr[26494]= 1415215352;
assign addr[26495]= 1296660098;
assign addr[26496]= 1171527280;
assign addr[26497]= 1040451659;
assign addr[26498]= 904098143;
assign addr[26499]= 763158411;
assign addr[26500]= 618347408;
assign addr[26501]= 470399716;
assign addr[26502]= 320065829;
assign addr[26503]= 168108346;
assign addr[26504]= 15298099;
assign addr[26505]= -137589750;
assign addr[26506]= -289779648;
assign addr[26507]= -440499581;
assign addr[26508]= -588984994;
assign addr[26509]= -734482665;
assign addr[26510]= -876254528;
assign addr[26511]= -1013581418;
assign addr[26512]= -1145766716;
assign addr[26513]= -1272139887;
assign addr[26514]= -1392059879;
assign addr[26515]= -1504918373;
assign addr[26516]= -1610142873;
assign addr[26517]= -1707199606;
assign addr[26518]= -1795596234;
assign addr[26519]= -1874884346;
assign addr[26520]= -1944661739;
assign addr[26521]= -2004574453;
assign addr[26522]= -2054318569;
assign addr[26523]= -2093641749;
assign addr[26524]= -2122344521;
assign addr[26525]= -2140281282;
assign addr[26526]= -2147361045;
assign addr[26527]= -2143547897;
assign addr[26528]= -2128861181;
assign addr[26529]= -2103375398;
assign addr[26530]= -2067219829;
assign addr[26531]= -2020577882;
assign addr[26532]= -1963686155;
assign addr[26533]= -1896833245;
assign addr[26534]= -1820358275;
assign addr[26535]= -1734649179;
assign addr[26536]= -1640140734;
assign addr[26537]= -1537312353;
assign addr[26538]= -1426685652;
assign addr[26539]= -1308821808;
assign addr[26540]= -1184318708;
assign addr[26541]= -1053807919;
assign addr[26542]= -917951481;
assign addr[26543]= -777438554;
assign addr[26544]= -632981917;
assign addr[26545]= -485314355;
assign addr[26546]= -335184940;
assign addr[26547]= -183355234;
assign addr[26548]= -30595422;
assign addr[26549]= 122319591;
assign addr[26550]= 274614114;
assign addr[26551]= 425515602;
assign addr[26552]= 574258580;
assign addr[26553]= 720088517;
assign addr[26554]= 862265664;
assign addr[26555]= 1000068799;
assign addr[26556]= 1132798888;
assign addr[26557]= 1259782632;
assign addr[26558]= 1380375881;
assign addr[26559]= 1493966902;
assign addr[26560]= 1599979481;
assign addr[26561]= 1697875851;
assign addr[26562]= 1787159411;
assign addr[26563]= 1867377253;
assign addr[26564]= 1938122457;
assign addr[26565]= 1999036154;
assign addr[26566]= 2049809346;
assign addr[26567]= 2090184478;
assign addr[26568]= 2119956737;
assign addr[26569]= 2138975100;
assign addr[26570]= 2147143090;
assign addr[26571]= 2144419275;
assign addr[26572]= 2130817471;
assign addr[26573]= 2106406677;
assign addr[26574]= 2071310720;
assign addr[26575]= 2025707632;
assign addr[26576]= 1969828744;
assign addr[26577]= 1903957513;
assign addr[26578]= 1828428082;
assign addr[26579]= 1743623590;
assign addr[26580]= 1649974225;
assign addr[26581]= 1547955041;
assign addr[26582]= 1438083551;
assign addr[26583]= 1320917099;
assign addr[26584]= 1197050035;
assign addr[26585]= 1067110699;
assign addr[26586]= 931758235;
assign addr[26587]= 791679244;
assign addr[26588]= 647584304;
assign addr[26589]= 500204365;
assign addr[26590]= 350287041;
assign addr[26591]= 198592817;
assign addr[26592]= 45891193;
assign addr[26593]= -107043224;
assign addr[26594]= -259434643;
assign addr[26595]= -410510029;
assign addr[26596]= -559503022;
assign addr[26597]= -705657826;
assign addr[26598]= -848233042;
assign addr[26599]= -986505429;
assign addr[26600]= -1119773573;
assign addr[26601]= -1247361445;
assign addr[26602]= -1368621831;
assign addr[26603]= -1482939614;
assign addr[26604]= -1589734894;
assign addr[26605]= -1688465931;
assign addr[26606]= -1778631892;
assign addr[26607]= -1859775393;
assign addr[26608]= -1931484818;
assign addr[26609]= -1993396407;
assign addr[26610]= -2045196100;
assign addr[26611]= -2086621133;
assign addr[26612]= -2117461370;
assign addr[26613]= -2137560369;
assign addr[26614]= -2146816171;
assign addr[26615]= -2145181827;
assign addr[26616]= -2132665626;
assign addr[26617]= -2109331059;
assign addr[26618]= -2075296495;
assign addr[26619]= -2030734582;
assign addr[26620]= -1975871368;
assign addr[26621]= -1910985158;
assign addr[26622]= -1836405100;
assign addr[26623]= -1752509516;
assign addr[26624]= -1659723983;
assign addr[26625]= -1558519173;
assign addr[26626]= -1449408469;
assign addr[26627]= -1332945355;
assign addr[26628]= -1209720613;
assign addr[26629]= -1080359326;
assign addr[26630]= -945517704;
assign addr[26631]= -805879757;
assign addr[26632]= -662153826;
assign addr[26633]= -515068990;
assign addr[26634]= -365371365;
assign addr[26635]= -213820322;
assign addr[26636]= -61184634;
assign addr[26637]= 91761426;
assign addr[26638]= 244242007;
assign addr[26639]= 395483624;
assign addr[26640]= 544719071;
assign addr[26641]= 691191324;
assign addr[26642]= 834157373;
assign addr[26643]= 972891995;
assign addr[26644]= 1106691431;
assign addr[26645]= 1234876957;
assign addr[26646]= 1356798326;
assign addr[26647]= 1471837070;
assign addr[26648]= 1579409630;
assign addr[26649]= 1678970324;
assign addr[26650]= 1770014111;
assign addr[26651]= 1852079154;
assign addr[26652]= 1924749160;
assign addr[26653]= 1987655498;
assign addr[26654]= 2040479063;
assign addr[26655]= 2082951896;
assign addr[26656]= 2114858546;
assign addr[26657]= 2136037160;
assign addr[26658]= 2146380306;
assign addr[26659]= 2145835515;
assign addr[26660]= 2134405552;
assign addr[26661]= 2112148396;
assign addr[26662]= 2079176953;
assign addr[26663]= 2035658475;
assign addr[26664]= 1981813720;
assign addr[26665]= 1917915825;
assign addr[26666]= 1844288924;
assign addr[26667]= 1761306505;
assign addr[26668]= 1669389513;
assign addr[26669]= 1569004214;
assign addr[26670]= 1460659832;
assign addr[26671]= 1344905966;
assign addr[26672]= 1222329801;
assign addr[26673]= 1093553126;
assign addr[26674]= 959229189;
assign addr[26675]= 820039373;
assign addr[26676]= 676689746;
assign addr[26677]= 529907477;
assign addr[26678]= 380437148;
assign addr[26679]= 229036977;
assign addr[26680]= 76474970;
assign addr[26681]= -76474970;
assign addr[26682]= -229036977;
assign addr[26683]= -380437148;
assign addr[26684]= -529907477;
assign addr[26685]= -676689746;
assign addr[26686]= -820039373;
assign addr[26687]= -959229189;
assign addr[26688]= -1093553126;
assign addr[26689]= -1222329801;
assign addr[26690]= -1344905966;
assign addr[26691]= -1460659832;
assign addr[26692]= -1569004214;
assign addr[26693]= -1669389513;
assign addr[26694]= -1761306505;
assign addr[26695]= -1844288924;
assign addr[26696]= -1917915825;
assign addr[26697]= -1981813720;
assign addr[26698]= -2035658475;
assign addr[26699]= -2079176953;
assign addr[26700]= -2112148396;
assign addr[26701]= -2134405552;
assign addr[26702]= -2145835515;
assign addr[26703]= -2146380306;
assign addr[26704]= -2136037160;
assign addr[26705]= -2114858546;
assign addr[26706]= -2082951896;
assign addr[26707]= -2040479063;
assign addr[26708]= -1987655498;
assign addr[26709]= -1924749160;
assign addr[26710]= -1852079154;
assign addr[26711]= -1770014111;
assign addr[26712]= -1678970324;
assign addr[26713]= -1579409630;
assign addr[26714]= -1471837070;
assign addr[26715]= -1356798326;
assign addr[26716]= -1234876957;
assign addr[26717]= -1106691431;
assign addr[26718]= -972891995;
assign addr[26719]= -834157373;
assign addr[26720]= -691191324;
assign addr[26721]= -544719071;
assign addr[26722]= -395483624;
assign addr[26723]= -244242007;
assign addr[26724]= -91761426;
assign addr[26725]= 61184634;
assign addr[26726]= 213820322;
assign addr[26727]= 365371365;
assign addr[26728]= 515068990;
assign addr[26729]= 662153826;
assign addr[26730]= 805879757;
assign addr[26731]= 945517704;
assign addr[26732]= 1080359326;
assign addr[26733]= 1209720613;
assign addr[26734]= 1332945355;
assign addr[26735]= 1449408469;
assign addr[26736]= 1558519173;
assign addr[26737]= 1659723983;
assign addr[26738]= 1752509516;
assign addr[26739]= 1836405100;
assign addr[26740]= 1910985158;
assign addr[26741]= 1975871368;
assign addr[26742]= 2030734582;
assign addr[26743]= 2075296495;
assign addr[26744]= 2109331059;
assign addr[26745]= 2132665626;
assign addr[26746]= 2145181827;
assign addr[26747]= 2146816171;
assign addr[26748]= 2137560369;
assign addr[26749]= 2117461370;
assign addr[26750]= 2086621133;
assign addr[26751]= 2045196100;
assign addr[26752]= 1993396407;
assign addr[26753]= 1931484818;
assign addr[26754]= 1859775393;
assign addr[26755]= 1778631892;
assign addr[26756]= 1688465931;
assign addr[26757]= 1589734894;
assign addr[26758]= 1482939614;
assign addr[26759]= 1368621831;
assign addr[26760]= 1247361445;
assign addr[26761]= 1119773573;
assign addr[26762]= 986505429;
assign addr[26763]= 848233042;
assign addr[26764]= 705657826;
assign addr[26765]= 559503022;
assign addr[26766]= 410510029;
assign addr[26767]= 259434643;
assign addr[26768]= 107043224;
assign addr[26769]= -45891193;
assign addr[26770]= -198592817;
assign addr[26771]= -350287041;
assign addr[26772]= -500204365;
assign addr[26773]= -647584304;
assign addr[26774]= -791679244;
assign addr[26775]= -931758235;
assign addr[26776]= -1067110699;
assign addr[26777]= -1197050035;
assign addr[26778]= -1320917099;
assign addr[26779]= -1438083551;
assign addr[26780]= -1547955041;
assign addr[26781]= -1649974225;
assign addr[26782]= -1743623590;
assign addr[26783]= -1828428082;
assign addr[26784]= -1903957513;
assign addr[26785]= -1969828744;
assign addr[26786]= -2025707632;
assign addr[26787]= -2071310720;
assign addr[26788]= -2106406677;
assign addr[26789]= -2130817471;
assign addr[26790]= -2144419275;
assign addr[26791]= -2147143090;
assign addr[26792]= -2138975100;
assign addr[26793]= -2119956737;
assign addr[26794]= -2090184478;
assign addr[26795]= -2049809346;
assign addr[26796]= -1999036154;
assign addr[26797]= -1938122457;
assign addr[26798]= -1867377253;
assign addr[26799]= -1787159411;
assign addr[26800]= -1697875851;
assign addr[26801]= -1599979481;
assign addr[26802]= -1493966902;
assign addr[26803]= -1380375881;
assign addr[26804]= -1259782632;
assign addr[26805]= -1132798888;
assign addr[26806]= -1000068799;
assign addr[26807]= -862265664;
assign addr[26808]= -720088517;
assign addr[26809]= -574258580;
assign addr[26810]= -425515602;
assign addr[26811]= -274614114;
assign addr[26812]= -122319591;
assign addr[26813]= 30595422;
assign addr[26814]= 183355234;
assign addr[26815]= 335184940;
assign addr[26816]= 485314355;
assign addr[26817]= 632981917;
assign addr[26818]= 777438554;
assign addr[26819]= 917951481;
assign addr[26820]= 1053807919;
assign addr[26821]= 1184318708;
assign addr[26822]= 1308821808;
assign addr[26823]= 1426685652;
assign addr[26824]= 1537312353;
assign addr[26825]= 1640140734;
assign addr[26826]= 1734649179;
assign addr[26827]= 1820358275;
assign addr[26828]= 1896833245;
assign addr[26829]= 1963686155;
assign addr[26830]= 2020577882;
assign addr[26831]= 2067219829;
assign addr[26832]= 2103375398;
assign addr[26833]= 2128861181;
assign addr[26834]= 2143547897;
assign addr[26835]= 2147361045;
assign addr[26836]= 2140281282;
assign addr[26837]= 2122344521;
assign addr[26838]= 2093641749;
assign addr[26839]= 2054318569;
assign addr[26840]= 2004574453;
assign addr[26841]= 1944661739;
assign addr[26842]= 1874884346;
assign addr[26843]= 1795596234;
assign addr[26844]= 1707199606;
assign addr[26845]= 1610142873;
assign addr[26846]= 1504918373;
assign addr[26847]= 1392059879;
assign addr[26848]= 1272139887;
assign addr[26849]= 1145766716;
assign addr[26850]= 1013581418;
assign addr[26851]= 876254528;
assign addr[26852]= 734482665;
assign addr[26853]= 588984994;
assign addr[26854]= 440499581;
assign addr[26855]= 289779648;
assign addr[26856]= 137589750;
assign addr[26857]= -15298099;
assign addr[26858]= -168108346;
assign addr[26859]= -320065829;
assign addr[26860]= -470399716;
assign addr[26861]= -618347408;
assign addr[26862]= -763158411;
assign addr[26863]= -904098143;
assign addr[26864]= -1040451659;
assign addr[26865]= -1171527280;
assign addr[26866]= -1296660098;
assign addr[26867]= -1415215352;
assign addr[26868]= -1526591649;
assign addr[26869]= -1630224009;
assign addr[26870]= -1725586737;
assign addr[26871]= -1812196087;
assign addr[26872]= -1889612716;
assign addr[26873]= -1957443913;
assign addr[26874]= -2015345591;
assign addr[26875]= -2063024031;
assign addr[26876]= -2100237377;
assign addr[26877]= -2126796855;
assign addr[26878]= -2142567738;
assign addr[26879]= -2147470025;
assign addr[26880]= -2141478848;
assign addr[26881]= -2124624598;
assign addr[26882]= -2096992772;
assign addr[26883]= -2058723538;
assign addr[26884]= -2010011024;
assign addr[26885]= -1951102334;
assign addr[26886]= -1882296293;
assign addr[26887]= -1803941934;
assign addr[26888]= -1716436725;
assign addr[26889]= -1620224553;
assign addr[26890]= -1515793473;
assign addr[26891]= -1403673233;
assign addr[26892]= -1284432584;
assign addr[26893]= -1158676398;
assign addr[26894]= -1027042599;
assign addr[26895]= -890198924;
assign addr[26896]= -748839539;
assign addr[26897]= -603681519;
assign addr[26898]= -455461206;
assign addr[26899]= -304930476;
assign addr[26900]= -152852926;
assign addr[26901]= 0;
assign addr[26902]= 152852926;
assign addr[26903]= 304930476;
assign addr[26904]= 455461206;
assign addr[26905]= 603681519;
assign addr[26906]= 748839539;
assign addr[26907]= 890198924;
assign addr[26908]= 1027042599;
assign addr[26909]= 1158676398;
assign addr[26910]= 1284432584;
assign addr[26911]= 1403673233;
assign addr[26912]= 1515793473;
assign addr[26913]= 1620224553;
assign addr[26914]= 1716436725;
assign addr[26915]= 1803941934;
assign addr[26916]= 1882296293;
assign addr[26917]= 1951102334;
assign addr[26918]= 2010011024;
assign addr[26919]= 2058723538;
assign addr[26920]= 2096992772;
assign addr[26921]= 2124624598;
assign addr[26922]= 2141478848;
assign addr[26923]= 2147470025;
assign addr[26924]= 2142567738;
assign addr[26925]= 2126796855;
assign addr[26926]= 2100237377;
assign addr[26927]= 2063024031;
assign addr[26928]= 2015345591;
assign addr[26929]= 1957443913;
assign addr[26930]= 1889612716;
assign addr[26931]= 1812196087;
assign addr[26932]= 1725586737;
assign addr[26933]= 1630224009;
assign addr[26934]= 1526591649;
assign addr[26935]= 1415215352;
assign addr[26936]= 1296660098;
assign addr[26937]= 1171527280;
assign addr[26938]= 1040451659;
assign addr[26939]= 904098143;
assign addr[26940]= 763158411;
assign addr[26941]= 618347408;
assign addr[26942]= 470399716;
assign addr[26943]= 320065829;
assign addr[26944]= 168108346;
assign addr[26945]= 15298099;
assign addr[26946]= -137589750;
assign addr[26947]= -289779648;
assign addr[26948]= -440499581;
assign addr[26949]= -588984994;
assign addr[26950]= -734482665;
assign addr[26951]= -876254528;
assign addr[26952]= -1013581418;
assign addr[26953]= -1145766716;
assign addr[26954]= -1272139887;
assign addr[26955]= -1392059879;
assign addr[26956]= -1504918373;
assign addr[26957]= -1610142873;
assign addr[26958]= -1707199606;
assign addr[26959]= -1795596234;
assign addr[26960]= -1874884346;
assign addr[26961]= -1944661739;
assign addr[26962]= -2004574453;
assign addr[26963]= -2054318569;
assign addr[26964]= -2093641749;
assign addr[26965]= -2122344521;
assign addr[26966]= -2140281282;
assign addr[26967]= -2147361045;
assign addr[26968]= -2143547897;
assign addr[26969]= -2128861181;
assign addr[26970]= -2103375398;
assign addr[26971]= -2067219829;
assign addr[26972]= -2020577882;
assign addr[26973]= -1963686155;
assign addr[26974]= -1896833245;
assign addr[26975]= -1820358275;
assign addr[26976]= -1734649179;
assign addr[26977]= -1640140734;
assign addr[26978]= -1537312353;
assign addr[26979]= -1426685652;
assign addr[26980]= -1308821808;
assign addr[26981]= -1184318708;
assign addr[26982]= -1053807919;
assign addr[26983]= -917951481;
assign addr[26984]= -777438554;
assign addr[26985]= -632981917;
assign addr[26986]= -485314355;
assign addr[26987]= -335184940;
assign addr[26988]= -183355234;
assign addr[26989]= -30595422;
assign addr[26990]= 122319591;
assign addr[26991]= 274614114;
assign addr[26992]= 425515602;
assign addr[26993]= 574258580;
assign addr[26994]= 720088517;
assign addr[26995]= 862265664;
assign addr[26996]= 1000068799;
assign addr[26997]= 1132798888;
assign addr[26998]= 1259782632;
assign addr[26999]= 1380375881;
assign addr[27000]= 1493966902;
assign addr[27001]= 1599979481;
assign addr[27002]= 1697875851;
assign addr[27003]= 1787159411;
assign addr[27004]= 1867377253;
assign addr[27005]= 1938122457;
assign addr[27006]= 1999036154;
assign addr[27007]= 2049809346;
assign addr[27008]= 2090184478;
assign addr[27009]= 2119956737;
assign addr[27010]= 2138975100;
assign addr[27011]= 2147143090;
assign addr[27012]= 2144419275;
assign addr[27013]= 2130817471;
assign addr[27014]= 2106406677;
assign addr[27015]= 2071310720;
assign addr[27016]= 2025707632;
assign addr[27017]= 1969828744;
assign addr[27018]= 1903957513;
assign addr[27019]= 1828428082;
assign addr[27020]= 1743623590;
assign addr[27021]= 1649974225;
assign addr[27022]= 1547955041;
assign addr[27023]= 1438083551;
assign addr[27024]= 1320917099;
assign addr[27025]= 1197050035;
assign addr[27026]= 1067110699;
assign addr[27027]= 931758235;
assign addr[27028]= 791679244;
assign addr[27029]= 647584304;
assign addr[27030]= 500204365;
assign addr[27031]= 350287041;
assign addr[27032]= 198592817;
assign addr[27033]= 45891193;
assign addr[27034]= -107043224;
assign addr[27035]= -259434643;
assign addr[27036]= -410510029;
assign addr[27037]= -559503022;
assign addr[27038]= -705657826;
assign addr[27039]= -848233042;
assign addr[27040]= -986505429;
assign addr[27041]= -1119773573;
assign addr[27042]= -1247361445;
assign addr[27043]= -1368621831;
assign addr[27044]= -1482939614;
assign addr[27045]= -1589734894;
assign addr[27046]= -1688465931;
assign addr[27047]= -1778631892;
assign addr[27048]= -1859775393;
assign addr[27049]= -1931484818;
assign addr[27050]= -1993396407;
assign addr[27051]= -2045196100;
assign addr[27052]= -2086621133;
assign addr[27053]= -2117461370;
assign addr[27054]= -2137560369;
assign addr[27055]= -2146816171;
assign addr[27056]= -2145181827;
assign addr[27057]= -2132665626;
assign addr[27058]= -2109331059;
assign addr[27059]= -2075296495;
assign addr[27060]= -2030734582;
assign addr[27061]= -1975871368;
assign addr[27062]= -1910985158;
assign addr[27063]= -1836405100;
assign addr[27064]= -1752509516;
assign addr[27065]= -1659723983;
assign addr[27066]= -1558519173;
assign addr[27067]= -1449408469;
assign addr[27068]= -1332945355;
assign addr[27069]= -1209720613;
assign addr[27070]= -1080359326;
assign addr[27071]= -945517704;
assign addr[27072]= -805879757;
assign addr[27073]= -662153826;
assign addr[27074]= -515068990;
assign addr[27075]= -365371365;
assign addr[27076]= -213820322;
assign addr[27077]= -61184634;
assign addr[27078]= 91761426;
assign addr[27079]= 244242007;
assign addr[27080]= 395483624;
assign addr[27081]= 544719071;
assign addr[27082]= 691191324;
assign addr[27083]= 834157373;
assign addr[27084]= 972891995;
assign addr[27085]= 1106691431;
assign addr[27086]= 1234876957;
assign addr[27087]= 1356798326;
assign addr[27088]= 1471837070;
assign addr[27089]= 1579409630;
assign addr[27090]= 1678970324;
assign addr[27091]= 1770014111;
assign addr[27092]= 1852079154;
assign addr[27093]= 1924749160;
assign addr[27094]= 1987655498;
assign addr[27095]= 2040479063;
assign addr[27096]= 2082951896;
assign addr[27097]= 2114858546;
assign addr[27098]= 2136037160;
assign addr[27099]= 2146380306;
assign addr[27100]= 2145835515;
assign addr[27101]= 2134405552;
assign addr[27102]= 2112148396;
assign addr[27103]= 2079176953;
assign addr[27104]= 2035658475;
assign addr[27105]= 1981813720;
assign addr[27106]= 1917915825;
assign addr[27107]= 1844288924;
assign addr[27108]= 1761306505;
assign addr[27109]= 1669389513;
assign addr[27110]= 1569004214;
assign addr[27111]= 1460659832;
assign addr[27112]= 1344905966;
assign addr[27113]= 1222329801;
assign addr[27114]= 1093553126;
assign addr[27115]= 959229189;
assign addr[27116]= 820039373;
assign addr[27117]= 676689746;
assign addr[27118]= 529907477;
assign addr[27119]= 380437148;
assign addr[27120]= 229036977;
assign addr[27121]= 76474970;
assign addr[27122]= -76474970;
assign addr[27123]= -229036977;
assign addr[27124]= -380437148;
assign addr[27125]= -529907477;
assign addr[27126]= -676689746;
assign addr[27127]= -820039373;
assign addr[27128]= -959229189;
assign addr[27129]= -1093553126;
assign addr[27130]= -1222329801;
assign addr[27131]= -1344905966;
assign addr[27132]= -1460659832;
assign addr[27133]= -1569004214;
assign addr[27134]= -1669389513;
assign addr[27135]= -1761306505;
assign addr[27136]= -1844288924;
assign addr[27137]= -1917915825;
assign addr[27138]= -1981813720;
assign addr[27139]= -2035658475;
assign addr[27140]= -2079176953;
assign addr[27141]= -2112148396;
assign addr[27142]= -2134405552;
assign addr[27143]= -2145835515;
assign addr[27144]= -2146380306;
assign addr[27145]= -2136037160;
assign addr[27146]= -2114858546;
assign addr[27147]= -2082951896;
assign addr[27148]= -2040479063;
assign addr[27149]= -1987655498;
assign addr[27150]= -1924749160;
assign addr[27151]= -1852079154;
assign addr[27152]= -1770014111;
assign addr[27153]= -1678970324;
assign addr[27154]= -1579409630;
assign addr[27155]= -1471837070;
assign addr[27156]= -1356798326;
assign addr[27157]= -1234876957;
assign addr[27158]= -1106691431;
assign addr[27159]= -972891995;
assign addr[27160]= -834157373;
assign addr[27161]= -691191324;
assign addr[27162]= -544719071;
assign addr[27163]= -395483624;
assign addr[27164]= -244242007;
assign addr[27165]= -91761426;
assign addr[27166]= 61184634;
assign addr[27167]= 213820322;
assign addr[27168]= 365371365;
assign addr[27169]= 515068990;
assign addr[27170]= 662153826;
assign addr[27171]= 805879757;
assign addr[27172]= 945517704;
assign addr[27173]= 1080359326;
assign addr[27174]= 1209720613;
assign addr[27175]= 1332945355;
assign addr[27176]= 1449408469;
assign addr[27177]= 1558519173;
assign addr[27178]= 1659723983;
assign addr[27179]= 1752509516;
assign addr[27180]= 1836405100;
assign addr[27181]= 1910985158;
assign addr[27182]= 1975871368;
assign addr[27183]= 2030734582;
assign addr[27184]= 2075296495;
assign addr[27185]= 2109331059;
assign addr[27186]= 2132665626;
assign addr[27187]= 2145181827;
assign addr[27188]= 2146816171;
assign addr[27189]= 2137560369;
assign addr[27190]= 2117461370;
assign addr[27191]= 2086621133;
assign addr[27192]= 2045196100;
assign addr[27193]= 1993396407;
assign addr[27194]= 1931484818;
assign addr[27195]= 1859775393;
assign addr[27196]= 1778631892;
assign addr[27197]= 1688465931;
assign addr[27198]= 1589734894;
assign addr[27199]= 1482939614;
assign addr[27200]= 1368621831;
assign addr[27201]= 1247361445;
assign addr[27202]= 1119773573;
assign addr[27203]= 986505429;
assign addr[27204]= 848233042;
assign addr[27205]= 705657826;
assign addr[27206]= 559503022;
assign addr[27207]= 410510029;
assign addr[27208]= 259434643;
assign addr[27209]= 107043224;
assign addr[27210]= -45891193;
assign addr[27211]= -198592817;
assign addr[27212]= -350287041;
assign addr[27213]= -500204365;
assign addr[27214]= -647584304;
assign addr[27215]= -791679244;
assign addr[27216]= -931758235;
assign addr[27217]= -1067110699;
assign addr[27218]= -1197050035;
assign addr[27219]= -1320917099;
assign addr[27220]= -1438083551;
assign addr[27221]= -1547955041;
assign addr[27222]= -1649974225;
assign addr[27223]= -1743623590;
assign addr[27224]= -1828428082;
assign addr[27225]= -1903957513;
assign addr[27226]= -1969828744;
assign addr[27227]= -2025707632;
assign addr[27228]= -2071310720;
assign addr[27229]= -2106406677;
assign addr[27230]= -2130817471;
assign addr[27231]= -2144419275;
assign addr[27232]= -2147143090;
assign addr[27233]= -2138975100;
assign addr[27234]= -2119956737;
assign addr[27235]= -2090184478;
assign addr[27236]= -2049809346;
assign addr[27237]= -1999036154;
assign addr[27238]= -1938122457;
assign addr[27239]= -1867377253;
assign addr[27240]= -1787159411;
assign addr[27241]= -1697875851;
assign addr[27242]= -1599979481;
assign addr[27243]= -1493966902;
assign addr[27244]= -1380375881;
assign addr[27245]= -1259782632;
assign addr[27246]= -1132798888;
assign addr[27247]= -1000068799;
assign addr[27248]= -862265664;
assign addr[27249]= -720088517;
assign addr[27250]= -574258580;
assign addr[27251]= -425515602;
assign addr[27252]= -274614114;
assign addr[27253]= -122319591;
assign addr[27254]= 30595422;
assign addr[27255]= 183355234;
assign addr[27256]= 335184940;
assign addr[27257]= 485314355;
assign addr[27258]= 632981917;
assign addr[27259]= 777438554;
assign addr[27260]= 917951481;
assign addr[27261]= 1053807919;
assign addr[27262]= 1184318708;
assign addr[27263]= 1308821808;
assign addr[27264]= 1426685652;
assign addr[27265]= 1537312353;
assign addr[27266]= 1640140734;
assign addr[27267]= 1734649179;
assign addr[27268]= 1820358275;
assign addr[27269]= 1896833245;
assign addr[27270]= 1963686155;
assign addr[27271]= 2020577882;
assign addr[27272]= 2067219829;
assign addr[27273]= 2103375398;
assign addr[27274]= 2128861181;
assign addr[27275]= 2143547897;
assign addr[27276]= 2147361045;
assign addr[27277]= 2140281282;
assign addr[27278]= 2122344521;
assign addr[27279]= 2093641749;
assign addr[27280]= 2054318569;
assign addr[27281]= 2004574453;
assign addr[27282]= 1944661739;
assign addr[27283]= 1874884346;
assign addr[27284]= 1795596234;
assign addr[27285]= 1707199606;
assign addr[27286]= 1610142873;
assign addr[27287]= 1504918373;
assign addr[27288]= 1392059879;
assign addr[27289]= 1272139887;
assign addr[27290]= 1145766716;
assign addr[27291]= 1013581418;
assign addr[27292]= 876254528;
assign addr[27293]= 734482665;
assign addr[27294]= 588984994;
assign addr[27295]= 440499581;
assign addr[27296]= 289779648;
assign addr[27297]= 137589750;
assign addr[27298]= -15298099;
assign addr[27299]= -168108346;
assign addr[27300]= -320065829;
assign addr[27301]= -470399716;
assign addr[27302]= -618347408;
assign addr[27303]= -763158411;
assign addr[27304]= -904098143;
assign addr[27305]= -1040451659;
assign addr[27306]= -1171527280;
assign addr[27307]= -1296660098;
assign addr[27308]= -1415215352;
assign addr[27309]= -1526591649;
assign addr[27310]= -1630224009;
assign addr[27311]= -1725586737;
assign addr[27312]= -1812196087;
assign addr[27313]= -1889612716;
assign addr[27314]= -1957443913;
assign addr[27315]= -2015345591;
assign addr[27316]= -2063024031;
assign addr[27317]= -2100237377;
assign addr[27318]= -2126796855;
assign addr[27319]= -2142567738;
assign addr[27320]= -2147470025;
assign addr[27321]= -2141478848;
assign addr[27322]= -2124624598;
assign addr[27323]= -2096992772;
assign addr[27324]= -2058723538;
assign addr[27325]= -2010011024;
assign addr[27326]= -1951102334;
assign addr[27327]= -1882296293;
assign addr[27328]= -1803941934;
assign addr[27329]= -1716436725;
assign addr[27330]= -1620224553;
assign addr[27331]= -1515793473;
assign addr[27332]= -1403673233;
assign addr[27333]= -1284432584;
assign addr[27334]= -1158676398;
assign addr[27335]= -1027042599;
assign addr[27336]= -890198924;
assign addr[27337]= -748839539;
assign addr[27338]= -603681519;
assign addr[27339]= -455461206;
assign addr[27340]= -304930476;
assign addr[27341]= -152852926;
assign addr[27342]= 0;
assign addr[27343]= 152852926;
assign addr[27344]= 304930476;
assign addr[27345]= 455461206;
assign addr[27346]= 603681519;
assign addr[27347]= 748839539;
assign addr[27348]= 890198924;
assign addr[27349]= 1027042599;
assign addr[27350]= 1158676398;
assign addr[27351]= 1284432584;
assign addr[27352]= 1403673233;
assign addr[27353]= 1515793473;
assign addr[27354]= 1620224553;
assign addr[27355]= 1716436725;
assign addr[27356]= 1803941934;
assign addr[27357]= 1882296293;
assign addr[27358]= 1951102334;
assign addr[27359]= 2010011024;
assign addr[27360]= 2058723538;
assign addr[27361]= 2096992772;
assign addr[27362]= 2124624598;
assign addr[27363]= 2141478848;
assign addr[27364]= 2147470025;
assign addr[27365]= 2142567738;
assign addr[27366]= 2126796855;
assign addr[27367]= 2100237377;
assign addr[27368]= 2063024031;
assign addr[27369]= 2015345591;
assign addr[27370]= 1957443913;
assign addr[27371]= 1889612716;
assign addr[27372]= 1812196087;
assign addr[27373]= 1725586737;
assign addr[27374]= 1630224009;
assign addr[27375]= 1526591649;
assign addr[27376]= 1415215352;
assign addr[27377]= 1296660098;
assign addr[27378]= 1171527280;
assign addr[27379]= 1040451659;
assign addr[27380]= 904098143;
assign addr[27381]= 763158411;
assign addr[27382]= 618347408;
assign addr[27383]= 470399716;
assign addr[27384]= 320065829;
assign addr[27385]= 168108346;
assign addr[27386]= 15298099;
assign addr[27387]= -137589750;
assign addr[27388]= -289779648;
assign addr[27389]= -440499581;
assign addr[27390]= -588984994;
assign addr[27391]= -734482665;
assign addr[27392]= -876254528;
assign addr[27393]= -1013581418;
assign addr[27394]= -1145766716;
assign addr[27395]= -1272139887;
assign addr[27396]= -1392059879;
assign addr[27397]= -1504918373;
assign addr[27398]= -1610142873;
assign addr[27399]= -1707199606;
assign addr[27400]= -1795596234;
assign addr[27401]= -1874884346;
assign addr[27402]= -1944661739;
assign addr[27403]= -2004574453;
assign addr[27404]= -2054318569;
assign addr[27405]= -2093641749;
assign addr[27406]= -2122344521;
assign addr[27407]= -2140281282;
assign addr[27408]= -2147361045;
assign addr[27409]= -2143547897;
assign addr[27410]= -2128861181;
assign addr[27411]= -2103375398;
assign addr[27412]= -2067219829;
assign addr[27413]= -2020577882;
assign addr[27414]= -1963686155;
assign addr[27415]= -1896833245;
assign addr[27416]= -1820358275;
assign addr[27417]= -1734649179;
assign addr[27418]= -1640140734;
assign addr[27419]= -1537312353;
assign addr[27420]= -1426685652;
assign addr[27421]= -1308821808;
assign addr[27422]= -1184318708;
assign addr[27423]= -1053807919;
assign addr[27424]= -917951481;
assign addr[27425]= -777438554;
assign addr[27426]= -632981917;
assign addr[27427]= -485314355;
assign addr[27428]= -335184940;
assign addr[27429]= -183355234;
assign addr[27430]= -30595422;
assign addr[27431]= 122319591;
assign addr[27432]= 274614114;
assign addr[27433]= 425515602;
assign addr[27434]= 574258580;
assign addr[27435]= 720088517;
assign addr[27436]= 862265664;
assign addr[27437]= 1000068799;
assign addr[27438]= 1132798888;
assign addr[27439]= 1259782632;
assign addr[27440]= 1380375881;
assign addr[27441]= 1493966902;
assign addr[27442]= 1599979481;
assign addr[27443]= 1697875851;
assign addr[27444]= 1787159411;
assign addr[27445]= 1867377253;
assign addr[27446]= 1938122457;
assign addr[27447]= 1999036154;
assign addr[27448]= 2049809346;
assign addr[27449]= 2090184478;
assign addr[27450]= 2119956737;
assign addr[27451]= 2138975100;
assign addr[27452]= 2147143090;
assign addr[27453]= 2144419275;
assign addr[27454]= 2130817471;
assign addr[27455]= 2106406677;
assign addr[27456]= 2071310720;
assign addr[27457]= 2025707632;
assign addr[27458]= 1969828744;
assign addr[27459]= 1903957513;
assign addr[27460]= 1828428082;
assign addr[27461]= 1743623590;
assign addr[27462]= 1649974225;
assign addr[27463]= 1547955041;
assign addr[27464]= 1438083551;
assign addr[27465]= 1320917099;
assign addr[27466]= 1197050035;
assign addr[27467]= 1067110699;
assign addr[27468]= 931758235;
assign addr[27469]= 791679244;
assign addr[27470]= 647584304;
assign addr[27471]= 500204365;
assign addr[27472]= 350287041;
assign addr[27473]= 198592817;
assign addr[27474]= 45891193;
assign addr[27475]= -107043224;
assign addr[27476]= -259434643;
assign addr[27477]= -410510029;
assign addr[27478]= -559503022;
assign addr[27479]= -705657826;
assign addr[27480]= -848233042;
assign addr[27481]= -986505429;
assign addr[27482]= -1119773573;
assign addr[27483]= -1247361445;
assign addr[27484]= -1368621831;
assign addr[27485]= -1482939614;
assign addr[27486]= -1589734894;
assign addr[27487]= -1688465931;
assign addr[27488]= -1778631892;
assign addr[27489]= -1859775393;
assign addr[27490]= -1931484818;
assign addr[27491]= -1993396407;
assign addr[27492]= -2045196100;
assign addr[27493]= -2086621133;
assign addr[27494]= -2117461370;
assign addr[27495]= -2137560369;
assign addr[27496]= -2146816171;
assign addr[27497]= -2145181827;
assign addr[27498]= -2132665626;
assign addr[27499]= -2109331059;
assign addr[27500]= -2075296495;
assign addr[27501]= -2030734582;
assign addr[27502]= -1975871368;
assign addr[27503]= -1910985158;
assign addr[27504]= -1836405100;
assign addr[27505]= -1752509516;
assign addr[27506]= -1659723983;
assign addr[27507]= -1558519173;
assign addr[27508]= -1449408469;
assign addr[27509]= -1332945355;
assign addr[27510]= -1209720613;
assign addr[27511]= -1080359326;
assign addr[27512]= -945517704;
assign addr[27513]= -805879757;
assign addr[27514]= -662153826;
assign addr[27515]= -515068990;
assign addr[27516]= -365371365;
assign addr[27517]= -213820322;
assign addr[27518]= -61184634;
assign addr[27519]= 91761426;
assign addr[27520]= 244242007;
assign addr[27521]= 395483624;
assign addr[27522]= 544719071;
assign addr[27523]= 691191324;
assign addr[27524]= 834157373;
assign addr[27525]= 972891995;
assign addr[27526]= 1106691431;
assign addr[27527]= 1234876957;
assign addr[27528]= 1356798326;
assign addr[27529]= 1471837070;
assign addr[27530]= 1579409630;
assign addr[27531]= 1678970324;
assign addr[27532]= 1770014111;
assign addr[27533]= 1852079154;
assign addr[27534]= 1924749160;
assign addr[27535]= 1987655498;
assign addr[27536]= 2040479063;
assign addr[27537]= 2082951896;
assign addr[27538]= 2114858546;
assign addr[27539]= 2136037160;
assign addr[27540]= 2146380306;
assign addr[27541]= 2145835515;
assign addr[27542]= 2134405552;
assign addr[27543]= 2112148396;
assign addr[27544]= 2079176953;
assign addr[27545]= 2035658475;
assign addr[27546]= 1981813720;
assign addr[27547]= 1917915825;
assign addr[27548]= 1844288924;
assign addr[27549]= 1761306505;
assign addr[27550]= 1669389513;
assign addr[27551]= 1569004214;
assign addr[27552]= 1460659832;
assign addr[27553]= 1344905966;
assign addr[27554]= 1222329801;
assign addr[27555]= 1093553126;
assign addr[27556]= 959229189;
assign addr[27557]= 820039373;
assign addr[27558]= 676689746;
assign addr[27559]= 529907477;
assign addr[27560]= 380437148;
assign addr[27561]= 229036977;
assign addr[27562]= 76474970;
assign addr[27563]= -76474970;
assign addr[27564]= -229036977;
assign addr[27565]= -380437148;
assign addr[27566]= -529907477;
assign addr[27567]= -676689746;
assign addr[27568]= -820039373;
assign addr[27569]= -959229189;
assign addr[27570]= -1093553126;
assign addr[27571]= -1222329801;
assign addr[27572]= -1344905966;
assign addr[27573]= -1460659832;
assign addr[27574]= -1569004214;
assign addr[27575]= -1669389513;
assign addr[27576]= -1761306505;
assign addr[27577]= -1844288924;
assign addr[27578]= -1917915825;
assign addr[27579]= -1981813720;
assign addr[27580]= -2035658475;
assign addr[27581]= -2079176953;
assign addr[27582]= -2112148396;
assign addr[27583]= -2134405552;
assign addr[27584]= -2145835515;
assign addr[27585]= -2146380306;
assign addr[27586]= -2136037160;
assign addr[27587]= -2114858546;
assign addr[27588]= -2082951896;
assign addr[27589]= -2040479063;
assign addr[27590]= -1987655498;
assign addr[27591]= -1924749160;
assign addr[27592]= -1852079154;
assign addr[27593]= -1770014111;
assign addr[27594]= -1678970324;
assign addr[27595]= -1579409630;
assign addr[27596]= -1471837070;
assign addr[27597]= -1356798326;
assign addr[27598]= -1234876957;
assign addr[27599]= -1106691431;
assign addr[27600]= -972891995;
assign addr[27601]= -834157373;
assign addr[27602]= -691191324;
assign addr[27603]= -544719071;
assign addr[27604]= -395483624;
assign addr[27605]= -244242007;
assign addr[27606]= -91761426;
assign addr[27607]= 61184634;
assign addr[27608]= 213820322;
assign addr[27609]= 365371365;
assign addr[27610]= 515068990;
assign addr[27611]= 662153826;
assign addr[27612]= 805879757;
assign addr[27613]= 945517704;
assign addr[27614]= 1080359326;
assign addr[27615]= 1209720613;
assign addr[27616]= 1332945355;
assign addr[27617]= 1449408469;
assign addr[27618]= 1558519173;
assign addr[27619]= 1659723983;
assign addr[27620]= 1752509516;
assign addr[27621]= 1836405100;
assign addr[27622]= 1910985158;
assign addr[27623]= 1975871368;
assign addr[27624]= 2030734582;
assign addr[27625]= 2075296495;
assign addr[27626]= 2109331059;
assign addr[27627]= 2132665626;
assign addr[27628]= 2145181827;
assign addr[27629]= 2146816171;
assign addr[27630]= 2137560369;
assign addr[27631]= 2117461370;
assign addr[27632]= 2086621133;
assign addr[27633]= 2045196100;
assign addr[27634]= 1993396407;
assign addr[27635]= 1931484818;
assign addr[27636]= 1859775393;
assign addr[27637]= 1778631892;
assign addr[27638]= 1688465931;
assign addr[27639]= 1589734894;
assign addr[27640]= 1482939614;
assign addr[27641]= 1368621831;
assign addr[27642]= 1247361445;
assign addr[27643]= 1119773573;
assign addr[27644]= 986505429;
assign addr[27645]= 848233042;
assign addr[27646]= 705657826;
assign addr[27647]= 559503022;
assign addr[27648]= 410510029;
assign addr[27649]= 259434643;
assign addr[27650]= 107043224;
assign addr[27651]= -45891193;
assign addr[27652]= -198592817;
assign addr[27653]= -350287041;
assign addr[27654]= -500204365;
assign addr[27655]= -647584304;
assign addr[27656]= -791679244;
assign addr[27657]= -931758235;
assign addr[27658]= -1067110699;
assign addr[27659]= -1197050035;
assign addr[27660]= -1320917099;
assign addr[27661]= -1438083551;
assign addr[27662]= -1547955041;
assign addr[27663]= -1649974225;
assign addr[27664]= -1743623590;
assign addr[27665]= -1828428082;
assign addr[27666]= -1903957513;
assign addr[27667]= -1969828744;
assign addr[27668]= -2025707632;
assign addr[27669]= -2071310720;
assign addr[27670]= -2106406677;
assign addr[27671]= -2130817471;
assign addr[27672]= -2144419275;
assign addr[27673]= -2147143090;
assign addr[27674]= -2138975100;
assign addr[27675]= -2119956737;
assign addr[27676]= -2090184478;
assign addr[27677]= -2049809346;
assign addr[27678]= -1999036154;
assign addr[27679]= -1938122457;
assign addr[27680]= -1867377253;
assign addr[27681]= -1787159411;
assign addr[27682]= -1697875851;
assign addr[27683]= -1599979481;
assign addr[27684]= -1493966902;
assign addr[27685]= -1380375881;
assign addr[27686]= -1259782632;
assign addr[27687]= -1132798888;
assign addr[27688]= -1000068799;
assign addr[27689]= -862265664;
assign addr[27690]= -720088517;
assign addr[27691]= -574258580;
assign addr[27692]= -425515602;
assign addr[27693]= -274614114;
assign addr[27694]= -122319591;
assign addr[27695]= 30595422;
assign addr[27696]= 183355234;
assign addr[27697]= 335184940;
assign addr[27698]= 485314355;
assign addr[27699]= 632981917;
assign addr[27700]= 777438554;
assign addr[27701]= 917951481;
assign addr[27702]= 1053807919;
assign addr[27703]= 1184318708;
assign addr[27704]= 1308821808;
assign addr[27705]= 1426685652;
assign addr[27706]= 1537312353;
assign addr[27707]= 1640140734;
assign addr[27708]= 1734649179;
assign addr[27709]= 1820358275;
assign addr[27710]= 1896833245;
assign addr[27711]= 1963686155;
assign addr[27712]= 2020577882;
assign addr[27713]= 2067219829;
assign addr[27714]= 2103375398;
assign addr[27715]= 2128861181;
assign addr[27716]= 2143547897;
assign addr[27717]= 2147361045;
assign addr[27718]= 2140281282;
assign addr[27719]= 2122344521;
assign addr[27720]= 2093641749;
assign addr[27721]= 2054318569;
assign addr[27722]= 2004574453;
assign addr[27723]= 1944661739;
assign addr[27724]= 1874884346;
assign addr[27725]= 1795596234;
assign addr[27726]= 1707199606;
assign addr[27727]= 1610142873;
assign addr[27728]= 1504918373;
assign addr[27729]= 1392059879;
assign addr[27730]= 1272139887;
assign addr[27731]= 1145766716;
assign addr[27732]= 1013581418;
assign addr[27733]= 876254528;
assign addr[27734]= 734482665;
assign addr[27735]= 588984994;
assign addr[27736]= 440499581;
assign addr[27737]= 289779648;
assign addr[27738]= 137589750;
assign addr[27739]= -15298099;
assign addr[27740]= -168108346;
assign addr[27741]= -320065829;
assign addr[27742]= -470399716;
assign addr[27743]= -618347408;
assign addr[27744]= -763158411;
assign addr[27745]= -904098143;
assign addr[27746]= -1040451659;
assign addr[27747]= -1171527280;
assign addr[27748]= -1296660098;
assign addr[27749]= -1415215352;
assign addr[27750]= -1526591649;
assign addr[27751]= -1630224009;
assign addr[27752]= -1725586737;
assign addr[27753]= -1812196087;
assign addr[27754]= -1889612716;
assign addr[27755]= -1957443913;
assign addr[27756]= -2015345591;
assign addr[27757]= -2063024031;
assign addr[27758]= -2100237377;
assign addr[27759]= -2126796855;
assign addr[27760]= -2142567738;
assign addr[27761]= -2147470025;
assign addr[27762]= -2141478848;
assign addr[27763]= -2124624598;
assign addr[27764]= -2096992772;
assign addr[27765]= -2058723538;
assign addr[27766]= -2010011024;
assign addr[27767]= -1951102334;
assign addr[27768]= -1882296293;
assign addr[27769]= -1803941934;
assign addr[27770]= -1716436725;
assign addr[27771]= -1620224553;
assign addr[27772]= -1515793473;
assign addr[27773]= -1403673233;
assign addr[27774]= -1284432584;
assign addr[27775]= -1158676398;
assign addr[27776]= -1027042599;
assign addr[27777]= -890198924;
assign addr[27778]= -748839539;
assign addr[27779]= -603681519;
assign addr[27780]= -455461206;
assign addr[27781]= -304930476;
assign addr[27782]= -152852926;
assign addr[27783]= 0;
assign addr[27784]= 152852926;
assign addr[27785]= 304930476;
assign addr[27786]= 455461206;
assign addr[27787]= 603681519;
assign addr[27788]= 748839539;
assign addr[27789]= 890198924;
assign addr[27790]= 1027042599;
assign addr[27791]= 1158676398;
assign addr[27792]= 1284432584;
assign addr[27793]= 1403673233;
assign addr[27794]= 1515793473;
assign addr[27795]= 1620224553;
assign addr[27796]= 1716436725;
assign addr[27797]= 1803941934;
assign addr[27798]= 1882296293;
assign addr[27799]= 1951102334;
assign addr[27800]= 2010011024;
assign addr[27801]= 2058723538;
assign addr[27802]= 2096992772;
assign addr[27803]= 2124624598;
assign addr[27804]= 2141478848;
assign addr[27805]= 2147470025;
assign addr[27806]= 2142567738;
assign addr[27807]= 2126796855;
assign addr[27808]= 2100237377;
assign addr[27809]= 2063024031;
assign addr[27810]= 2015345591;
assign addr[27811]= 1957443913;
assign addr[27812]= 1889612716;
assign addr[27813]= 1812196087;
assign addr[27814]= 1725586737;
assign addr[27815]= 1630224009;
assign addr[27816]= 1526591649;
assign addr[27817]= 1415215352;
assign addr[27818]= 1296660098;
assign addr[27819]= 1171527280;
assign addr[27820]= 1040451659;
assign addr[27821]= 904098143;
assign addr[27822]= 763158411;
assign addr[27823]= 618347408;
assign addr[27824]= 470399716;
assign addr[27825]= 320065829;
assign addr[27826]= 168108346;
assign addr[27827]= 15298099;
assign addr[27828]= -137589750;
assign addr[27829]= -289779648;
assign addr[27830]= -440499581;
assign addr[27831]= -588984994;
assign addr[27832]= -734482665;
assign addr[27833]= -876254528;
assign addr[27834]= -1013581418;
assign addr[27835]= -1145766716;
assign addr[27836]= -1272139887;
assign addr[27837]= -1392059879;
assign addr[27838]= -1504918373;
assign addr[27839]= -1610142873;
assign addr[27840]= -1707199606;
assign addr[27841]= -1795596234;
assign addr[27842]= -1874884346;
assign addr[27843]= -1944661739;
assign addr[27844]= -2004574453;
assign addr[27845]= -2054318569;
assign addr[27846]= -2093641749;
assign addr[27847]= -2122344521;
assign addr[27848]= -2140281282;
assign addr[27849]= -2147361045;
assign addr[27850]= -2143547897;
assign addr[27851]= -2128861181;
assign addr[27852]= -2103375398;
assign addr[27853]= -2067219829;
assign addr[27854]= -2020577882;
assign addr[27855]= -1963686155;
assign addr[27856]= -1896833245;
assign addr[27857]= -1820358275;
assign addr[27858]= -1734649179;
assign addr[27859]= -1640140734;
assign addr[27860]= -1537312353;
assign addr[27861]= -1426685652;
assign addr[27862]= -1308821808;
assign addr[27863]= -1184318708;
assign addr[27864]= -1053807919;
assign addr[27865]= -917951481;
assign addr[27866]= -777438554;
assign addr[27867]= -632981917;
assign addr[27868]= -485314355;
assign addr[27869]= -335184940;
assign addr[27870]= -183355234;
assign addr[27871]= -30595422;
assign addr[27872]= 122319591;
assign addr[27873]= 274614114;
assign addr[27874]= 425515602;
assign addr[27875]= 574258580;
assign addr[27876]= 720088517;
assign addr[27877]= 862265664;
assign addr[27878]= 1000068799;
assign addr[27879]= 1132798888;
assign addr[27880]= 1259782632;
assign addr[27881]= 1380375881;
assign addr[27882]= 1493966902;
assign addr[27883]= 1599979481;
assign addr[27884]= 1697875851;
assign addr[27885]= 1787159411;
assign addr[27886]= 1867377253;
assign addr[27887]= 1938122457;
assign addr[27888]= 1999036154;
assign addr[27889]= 2049809346;
assign addr[27890]= 2090184478;
assign addr[27891]= 2119956737;
assign addr[27892]= 2138975100;
assign addr[27893]= 2147143090;
assign addr[27894]= 2144419275;
assign addr[27895]= 2130817471;
assign addr[27896]= 2106406677;
assign addr[27897]= 2071310720;
assign addr[27898]= 2025707632;
assign addr[27899]= 1969828744;
assign addr[27900]= 1903957513;
assign addr[27901]= 1828428082;
assign addr[27902]= 1743623590;
assign addr[27903]= 1649974225;
assign addr[27904]= 1547955041;
assign addr[27905]= 1438083551;
assign addr[27906]= 1320917099;
assign addr[27907]= 1197050035;
assign addr[27908]= 1067110699;
assign addr[27909]= 931758235;
assign addr[27910]= 791679244;
assign addr[27911]= 647584304;
assign addr[27912]= 500204365;
assign addr[27913]= 350287041;
assign addr[27914]= 198592817;
assign addr[27915]= 45891193;
assign addr[27916]= -107043224;
assign addr[27917]= -259434643;
assign addr[27918]= -410510029;
assign addr[27919]= -559503022;
assign addr[27920]= -705657826;
assign addr[27921]= -848233042;
assign addr[27922]= -986505429;
assign addr[27923]= -1119773573;
assign addr[27924]= -1247361445;
assign addr[27925]= -1368621831;
assign addr[27926]= -1482939614;
assign addr[27927]= -1589734894;
assign addr[27928]= -1688465931;
assign addr[27929]= -1778631892;
assign addr[27930]= -1859775393;
assign addr[27931]= -1931484818;
assign addr[27932]= -1993396407;
assign addr[27933]= -2045196100;
assign addr[27934]= -2086621133;
assign addr[27935]= -2117461370;
assign addr[27936]= -2137560369;
assign addr[27937]= -2146816171;
assign addr[27938]= -2145181827;
assign addr[27939]= -2132665626;
assign addr[27940]= -2109331059;
assign addr[27941]= -2075296495;
assign addr[27942]= -2030734582;
assign addr[27943]= -1975871368;
assign addr[27944]= -1910985158;
assign addr[27945]= -1836405100;
assign addr[27946]= -1752509516;
assign addr[27947]= -1659723983;
assign addr[27948]= -1558519173;
assign addr[27949]= -1449408469;
assign addr[27950]= -1332945355;
assign addr[27951]= -1209720613;
assign addr[27952]= -1080359326;
assign addr[27953]= -945517704;
assign addr[27954]= -805879757;
assign addr[27955]= -662153826;
assign addr[27956]= -515068990;
assign addr[27957]= -365371365;
assign addr[27958]= -213820322;
assign addr[27959]= -61184634;
assign addr[27960]= 91761426;
assign addr[27961]= 244242007;
assign addr[27962]= 395483624;
assign addr[27963]= 544719071;
assign addr[27964]= 691191324;
assign addr[27965]= 834157373;
assign addr[27966]= 972891995;
assign addr[27967]= 1106691431;
assign addr[27968]= 1234876957;
assign addr[27969]= 1356798326;
assign addr[27970]= 1471837070;
assign addr[27971]= 1579409630;
assign addr[27972]= 1678970324;
assign addr[27973]= 1770014111;
assign addr[27974]= 1852079154;
assign addr[27975]= 1924749160;
assign addr[27976]= 1987655498;
assign addr[27977]= 2040479063;
assign addr[27978]= 2082951896;
assign addr[27979]= 2114858546;
assign addr[27980]= 2136037160;
assign addr[27981]= 2146380306;
assign addr[27982]= 2145835515;
assign addr[27983]= 2134405552;
assign addr[27984]= 2112148396;
assign addr[27985]= 2079176953;
assign addr[27986]= 2035658475;
assign addr[27987]= 1981813720;
assign addr[27988]= 1917915825;
assign addr[27989]= 1844288924;
assign addr[27990]= 1761306505;
assign addr[27991]= 1669389513;
assign addr[27992]= 1569004214;
assign addr[27993]= 1460659832;
assign addr[27994]= 1344905966;
assign addr[27995]= 1222329801;
assign addr[27996]= 1093553126;
assign addr[27997]= 959229189;
assign addr[27998]= 820039373;
assign addr[27999]= 676689746;
assign addr[28000]= 529907477;
assign addr[28001]= 380437148;
assign addr[28002]= 229036977;
assign addr[28003]= 76474970;
assign addr[28004]= -76474970;
assign addr[28005]= -229036977;
assign addr[28006]= -380437148;
assign addr[28007]= -529907477;
assign addr[28008]= -676689746;
assign addr[28009]= -820039373;
assign addr[28010]= -959229189;
assign addr[28011]= -1093553126;
assign addr[28012]= -1222329801;
assign addr[28013]= -1344905966;
assign addr[28014]= -1460659832;
assign addr[28015]= -1569004214;
assign addr[28016]= -1669389513;
assign addr[28017]= -1761306505;
assign addr[28018]= -1844288924;
assign addr[28019]= -1917915825;
assign addr[28020]= -1981813720;
assign addr[28021]= -2035658475;
assign addr[28022]= -2079176953;
assign addr[28023]= -2112148396;
assign addr[28024]= -2134405552;
assign addr[28025]= -2145835515;
assign addr[28026]= -2146380306;
assign addr[28027]= -2136037160;
assign addr[28028]= -2114858546;
assign addr[28029]= -2082951896;
assign addr[28030]= -2040479063;
assign addr[28031]= -1987655498;
assign addr[28032]= -1924749160;
assign addr[28033]= -1852079154;
assign addr[28034]= -1770014111;
assign addr[28035]= -1678970324;
assign addr[28036]= -1579409630;
assign addr[28037]= -1471837070;
assign addr[28038]= -1356798326;
assign addr[28039]= -1234876957;
assign addr[28040]= -1106691431;
assign addr[28041]= -972891995;
assign addr[28042]= -834157373;
assign addr[28043]= -691191324;
assign addr[28044]= -544719071;
assign addr[28045]= -395483624;
assign addr[28046]= -244242007;
assign addr[28047]= -91761426;
assign addr[28048]= 61184634;
assign addr[28049]= 213820322;
assign addr[28050]= 365371365;
assign addr[28051]= 515068990;
assign addr[28052]= 662153826;
assign addr[28053]= 805879757;
assign addr[28054]= 945517704;
assign addr[28055]= 1080359326;
assign addr[28056]= 1209720613;
assign addr[28057]= 1332945355;
assign addr[28058]= 1449408469;
assign addr[28059]= 1558519173;
assign addr[28060]= 1659723983;
assign addr[28061]= 1752509516;
assign addr[28062]= 1836405100;
assign addr[28063]= 1910985158;
assign addr[28064]= 1975871368;
assign addr[28065]= 2030734582;
assign addr[28066]= 2075296495;
assign addr[28067]= 2109331059;
assign addr[28068]= 2132665626;
assign addr[28069]= 2145181827;
assign addr[28070]= 2146816171;
assign addr[28071]= 2137560369;
assign addr[28072]= 2117461370;
assign addr[28073]= 2086621133;
assign addr[28074]= 2045196100;
assign addr[28075]= 1993396407;
assign addr[28076]= 1931484818;
assign addr[28077]= 1859775393;
assign addr[28078]= 1778631892;
assign addr[28079]= 1688465931;
assign addr[28080]= 1589734894;
assign addr[28081]= 1482939614;
assign addr[28082]= 1368621831;
assign addr[28083]= 1247361445;
assign addr[28084]= 1119773573;
assign addr[28085]= 986505429;
assign addr[28086]= 848233042;
assign addr[28087]= 705657826;
assign addr[28088]= 559503022;
assign addr[28089]= 410510029;
assign addr[28090]= 259434643;
assign addr[28091]= 107043224;
assign addr[28092]= -45891193;
assign addr[28093]= -198592817;
assign addr[28094]= -350287041;
assign addr[28095]= -500204365;
assign addr[28096]= -647584304;
assign addr[28097]= -791679244;
assign addr[28098]= -931758235;
assign addr[28099]= -1067110699;
assign addr[28100]= -1197050035;
assign addr[28101]= -1320917099;
assign addr[28102]= -1438083551;
assign addr[28103]= -1547955041;
assign addr[28104]= -1649974225;
assign addr[28105]= -1743623590;
assign addr[28106]= -1828428082;
assign addr[28107]= -1903957513;
assign addr[28108]= -1969828744;
assign addr[28109]= -2025707632;
assign addr[28110]= -2071310720;
assign addr[28111]= -2106406677;
assign addr[28112]= -2130817471;
assign addr[28113]= -2144419275;
assign addr[28114]= -2147143090;
assign addr[28115]= -2138975100;
assign addr[28116]= -2119956737;
assign addr[28117]= -2090184478;
assign addr[28118]= -2049809346;
assign addr[28119]= -1999036154;
assign addr[28120]= -1938122457;
assign addr[28121]= -1867377253;
assign addr[28122]= -1787159411;
assign addr[28123]= -1697875851;
assign addr[28124]= -1599979481;
assign addr[28125]= -1493966902;
assign addr[28126]= -1380375881;
assign addr[28127]= -1259782632;
assign addr[28128]= -1132798888;
assign addr[28129]= -1000068799;
assign addr[28130]= -862265664;
assign addr[28131]= -720088517;
assign addr[28132]= -574258580;
assign addr[28133]= -425515602;
assign addr[28134]= -274614114;
assign addr[28135]= -122319591;
assign addr[28136]= 30595422;
assign addr[28137]= 183355234;
assign addr[28138]= 335184940;
assign addr[28139]= 485314355;
assign addr[28140]= 632981917;
assign addr[28141]= 777438554;
assign addr[28142]= 917951481;
assign addr[28143]= 1053807919;
assign addr[28144]= 1184318708;
assign addr[28145]= 1308821808;
assign addr[28146]= 1426685652;
assign addr[28147]= 1537312353;
assign addr[28148]= 1640140734;
assign addr[28149]= 1734649179;
assign addr[28150]= 1820358275;
assign addr[28151]= 1896833245;
assign addr[28152]= 1963686155;
assign addr[28153]= 2020577882;
assign addr[28154]= 2067219829;
assign addr[28155]= 2103375398;
assign addr[28156]= 2128861181;
assign addr[28157]= 2143547897;
assign addr[28158]= 2147361045;
assign addr[28159]= 2140281282;
assign addr[28160]= 2122344521;
assign addr[28161]= 2093641749;
assign addr[28162]= 2054318569;
assign addr[28163]= 2004574453;
assign addr[28164]= 1944661739;
assign addr[28165]= 1874884346;
assign addr[28166]= 1795596234;
assign addr[28167]= 1707199606;
assign addr[28168]= 1610142873;
assign addr[28169]= 1504918373;
assign addr[28170]= 1392059879;
assign addr[28171]= 1272139887;
assign addr[28172]= 1145766716;
assign addr[28173]= 1013581418;
assign addr[28174]= 876254528;
assign addr[28175]= 734482665;
assign addr[28176]= 588984994;
assign addr[28177]= 440499581;
assign addr[28178]= 289779648;
assign addr[28179]= 137589750;
assign addr[28180]= -15298099;
assign addr[28181]= -168108346;
assign addr[28182]= -320065829;
assign addr[28183]= -470399716;
assign addr[28184]= -618347408;
assign addr[28185]= -763158411;
assign addr[28186]= -904098143;
assign addr[28187]= -1040451659;
assign addr[28188]= -1171527280;
assign addr[28189]= -1296660098;
assign addr[28190]= -1415215352;
assign addr[28191]= -1526591649;
assign addr[28192]= -1630224009;
assign addr[28193]= -1725586737;
assign addr[28194]= -1812196087;
assign addr[28195]= -1889612716;
assign addr[28196]= -1957443913;
assign addr[28197]= -2015345591;
assign addr[28198]= -2063024031;
assign addr[28199]= -2100237377;
assign addr[28200]= -2126796855;
assign addr[28201]= -2142567738;
assign addr[28202]= -2147470025;
assign addr[28203]= -2141478848;
assign addr[28204]= -2124624598;
assign addr[28205]= -2096992772;
assign addr[28206]= -2058723538;
assign addr[28207]= -2010011024;
assign addr[28208]= -1951102334;
assign addr[28209]= -1882296293;
assign addr[28210]= -1803941934;
assign addr[28211]= -1716436725;
assign addr[28212]= -1620224553;
assign addr[28213]= -1515793473;
assign addr[28214]= -1403673233;
assign addr[28215]= -1284432584;
assign addr[28216]= -1158676398;
assign addr[28217]= -1027042599;
assign addr[28218]= -890198924;
assign addr[28219]= -748839539;
assign addr[28220]= -603681519;
assign addr[28221]= -455461206;
assign addr[28222]= -304930476;
assign addr[28223]= -152852926;
assign addr[28224]= 0;
assign addr[28225]= 152852926;
assign addr[28226]= 304930476;
assign addr[28227]= 455461206;
assign addr[28228]= 603681519;
assign addr[28229]= 748839539;
assign addr[28230]= 890198924;
assign addr[28231]= 1027042599;
assign addr[28232]= 1158676398;
assign addr[28233]= 1284432584;
assign addr[28234]= 1403673233;
assign addr[28235]= 1515793473;
assign addr[28236]= 1620224553;
assign addr[28237]= 1716436725;
assign addr[28238]= 1803941934;
assign addr[28239]= 1882296293;
assign addr[28240]= 1951102334;
assign addr[28241]= 2010011024;
assign addr[28242]= 2058723538;
assign addr[28243]= 2096992772;
assign addr[28244]= 2124624598;
assign addr[28245]= 2141478848;
assign addr[28246]= 2147470025;
assign addr[28247]= 2142567738;
assign addr[28248]= 2126796855;
assign addr[28249]= 2100237377;
assign addr[28250]= 2063024031;
assign addr[28251]= 2015345591;
assign addr[28252]= 1957443913;
assign addr[28253]= 1889612716;
assign addr[28254]= 1812196087;
assign addr[28255]= 1725586737;
assign addr[28256]= 1630224009;
assign addr[28257]= 1526591649;
assign addr[28258]= 1415215352;
assign addr[28259]= 1296660098;
assign addr[28260]= 1171527280;
assign addr[28261]= 1040451659;
assign addr[28262]= 904098143;
assign addr[28263]= 763158411;
assign addr[28264]= 618347408;
assign addr[28265]= 470399716;
assign addr[28266]= 320065829;
assign addr[28267]= 168108346;
assign addr[28268]= 15298099;
assign addr[28269]= -137589750;
assign addr[28270]= -289779648;
assign addr[28271]= -440499581;
assign addr[28272]= -588984994;
assign addr[28273]= -734482665;
assign addr[28274]= -876254528;
assign addr[28275]= -1013581418;
assign addr[28276]= -1145766716;
assign addr[28277]= -1272139887;
assign addr[28278]= -1392059879;
assign addr[28279]= -1504918373;
assign addr[28280]= -1610142873;
assign addr[28281]= -1707199606;
assign addr[28282]= -1795596234;
assign addr[28283]= -1874884346;
assign addr[28284]= -1944661739;
assign addr[28285]= -2004574453;
assign addr[28286]= -2054318569;
assign addr[28287]= -2093641749;
assign addr[28288]= -2122344521;
assign addr[28289]= -2140281282;
assign addr[28290]= -2147361045;
assign addr[28291]= -2143547897;
assign addr[28292]= -2128861181;
assign addr[28293]= -2103375398;
assign addr[28294]= -2067219829;
assign addr[28295]= -2020577882;
assign addr[28296]= -1963686155;
assign addr[28297]= -1896833245;
assign addr[28298]= -1820358275;
assign addr[28299]= -1734649179;
assign addr[28300]= -1640140734;
assign addr[28301]= -1537312353;
assign addr[28302]= -1426685652;
assign addr[28303]= -1308821808;
assign addr[28304]= -1184318708;
assign addr[28305]= -1053807919;
assign addr[28306]= -917951481;
assign addr[28307]= -777438554;
assign addr[28308]= -632981917;
assign addr[28309]= -485314355;
assign addr[28310]= -335184940;
assign addr[28311]= -183355234;
assign addr[28312]= -30595422;
assign addr[28313]= 122319591;
assign addr[28314]= 274614114;
assign addr[28315]= 425515602;
assign addr[28316]= 574258580;
assign addr[28317]= 720088517;
assign addr[28318]= 862265664;
assign addr[28319]= 1000068799;
assign addr[28320]= 1132798888;
assign addr[28321]= 1259782632;
assign addr[28322]= 1380375881;
assign addr[28323]= 1493966902;
assign addr[28324]= 1599979481;
assign addr[28325]= 1697875851;
assign addr[28326]= 1787159411;
assign addr[28327]= 1867377253;
assign addr[28328]= 1938122457;
assign addr[28329]= 1999036154;
assign addr[28330]= 2049809346;
assign addr[28331]= 2090184478;
assign addr[28332]= 2119956737;
assign addr[28333]= 2138975100;
assign addr[28334]= 2147143090;
assign addr[28335]= 2144419275;
assign addr[28336]= 2130817471;
assign addr[28337]= 2106406677;
assign addr[28338]= 2071310720;
assign addr[28339]= 2025707632;
assign addr[28340]= 1969828744;
assign addr[28341]= 1903957513;
assign addr[28342]= 1828428082;
assign addr[28343]= 1743623590;
assign addr[28344]= 1649974225;
assign addr[28345]= 1547955041;
assign addr[28346]= 1438083551;
assign addr[28347]= 1320917099;
assign addr[28348]= 1197050035;
assign addr[28349]= 1067110699;
assign addr[28350]= 931758235;
assign addr[28351]= 791679244;
assign addr[28352]= 647584304;
assign addr[28353]= 500204365;
assign addr[28354]= 350287041;
assign addr[28355]= 198592817;
assign addr[28356]= 45891193;
assign addr[28357]= -107043224;
assign addr[28358]= -259434643;
assign addr[28359]= -410510029;
assign addr[28360]= -559503022;
assign addr[28361]= -705657826;
assign addr[28362]= -848233042;
assign addr[28363]= -986505429;
assign addr[28364]= -1119773573;
assign addr[28365]= -1247361445;
assign addr[28366]= -1368621831;
assign addr[28367]= -1482939614;
assign addr[28368]= -1589734894;
assign addr[28369]= -1688465931;
assign addr[28370]= -1778631892;
assign addr[28371]= -1859775393;
assign addr[28372]= -1931484818;
assign addr[28373]= -1993396407;
assign addr[28374]= -2045196100;
assign addr[28375]= -2086621133;
assign addr[28376]= -2117461370;
assign addr[28377]= -2137560369;
assign addr[28378]= -2146816171;
assign addr[28379]= -2145181827;
assign addr[28380]= -2132665626;
assign addr[28381]= -2109331059;
assign addr[28382]= -2075296495;
assign addr[28383]= -2030734582;
assign addr[28384]= -1975871368;
assign addr[28385]= -1910985158;
assign addr[28386]= -1836405100;
assign addr[28387]= -1752509516;
assign addr[28388]= -1659723983;
assign addr[28389]= -1558519173;
assign addr[28390]= -1449408469;
assign addr[28391]= -1332945355;
assign addr[28392]= -1209720613;
assign addr[28393]= -1080359326;
assign addr[28394]= -945517704;
assign addr[28395]= -805879757;
assign addr[28396]= -662153826;
assign addr[28397]= -515068990;
assign addr[28398]= -365371365;
assign addr[28399]= -213820322;
assign addr[28400]= -61184634;
assign addr[28401]= 91761426;
assign addr[28402]= 244242007;
assign addr[28403]= 395483624;
assign addr[28404]= 544719071;
assign addr[28405]= 691191324;
assign addr[28406]= 834157373;
assign addr[28407]= 972891995;
assign addr[28408]= 1106691431;
assign addr[28409]= 1234876957;
assign addr[28410]= 1356798326;
assign addr[28411]= 1471837070;
assign addr[28412]= 1579409630;
assign addr[28413]= 1678970324;
assign addr[28414]= 1770014111;
assign addr[28415]= 1852079154;
assign addr[28416]= 1924749160;
assign addr[28417]= 1987655498;
assign addr[28418]= 2040479063;
assign addr[28419]= 2082951896;
assign addr[28420]= 2114858546;
assign addr[28421]= 2136037160;
assign addr[28422]= 2146380306;
assign addr[28423]= 2145835515;
assign addr[28424]= 2134405552;
assign addr[28425]= 2112148396;
assign addr[28426]= 2079176953;
assign addr[28427]= 2035658475;
assign addr[28428]= 1981813720;
assign addr[28429]= 1917915825;
assign addr[28430]= 1844288924;
assign addr[28431]= 1761306505;
assign addr[28432]= 1669389513;
assign addr[28433]= 1569004214;
assign addr[28434]= 1460659832;
assign addr[28435]= 1344905966;
assign addr[28436]= 1222329801;
assign addr[28437]= 1093553126;
assign addr[28438]= 959229189;
assign addr[28439]= 820039373;
assign addr[28440]= 676689746;
assign addr[28441]= 529907477;
assign addr[28442]= 380437148;
assign addr[28443]= 229036977;
assign addr[28444]= 76474970;
assign addr[28445]= -76474970;
assign addr[28446]= -229036977;
assign addr[28447]= -380437148;
assign addr[28448]= -529907477;
assign addr[28449]= -676689746;
assign addr[28450]= -820039373;
assign addr[28451]= -959229189;
assign addr[28452]= -1093553126;
assign addr[28453]= -1222329801;
assign addr[28454]= -1344905966;
assign addr[28455]= -1460659832;
assign addr[28456]= -1569004214;
assign addr[28457]= -1669389513;
assign addr[28458]= -1761306505;
assign addr[28459]= -1844288924;
assign addr[28460]= -1917915825;
assign addr[28461]= -1981813720;
assign addr[28462]= -2035658475;
assign addr[28463]= -2079176953;
assign addr[28464]= -2112148396;
assign addr[28465]= -2134405552;
assign addr[28466]= -2145835515;
assign addr[28467]= -2146380306;
assign addr[28468]= -2136037160;
assign addr[28469]= -2114858546;
assign addr[28470]= -2082951896;
assign addr[28471]= -2040479063;
assign addr[28472]= -1987655498;
assign addr[28473]= -1924749160;
assign addr[28474]= -1852079154;
assign addr[28475]= -1770014111;
assign addr[28476]= -1678970324;
assign addr[28477]= -1579409630;
assign addr[28478]= -1471837070;
assign addr[28479]= -1356798326;
assign addr[28480]= -1234876957;
assign addr[28481]= -1106691431;
assign addr[28482]= -972891995;
assign addr[28483]= -834157373;
assign addr[28484]= -691191324;
assign addr[28485]= -544719071;
assign addr[28486]= -395483624;
assign addr[28487]= -244242007;
assign addr[28488]= -91761426;
assign addr[28489]= 61184634;
assign addr[28490]= 213820322;
assign addr[28491]= 365371365;
assign addr[28492]= 515068990;
assign addr[28493]= 662153826;
assign addr[28494]= 805879757;
assign addr[28495]= 945517704;
assign addr[28496]= 1080359326;
assign addr[28497]= 1209720613;
assign addr[28498]= 1332945355;
assign addr[28499]= 1449408469;
assign addr[28500]= 1558519173;
assign addr[28501]= 1659723983;
assign addr[28502]= 1752509516;
assign addr[28503]= 1836405100;
assign addr[28504]= 1910985158;
assign addr[28505]= 1975871368;
assign addr[28506]= 2030734582;
assign addr[28507]= 2075296495;
assign addr[28508]= 2109331059;
assign addr[28509]= 2132665626;
assign addr[28510]= 2145181827;
assign addr[28511]= 2146816171;
assign addr[28512]= 2137560369;
assign addr[28513]= 2117461370;
assign addr[28514]= 2086621133;
assign addr[28515]= 2045196100;
assign addr[28516]= 1993396407;
assign addr[28517]= 1931484818;
assign addr[28518]= 1859775393;
assign addr[28519]= 1778631892;
assign addr[28520]= 1688465931;
assign addr[28521]= 1589734894;
assign addr[28522]= 1482939614;
assign addr[28523]= 1368621831;
assign addr[28524]= 1247361445;
assign addr[28525]= 1119773573;
assign addr[28526]= 986505429;
assign addr[28527]= 848233042;
assign addr[28528]= 705657826;
assign addr[28529]= 559503022;
assign addr[28530]= 410510029;
assign addr[28531]= 259434643;
assign addr[28532]= 107043224;
assign addr[28533]= -45891193;
assign addr[28534]= -198592817;
assign addr[28535]= -350287041;
assign addr[28536]= -500204365;
assign addr[28537]= -647584304;
assign addr[28538]= -791679244;
assign addr[28539]= -931758235;
assign addr[28540]= -1067110699;
assign addr[28541]= -1197050035;
assign addr[28542]= -1320917099;
assign addr[28543]= -1438083551;
assign addr[28544]= -1547955041;
assign addr[28545]= -1649974225;
assign addr[28546]= -1743623590;
assign addr[28547]= -1828428082;
assign addr[28548]= -1903957513;
assign addr[28549]= -1969828744;
assign addr[28550]= -2025707632;
assign addr[28551]= -2071310720;
assign addr[28552]= -2106406677;
assign addr[28553]= -2130817471;
assign addr[28554]= -2144419275;
assign addr[28555]= -2147143090;
assign addr[28556]= -2138975100;
assign addr[28557]= -2119956737;
assign addr[28558]= -2090184478;
assign addr[28559]= -2049809346;
assign addr[28560]= -1999036154;
assign addr[28561]= -1938122457;
assign addr[28562]= -1867377253;
assign addr[28563]= -1787159411;
assign addr[28564]= -1697875851;
assign addr[28565]= -1599979481;
assign addr[28566]= -1493966902;
assign addr[28567]= -1380375881;
assign addr[28568]= -1259782632;
assign addr[28569]= -1132798888;
assign addr[28570]= -1000068799;
assign addr[28571]= -862265664;
assign addr[28572]= -720088517;
assign addr[28573]= -574258580;
assign addr[28574]= -425515602;
assign addr[28575]= -274614114;
assign addr[28576]= -122319591;
assign addr[28577]= 30595422;
assign addr[28578]= 183355234;
assign addr[28579]= 335184940;
assign addr[28580]= 485314355;
assign addr[28581]= 632981917;
assign addr[28582]= 777438554;
assign addr[28583]= 917951481;
assign addr[28584]= 1053807919;
assign addr[28585]= 1184318708;
assign addr[28586]= 1308821808;
assign addr[28587]= 1426685652;
assign addr[28588]= 1537312353;
assign addr[28589]= 1640140734;
assign addr[28590]= 1734649179;
assign addr[28591]= 1820358275;
assign addr[28592]= 1896833245;
assign addr[28593]= 1963686155;
assign addr[28594]= 2020577882;
assign addr[28595]= 2067219829;
assign addr[28596]= 2103375398;
assign addr[28597]= 2128861181;
assign addr[28598]= 2143547897;
assign addr[28599]= 2147361045;
assign addr[28600]= 2140281282;
assign addr[28601]= 2122344521;
assign addr[28602]= 2093641749;
assign addr[28603]= 2054318569;
assign addr[28604]= 2004574453;
assign addr[28605]= 1944661739;
assign addr[28606]= 1874884346;
assign addr[28607]= 1795596234;
assign addr[28608]= 1707199606;
assign addr[28609]= 1610142873;
assign addr[28610]= 1504918373;
assign addr[28611]= 1392059879;
assign addr[28612]= 1272139887;
assign addr[28613]= 1145766716;
assign addr[28614]= 1013581418;
assign addr[28615]= 876254528;
assign addr[28616]= 734482665;
assign addr[28617]= 588984994;
assign addr[28618]= 440499581;
assign addr[28619]= 289779648;
assign addr[28620]= 137589750;
assign addr[28621]= -15298099;
assign addr[28622]= -168108346;
assign addr[28623]= -320065829;
assign addr[28624]= -470399716;
assign addr[28625]= -618347408;
assign addr[28626]= -763158411;
assign addr[28627]= -904098143;
assign addr[28628]= -1040451659;
assign addr[28629]= -1171527280;
assign addr[28630]= -1296660098;
assign addr[28631]= -1415215352;
assign addr[28632]= -1526591649;
assign addr[28633]= -1630224009;
assign addr[28634]= -1725586737;
assign addr[28635]= -1812196087;
assign addr[28636]= -1889612716;
assign addr[28637]= -1957443913;
assign addr[28638]= -2015345591;
assign addr[28639]= -2063024031;
assign addr[28640]= -2100237377;
assign addr[28641]= -2126796855;
assign addr[28642]= -2142567738;
assign addr[28643]= -2147470025;
assign addr[28644]= -2141478848;
assign addr[28645]= -2124624598;
assign addr[28646]= -2096992772;
assign addr[28647]= -2058723538;
assign addr[28648]= -2010011024;
assign addr[28649]= -1951102334;
assign addr[28650]= -1882296293;
assign addr[28651]= -1803941934;
assign addr[28652]= -1716436725;
assign addr[28653]= -1620224553;
assign addr[28654]= -1515793473;
assign addr[28655]= -1403673233;
assign addr[28656]= -1284432584;
assign addr[28657]= -1158676398;
assign addr[28658]= -1027042599;
assign addr[28659]= -890198924;
assign addr[28660]= -748839539;
assign addr[28661]= -603681519;
assign addr[28662]= -455461206;
assign addr[28663]= -304930476;
assign addr[28664]= -152852926;
assign addr[28665]= 0;
assign addr[28666]= 152852926;
assign addr[28667]= 304930476;
assign addr[28668]= 455461206;
assign addr[28669]= 603681519;
assign addr[28670]= 748839539;
assign addr[28671]= 890198924;
assign addr[28672]= 1027042599;
assign addr[28673]= 1158676398;
assign addr[28674]= 1284432584;
assign addr[28675]= 1403673233;
assign addr[28676]= 1515793473;
assign addr[28677]= 1620224553;
assign addr[28678]= 1716436725;
assign addr[28679]= 1803941934;
assign addr[28680]= 1882296293;
assign addr[28681]= 1951102334;
assign addr[28682]= 2010011024;
assign addr[28683]= 2058723538;
assign addr[28684]= 2096992772;
assign addr[28685]= 2124624598;
assign addr[28686]= 2141478848;
assign addr[28687]= 2147470025;
assign addr[28688]= 2142567738;
assign addr[28689]= 2126796855;
assign addr[28690]= 2100237377;
assign addr[28691]= 2063024031;
assign addr[28692]= 2015345591;
assign addr[28693]= 1957443913;
assign addr[28694]= 1889612716;
assign addr[28695]= 1812196087;
assign addr[28696]= 1725586737;
assign addr[28697]= 1630224009;
assign addr[28698]= 1526591649;
assign addr[28699]= 1415215352;
assign addr[28700]= 1296660098;
assign addr[28701]= 1171527280;
assign addr[28702]= 1040451659;
assign addr[28703]= 904098143;
assign addr[28704]= 763158411;
assign addr[28705]= 618347408;
assign addr[28706]= 470399716;
assign addr[28707]= 320065829;
assign addr[28708]= 168108346;
assign addr[28709]= 15298099;
assign addr[28710]= -137589750;
assign addr[28711]= -289779648;
assign addr[28712]= -440499581;
assign addr[28713]= -588984994;
assign addr[28714]= -734482665;
assign addr[28715]= -876254528;
assign addr[28716]= -1013581418;
assign addr[28717]= -1145766716;
assign addr[28718]= -1272139887;
assign addr[28719]= -1392059879;
assign addr[28720]= -1504918373;
assign addr[28721]= -1610142873;
assign addr[28722]= -1707199606;
assign addr[28723]= -1795596234;
assign addr[28724]= -1874884346;
assign addr[28725]= -1944661739;
assign addr[28726]= -2004574453;
assign addr[28727]= -2054318569;
assign addr[28728]= -2093641749;
assign addr[28729]= -2122344521;
assign addr[28730]= -2140281282;
assign addr[28731]= -2147361045;
assign addr[28732]= -2143547897;
assign addr[28733]= -2128861181;
assign addr[28734]= -2103375398;
assign addr[28735]= -2067219829;
assign addr[28736]= -2020577882;
assign addr[28737]= -1963686155;
assign addr[28738]= -1896833245;
assign addr[28739]= -1820358275;
assign addr[28740]= -1734649179;
assign addr[28741]= -1640140734;
assign addr[28742]= -1537312353;
assign addr[28743]= -1426685652;
assign addr[28744]= -1308821808;
assign addr[28745]= -1184318708;
assign addr[28746]= -1053807919;
assign addr[28747]= -917951481;
assign addr[28748]= -777438554;
assign addr[28749]= -632981917;
assign addr[28750]= -485314355;
assign addr[28751]= -335184940;
assign addr[28752]= -183355234;
assign addr[28753]= -30595422;
assign addr[28754]= 122319591;
assign addr[28755]= 274614114;
assign addr[28756]= 425515602;
assign addr[28757]= 574258580;
assign addr[28758]= 720088517;
assign addr[28759]= 862265664;
assign addr[28760]= 1000068799;
assign addr[28761]= 1132798888;
assign addr[28762]= 1259782632;
assign addr[28763]= 1380375881;
assign addr[28764]= 1493966902;
assign addr[28765]= 1599979481;
assign addr[28766]= 1697875851;
assign addr[28767]= 1787159411;
assign addr[28768]= 1867377253;
assign addr[28769]= 1938122457;
assign addr[28770]= 1999036154;
assign addr[28771]= 2049809346;
assign addr[28772]= 2090184478;
assign addr[28773]= 2119956737;
assign addr[28774]= 2138975100;
assign addr[28775]= 2147143090;
assign addr[28776]= 2144419275;
assign addr[28777]= 2130817471;
assign addr[28778]= 2106406677;
assign addr[28779]= 2071310720;
assign addr[28780]= 2025707632;
assign addr[28781]= 1969828744;
assign addr[28782]= 1903957513;
assign addr[28783]= 1828428082;
assign addr[28784]= 1743623590;
assign addr[28785]= 1649974225;
assign addr[28786]= 1547955041;
assign addr[28787]= 1438083551;
assign addr[28788]= 1320917099;
assign addr[28789]= 1197050035;
assign addr[28790]= 1067110699;
assign addr[28791]= 931758235;
assign addr[28792]= 791679244;
assign addr[28793]= 647584304;
assign addr[28794]= 500204365;
assign addr[28795]= 350287041;
assign addr[28796]= 198592817;
assign addr[28797]= 45891193;
assign addr[28798]= -107043224;
assign addr[28799]= -259434643;
assign addr[28800]= -410510029;
assign addr[28801]= -559503022;
assign addr[28802]= -705657826;
assign addr[28803]= -848233042;
assign addr[28804]= -986505429;
assign addr[28805]= -1119773573;
assign addr[28806]= -1247361445;
assign addr[28807]= -1368621831;
assign addr[28808]= -1482939614;
assign addr[28809]= -1589734894;
assign addr[28810]= -1688465931;
assign addr[28811]= -1778631892;
assign addr[28812]= -1859775393;
assign addr[28813]= -1931484818;
assign addr[28814]= -1993396407;
assign addr[28815]= -2045196100;
assign addr[28816]= -2086621133;
assign addr[28817]= -2117461370;
assign addr[28818]= -2137560369;
assign addr[28819]= -2146816171;
assign addr[28820]= -2145181827;
assign addr[28821]= -2132665626;
assign addr[28822]= -2109331059;
assign addr[28823]= -2075296495;
assign addr[28824]= -2030734582;
assign addr[28825]= -1975871368;
assign addr[28826]= -1910985158;
assign addr[28827]= -1836405100;
assign addr[28828]= -1752509516;
assign addr[28829]= -1659723983;
assign addr[28830]= -1558519173;
assign addr[28831]= -1449408469;
assign addr[28832]= -1332945355;
assign addr[28833]= -1209720613;
assign addr[28834]= -1080359326;
assign addr[28835]= -945517704;
assign addr[28836]= -805879757;
assign addr[28837]= -662153826;
assign addr[28838]= -515068990;
assign addr[28839]= -365371365;
assign addr[28840]= -213820322;
assign addr[28841]= -61184634;
assign addr[28842]= 91761426;
assign addr[28843]= 244242007;
assign addr[28844]= 395483624;
assign addr[28845]= 544719071;
assign addr[28846]= 691191324;
assign addr[28847]= 834157373;
assign addr[28848]= 972891995;
assign addr[28849]= 1106691431;
assign addr[28850]= 1234876957;
assign addr[28851]= 1356798326;
assign addr[28852]= 1471837070;
assign addr[28853]= 1579409630;
assign addr[28854]= 1678970324;
assign addr[28855]= 1770014111;
assign addr[28856]= 1852079154;
assign addr[28857]= 1924749160;
assign addr[28858]= 1987655498;
assign addr[28859]= 2040479063;
assign addr[28860]= 2082951896;
assign addr[28861]= 2114858546;
assign addr[28862]= 2136037160;
assign addr[28863]= 2146380306;
assign addr[28864]= 2145835515;
assign addr[28865]= 2134405552;
assign addr[28866]= 2112148396;
assign addr[28867]= 2079176953;
assign addr[28868]= 2035658475;
assign addr[28869]= 1981813720;
assign addr[28870]= 1917915825;
assign addr[28871]= 1844288924;
assign addr[28872]= 1761306505;
assign addr[28873]= 1669389513;
assign addr[28874]= 1569004214;
assign addr[28875]= 1460659832;
assign addr[28876]= 1344905966;
assign addr[28877]= 1222329801;
assign addr[28878]= 1093553126;
assign addr[28879]= 959229189;
assign addr[28880]= 820039373;
assign addr[28881]= 676689746;
assign addr[28882]= 529907477;
assign addr[28883]= 380437148;
assign addr[28884]= 229036977;
assign addr[28885]= 76474970;
assign addr[28886]= -76474970;
assign addr[28887]= -229036977;
assign addr[28888]= -380437148;
assign addr[28889]= -529907477;
assign addr[28890]= -676689746;
assign addr[28891]= -820039373;
assign addr[28892]= -959229189;
assign addr[28893]= -1093553126;
assign addr[28894]= -1222329801;
assign addr[28895]= -1344905966;
assign addr[28896]= -1460659832;
assign addr[28897]= -1569004214;
assign addr[28898]= -1669389513;
assign addr[28899]= -1761306505;
assign addr[28900]= -1844288924;
assign addr[28901]= -1917915825;
assign addr[28902]= -1981813720;
assign addr[28903]= -2035658475;
assign addr[28904]= -2079176953;
assign addr[28905]= -2112148396;
assign addr[28906]= -2134405552;
assign addr[28907]= -2145835515;
assign addr[28908]= -2146380306;
assign addr[28909]= -2136037160;
assign addr[28910]= -2114858546;
assign addr[28911]= -2082951896;
assign addr[28912]= -2040479063;
assign addr[28913]= -1987655498;
assign addr[28914]= -1924749160;
assign addr[28915]= -1852079154;
assign addr[28916]= -1770014111;
assign addr[28917]= -1678970324;
assign addr[28918]= -1579409630;
assign addr[28919]= -1471837070;
assign addr[28920]= -1356798326;
assign addr[28921]= -1234876957;
assign addr[28922]= -1106691431;
assign addr[28923]= -972891995;
assign addr[28924]= -834157373;
assign addr[28925]= -691191324;
assign addr[28926]= -544719071;
assign addr[28927]= -395483624;
assign addr[28928]= -244242007;
assign addr[28929]= -91761426;
assign addr[28930]= 61184634;
assign addr[28931]= 213820322;
assign addr[28932]= 365371365;
assign addr[28933]= 515068990;
assign addr[28934]= 662153826;
assign addr[28935]= 805879757;
assign addr[28936]= 945517704;
assign addr[28937]= 1080359326;
assign addr[28938]= 1209720613;
assign addr[28939]= 1332945355;
assign addr[28940]= 1449408469;
assign addr[28941]= 1558519173;
assign addr[28942]= 1659723983;
assign addr[28943]= 1752509516;
assign addr[28944]= 1836405100;
assign addr[28945]= 1910985158;
assign addr[28946]= 1975871368;
assign addr[28947]= 2030734582;
assign addr[28948]= 2075296495;
assign addr[28949]= 2109331059;
assign addr[28950]= 2132665626;
assign addr[28951]= 2145181827;
assign addr[28952]= 2146816171;
assign addr[28953]= 2137560369;
assign addr[28954]= 2117461370;
assign addr[28955]= 2086621133;
assign addr[28956]= 2045196100;
assign addr[28957]= 1993396407;
assign addr[28958]= 1931484818;
assign addr[28959]= 1859775393;
assign addr[28960]= 1778631892;
assign addr[28961]= 1688465931;
assign addr[28962]= 1589734894;
assign addr[28963]= 1482939614;
assign addr[28964]= 1368621831;
assign addr[28965]= 1247361445;
assign addr[28966]= 1119773573;
assign addr[28967]= 986505429;
assign addr[28968]= 848233042;
assign addr[28969]= 705657826;
assign addr[28970]= 559503022;
assign addr[28971]= 410510029;
assign addr[28972]= 259434643;
assign addr[28973]= 107043224;
assign addr[28974]= -45891193;
assign addr[28975]= -198592817;
assign addr[28976]= -350287041;
assign addr[28977]= -500204365;
assign addr[28978]= -647584304;
assign addr[28979]= -791679244;
assign addr[28980]= -931758235;
assign addr[28981]= -1067110699;
assign addr[28982]= -1197050035;
assign addr[28983]= -1320917099;
assign addr[28984]= -1438083551;
assign addr[28985]= -1547955041;
assign addr[28986]= -1649974225;
assign addr[28987]= -1743623590;
assign addr[28988]= -1828428082;
assign addr[28989]= -1903957513;
assign addr[28990]= -1969828744;
assign addr[28991]= -2025707632;
assign addr[28992]= -2071310720;
assign addr[28993]= -2106406677;
assign addr[28994]= -2130817471;
assign addr[28995]= -2144419275;
assign addr[28996]= -2147143090;
assign addr[28997]= -2138975100;
assign addr[28998]= -2119956737;
assign addr[28999]= -2090184478;
assign addr[29000]= -2049809346;
assign addr[29001]= -1999036154;
assign addr[29002]= -1938122457;
assign addr[29003]= -1867377253;
assign addr[29004]= -1787159411;
assign addr[29005]= -1697875851;
assign addr[29006]= -1599979481;
assign addr[29007]= -1493966902;
assign addr[29008]= -1380375881;
assign addr[29009]= -1259782632;
assign addr[29010]= -1132798888;
assign addr[29011]= -1000068799;
assign addr[29012]= -862265664;
assign addr[29013]= -720088517;
assign addr[29014]= -574258580;
assign addr[29015]= -425515602;
assign addr[29016]= -274614114;
assign addr[29017]= -122319591;
assign addr[29018]= 30595422;
assign addr[29019]= 183355234;
assign addr[29020]= 335184940;
assign addr[29021]= 485314355;
assign addr[29022]= 632981917;
assign addr[29023]= 777438554;
assign addr[29024]= 917951481;
assign addr[29025]= 1053807919;
assign addr[29026]= 1184318708;
assign addr[29027]= 1308821808;
assign addr[29028]= 1426685652;
assign addr[29029]= 1537312353;
assign addr[29030]= 1640140734;
assign addr[29031]= 1734649179;
assign addr[29032]= 1820358275;
assign addr[29033]= 1896833245;
assign addr[29034]= 1963686155;
assign addr[29035]= 2020577882;
assign addr[29036]= 2067219829;
assign addr[29037]= 2103375398;
assign addr[29038]= 2128861181;
assign addr[29039]= 2143547897;
assign addr[29040]= 2147361045;
assign addr[29041]= 2140281282;
assign addr[29042]= 2122344521;
assign addr[29043]= 2093641749;
assign addr[29044]= 2054318569;
assign addr[29045]= 2004574453;
assign addr[29046]= 1944661739;
assign addr[29047]= 1874884346;
assign addr[29048]= 1795596234;
assign addr[29049]= 1707199606;
assign addr[29050]= 1610142873;
assign addr[29051]= 1504918373;
assign addr[29052]= 1392059879;
assign addr[29053]= 1272139887;
assign addr[29054]= 1145766716;
assign addr[29055]= 1013581418;
assign addr[29056]= 876254528;
assign addr[29057]= 734482665;
assign addr[29058]= 588984994;
assign addr[29059]= 440499581;
assign addr[29060]= 289779648;
assign addr[29061]= 137589750;
assign addr[29062]= -15298099;
assign addr[29063]= -168108346;
assign addr[29064]= -320065829;
assign addr[29065]= -470399716;
assign addr[29066]= -618347408;
assign addr[29067]= -763158411;
assign addr[29068]= -904098143;
assign addr[29069]= -1040451659;
assign addr[29070]= -1171527280;
assign addr[29071]= -1296660098;
assign addr[29072]= -1415215352;
assign addr[29073]= -1526591649;
assign addr[29074]= -1630224009;
assign addr[29075]= -1725586737;
assign addr[29076]= -1812196087;
assign addr[29077]= -1889612716;
assign addr[29078]= -1957443913;
assign addr[29079]= -2015345591;
assign addr[29080]= -2063024031;
assign addr[29081]= -2100237377;
assign addr[29082]= -2126796855;
assign addr[29083]= -2142567738;
assign addr[29084]= -2147470025;
assign addr[29085]= -2141478848;
assign addr[29086]= -2124624598;
assign addr[29087]= -2096992772;
assign addr[29088]= -2058723538;
assign addr[29089]= -2010011024;
assign addr[29090]= -1951102334;
assign addr[29091]= -1882296293;
assign addr[29092]= -1803941934;
assign addr[29093]= -1716436725;
assign addr[29094]= -1620224553;
assign addr[29095]= -1515793473;
assign addr[29096]= -1403673233;
assign addr[29097]= -1284432584;
assign addr[29098]= -1158676398;
assign addr[29099]= -1027042599;
assign addr[29100]= -890198924;
assign addr[29101]= -748839539;
assign addr[29102]= -603681519;
assign addr[29103]= -455461206;
assign addr[29104]= -304930476;
assign addr[29105]= -152852926;
assign addr[29106]= 0;
assign addr[29107]= 152852926;
assign addr[29108]= 304930476;
assign addr[29109]= 455461206;
assign addr[29110]= 603681519;
assign addr[29111]= 748839539;
assign addr[29112]= 890198924;
assign addr[29113]= 1027042599;
assign addr[29114]= 1158676398;
assign addr[29115]= 1284432584;
assign addr[29116]= 1403673233;
assign addr[29117]= 1515793473;
assign addr[29118]= 1620224553;
assign addr[29119]= 1716436725;
assign addr[29120]= 1803941934;
assign addr[29121]= 1882296293;
assign addr[29122]= 1951102334;
assign addr[29123]= 2010011024;
assign addr[29124]= 2058723538;
assign addr[29125]= 2096992772;
assign addr[29126]= 2124624598;
assign addr[29127]= 2141478848;
assign addr[29128]= 2147470025;
assign addr[29129]= 2142567738;
assign addr[29130]= 2126796855;
assign addr[29131]= 2100237377;
assign addr[29132]= 2063024031;
assign addr[29133]= 2015345591;
assign addr[29134]= 1957443913;
assign addr[29135]= 1889612716;
assign addr[29136]= 1812196087;
assign addr[29137]= 1725586737;
assign addr[29138]= 1630224009;
assign addr[29139]= 1526591649;
assign addr[29140]= 1415215352;
assign addr[29141]= 1296660098;
assign addr[29142]= 1171527280;
assign addr[29143]= 1040451659;
assign addr[29144]= 904098143;
assign addr[29145]= 763158411;
assign addr[29146]= 618347408;
assign addr[29147]= 470399716;
assign addr[29148]= 320065829;
assign addr[29149]= 168108346;
assign addr[29150]= 15298099;
assign addr[29151]= -137589750;
assign addr[29152]= -289779648;
assign addr[29153]= -440499581;
assign addr[29154]= -588984994;
assign addr[29155]= -734482665;
assign addr[29156]= -876254528;
assign addr[29157]= -1013581418;
assign addr[29158]= -1145766716;
assign addr[29159]= -1272139887;
assign addr[29160]= -1392059879;
assign addr[29161]= -1504918373;
assign addr[29162]= -1610142873;
assign addr[29163]= -1707199606;
assign addr[29164]= -1795596234;
assign addr[29165]= -1874884346;
assign addr[29166]= -1944661739;
assign addr[29167]= -2004574453;
assign addr[29168]= -2054318569;
assign addr[29169]= -2093641749;
assign addr[29170]= -2122344521;
assign addr[29171]= -2140281282;
assign addr[29172]= -2147361045;
assign addr[29173]= -2143547897;
assign addr[29174]= -2128861181;
assign addr[29175]= -2103375398;
assign addr[29176]= -2067219829;
assign addr[29177]= -2020577882;
assign addr[29178]= -1963686155;
assign addr[29179]= -1896833245;
assign addr[29180]= -1820358275;
assign addr[29181]= -1734649179;
assign addr[29182]= -1640140734;
assign addr[29183]= -1537312353;
assign addr[29184]= -1426685652;
assign addr[29185]= -1308821808;
assign addr[29186]= -1184318708;
assign addr[29187]= -1053807919;
assign addr[29188]= -917951481;
assign addr[29189]= -777438554;
assign addr[29190]= -632981917;
assign addr[29191]= -485314355;
assign addr[29192]= -335184940;
assign addr[29193]= -183355234;
assign addr[29194]= -30595422;
assign addr[29195]= 122319591;
assign addr[29196]= 274614114;
assign addr[29197]= 425515602;
assign addr[29198]= 574258580;
assign addr[29199]= 720088517;
assign addr[29200]= 862265664;
assign addr[29201]= 1000068799;
assign addr[29202]= 1132798888;
assign addr[29203]= 1259782632;
assign addr[29204]= 1380375881;
assign addr[29205]= 1493966902;
assign addr[29206]= 1599979481;
assign addr[29207]= 1697875851;
assign addr[29208]= 1787159411;
assign addr[29209]= 1867377253;
assign addr[29210]= 1938122457;
assign addr[29211]= 1999036154;
assign addr[29212]= 2049809346;
assign addr[29213]= 2090184478;
assign addr[29214]= 2119956737;
assign addr[29215]= 2138975100;
assign addr[29216]= 2147143090;
assign addr[29217]= 2144419275;
assign addr[29218]= 2130817471;
assign addr[29219]= 2106406677;
assign addr[29220]= 2071310720;
assign addr[29221]= 2025707632;
assign addr[29222]= 1969828744;
assign addr[29223]= 1903957513;
assign addr[29224]= 1828428082;
assign addr[29225]= 1743623590;
assign addr[29226]= 1649974225;
assign addr[29227]= 1547955041;
assign addr[29228]= 1438083551;
assign addr[29229]= 1320917099;
assign addr[29230]= 1197050035;
assign addr[29231]= 1067110699;
assign addr[29232]= 931758235;
assign addr[29233]= 791679244;
assign addr[29234]= 647584304;
assign addr[29235]= 500204365;
assign addr[29236]= 350287041;
assign addr[29237]= 198592817;
assign addr[29238]= 45891193;
assign addr[29239]= -107043224;
assign addr[29240]= -259434643;
assign addr[29241]= -410510029;
assign addr[29242]= -559503022;
assign addr[29243]= -705657826;
assign addr[29244]= -848233042;
assign addr[29245]= -986505429;
assign addr[29246]= -1119773573;
assign addr[29247]= -1247361445;
assign addr[29248]= -1368621831;
assign addr[29249]= -1482939614;
assign addr[29250]= -1589734894;
assign addr[29251]= -1688465931;
assign addr[29252]= -1778631892;
assign addr[29253]= -1859775393;
assign addr[29254]= -1931484818;
assign addr[29255]= -1993396407;
assign addr[29256]= -2045196100;
assign addr[29257]= -2086621133;
assign addr[29258]= -2117461370;
assign addr[29259]= -2137560369;
assign addr[29260]= -2146816171;
assign addr[29261]= -2145181827;
assign addr[29262]= -2132665626;
assign addr[29263]= -2109331059;
assign addr[29264]= -2075296495;
assign addr[29265]= -2030734582;
assign addr[29266]= -1975871368;
assign addr[29267]= -1910985158;
assign addr[29268]= -1836405100;
assign addr[29269]= -1752509516;
assign addr[29270]= -1659723983;
assign addr[29271]= -1558519173;
assign addr[29272]= -1449408469;
assign addr[29273]= -1332945355;
assign addr[29274]= -1209720613;
assign addr[29275]= -1080359326;
assign addr[29276]= -945517704;
assign addr[29277]= -805879757;
assign addr[29278]= -662153826;
assign addr[29279]= -515068990;
assign addr[29280]= -365371365;
assign addr[29281]= -213820322;
assign addr[29282]= -61184634;
assign addr[29283]= 91761426;
assign addr[29284]= 244242007;
assign addr[29285]= 395483624;
assign addr[29286]= 544719071;
assign addr[29287]= 691191324;
assign addr[29288]= 834157373;
assign addr[29289]= 972891995;
assign addr[29290]= 1106691431;
assign addr[29291]= 1234876957;
assign addr[29292]= 1356798326;
assign addr[29293]= 1471837070;
assign addr[29294]= 1579409630;
assign addr[29295]= 1678970324;
assign addr[29296]= 1770014111;
assign addr[29297]= 1852079154;
assign addr[29298]= 1924749160;
assign addr[29299]= 1987655498;
assign addr[29300]= 2040479063;
assign addr[29301]= 2082951896;
assign addr[29302]= 2114858546;
assign addr[29303]= 2136037160;
assign addr[29304]= 2146380306;
assign addr[29305]= 2145835515;
assign addr[29306]= 2134405552;
assign addr[29307]= 2112148396;
assign addr[29308]= 2079176953;
assign addr[29309]= 2035658475;
assign addr[29310]= 1981813720;
assign addr[29311]= 1917915825;
assign addr[29312]= 1844288924;
assign addr[29313]= 1761306505;
assign addr[29314]= 1669389513;
assign addr[29315]= 1569004214;
assign addr[29316]= 1460659832;
assign addr[29317]= 1344905966;
assign addr[29318]= 1222329801;
assign addr[29319]= 1093553126;
assign addr[29320]= 959229189;
assign addr[29321]= 820039373;
assign addr[29322]= 676689746;
assign addr[29323]= 529907477;
assign addr[29324]= 380437148;
assign addr[29325]= 229036977;
assign addr[29326]= 76474970;
assign addr[29327]= -76474970;
assign addr[29328]= -229036977;
assign addr[29329]= -380437148;
assign addr[29330]= -529907477;
assign addr[29331]= -676689746;
assign addr[29332]= -820039373;
assign addr[29333]= -959229189;
assign addr[29334]= -1093553126;
assign addr[29335]= -1222329801;
assign addr[29336]= -1344905966;
assign addr[29337]= -1460659832;
assign addr[29338]= -1569004214;
assign addr[29339]= -1669389513;
assign addr[29340]= -1761306505;
assign addr[29341]= -1844288924;
assign addr[29342]= -1917915825;
assign addr[29343]= -1981813720;
assign addr[29344]= -2035658475;
assign addr[29345]= -2079176953;
assign addr[29346]= -2112148396;
assign addr[29347]= -2134405552;
assign addr[29348]= -2145835515;
assign addr[29349]= -2146380306;
assign addr[29350]= -2136037160;
assign addr[29351]= -2114858546;
assign addr[29352]= -2082951896;
assign addr[29353]= -2040479063;
assign addr[29354]= -1987655498;
assign addr[29355]= -1924749160;
assign addr[29356]= -1852079154;
assign addr[29357]= -1770014111;
assign addr[29358]= -1678970324;
assign addr[29359]= -1579409630;
assign addr[29360]= -1471837070;
assign addr[29361]= -1356798326;
assign addr[29362]= -1234876957;
assign addr[29363]= -1106691431;
assign addr[29364]= -972891995;
assign addr[29365]= -834157373;
assign addr[29366]= -691191324;
assign addr[29367]= -544719071;
assign addr[29368]= -395483624;
assign addr[29369]= -244242007;
assign addr[29370]= -91761426;
assign addr[29371]= 61184634;
assign addr[29372]= 213820322;
assign addr[29373]= 365371365;
assign addr[29374]= 515068990;
assign addr[29375]= 662153826;
assign addr[29376]= 805879757;
assign addr[29377]= 945517704;
assign addr[29378]= 1080359326;
assign addr[29379]= 1209720613;
assign addr[29380]= 1332945355;
assign addr[29381]= 1449408469;
assign addr[29382]= 1558519173;
assign addr[29383]= 1659723983;
assign addr[29384]= 1752509516;
assign addr[29385]= 1836405100;
assign addr[29386]= 1910985158;
assign addr[29387]= 1975871368;
assign addr[29388]= 2030734582;
assign addr[29389]= 2075296495;
assign addr[29390]= 2109331059;
assign addr[29391]= 2132665626;
assign addr[29392]= 2145181827;
assign addr[29393]= 2146816171;
assign addr[29394]= 2137560369;
assign addr[29395]= 2117461370;
assign addr[29396]= 2086621133;
assign addr[29397]= 2045196100;
assign addr[29398]= 1993396407;
assign addr[29399]= 1931484818;
assign addr[29400]= 1859775393;
assign addr[29401]= 1778631892;
assign addr[29402]= 1688465931;
assign addr[29403]= 1589734894;
assign addr[29404]= 1482939614;
assign addr[29405]= 1368621831;
assign addr[29406]= 1247361445;
assign addr[29407]= 1119773573;
assign addr[29408]= 986505429;
assign addr[29409]= 848233042;
assign addr[29410]= 705657826;
assign addr[29411]= 559503022;
assign addr[29412]= 410510029;
assign addr[29413]= 259434643;
assign addr[29414]= 107043224;
assign addr[29415]= -45891193;
assign addr[29416]= -198592817;
assign addr[29417]= -350287041;
assign addr[29418]= -500204365;
assign addr[29419]= -647584304;
assign addr[29420]= -791679244;
assign addr[29421]= -931758235;
assign addr[29422]= -1067110699;
assign addr[29423]= -1197050035;
assign addr[29424]= -1320917099;
assign addr[29425]= -1438083551;
assign addr[29426]= -1547955041;
assign addr[29427]= -1649974225;
assign addr[29428]= -1743623590;
assign addr[29429]= -1828428082;
assign addr[29430]= -1903957513;
assign addr[29431]= -1969828744;
assign addr[29432]= -2025707632;
assign addr[29433]= -2071310720;
assign addr[29434]= -2106406677;
assign addr[29435]= -2130817471;
assign addr[29436]= -2144419275;
assign addr[29437]= -2147143090;
assign addr[29438]= -2138975100;
assign addr[29439]= -2119956737;
assign addr[29440]= -2090184478;
assign addr[29441]= -2049809346;
assign addr[29442]= -1999036154;
assign addr[29443]= -1938122457;
assign addr[29444]= -1867377253;
assign addr[29445]= -1787159411;
assign addr[29446]= -1697875851;
assign addr[29447]= -1599979481;
assign addr[29448]= -1493966902;
assign addr[29449]= -1380375881;
assign addr[29450]= -1259782632;
assign addr[29451]= -1132798888;
assign addr[29452]= -1000068799;
assign addr[29453]= -862265664;
assign addr[29454]= -720088517;
assign addr[29455]= -574258580;
assign addr[29456]= -425515602;
assign addr[29457]= -274614114;
assign addr[29458]= -122319591;
assign addr[29459]= 30595422;
assign addr[29460]= 183355234;
assign addr[29461]= 335184940;
assign addr[29462]= 485314355;
assign addr[29463]= 632981917;
assign addr[29464]= 777438554;
assign addr[29465]= 917951481;
assign addr[29466]= 1053807919;
assign addr[29467]= 1184318708;
assign addr[29468]= 1308821808;
assign addr[29469]= 1426685652;
assign addr[29470]= 1537312353;
assign addr[29471]= 1640140734;
assign addr[29472]= 1734649179;
assign addr[29473]= 1820358275;
assign addr[29474]= 1896833245;
assign addr[29475]= 1963686155;
assign addr[29476]= 2020577882;
assign addr[29477]= 2067219829;
assign addr[29478]= 2103375398;
assign addr[29479]= 2128861181;
assign addr[29480]= 2143547897;
assign addr[29481]= 2147361045;
assign addr[29482]= 2140281282;
assign addr[29483]= 2122344521;
assign addr[29484]= 2093641749;
assign addr[29485]= 2054318569;
assign addr[29486]= 2004574453;
assign addr[29487]= 1944661739;
assign addr[29488]= 1874884346;
assign addr[29489]= 1795596234;
assign addr[29490]= 1707199606;
assign addr[29491]= 1610142873;
assign addr[29492]= 1504918373;
assign addr[29493]= 1392059879;
assign addr[29494]= 1272139887;
assign addr[29495]= 1145766716;
assign addr[29496]= 1013581418;
assign addr[29497]= 876254528;
assign addr[29498]= 734482665;
assign addr[29499]= 588984994;
assign addr[29500]= 440499581;
assign addr[29501]= 289779648;
assign addr[29502]= 137589750;
assign addr[29503]= -15298099;
assign addr[29504]= -168108346;
assign addr[29505]= -320065829;
assign addr[29506]= -470399716;
assign addr[29507]= -618347408;
assign addr[29508]= -763158411;
assign addr[29509]= -904098143;
assign addr[29510]= -1040451659;
assign addr[29511]= -1171527280;
assign addr[29512]= -1296660098;
assign addr[29513]= -1415215352;
assign addr[29514]= -1526591649;
assign addr[29515]= -1630224009;
assign addr[29516]= -1725586737;
assign addr[29517]= -1812196087;
assign addr[29518]= -1889612716;
assign addr[29519]= -1957443913;
assign addr[29520]= -2015345591;
assign addr[29521]= -2063024031;
assign addr[29522]= -2100237377;
assign addr[29523]= -2126796855;
assign addr[29524]= -2142567738;
assign addr[29525]= -2147470025;
assign addr[29526]= -2141478848;
assign addr[29527]= -2124624598;
assign addr[29528]= -2096992772;
assign addr[29529]= -2058723538;
assign addr[29530]= -2010011024;
assign addr[29531]= -1951102334;
assign addr[29532]= -1882296293;
assign addr[29533]= -1803941934;
assign addr[29534]= -1716436725;
assign addr[29535]= -1620224553;
assign addr[29536]= -1515793473;
assign addr[29537]= -1403673233;
assign addr[29538]= -1284432584;
assign addr[29539]= -1158676398;
assign addr[29540]= -1027042599;
assign addr[29541]= -890198924;
assign addr[29542]= -748839539;
assign addr[29543]= -603681519;
assign addr[29544]= -455461206;
assign addr[29545]= -304930476;
assign addr[29546]= -152852926;
assign addr[29547]= 0;
assign addr[29548]= 152852926;
assign addr[29549]= 304930476;
assign addr[29550]= 455461206;
assign addr[29551]= 603681519;
assign addr[29552]= 748839539;
assign addr[29553]= 890198924;
assign addr[29554]= 1027042599;
assign addr[29555]= 1158676398;
assign addr[29556]= 1284432584;
assign addr[29557]= 1403673233;
assign addr[29558]= 1515793473;
assign addr[29559]= 1620224553;
assign addr[29560]= 1716436725;
assign addr[29561]= 1803941934;
assign addr[29562]= 1882296293;
assign addr[29563]= 1951102334;
assign addr[29564]= 2010011024;
assign addr[29565]= 2058723538;
assign addr[29566]= 2096992772;
assign addr[29567]= 2124624598;
assign addr[29568]= 2141478848;
assign addr[29569]= 2147470025;
assign addr[29570]= 2142567738;
assign addr[29571]= 2126796855;
assign addr[29572]= 2100237377;
assign addr[29573]= 2063024031;
assign addr[29574]= 2015345591;
assign addr[29575]= 1957443913;
assign addr[29576]= 1889612716;
assign addr[29577]= 1812196087;
assign addr[29578]= 1725586737;
assign addr[29579]= 1630224009;
assign addr[29580]= 1526591649;
assign addr[29581]= 1415215352;
assign addr[29582]= 1296660098;
assign addr[29583]= 1171527280;
assign addr[29584]= 1040451659;
assign addr[29585]= 904098143;
assign addr[29586]= 763158411;
assign addr[29587]= 618347408;
assign addr[29588]= 470399716;
assign addr[29589]= 320065829;
assign addr[29590]= 168108346;
assign addr[29591]= 15298099;
assign addr[29592]= -137589750;
assign addr[29593]= -289779648;
assign addr[29594]= -440499581;
assign addr[29595]= -588984994;
assign addr[29596]= -734482665;
assign addr[29597]= -876254528;
assign addr[29598]= -1013581418;
assign addr[29599]= -1145766716;
assign addr[29600]= -1272139887;
assign addr[29601]= -1392059879;
assign addr[29602]= -1504918373;
assign addr[29603]= -1610142873;
assign addr[29604]= -1707199606;
assign addr[29605]= -1795596234;
assign addr[29606]= -1874884346;
assign addr[29607]= -1944661739;
assign addr[29608]= -2004574453;
assign addr[29609]= -2054318569;
assign addr[29610]= -2093641749;
assign addr[29611]= -2122344521;
assign addr[29612]= -2140281282;
assign addr[29613]= -2147361045;
assign addr[29614]= -2143547897;
assign addr[29615]= -2128861181;
assign addr[29616]= -2103375398;
assign addr[29617]= -2067219829;
assign addr[29618]= -2020577882;
assign addr[29619]= -1963686155;
assign addr[29620]= -1896833245;
assign addr[29621]= -1820358275;
assign addr[29622]= -1734649179;
assign addr[29623]= -1640140734;
assign addr[29624]= -1537312353;
assign addr[29625]= -1426685652;
assign addr[29626]= -1308821808;
assign addr[29627]= -1184318708;
assign addr[29628]= -1053807919;
assign addr[29629]= -917951481;
assign addr[29630]= -777438554;
assign addr[29631]= -632981917;
assign addr[29632]= -485314355;
assign addr[29633]= -335184940;
assign addr[29634]= -183355234;
assign addr[29635]= -30595422;
assign addr[29636]= 122319591;
assign addr[29637]= 274614114;
assign addr[29638]= 425515602;
assign addr[29639]= 574258580;
assign addr[29640]= 720088517;
assign addr[29641]= 862265664;
assign addr[29642]= 1000068799;
assign addr[29643]= 1132798888;
assign addr[29644]= 1259782632;
assign addr[29645]= 1380375881;
assign addr[29646]= 1493966902;
assign addr[29647]= 1599979481;
assign addr[29648]= 1697875851;
assign addr[29649]= 1787159411;
assign addr[29650]= 1867377253;
assign addr[29651]= 1938122457;
assign addr[29652]= 1999036154;
assign addr[29653]= 2049809346;
assign addr[29654]= 2090184478;
assign addr[29655]= 2119956737;
assign addr[29656]= 2138975100;
assign addr[29657]= 2147143090;
assign addr[29658]= 2144419275;
assign addr[29659]= 2130817471;
assign addr[29660]= 2106406677;
assign addr[29661]= 2071310720;
assign addr[29662]= 2025707632;
assign addr[29663]= 1969828744;
assign addr[29664]= 1903957513;
assign addr[29665]= 1828428082;
assign addr[29666]= 1743623590;
assign addr[29667]= 1649974225;
assign addr[29668]= 1547955041;
assign addr[29669]= 1438083551;
assign addr[29670]= 1320917099;
assign addr[29671]= 1197050035;
assign addr[29672]= 1067110699;
assign addr[29673]= 931758235;
assign addr[29674]= 791679244;
assign addr[29675]= 647584304;
assign addr[29676]= 500204365;
assign addr[29677]= 350287041;
assign addr[29678]= 198592817;
assign addr[29679]= 45891193;
assign addr[29680]= -107043224;
assign addr[29681]= -259434643;
assign addr[29682]= -410510029;
assign addr[29683]= -559503022;
assign addr[29684]= -705657826;
assign addr[29685]= -848233042;
assign addr[29686]= -986505429;
assign addr[29687]= -1119773573;
assign addr[29688]= -1247361445;
assign addr[29689]= -1368621831;
assign addr[29690]= -1482939614;
assign addr[29691]= -1589734894;
assign addr[29692]= -1688465931;
assign addr[29693]= -1778631892;
assign addr[29694]= -1859775393;
assign addr[29695]= -1931484818;
assign addr[29696]= -1993396407;
assign addr[29697]= -2045196100;
assign addr[29698]= -2086621133;
assign addr[29699]= -2117461370;
assign addr[29700]= -2137560369;
assign addr[29701]= -2146816171;
assign addr[29702]= -2145181827;
assign addr[29703]= -2132665626;
assign addr[29704]= -2109331059;
assign addr[29705]= -2075296495;
assign addr[29706]= -2030734582;
assign addr[29707]= -1975871368;
assign addr[29708]= -1910985158;
assign addr[29709]= -1836405100;
assign addr[29710]= -1752509516;
assign addr[29711]= -1659723983;
assign addr[29712]= -1558519173;
assign addr[29713]= -1449408469;
assign addr[29714]= -1332945355;
assign addr[29715]= -1209720613;
assign addr[29716]= -1080359326;
assign addr[29717]= -945517704;
assign addr[29718]= -805879757;
assign addr[29719]= -662153826;
assign addr[29720]= -515068990;
assign addr[29721]= -365371365;
assign addr[29722]= -213820322;
assign addr[29723]= -61184634;
assign addr[29724]= 91761426;
assign addr[29725]= 244242007;
assign addr[29726]= 395483624;
assign addr[29727]= 544719071;
assign addr[29728]= 691191324;
assign addr[29729]= 834157373;
assign addr[29730]= 972891995;
assign addr[29731]= 1106691431;
assign addr[29732]= 1234876957;
assign addr[29733]= 1356798326;
assign addr[29734]= 1471837070;
assign addr[29735]= 1579409630;
assign addr[29736]= 1678970324;
assign addr[29737]= 1770014111;
assign addr[29738]= 1852079154;
assign addr[29739]= 1924749160;
assign addr[29740]= 1987655498;
assign addr[29741]= 2040479063;
assign addr[29742]= 2082951896;
assign addr[29743]= 2114858546;
assign addr[29744]= 2136037160;
assign addr[29745]= 2146380306;
assign addr[29746]= 2145835515;
assign addr[29747]= 2134405552;
assign addr[29748]= 2112148396;
assign addr[29749]= 2079176953;
assign addr[29750]= 2035658475;
assign addr[29751]= 1981813720;
assign addr[29752]= 1917915825;
assign addr[29753]= 1844288924;
assign addr[29754]= 1761306505;
assign addr[29755]= 1669389513;
assign addr[29756]= 1569004214;
assign addr[29757]= 1460659832;
assign addr[29758]= 1344905966;
assign addr[29759]= 1222329801;
assign addr[29760]= 1093553126;
assign addr[29761]= 959229189;
assign addr[29762]= 820039373;
assign addr[29763]= 676689746;
assign addr[29764]= 529907477;
assign addr[29765]= 380437148;
assign addr[29766]= 229036977;
assign addr[29767]= 76474970;
assign addr[29768]= -76474970;
assign addr[29769]= -229036977;
assign addr[29770]= -380437148;
assign addr[29771]= -529907477;
assign addr[29772]= -676689746;
assign addr[29773]= -820039373;
assign addr[29774]= -959229189;
assign addr[29775]= -1093553126;
assign addr[29776]= -1222329801;
assign addr[29777]= -1344905966;
assign addr[29778]= -1460659832;
assign addr[29779]= -1569004214;
assign addr[29780]= -1669389513;
assign addr[29781]= -1761306505;
assign addr[29782]= -1844288924;
assign addr[29783]= -1917915825;
assign addr[29784]= -1981813720;
assign addr[29785]= -2035658475;
assign addr[29786]= -2079176953;
assign addr[29787]= -2112148396;
assign addr[29788]= -2134405552;
assign addr[29789]= -2145835515;
assign addr[29790]= -2146380306;
assign addr[29791]= -2136037160;
assign addr[29792]= -2114858546;
assign addr[29793]= -2082951896;
assign addr[29794]= -2040479063;
assign addr[29795]= -1987655498;
assign addr[29796]= -1924749160;
assign addr[29797]= -1852079154;
assign addr[29798]= -1770014111;
assign addr[29799]= -1678970324;
assign addr[29800]= -1579409630;
assign addr[29801]= -1471837070;
assign addr[29802]= -1356798326;
assign addr[29803]= -1234876957;
assign addr[29804]= -1106691431;
assign addr[29805]= -972891995;
assign addr[29806]= -834157373;
assign addr[29807]= -691191324;
assign addr[29808]= -544719071;
assign addr[29809]= -395483624;
assign addr[29810]= -244242007;
assign addr[29811]= -91761426;
assign addr[29812]= 61184634;
assign addr[29813]= 213820322;
assign addr[29814]= 365371365;
assign addr[29815]= 515068990;
assign addr[29816]= 662153826;
assign addr[29817]= 805879757;
assign addr[29818]= 945517704;
assign addr[29819]= 1080359326;
assign addr[29820]= 1209720613;
assign addr[29821]= 1332945355;
assign addr[29822]= 1449408469;
assign addr[29823]= 1558519173;
assign addr[29824]= 1659723983;
assign addr[29825]= 1752509516;
assign addr[29826]= 1836405100;
assign addr[29827]= 1910985158;
assign addr[29828]= 1975871368;
assign addr[29829]= 2030734582;
assign addr[29830]= 2075296495;
assign addr[29831]= 2109331059;
assign addr[29832]= 2132665626;
assign addr[29833]= 2145181827;
assign addr[29834]= 2146816171;
assign addr[29835]= 2137560369;
assign addr[29836]= 2117461370;
assign addr[29837]= 2086621133;
assign addr[29838]= 2045196100;
assign addr[29839]= 1993396407;
assign addr[29840]= 1931484818;
assign addr[29841]= 1859775393;
assign addr[29842]= 1778631892;
assign addr[29843]= 1688465931;
assign addr[29844]= 1589734894;
assign addr[29845]= 1482939614;
assign addr[29846]= 1368621831;
assign addr[29847]= 1247361445;
assign addr[29848]= 1119773573;
assign addr[29849]= 986505429;
assign addr[29850]= 848233042;
assign addr[29851]= 705657826;
assign addr[29852]= 559503022;
assign addr[29853]= 410510029;
assign addr[29854]= 259434643;
assign addr[29855]= 107043224;
assign addr[29856]= -45891193;
assign addr[29857]= -198592817;
assign addr[29858]= -350287041;
assign addr[29859]= -500204365;
assign addr[29860]= -647584304;
assign addr[29861]= -791679244;
assign addr[29862]= -931758235;
assign addr[29863]= -1067110699;
assign addr[29864]= -1197050035;
assign addr[29865]= -1320917099;
assign addr[29866]= -1438083551;
assign addr[29867]= -1547955041;
assign addr[29868]= -1649974225;
assign addr[29869]= -1743623590;
assign addr[29870]= -1828428082;
assign addr[29871]= -1903957513;
assign addr[29872]= -1969828744;
assign addr[29873]= -2025707632;
assign addr[29874]= -2071310720;
assign addr[29875]= -2106406677;
assign addr[29876]= -2130817471;
assign addr[29877]= -2144419275;
assign addr[29878]= -2147143090;
assign addr[29879]= -2138975100;
assign addr[29880]= -2119956737;
assign addr[29881]= -2090184478;
assign addr[29882]= -2049809346;
assign addr[29883]= -1999036154;
assign addr[29884]= -1938122457;
assign addr[29885]= -1867377253;
assign addr[29886]= -1787159411;
assign addr[29887]= -1697875851;
assign addr[29888]= -1599979481;
assign addr[29889]= -1493966902;
assign addr[29890]= -1380375881;
assign addr[29891]= -1259782632;
assign addr[29892]= -1132798888;
assign addr[29893]= -1000068799;
assign addr[29894]= -862265664;
assign addr[29895]= -720088517;
assign addr[29896]= -574258580;
assign addr[29897]= -425515602;
assign addr[29898]= -274614114;
assign addr[29899]= -122319591;
assign addr[29900]= 30595422;
assign addr[29901]= 183355234;
assign addr[29902]= 335184940;
assign addr[29903]= 485314355;
assign addr[29904]= 632981917;
assign addr[29905]= 777438554;
assign addr[29906]= 917951481;
assign addr[29907]= 1053807919;
assign addr[29908]= 1184318708;
assign addr[29909]= 1308821808;
assign addr[29910]= 1426685652;
assign addr[29911]= 1537312353;
assign addr[29912]= 1640140734;
assign addr[29913]= 1734649179;
assign addr[29914]= 1820358275;
assign addr[29915]= 1896833245;
assign addr[29916]= 1963686155;
assign addr[29917]= 2020577882;
assign addr[29918]= 2067219829;
assign addr[29919]= 2103375398;
assign addr[29920]= 2128861181;
assign addr[29921]= 2143547897;
assign addr[29922]= 2147361045;
assign addr[29923]= 2140281282;
assign addr[29924]= 2122344521;
assign addr[29925]= 2093641749;
assign addr[29926]= 2054318569;
assign addr[29927]= 2004574453;
assign addr[29928]= 1944661739;
assign addr[29929]= 1874884346;
assign addr[29930]= 1795596234;
assign addr[29931]= 1707199606;
assign addr[29932]= 1610142873;
assign addr[29933]= 1504918373;
assign addr[29934]= 1392059879;
assign addr[29935]= 1272139887;
assign addr[29936]= 1145766716;
assign addr[29937]= 1013581418;
assign addr[29938]= 876254528;
assign addr[29939]= 734482665;
assign addr[29940]= 588984994;
assign addr[29941]= 440499581;
assign addr[29942]= 289779648;
assign addr[29943]= 137589750;
assign addr[29944]= -15298099;
assign addr[29945]= -168108346;
assign addr[29946]= -320065829;
assign addr[29947]= -470399716;
assign addr[29948]= -618347408;
assign addr[29949]= -763158411;
assign addr[29950]= -904098143;
assign addr[29951]= -1040451659;
assign addr[29952]= -1171527280;
assign addr[29953]= -1296660098;
assign addr[29954]= -1415215352;
assign addr[29955]= -1526591649;
assign addr[29956]= -1630224009;
assign addr[29957]= -1725586737;
assign addr[29958]= -1812196087;
assign addr[29959]= -1889612716;
assign addr[29960]= -1957443913;
assign addr[29961]= -2015345591;
assign addr[29962]= -2063024031;
assign addr[29963]= -2100237377;
assign addr[29964]= -2126796855;
assign addr[29965]= -2142567738;
assign addr[29966]= -2147470025;
assign addr[29967]= -2141478848;
assign addr[29968]= -2124624598;
assign addr[29969]= -2096992772;
assign addr[29970]= -2058723538;
assign addr[29971]= -2010011024;
assign addr[29972]= -1951102334;
assign addr[29973]= -1882296293;
assign addr[29974]= -1803941934;
assign addr[29975]= -1716436725;
assign addr[29976]= -1620224553;
assign addr[29977]= -1515793473;
assign addr[29978]= -1403673233;
assign addr[29979]= -1284432584;
assign addr[29980]= -1158676398;
assign addr[29981]= -1027042599;
assign addr[29982]= -890198924;
assign addr[29983]= -748839539;
assign addr[29984]= -603681519;
assign addr[29985]= -455461206;
assign addr[29986]= -304930476;
assign addr[29987]= -152852926;
assign addr[29988]= 0;
assign addr[29989]= 152852926;
assign addr[29990]= 304930476;
assign addr[29991]= 455461206;
assign addr[29992]= 603681519;
assign addr[29993]= 748839539;
assign addr[29994]= 890198924;
assign addr[29995]= 1027042599;
assign addr[29996]= 1158676398;
assign addr[29997]= 1284432584;
assign addr[29998]= 1403673233;
assign addr[29999]= 1515793473;
assign addr[30000]= 1620224553;
assign addr[30001]= 1716436725;
assign addr[30002]= 1803941934;
assign addr[30003]= 1882296293;
assign addr[30004]= 1951102334;
assign addr[30005]= 2010011024;
assign addr[30006]= 2058723538;
assign addr[30007]= 2096992772;
assign addr[30008]= 2124624598;
assign addr[30009]= 2141478848;
assign addr[30010]= 2147470025;
assign addr[30011]= 2142567738;
assign addr[30012]= 2126796855;
assign addr[30013]= 2100237377;
assign addr[30014]= 2063024031;
assign addr[30015]= 2015345591;
assign addr[30016]= 1957443913;
assign addr[30017]= 1889612716;
assign addr[30018]= 1812196087;
assign addr[30019]= 1725586737;
assign addr[30020]= 1630224009;
assign addr[30021]= 1526591649;
assign addr[30022]= 1415215352;
assign addr[30023]= 1296660098;
assign addr[30024]= 1171527280;
assign addr[30025]= 1040451659;
assign addr[30026]= 904098143;
assign addr[30027]= 763158411;
assign addr[30028]= 618347408;
assign addr[30029]= 470399716;
assign addr[30030]= 320065829;
assign addr[30031]= 168108346;
assign addr[30032]= 15298099;
assign addr[30033]= -137589750;
assign addr[30034]= -289779648;
assign addr[30035]= -440499581;
assign addr[30036]= -588984994;
assign addr[30037]= -734482665;
assign addr[30038]= -876254528;
assign addr[30039]= -1013581418;
assign addr[30040]= -1145766716;
assign addr[30041]= -1272139887;
assign addr[30042]= -1392059879;
assign addr[30043]= -1504918373;
assign addr[30044]= -1610142873;
assign addr[30045]= -1707199606;
assign addr[30046]= -1795596234;
assign addr[30047]= -1874884346;
assign addr[30048]= -1944661739;
assign addr[30049]= -2004574453;
assign addr[30050]= -2054318569;
assign addr[30051]= -2093641749;
assign addr[30052]= -2122344521;
assign addr[30053]= -2140281282;
assign addr[30054]= -2147361045;
assign addr[30055]= -2143547897;
assign addr[30056]= -2128861181;
assign addr[30057]= -2103375398;
assign addr[30058]= -2067219829;
assign addr[30059]= -2020577882;
assign addr[30060]= -1963686155;
assign addr[30061]= -1896833245;
assign addr[30062]= -1820358275;
assign addr[30063]= -1734649179;
assign addr[30064]= -1640140734;
assign addr[30065]= -1537312353;
assign addr[30066]= -1426685652;
assign addr[30067]= -1308821808;
assign addr[30068]= -1184318708;
assign addr[30069]= -1053807919;
assign addr[30070]= -917951481;
assign addr[30071]= -777438554;
assign addr[30072]= -632981917;
assign addr[30073]= -485314355;
assign addr[30074]= -335184940;
assign addr[30075]= -183355234;
assign addr[30076]= -30595422;
assign addr[30077]= 122319591;
assign addr[30078]= 274614114;
assign addr[30079]= 425515602;
assign addr[30080]= 574258580;
assign addr[30081]= 720088517;
assign addr[30082]= 862265664;
assign addr[30083]= 1000068799;
assign addr[30084]= 1132798888;
assign addr[30085]= 1259782632;
assign addr[30086]= 1380375881;
assign addr[30087]= 1493966902;
assign addr[30088]= 1599979481;
assign addr[30089]= 1697875851;
assign addr[30090]= 1787159411;
assign addr[30091]= 1867377253;
assign addr[30092]= 1938122457;
assign addr[30093]= 1999036154;
assign addr[30094]= 2049809346;
assign addr[30095]= 2090184478;
assign addr[30096]= 2119956737;
assign addr[30097]= 2138975100;
assign addr[30098]= 2147143090;
assign addr[30099]= 2144419275;
assign addr[30100]= 2130817471;
assign addr[30101]= 2106406677;
assign addr[30102]= 2071310720;
assign addr[30103]= 2025707632;
assign addr[30104]= 1969828744;
assign addr[30105]= 1903957513;
assign addr[30106]= 1828428082;
assign addr[30107]= 1743623590;
assign addr[30108]= 1649974225;
assign addr[30109]= 1547955041;
assign addr[30110]= 1438083551;
assign addr[30111]= 1320917099;
assign addr[30112]= 1197050035;
assign addr[30113]= 1067110699;
assign addr[30114]= 931758235;
assign addr[30115]= 791679244;
assign addr[30116]= 647584304;
assign addr[30117]= 500204365;
assign addr[30118]= 350287041;
assign addr[30119]= 198592817;
assign addr[30120]= 45891193;
assign addr[30121]= -107043224;
assign addr[30122]= -259434643;
assign addr[30123]= -410510029;
assign addr[30124]= -559503022;
assign addr[30125]= -705657826;
assign addr[30126]= -848233042;
assign addr[30127]= -986505429;
assign addr[30128]= -1119773573;
assign addr[30129]= -1247361445;
assign addr[30130]= -1368621831;
assign addr[30131]= -1482939614;
assign addr[30132]= -1589734894;
assign addr[30133]= -1688465931;
assign addr[30134]= -1778631892;
assign addr[30135]= -1859775393;
assign addr[30136]= -1931484818;
assign addr[30137]= -1993396407;
assign addr[30138]= -2045196100;
assign addr[30139]= -2086621133;
assign addr[30140]= -2117461370;
assign addr[30141]= -2137560369;
assign addr[30142]= -2146816171;
assign addr[30143]= -2145181827;
assign addr[30144]= -2132665626;
assign addr[30145]= -2109331059;
assign addr[30146]= -2075296495;
assign addr[30147]= -2030734582;
assign addr[30148]= -1975871368;
assign addr[30149]= -1910985158;
assign addr[30150]= -1836405100;
assign addr[30151]= -1752509516;
assign addr[30152]= -1659723983;
assign addr[30153]= -1558519173;
assign addr[30154]= -1449408469;
assign addr[30155]= -1332945355;
assign addr[30156]= -1209720613;
assign addr[30157]= -1080359326;
assign addr[30158]= -945517704;
assign addr[30159]= -805879757;
assign addr[30160]= -662153826;
assign addr[30161]= -515068990;
assign addr[30162]= -365371365;
assign addr[30163]= -213820322;
assign addr[30164]= -61184634;
assign addr[30165]= 91761426;
assign addr[30166]= 244242007;
assign addr[30167]= 395483624;
assign addr[30168]= 544719071;
assign addr[30169]= 691191324;
assign addr[30170]= 834157373;
assign addr[30171]= 972891995;
assign addr[30172]= 1106691431;
assign addr[30173]= 1234876957;
assign addr[30174]= 1356798326;
assign addr[30175]= 1471837070;
assign addr[30176]= 1579409630;
assign addr[30177]= 1678970324;
assign addr[30178]= 1770014111;
assign addr[30179]= 1852079154;
assign addr[30180]= 1924749160;
assign addr[30181]= 1987655498;
assign addr[30182]= 2040479063;
assign addr[30183]= 2082951896;
assign addr[30184]= 2114858546;
assign addr[30185]= 2136037160;
assign addr[30186]= 2146380306;
assign addr[30187]= 2145835515;
assign addr[30188]= 2134405552;
assign addr[30189]= 2112148396;
assign addr[30190]= 2079176953;
assign addr[30191]= 2035658475;
assign addr[30192]= 1981813720;
assign addr[30193]= 1917915825;
assign addr[30194]= 1844288924;
assign addr[30195]= 1761306505;
assign addr[30196]= 1669389513;
assign addr[30197]= 1569004214;
assign addr[30198]= 1460659832;
assign addr[30199]= 1344905966;
assign addr[30200]= 1222329801;
assign addr[30201]= 1093553126;
assign addr[30202]= 959229189;
assign addr[30203]= 820039373;
assign addr[30204]= 676689746;
assign addr[30205]= 529907477;
assign addr[30206]= 380437148;
assign addr[30207]= 229036977;
assign addr[30208]= 76474970;
assign addr[30209]= -76474970;
assign addr[30210]= -229036977;
assign addr[30211]= -380437148;
assign addr[30212]= -529907477;
assign addr[30213]= -676689746;
assign addr[30214]= -820039373;
assign addr[30215]= -959229189;
assign addr[30216]= -1093553126;
assign addr[30217]= -1222329801;
assign addr[30218]= -1344905966;
assign addr[30219]= -1460659832;
assign addr[30220]= -1569004214;
assign addr[30221]= -1669389513;
assign addr[30222]= -1761306505;
assign addr[30223]= -1844288924;
assign addr[30224]= -1917915825;
assign addr[30225]= -1981813720;
assign addr[30226]= -2035658475;
assign addr[30227]= -2079176953;
assign addr[30228]= -2112148396;
assign addr[30229]= -2134405552;
assign addr[30230]= -2145835515;
assign addr[30231]= -2146380306;
assign addr[30232]= -2136037160;
assign addr[30233]= -2114858546;
assign addr[30234]= -2082951896;
assign addr[30235]= -2040479063;
assign addr[30236]= -1987655498;
assign addr[30237]= -1924749160;
assign addr[30238]= -1852079154;
assign addr[30239]= -1770014111;
assign addr[30240]= -1678970324;
assign addr[30241]= -1579409630;
assign addr[30242]= -1471837070;
assign addr[30243]= -1356798326;
assign addr[30244]= -1234876957;
assign addr[30245]= -1106691431;
assign addr[30246]= -972891995;
assign addr[30247]= -834157373;
assign addr[30248]= -691191324;
assign addr[30249]= -544719071;
assign addr[30250]= -395483624;
assign addr[30251]= -244242007;
assign addr[30252]= -91761426;
assign addr[30253]= 61184634;
assign addr[30254]= 213820322;
assign addr[30255]= 365371365;
assign addr[30256]= 515068990;
assign addr[30257]= 662153826;
assign addr[30258]= 805879757;
assign addr[30259]= 945517704;
assign addr[30260]= 1080359326;
assign addr[30261]= 1209720613;
assign addr[30262]= 1332945355;
assign addr[30263]= 1449408469;
assign addr[30264]= 1558519173;
assign addr[30265]= 1659723983;
assign addr[30266]= 1752509516;
assign addr[30267]= 1836405100;
assign addr[30268]= 1910985158;
assign addr[30269]= 1975871368;
assign addr[30270]= 2030734582;
assign addr[30271]= 2075296495;
assign addr[30272]= 2109331059;
assign addr[30273]= 2132665626;
assign addr[30274]= 2145181827;
assign addr[30275]= 2146816171;
assign addr[30276]= 2137560369;
assign addr[30277]= 2117461370;
assign addr[30278]= 2086621133;
assign addr[30279]= 2045196100;
assign addr[30280]= 1993396407;
assign addr[30281]= 1931484818;
assign addr[30282]= 1859775393;
assign addr[30283]= 1778631892;
assign addr[30284]= 1688465931;
assign addr[30285]= 1589734894;
assign addr[30286]= 1482939614;
assign addr[30287]= 1368621831;
assign addr[30288]= 1247361445;
assign addr[30289]= 1119773573;
assign addr[30290]= 986505429;
assign addr[30291]= 848233042;
assign addr[30292]= 705657826;
assign addr[30293]= 559503022;
assign addr[30294]= 410510029;
assign addr[30295]= 259434643;
assign addr[30296]= 107043224;
assign addr[30297]= -45891193;
assign addr[30298]= -198592817;
assign addr[30299]= -350287041;
assign addr[30300]= -500204365;
assign addr[30301]= -647584304;
assign addr[30302]= -791679244;
assign addr[30303]= -931758235;
assign addr[30304]= -1067110699;
assign addr[30305]= -1197050035;
assign addr[30306]= -1320917099;
assign addr[30307]= -1438083551;
assign addr[30308]= -1547955041;
assign addr[30309]= -1649974225;
assign addr[30310]= -1743623590;
assign addr[30311]= -1828428082;
assign addr[30312]= -1903957513;
assign addr[30313]= -1969828744;
assign addr[30314]= -2025707632;
assign addr[30315]= -2071310720;
assign addr[30316]= -2106406677;
assign addr[30317]= -2130817471;
assign addr[30318]= -2144419275;
assign addr[30319]= -2147143090;
assign addr[30320]= -2138975100;
assign addr[30321]= -2119956737;
assign addr[30322]= -2090184478;
assign addr[30323]= -2049809346;
assign addr[30324]= -1999036154;
assign addr[30325]= -1938122457;
assign addr[30326]= -1867377253;
assign addr[30327]= -1787159411;
assign addr[30328]= -1697875851;
assign addr[30329]= -1599979481;
assign addr[30330]= -1493966902;
assign addr[30331]= -1380375881;
assign addr[30332]= -1259782632;
assign addr[30333]= -1132798888;
assign addr[30334]= -1000068799;
assign addr[30335]= -862265664;
assign addr[30336]= -720088517;
assign addr[30337]= -574258580;
assign addr[30338]= -425515602;
assign addr[30339]= -274614114;
assign addr[30340]= -122319591;
assign addr[30341]= 30595422;
assign addr[30342]= 183355234;
assign addr[30343]= 335184940;
assign addr[30344]= 485314355;
assign addr[30345]= 632981917;
assign addr[30346]= 777438554;
assign addr[30347]= 917951481;
assign addr[30348]= 1053807919;
assign addr[30349]= 1184318708;
assign addr[30350]= 1308821808;
assign addr[30351]= 1426685652;
assign addr[30352]= 1537312353;
assign addr[30353]= 1640140734;
assign addr[30354]= 1734649179;
assign addr[30355]= 1820358275;
assign addr[30356]= 1896833245;
assign addr[30357]= 1963686155;
assign addr[30358]= 2020577882;
assign addr[30359]= 2067219829;
assign addr[30360]= 2103375398;
assign addr[30361]= 2128861181;
assign addr[30362]= 2143547897;
assign addr[30363]= 2147361045;
assign addr[30364]= 2140281282;
assign addr[30365]= 2122344521;
assign addr[30366]= 2093641749;
assign addr[30367]= 2054318569;
assign addr[30368]= 2004574453;
assign addr[30369]= 1944661739;
assign addr[30370]= 1874884346;
assign addr[30371]= 1795596234;
assign addr[30372]= 1707199606;
assign addr[30373]= 1610142873;
assign addr[30374]= 1504918373;
assign addr[30375]= 1392059879;
assign addr[30376]= 1272139887;
assign addr[30377]= 1145766716;
assign addr[30378]= 1013581418;
assign addr[30379]= 876254528;
assign addr[30380]= 734482665;
assign addr[30381]= 588984994;
assign addr[30382]= 440499581;
assign addr[30383]= 289779648;
assign addr[30384]= 137589750;
assign addr[30385]= -15298099;
assign addr[30386]= -168108346;
assign addr[30387]= -320065829;
assign addr[30388]= -470399716;
assign addr[30389]= -618347408;
assign addr[30390]= -763158411;
assign addr[30391]= -904098143;
assign addr[30392]= -1040451659;
assign addr[30393]= -1171527280;
assign addr[30394]= -1296660098;
assign addr[30395]= -1415215352;
assign addr[30396]= -1526591649;
assign addr[30397]= -1630224009;
assign addr[30398]= -1725586737;
assign addr[30399]= -1812196087;
assign addr[30400]= -1889612716;
assign addr[30401]= -1957443913;
assign addr[30402]= -2015345591;
assign addr[30403]= -2063024031;
assign addr[30404]= -2100237377;
assign addr[30405]= -2126796855;
assign addr[30406]= -2142567738;
assign addr[30407]= -2147470025;
assign addr[30408]= -2141478848;
assign addr[30409]= -2124624598;
assign addr[30410]= -2096992772;
assign addr[30411]= -2058723538;
assign addr[30412]= -2010011024;
assign addr[30413]= -1951102334;
assign addr[30414]= -1882296293;
assign addr[30415]= -1803941934;
assign addr[30416]= -1716436725;
assign addr[30417]= -1620224553;
assign addr[30418]= -1515793473;
assign addr[30419]= -1403673233;
assign addr[30420]= -1284432584;
assign addr[30421]= -1158676398;
assign addr[30422]= -1027042599;
assign addr[30423]= -890198924;
assign addr[30424]= -748839539;
assign addr[30425]= -603681519;
assign addr[30426]= -455461206;
assign addr[30427]= -304930476;
assign addr[30428]= -152852926;
assign addr[30429]= 0;
assign addr[30430]= 152852926;
assign addr[30431]= 304930476;
assign addr[30432]= 455461206;
assign addr[30433]= 603681519;
assign addr[30434]= 748839539;
assign addr[30435]= 890198924;
assign addr[30436]= 1027042599;
assign addr[30437]= 1158676398;
assign addr[30438]= 1284432584;
assign addr[30439]= 1403673233;
assign addr[30440]= 1515793473;
assign addr[30441]= 1620224553;
assign addr[30442]= 1716436725;
assign addr[30443]= 1803941934;
assign addr[30444]= 1882296293;
assign addr[30445]= 1951102334;
assign addr[30446]= 2010011024;
assign addr[30447]= 2058723538;
assign addr[30448]= 2096992772;
assign addr[30449]= 2124624598;
assign addr[30450]= 2141478848;
assign addr[30451]= 2147470025;
assign addr[30452]= 2142567738;
assign addr[30453]= 2126796855;
assign addr[30454]= 2100237377;
assign addr[30455]= 2063024031;
assign addr[30456]= 2015345591;
assign addr[30457]= 1957443913;
assign addr[30458]= 1889612716;
assign addr[30459]= 1812196087;
assign addr[30460]= 1725586737;
assign addr[30461]= 1630224009;
assign addr[30462]= 1526591649;
assign addr[30463]= 1415215352;
assign addr[30464]= 1296660098;
assign addr[30465]= 1171527280;
assign addr[30466]= 1040451659;
assign addr[30467]= 904098143;
assign addr[30468]= 763158411;
assign addr[30469]= 618347408;
assign addr[30470]= 470399716;
assign addr[30471]= 320065829;
assign addr[30472]= 168108346;
assign addr[30473]= 15298099;
assign addr[30474]= -137589750;
assign addr[30475]= -289779648;
assign addr[30476]= -440499581;
assign addr[30477]= -588984994;
assign addr[30478]= -734482665;
assign addr[30479]= -876254528;
assign addr[30480]= -1013581418;
assign addr[30481]= -1145766716;
assign addr[30482]= -1272139887;
assign addr[30483]= -1392059879;
assign addr[30484]= -1504918373;
assign addr[30485]= -1610142873;
assign addr[30486]= -1707199606;
assign addr[30487]= -1795596234;
assign addr[30488]= -1874884346;
assign addr[30489]= -1944661739;
assign addr[30490]= -2004574453;
assign addr[30491]= -2054318569;
assign addr[30492]= -2093641749;
assign addr[30493]= -2122344521;
assign addr[30494]= -2140281282;
assign addr[30495]= -2147361045;
assign addr[30496]= -2143547897;
assign addr[30497]= -2128861181;
assign addr[30498]= -2103375398;
assign addr[30499]= -2067219829;
assign addr[30500]= -2020577882;
assign addr[30501]= -1963686155;
assign addr[30502]= -1896833245;
assign addr[30503]= -1820358275;
assign addr[30504]= -1734649179;
assign addr[30505]= -1640140734;
assign addr[30506]= -1537312353;
assign addr[30507]= -1426685652;
assign addr[30508]= -1308821808;
assign addr[30509]= -1184318708;
assign addr[30510]= -1053807919;
assign addr[30511]= -917951481;
assign addr[30512]= -777438554;
assign addr[30513]= -632981917;
assign addr[30514]= -485314355;
assign addr[30515]= -335184940;
assign addr[30516]= -183355234;
assign addr[30517]= -30595422;
assign addr[30518]= 122319591;
assign addr[30519]= 274614114;
assign addr[30520]= 425515602;
assign addr[30521]= 574258580;
assign addr[30522]= 720088517;
assign addr[30523]= 862265664;
assign addr[30524]= 1000068799;
assign addr[30525]= 1132798888;
assign addr[30526]= 1259782632;
assign addr[30527]= 1380375881;
assign addr[30528]= 1493966902;
assign addr[30529]= 1599979481;
assign addr[30530]= 1697875851;
assign addr[30531]= 1787159411;
assign addr[30532]= 1867377253;
assign addr[30533]= 1938122457;
assign addr[30534]= 1999036154;
assign addr[30535]= 2049809346;
assign addr[30536]= 2090184478;
assign addr[30537]= 2119956737;
assign addr[30538]= 2138975100;
assign addr[30539]= 2147143090;
assign addr[30540]= 2144419275;
assign addr[30541]= 2130817471;
assign addr[30542]= 2106406677;
assign addr[30543]= 2071310720;
assign addr[30544]= 2025707632;
assign addr[30545]= 1969828744;
assign addr[30546]= 1903957513;
assign addr[30547]= 1828428082;
assign addr[30548]= 1743623590;
assign addr[30549]= 1649974225;
assign addr[30550]= 1547955041;
assign addr[30551]= 1438083551;
assign addr[30552]= 1320917099;
assign addr[30553]= 1197050035;
assign addr[30554]= 1067110699;
assign addr[30555]= 931758235;
assign addr[30556]= 791679244;
assign addr[30557]= 647584304;
assign addr[30558]= 500204365;
assign addr[30559]= 350287041;
assign addr[30560]= 198592817;
assign addr[30561]= 45891193;
assign addr[30562]= -107043224;
assign addr[30563]= -259434643;
assign addr[30564]= -410510029;
assign addr[30565]= -559503022;
assign addr[30566]= -705657826;
assign addr[30567]= -848233042;
assign addr[30568]= -986505429;
assign addr[30569]= -1119773573;
assign addr[30570]= -1247361445;
assign addr[30571]= -1368621831;
assign addr[30572]= -1482939614;
assign addr[30573]= -1589734894;
assign addr[30574]= -1688465931;
assign addr[30575]= -1778631892;
assign addr[30576]= -1859775393;
assign addr[30577]= -1931484818;
assign addr[30578]= -1993396407;
assign addr[30579]= -2045196100;
assign addr[30580]= -2086621133;
assign addr[30581]= -2117461370;
assign addr[30582]= -2137560369;
assign addr[30583]= -2146816171;
assign addr[30584]= -2145181827;
assign addr[30585]= -2132665626;
assign addr[30586]= -2109331059;
assign addr[30587]= -2075296495;
assign addr[30588]= -2030734582;
assign addr[30589]= -1975871368;
assign addr[30590]= -1910985158;
assign addr[30591]= -1836405100;
assign addr[30592]= -1752509516;
assign addr[30593]= -1659723983;
assign addr[30594]= -1558519173;
assign addr[30595]= -1449408469;
assign addr[30596]= -1332945355;
assign addr[30597]= -1209720613;
assign addr[30598]= -1080359326;
assign addr[30599]= -945517704;
assign addr[30600]= -805879757;
assign addr[30601]= -662153826;
assign addr[30602]= -515068990;
assign addr[30603]= -365371365;
assign addr[30604]= -213820322;
assign addr[30605]= -61184634;
assign addr[30606]= 91761426;
assign addr[30607]= 244242007;
assign addr[30608]= 395483624;
assign addr[30609]= 544719071;
assign addr[30610]= 691191324;
assign addr[30611]= 834157373;
assign addr[30612]= 972891995;
assign addr[30613]= 1106691431;
assign addr[30614]= 1234876957;
assign addr[30615]= 1356798326;
assign addr[30616]= 1471837070;
assign addr[30617]= 1579409630;
assign addr[30618]= 1678970324;
assign addr[30619]= 1770014111;
assign addr[30620]= 1852079154;
assign addr[30621]= 1924749160;
assign addr[30622]= 1987655498;
assign addr[30623]= 2040479063;
assign addr[30624]= 2082951896;
assign addr[30625]= 2114858546;
assign addr[30626]= 2136037160;
assign addr[30627]= 2146380306;
assign addr[30628]= 2145835515;
assign addr[30629]= 2134405552;
assign addr[30630]= 2112148396;
assign addr[30631]= 2079176953;
assign addr[30632]= 2035658475;
assign addr[30633]= 1981813720;
assign addr[30634]= 1917915825;
assign addr[30635]= 1844288924;
assign addr[30636]= 1761306505;
assign addr[30637]= 1669389513;
assign addr[30638]= 1569004214;
assign addr[30639]= 1460659832;
assign addr[30640]= 1344905966;
assign addr[30641]= 1222329801;
assign addr[30642]= 1093553126;
assign addr[30643]= 959229189;
assign addr[30644]= 820039373;
assign addr[30645]= 676689746;
assign addr[30646]= 529907477;
assign addr[30647]= 380437148;
assign addr[30648]= 229036977;
assign addr[30649]= 76474970;
assign addr[30650]= -76474970;
assign addr[30651]= -229036977;
assign addr[30652]= -380437148;
assign addr[30653]= -529907477;
assign addr[30654]= -676689746;
assign addr[30655]= -820039373;
assign addr[30656]= -959229189;
assign addr[30657]= -1093553126;
assign addr[30658]= -1222329801;
assign addr[30659]= -1344905966;
assign addr[30660]= -1460659832;
assign addr[30661]= -1569004214;
assign addr[30662]= -1669389513;
assign addr[30663]= -1761306505;
assign addr[30664]= -1844288924;
assign addr[30665]= -1917915825;
assign addr[30666]= -1981813720;
assign addr[30667]= -2035658475;
assign addr[30668]= -2079176953;
assign addr[30669]= -2112148396;
assign addr[30670]= -2134405552;
assign addr[30671]= -2145835515;
assign addr[30672]= -2146380306;
assign addr[30673]= -2136037160;
assign addr[30674]= -2114858546;
assign addr[30675]= -2082951896;
assign addr[30676]= -2040479063;
assign addr[30677]= -1987655498;
assign addr[30678]= -1924749160;
assign addr[30679]= -1852079154;
assign addr[30680]= -1770014111;
assign addr[30681]= -1678970324;
assign addr[30682]= -1579409630;
assign addr[30683]= -1471837070;
assign addr[30684]= -1356798326;
assign addr[30685]= -1234876957;
assign addr[30686]= -1106691431;
assign addr[30687]= -972891995;
assign addr[30688]= -834157373;
assign addr[30689]= -691191324;
assign addr[30690]= -544719071;
assign addr[30691]= -395483624;
assign addr[30692]= -244242007;
assign addr[30693]= -91761426;
assign addr[30694]= 61184634;
assign addr[30695]= 213820322;
assign addr[30696]= 365371365;
assign addr[30697]= 515068990;
assign addr[30698]= 662153826;
assign addr[30699]= 805879757;
assign addr[30700]= 945517704;
assign addr[30701]= 1080359326;
assign addr[30702]= 1209720613;
assign addr[30703]= 1332945355;
assign addr[30704]= 1449408469;
assign addr[30705]= 1558519173;
assign addr[30706]= 1659723983;
assign addr[30707]= 1752509516;
assign addr[30708]= 1836405100;
assign addr[30709]= 1910985158;
assign addr[30710]= 1975871368;
assign addr[30711]= 2030734582;
assign addr[30712]= 2075296495;
assign addr[30713]= 2109331059;
assign addr[30714]= 2132665626;
assign addr[30715]= 2145181827;
assign addr[30716]= 2146816171;
assign addr[30717]= 2137560369;
assign addr[30718]= 2117461370;
assign addr[30719]= 2086621133;
assign addr[30720]= 2045196100;
assign addr[30721]= 1993396407;
assign addr[30722]= 1931484818;
assign addr[30723]= 1859775393;
assign addr[30724]= 1778631892;
assign addr[30725]= 1688465931;
assign addr[30726]= 1589734894;
assign addr[30727]= 1482939614;
assign addr[30728]= 1368621831;
assign addr[30729]= 1247361445;
assign addr[30730]= 1119773573;
assign addr[30731]= 986505429;
assign addr[30732]= 848233042;
assign addr[30733]= 705657826;
assign addr[30734]= 559503022;
assign addr[30735]= 410510029;
assign addr[30736]= 259434643;
assign addr[30737]= 107043224;
assign addr[30738]= -45891193;
assign addr[30739]= -198592817;
assign addr[30740]= -350287041;
assign addr[30741]= -500204365;
assign addr[30742]= -647584304;
assign addr[30743]= -791679244;
assign addr[30744]= -931758235;
assign addr[30745]= -1067110699;
assign addr[30746]= -1197050035;
assign addr[30747]= -1320917099;
assign addr[30748]= -1438083551;
assign addr[30749]= -1547955041;
assign addr[30750]= -1649974225;
assign addr[30751]= -1743623590;
assign addr[30752]= -1828428082;
assign addr[30753]= -1903957513;
assign addr[30754]= -1969828744;
assign addr[30755]= -2025707632;
assign addr[30756]= -2071310720;
assign addr[30757]= -2106406677;
assign addr[30758]= -2130817471;
assign addr[30759]= -2144419275;
assign addr[30760]= -2147143090;
assign addr[30761]= -2138975100;
assign addr[30762]= -2119956737;
assign addr[30763]= -2090184478;
assign addr[30764]= -2049809346;
assign addr[30765]= -1999036154;
assign addr[30766]= -1938122457;
assign addr[30767]= -1867377253;
assign addr[30768]= -1787159411;
assign addr[30769]= -1697875851;
assign addr[30770]= -1599979481;
assign addr[30771]= -1493966902;
assign addr[30772]= -1380375881;
assign addr[30773]= -1259782632;
assign addr[30774]= -1132798888;
assign addr[30775]= -1000068799;
assign addr[30776]= -862265664;
assign addr[30777]= -720088517;
assign addr[30778]= -574258580;
assign addr[30779]= -425515602;
assign addr[30780]= -274614114;
assign addr[30781]= -122319591;
assign addr[30782]= 30595422;
assign addr[30783]= 183355234;
assign addr[30784]= 335184940;
assign addr[30785]= 485314355;
assign addr[30786]= 632981917;
assign addr[30787]= 777438554;
assign addr[30788]= 917951481;
assign addr[30789]= 1053807919;
assign addr[30790]= 1184318708;
assign addr[30791]= 1308821808;
assign addr[30792]= 1426685652;
assign addr[30793]= 1537312353;
assign addr[30794]= 1640140734;
assign addr[30795]= 1734649179;
assign addr[30796]= 1820358275;
assign addr[30797]= 1896833245;
assign addr[30798]= 1963686155;
assign addr[30799]= 2020577882;
assign addr[30800]= 2067219829;
assign addr[30801]= 2103375398;
assign addr[30802]= 2128861181;
assign addr[30803]= 2143547897;
assign addr[30804]= 2147361045;
assign addr[30805]= 2140281282;
assign addr[30806]= 2122344521;
assign addr[30807]= 2093641749;
assign addr[30808]= 2054318569;
assign addr[30809]= 2004574453;
assign addr[30810]= 1944661739;
assign addr[30811]= 1874884346;
assign addr[30812]= 1795596234;
assign addr[30813]= 1707199606;
assign addr[30814]= 1610142873;
assign addr[30815]= 1504918373;
assign addr[30816]= 1392059879;
assign addr[30817]= 1272139887;
assign addr[30818]= 1145766716;
assign addr[30819]= 1013581418;
assign addr[30820]= 876254528;
assign addr[30821]= 734482665;
assign addr[30822]= 588984994;
assign addr[30823]= 440499581;
assign addr[30824]= 289779648;
assign addr[30825]= 137589750;
assign addr[30826]= -15298099;
assign addr[30827]= -168108346;
assign addr[30828]= -320065829;
assign addr[30829]= -470399716;
assign addr[30830]= -618347408;
assign addr[30831]= -763158411;
assign addr[30832]= -904098143;
assign addr[30833]= -1040451659;
assign addr[30834]= -1171527280;
assign addr[30835]= -1296660098;
assign addr[30836]= -1415215352;
assign addr[30837]= -1526591649;
assign addr[30838]= -1630224009;
assign addr[30839]= -1725586737;
assign addr[30840]= -1812196087;
assign addr[30841]= -1889612716;
assign addr[30842]= -1957443913;
assign addr[30843]= -2015345591;
assign addr[30844]= -2063024031;
assign addr[30845]= -2100237377;
assign addr[30846]= -2126796855;
assign addr[30847]= -2142567738;
assign addr[30848]= -2147470025;
assign addr[30849]= -2141478848;
assign addr[30850]= -2124624598;
assign addr[30851]= -2096992772;
assign addr[30852]= -2058723538;
assign addr[30853]= -2010011024;
assign addr[30854]= -1951102334;
assign addr[30855]= -1882296293;
assign addr[30856]= -1803941934;
assign addr[30857]= -1716436725;
assign addr[30858]= -1620224553;
assign addr[30859]= -1515793473;
assign addr[30860]= -1403673233;
assign addr[30861]= -1284432584;
assign addr[30862]= -1158676398;
assign addr[30863]= -1027042599;
assign addr[30864]= -890198924;
assign addr[30865]= -748839539;
assign addr[30866]= -603681519;
assign addr[30867]= -455461206;
assign addr[30868]= -304930476;
assign addr[30869]= -152852926;
assign addr[30870]= 0;
assign addr[30871]= 152852926;
assign addr[30872]= 304930476;
assign addr[30873]= 455461206;
assign addr[30874]= 603681519;
assign addr[30875]= 748839539;
assign addr[30876]= 890198924;
assign addr[30877]= 1027042599;
assign addr[30878]= 1158676398;
assign addr[30879]= 1284432584;
assign addr[30880]= 1403673233;
assign addr[30881]= 1515793473;
assign addr[30882]= 1620224553;
assign addr[30883]= 1716436725;
assign addr[30884]= 1803941934;
assign addr[30885]= 1882296293;
assign addr[30886]= 1951102334;
assign addr[30887]= 2010011024;
assign addr[30888]= 2058723538;
assign addr[30889]= 2096992772;
assign addr[30890]= 2124624598;
assign addr[30891]= 2141478848;
assign addr[30892]= 2147470025;
assign addr[30893]= 2142567738;
assign addr[30894]= 2126796855;
assign addr[30895]= 2100237377;
assign addr[30896]= 2063024031;
assign addr[30897]= 2015345591;
assign addr[30898]= 1957443913;
assign addr[30899]= 1889612716;
assign addr[30900]= 1812196087;
assign addr[30901]= 1725586737;
assign addr[30902]= 1630224009;
assign addr[30903]= 1526591649;
assign addr[30904]= 1415215352;
assign addr[30905]= 1296660098;
assign addr[30906]= 1171527280;
assign addr[30907]= 1040451659;
assign addr[30908]= 904098143;
assign addr[30909]= 763158411;
assign addr[30910]= 618347408;
assign addr[30911]= 470399716;
assign addr[30912]= 320065829;
assign addr[30913]= 168108346;
assign addr[30914]= 15298099;
assign addr[30915]= -137589750;
assign addr[30916]= -289779648;
assign addr[30917]= -440499581;
assign addr[30918]= -588984994;
assign addr[30919]= -734482665;
assign addr[30920]= -876254528;
assign addr[30921]= -1013581418;
assign addr[30922]= -1145766716;
assign addr[30923]= -1272139887;
assign addr[30924]= -1392059879;
assign addr[30925]= -1504918373;
assign addr[30926]= -1610142873;
assign addr[30927]= -1707199606;
assign addr[30928]= -1795596234;
assign addr[30929]= -1874884346;
assign addr[30930]= -1944661739;
assign addr[30931]= -2004574453;
assign addr[30932]= -2054318569;
assign addr[30933]= -2093641749;
assign addr[30934]= -2122344521;
assign addr[30935]= -2140281282;
assign addr[30936]= -2147361045;
assign addr[30937]= -2143547897;
assign addr[30938]= -2128861181;
assign addr[30939]= -2103375398;
assign addr[30940]= -2067219829;
assign addr[30941]= -2020577882;
assign addr[30942]= -1963686155;
assign addr[30943]= -1896833245;
assign addr[30944]= -1820358275;
assign addr[30945]= -1734649179;
assign addr[30946]= -1640140734;
assign addr[30947]= -1537312353;
assign addr[30948]= -1426685652;
assign addr[30949]= -1308821808;
assign addr[30950]= -1184318708;
assign addr[30951]= -1053807919;
assign addr[30952]= -917951481;
assign addr[30953]= -777438554;
assign addr[30954]= -632981917;
assign addr[30955]= -485314355;
assign addr[30956]= -335184940;
assign addr[30957]= -183355234;
assign addr[30958]= -30595422;
assign addr[30959]= 122319591;
assign addr[30960]= 274614114;
assign addr[30961]= 425515602;
assign addr[30962]= 574258580;
assign addr[30963]= 720088517;
assign addr[30964]= 862265664;
assign addr[30965]= 1000068799;
assign addr[30966]= 1132798888;
assign addr[30967]= 1259782632;
assign addr[30968]= 1380375881;
assign addr[30969]= 1493966902;
assign addr[30970]= 1599979481;
assign addr[30971]= 1697875851;
assign addr[30972]= 1787159411;
assign addr[30973]= 1867377253;
assign addr[30974]= 1938122457;
assign addr[30975]= 1999036154;
assign addr[30976]= 2049809346;
assign addr[30977]= 2090184478;
assign addr[30978]= 2119956737;
assign addr[30979]= 2138975100;
assign addr[30980]= 2147143090;
assign addr[30981]= 2144419275;
assign addr[30982]= 2130817471;
assign addr[30983]= 2106406677;
assign addr[30984]= 2071310720;
assign addr[30985]= 2025707632;
assign addr[30986]= 1969828744;
assign addr[30987]= 1903957513;
assign addr[30988]= 1828428082;
assign addr[30989]= 1743623590;
assign addr[30990]= 1649974225;
assign addr[30991]= 1547955041;
assign addr[30992]= 1438083551;
assign addr[30993]= 1320917099;
assign addr[30994]= 1197050035;
assign addr[30995]= 1067110699;
assign addr[30996]= 931758235;
assign addr[30997]= 791679244;
assign addr[30998]= 647584304;
assign addr[30999]= 500204365;
assign addr[31000]= 350287041;
assign addr[31001]= 198592817;
assign addr[31002]= 45891193;
assign addr[31003]= -107043224;
assign addr[31004]= -259434643;
assign addr[31005]= -410510029;
assign addr[31006]= -559503022;
assign addr[31007]= -705657826;
assign addr[31008]= -848233042;
assign addr[31009]= -986505429;
assign addr[31010]= -1119773573;
assign addr[31011]= -1247361445;
assign addr[31012]= -1368621831;
assign addr[31013]= -1482939614;
assign addr[31014]= -1589734894;
assign addr[31015]= -1688465931;
assign addr[31016]= -1778631892;
assign addr[31017]= -1859775393;
assign addr[31018]= -1931484818;
assign addr[31019]= -1993396407;
assign addr[31020]= -2045196100;
assign addr[31021]= -2086621133;
assign addr[31022]= -2117461370;
assign addr[31023]= -2137560369;
assign addr[31024]= -2146816171;
assign addr[31025]= -2145181827;
assign addr[31026]= -2132665626;
assign addr[31027]= -2109331059;
assign addr[31028]= -2075296495;
assign addr[31029]= -2030734582;
assign addr[31030]= -1975871368;
assign addr[31031]= -1910985158;
assign addr[31032]= -1836405100;
assign addr[31033]= -1752509516;
assign addr[31034]= -1659723983;
assign addr[31035]= -1558519173;
assign addr[31036]= -1449408469;
assign addr[31037]= -1332945355;
assign addr[31038]= -1209720613;
assign addr[31039]= -1080359326;
assign addr[31040]= -945517704;
assign addr[31041]= -805879757;
assign addr[31042]= -662153826;
assign addr[31043]= -515068990;
assign addr[31044]= -365371365;
assign addr[31045]= -213820322;
assign addr[31046]= -61184634;
assign addr[31047]= 91761426;
assign addr[31048]= 244242007;
assign addr[31049]= 395483624;
assign addr[31050]= 544719071;
assign addr[31051]= 691191324;
assign addr[31052]= 834157373;
assign addr[31053]= 972891995;
assign addr[31054]= 1106691431;
assign addr[31055]= 1234876957;
assign addr[31056]= 1356798326;
assign addr[31057]= 1471837070;
assign addr[31058]= 1579409630;
assign addr[31059]= 1678970324;
assign addr[31060]= 1770014111;
assign addr[31061]= 1852079154;
assign addr[31062]= 1924749160;
assign addr[31063]= 1987655498;
assign addr[31064]= 2040479063;
assign addr[31065]= 2082951896;
assign addr[31066]= 2114858546;
assign addr[31067]= 2136037160;
assign addr[31068]= 2146380306;
assign addr[31069]= 2145835515;
assign addr[31070]= 2134405552;
assign addr[31071]= 2112148396;
assign addr[31072]= 2079176953;
assign addr[31073]= 2035658475;
assign addr[31074]= 1981813720;
assign addr[31075]= 1917915825;
assign addr[31076]= 1844288924;
assign addr[31077]= 1761306505;
assign addr[31078]= 1669389513;
assign addr[31079]= 1569004214;
assign addr[31080]= 1460659832;
assign addr[31081]= 1344905966;
assign addr[31082]= 1222329801;
assign addr[31083]= 1093553126;
assign addr[31084]= 959229189;
assign addr[31085]= 820039373;
assign addr[31086]= 676689746;
assign addr[31087]= 529907477;
assign addr[31088]= 380437148;
assign addr[31089]= 229036977;
assign addr[31090]= 76474970;
assign addr[31091]= -76474970;
assign addr[31092]= -229036977;
assign addr[31093]= -380437148;
assign addr[31094]= -529907477;
assign addr[31095]= -676689746;
assign addr[31096]= -820039373;
assign addr[31097]= -959229189;
assign addr[31098]= -1093553126;
assign addr[31099]= -1222329801;
assign addr[31100]= -1344905966;
assign addr[31101]= -1460659832;
assign addr[31102]= -1569004214;
assign addr[31103]= -1669389513;
assign addr[31104]= -1761306505;
assign addr[31105]= -1844288924;
assign addr[31106]= -1917915825;
assign addr[31107]= -1981813720;
assign addr[31108]= -2035658475;
assign addr[31109]= -2079176953;
assign addr[31110]= -2112148396;
assign addr[31111]= -2134405552;
assign addr[31112]= -2145835515;
assign addr[31113]= -2146380306;
assign addr[31114]= -2136037160;
assign addr[31115]= -2114858546;
assign addr[31116]= -2082951896;
assign addr[31117]= -2040479063;
assign addr[31118]= -1987655498;
assign addr[31119]= -1924749160;
assign addr[31120]= -1852079154;
assign addr[31121]= -1770014111;
assign addr[31122]= -1678970324;
assign addr[31123]= -1579409630;
assign addr[31124]= -1471837070;
assign addr[31125]= -1356798326;
assign addr[31126]= -1234876957;
assign addr[31127]= -1106691431;
assign addr[31128]= -972891995;
assign addr[31129]= -834157373;
assign addr[31130]= -691191324;
assign addr[31131]= -544719071;
assign addr[31132]= -395483624;
assign addr[31133]= -244242007;
assign addr[31134]= -91761426;
assign addr[31135]= 61184634;
assign addr[31136]= 213820322;
assign addr[31137]= 365371365;
assign addr[31138]= 515068990;
assign addr[31139]= 662153826;
assign addr[31140]= 805879757;
assign addr[31141]= 945517704;
assign addr[31142]= 1080359326;
assign addr[31143]= 1209720613;
assign addr[31144]= 1332945355;
assign addr[31145]= 1449408469;
assign addr[31146]= 1558519173;
assign addr[31147]= 1659723983;
assign addr[31148]= 1752509516;
assign addr[31149]= 1836405100;
assign addr[31150]= 1910985158;
assign addr[31151]= 1975871368;
assign addr[31152]= 2030734582;
assign addr[31153]= 2075296495;
assign addr[31154]= 2109331059;
assign addr[31155]= 2132665626;
assign addr[31156]= 2145181827;
assign addr[31157]= 2146816171;
assign addr[31158]= 2137560369;
assign addr[31159]= 2117461370;
assign addr[31160]= 2086621133;
assign addr[31161]= 2045196100;
assign addr[31162]= 1993396407;
assign addr[31163]= 1931484818;
assign addr[31164]= 1859775393;
assign addr[31165]= 1778631892;
assign addr[31166]= 1688465931;
assign addr[31167]= 1589734894;
assign addr[31168]= 1482939614;
assign addr[31169]= 1368621831;
assign addr[31170]= 1247361445;
assign addr[31171]= 1119773573;
assign addr[31172]= 986505429;
assign addr[31173]= 848233042;
assign addr[31174]= 705657826;
assign addr[31175]= 559503022;
assign addr[31176]= 410510029;
assign addr[31177]= 259434643;
assign addr[31178]= 107043224;
assign addr[31179]= -45891193;
assign addr[31180]= -198592817;
assign addr[31181]= -350287041;
assign addr[31182]= -500204365;
assign addr[31183]= -647584304;
assign addr[31184]= -791679244;
assign addr[31185]= -931758235;
assign addr[31186]= -1067110699;
assign addr[31187]= -1197050035;
assign addr[31188]= -1320917099;
assign addr[31189]= -1438083551;
assign addr[31190]= -1547955041;
assign addr[31191]= -1649974225;
assign addr[31192]= -1743623590;
assign addr[31193]= -1828428082;
assign addr[31194]= -1903957513;
assign addr[31195]= -1969828744;
assign addr[31196]= -2025707632;
assign addr[31197]= -2071310720;
assign addr[31198]= -2106406677;
assign addr[31199]= -2130817471;
assign addr[31200]= -2144419275;
assign addr[31201]= -2147143090;
assign addr[31202]= -2138975100;
assign addr[31203]= -2119956737;
assign addr[31204]= -2090184478;
assign addr[31205]= -2049809346;
assign addr[31206]= -1999036154;
assign addr[31207]= -1938122457;
assign addr[31208]= -1867377253;
assign addr[31209]= -1787159411;
assign addr[31210]= -1697875851;
assign addr[31211]= -1599979481;
assign addr[31212]= -1493966902;
assign addr[31213]= -1380375881;
assign addr[31214]= -1259782632;
assign addr[31215]= -1132798888;
assign addr[31216]= -1000068799;
assign addr[31217]= -862265664;
assign addr[31218]= -720088517;
assign addr[31219]= -574258580;
assign addr[31220]= -425515602;
assign addr[31221]= -274614114;
assign addr[31222]= -122319591;
assign addr[31223]= 30595422;
assign addr[31224]= 183355234;
assign addr[31225]= 335184940;
assign addr[31226]= 485314355;
assign addr[31227]= 632981917;
assign addr[31228]= 777438554;
assign addr[31229]= 917951481;
assign addr[31230]= 1053807919;
assign addr[31231]= 1184318708;
assign addr[31232]= 1308821808;
assign addr[31233]= 1426685652;
assign addr[31234]= 1537312353;
assign addr[31235]= 1640140734;
assign addr[31236]= 1734649179;
assign addr[31237]= 1820358275;
assign addr[31238]= 1896833245;
assign addr[31239]= 1963686155;
assign addr[31240]= 2020577882;
assign addr[31241]= 2067219829;
assign addr[31242]= 2103375398;
assign addr[31243]= 2128861181;
assign addr[31244]= 2143547897;
assign addr[31245]= 2147361045;
assign addr[31246]= 2140281282;
assign addr[31247]= 2122344521;
assign addr[31248]= 2093641749;
assign addr[31249]= 2054318569;
assign addr[31250]= 2004574453;
assign addr[31251]= 1944661739;
assign addr[31252]= 1874884346;
assign addr[31253]= 1795596234;
assign addr[31254]= 1707199606;
assign addr[31255]= 1610142873;
assign addr[31256]= 1504918373;
assign addr[31257]= 1392059879;
assign addr[31258]= 1272139887;
assign addr[31259]= 1145766716;
assign addr[31260]= 1013581418;
assign addr[31261]= 876254528;
assign addr[31262]= 734482665;
assign addr[31263]= 588984994;
assign addr[31264]= 440499581;
assign addr[31265]= 289779648;
assign addr[31266]= 137589750;
assign addr[31267]= -15298099;
assign addr[31268]= -168108346;
assign addr[31269]= -320065829;
assign addr[31270]= -470399716;
assign addr[31271]= -618347408;
assign addr[31272]= -763158411;
assign addr[31273]= -904098143;
assign addr[31274]= -1040451659;
assign addr[31275]= -1171527280;
assign addr[31276]= -1296660098;
assign addr[31277]= -1415215352;
assign addr[31278]= -1526591649;
assign addr[31279]= -1630224009;
assign addr[31280]= -1725586737;
assign addr[31281]= -1812196087;
assign addr[31282]= -1889612716;
assign addr[31283]= -1957443913;
assign addr[31284]= -2015345591;
assign addr[31285]= -2063024031;
assign addr[31286]= -2100237377;
assign addr[31287]= -2126796855;
assign addr[31288]= -2142567738;
assign addr[31289]= -2147470025;
assign addr[31290]= -2141478848;
assign addr[31291]= -2124624598;
assign addr[31292]= -2096992772;
assign addr[31293]= -2058723538;
assign addr[31294]= -2010011024;
assign addr[31295]= -1951102334;
assign addr[31296]= -1882296293;
assign addr[31297]= -1803941934;
assign addr[31298]= -1716436725;
assign addr[31299]= -1620224553;
assign addr[31300]= -1515793473;
assign addr[31301]= -1403673233;
assign addr[31302]= -1284432584;
assign addr[31303]= -1158676398;
assign addr[31304]= -1027042599;
assign addr[31305]= -890198924;
assign addr[31306]= -748839539;
assign addr[31307]= -603681519;
assign addr[31308]= -455461206;
assign addr[31309]= -304930476;
assign addr[31310]= -152852926;
assign addr[31311]= 0;
assign addr[31312]= 152852926;
assign addr[31313]= 304930476;
assign addr[31314]= 455461206;
assign addr[31315]= 603681519;
assign addr[31316]= 748839539;
assign addr[31317]= 890198924;
assign addr[31318]= 1027042599;
assign addr[31319]= 1158676398;
assign addr[31320]= 1284432584;
assign addr[31321]= 1403673233;
assign addr[31322]= 1515793473;
assign addr[31323]= 1620224553;
assign addr[31324]= 1716436725;
assign addr[31325]= 1803941934;
assign addr[31326]= 1882296293;
assign addr[31327]= 1951102334;
assign addr[31328]= 2010011024;
assign addr[31329]= 2058723538;
assign addr[31330]= 2096992772;
assign addr[31331]= 2124624598;
assign addr[31332]= 2141478848;
assign addr[31333]= 2147470025;
assign addr[31334]= 2142567738;
assign addr[31335]= 2126796855;
assign addr[31336]= 2100237377;
assign addr[31337]= 2063024031;
assign addr[31338]= 2015345591;
assign addr[31339]= 1957443913;
assign addr[31340]= 1889612716;
assign addr[31341]= 1812196087;
assign addr[31342]= 1725586737;
assign addr[31343]= 1630224009;
assign addr[31344]= 1526591649;
assign addr[31345]= 1415215352;
assign addr[31346]= 1296660098;
assign addr[31347]= 1171527280;
assign addr[31348]= 1040451659;
assign addr[31349]= 904098143;
assign addr[31350]= 763158411;
assign addr[31351]= 618347408;
assign addr[31352]= 470399716;
assign addr[31353]= 320065829;
assign addr[31354]= 168108346;
assign addr[31355]= 15298099;
assign addr[31356]= -137589750;
assign addr[31357]= -289779648;
assign addr[31358]= -440499581;
assign addr[31359]= -588984994;
assign addr[31360]= -734482665;
assign addr[31361]= -876254528;
assign addr[31362]= -1013581418;
assign addr[31363]= -1145766716;
assign addr[31364]= -1272139887;
assign addr[31365]= -1392059879;
assign addr[31366]= -1504918373;
assign addr[31367]= -1610142873;
assign addr[31368]= -1707199606;
assign addr[31369]= -1795596234;
assign addr[31370]= -1874884346;
assign addr[31371]= -1944661739;
assign addr[31372]= -2004574453;
assign addr[31373]= -2054318569;
assign addr[31374]= -2093641749;
assign addr[31375]= -2122344521;
assign addr[31376]= -2140281282;
assign addr[31377]= -2147361045;
assign addr[31378]= -2143547897;
assign addr[31379]= -2128861181;
assign addr[31380]= -2103375398;
assign addr[31381]= -2067219829;
assign addr[31382]= -2020577882;
assign addr[31383]= -1963686155;
assign addr[31384]= -1896833245;
assign addr[31385]= -1820358275;
assign addr[31386]= -1734649179;
assign addr[31387]= -1640140734;
assign addr[31388]= -1537312353;
assign addr[31389]= -1426685652;
assign addr[31390]= -1308821808;
assign addr[31391]= -1184318708;
assign addr[31392]= -1053807919;
assign addr[31393]= -917951481;
assign addr[31394]= -777438554;
assign addr[31395]= -632981917;
assign addr[31396]= -485314355;
assign addr[31397]= -335184940;
assign addr[31398]= -183355234;
assign addr[31399]= -30595422;
assign addr[31400]= 122319591;
assign addr[31401]= 274614114;
assign addr[31402]= 425515602;
assign addr[31403]= 574258580;
assign addr[31404]= 720088517;
assign addr[31405]= 862265664;
assign addr[31406]= 1000068799;
assign addr[31407]= 1132798888;
assign addr[31408]= 1259782632;
assign addr[31409]= 1380375881;
assign addr[31410]= 1493966902;
assign addr[31411]= 1599979481;
assign addr[31412]= 1697875851;
assign addr[31413]= 1787159411;
assign addr[31414]= 1867377253;
assign addr[31415]= 1938122457;
assign addr[31416]= 1999036154;
assign addr[31417]= 2049809346;
assign addr[31418]= 2090184478;
assign addr[31419]= 2119956737;
assign addr[31420]= 2138975100;
assign addr[31421]= 2147143090;
assign addr[31422]= 2144419275;
assign addr[31423]= 2130817471;
assign addr[31424]= 2106406677;
assign addr[31425]= 2071310720;
assign addr[31426]= 2025707632;
assign addr[31427]= 1969828744;
assign addr[31428]= 1903957513;
assign addr[31429]= 1828428082;
assign addr[31430]= 1743623590;
assign addr[31431]= 1649974225;
assign addr[31432]= 1547955041;
assign addr[31433]= 1438083551;
assign addr[31434]= 1320917099;
assign addr[31435]= 1197050035;
assign addr[31436]= 1067110699;
assign addr[31437]= 931758235;
assign addr[31438]= 791679244;
assign addr[31439]= 647584304;
assign addr[31440]= 500204365;
assign addr[31441]= 350287041;
assign addr[31442]= 198592817;
assign addr[31443]= 45891193;
assign addr[31444]= -107043224;
assign addr[31445]= -259434643;
assign addr[31446]= -410510029;
assign addr[31447]= -559503022;
assign addr[31448]= -705657826;
assign addr[31449]= -848233042;
assign addr[31450]= -986505429;
assign addr[31451]= -1119773573;
assign addr[31452]= -1247361445;
assign addr[31453]= -1368621831;
assign addr[31454]= -1482939614;
assign addr[31455]= -1589734894;
assign addr[31456]= -1688465931;
assign addr[31457]= -1778631892;
assign addr[31458]= -1859775393;
assign addr[31459]= -1931484818;
assign addr[31460]= -1993396407;
assign addr[31461]= -2045196100;
assign addr[31462]= -2086621133;
assign addr[31463]= -2117461370;
assign addr[31464]= -2137560369;
assign addr[31465]= -2146816171;
assign addr[31466]= -2145181827;
assign addr[31467]= -2132665626;
assign addr[31468]= -2109331059;
assign addr[31469]= -2075296495;
assign addr[31470]= -2030734582;
assign addr[31471]= -1975871368;
assign addr[31472]= -1910985158;
assign addr[31473]= -1836405100;
assign addr[31474]= -1752509516;
assign addr[31475]= -1659723983;
assign addr[31476]= -1558519173;
assign addr[31477]= -1449408469;
assign addr[31478]= -1332945355;
assign addr[31479]= -1209720613;
assign addr[31480]= -1080359326;
assign addr[31481]= -945517704;
assign addr[31482]= -805879757;
assign addr[31483]= -662153826;
assign addr[31484]= -515068990;
assign addr[31485]= -365371365;
assign addr[31486]= -213820322;
assign addr[31487]= -61184634;
assign addr[31488]= 91761426;
assign addr[31489]= 244242007;
assign addr[31490]= 395483624;
assign addr[31491]= 544719071;
assign addr[31492]= 691191324;
assign addr[31493]= 834157373;
assign addr[31494]= 972891995;
assign addr[31495]= 1106691431;
assign addr[31496]= 1234876957;
assign addr[31497]= 1356798326;
assign addr[31498]= 1471837070;
assign addr[31499]= 1579409630;
assign addr[31500]= 1678970324;
assign addr[31501]= 1770014111;
assign addr[31502]= 1852079154;
assign addr[31503]= 1924749160;
assign addr[31504]= 1987655498;
assign addr[31505]= 2040479063;
assign addr[31506]= 2082951896;
assign addr[31507]= 2114858546;
assign addr[31508]= 2136037160;
assign addr[31509]= 2146380306;
assign addr[31510]= 2145835515;
assign addr[31511]= 2134405552;
assign addr[31512]= 2112148396;
assign addr[31513]= 2079176953;
assign addr[31514]= 2035658475;
assign addr[31515]= 1981813720;
assign addr[31516]= 1917915825;
assign addr[31517]= 1844288924;
assign addr[31518]= 1761306505;
assign addr[31519]= 1669389513;
assign addr[31520]= 1569004214;
assign addr[31521]= 1460659832;
assign addr[31522]= 1344905966;
assign addr[31523]= 1222329801;
assign addr[31524]= 1093553126;
assign addr[31525]= 959229189;
assign addr[31526]= 820039373;
assign addr[31527]= 676689746;
assign addr[31528]= 529907477;
assign addr[31529]= 380437148;
assign addr[31530]= 229036977;
assign addr[31531]= 76474970;
assign addr[31532]= -76474970;
assign addr[31533]= -229036977;
assign addr[31534]= -380437148;
assign addr[31535]= -529907477;
assign addr[31536]= -676689746;
assign addr[31537]= -820039373;
assign addr[31538]= -959229189;
assign addr[31539]= -1093553126;
assign addr[31540]= -1222329801;
assign addr[31541]= -1344905966;
assign addr[31542]= -1460659832;
assign addr[31543]= -1569004214;
assign addr[31544]= -1669389513;
assign addr[31545]= -1761306505;
assign addr[31546]= -1844288924;
assign addr[31547]= -1917915825;
assign addr[31548]= -1981813720;
assign addr[31549]= -2035658475;
assign addr[31550]= -2079176953;
assign addr[31551]= -2112148396;
assign addr[31552]= -2134405552;
assign addr[31553]= -2145835515;
assign addr[31554]= -2146380306;
assign addr[31555]= -2136037160;
assign addr[31556]= -2114858546;
assign addr[31557]= -2082951896;
assign addr[31558]= -2040479063;
assign addr[31559]= -1987655498;
assign addr[31560]= -1924749160;
assign addr[31561]= -1852079154;
assign addr[31562]= -1770014111;
assign addr[31563]= -1678970324;
assign addr[31564]= -1579409630;
assign addr[31565]= -1471837070;
assign addr[31566]= -1356798326;
assign addr[31567]= -1234876957;
assign addr[31568]= -1106691431;
assign addr[31569]= -972891995;
assign addr[31570]= -834157373;
assign addr[31571]= -691191324;
assign addr[31572]= -544719071;
assign addr[31573]= -395483624;
assign addr[31574]= -244242007;
assign addr[31575]= -91761426;
assign addr[31576]= 61184634;
assign addr[31577]= 213820322;
assign addr[31578]= 365371365;
assign addr[31579]= 515068990;
assign addr[31580]= 662153826;
assign addr[31581]= 805879757;
assign addr[31582]= 945517704;
assign addr[31583]= 1080359326;
assign addr[31584]= 1209720613;
assign addr[31585]= 1332945355;
assign addr[31586]= 1449408469;
assign addr[31587]= 1558519173;
assign addr[31588]= 1659723983;
assign addr[31589]= 1752509516;
assign addr[31590]= 1836405100;
assign addr[31591]= 1910985158;
assign addr[31592]= 1975871368;
assign addr[31593]= 2030734582;
assign addr[31594]= 2075296495;
assign addr[31595]= 2109331059;
assign addr[31596]= 2132665626;
assign addr[31597]= 2145181827;
assign addr[31598]= 2146816171;
assign addr[31599]= 2137560369;
assign addr[31600]= 2117461370;
assign addr[31601]= 2086621133;
assign addr[31602]= 2045196100;
assign addr[31603]= 1993396407;
assign addr[31604]= 1931484818;
assign addr[31605]= 1859775393;
assign addr[31606]= 1778631892;
assign addr[31607]= 1688465931;
assign addr[31608]= 1589734894;
assign addr[31609]= 1482939614;
assign addr[31610]= 1368621831;
assign addr[31611]= 1247361445;
assign addr[31612]= 1119773573;
assign addr[31613]= 986505429;
assign addr[31614]= 848233042;
assign addr[31615]= 705657826;
assign addr[31616]= 559503022;
assign addr[31617]= 410510029;
assign addr[31618]= 259434643;
assign addr[31619]= 107043224;
assign addr[31620]= -45891193;
assign addr[31621]= -198592817;
assign addr[31622]= -350287041;
assign addr[31623]= -500204365;
assign addr[31624]= -647584304;
assign addr[31625]= -791679244;
assign addr[31626]= -931758235;
assign addr[31627]= -1067110699;
assign addr[31628]= -1197050035;
assign addr[31629]= -1320917099;
assign addr[31630]= -1438083551;
assign addr[31631]= -1547955041;
assign addr[31632]= -1649974225;
assign addr[31633]= -1743623590;
assign addr[31634]= -1828428082;
assign addr[31635]= -1903957513;
assign addr[31636]= -1969828744;
assign addr[31637]= -2025707632;
assign addr[31638]= -2071310720;
assign addr[31639]= -2106406677;
assign addr[31640]= -2130817471;
assign addr[31641]= -2144419275;
assign addr[31642]= -2147143090;
assign addr[31643]= -2138975100;
assign addr[31644]= -2119956737;
assign addr[31645]= -2090184478;
assign addr[31646]= -2049809346;
assign addr[31647]= -1999036154;
assign addr[31648]= -1938122457;
assign addr[31649]= -1867377253;
assign addr[31650]= -1787159411;
assign addr[31651]= -1697875851;
assign addr[31652]= -1599979481;
assign addr[31653]= -1493966902;
assign addr[31654]= -1380375881;
assign addr[31655]= -1259782632;
assign addr[31656]= -1132798888;
assign addr[31657]= -1000068799;
assign addr[31658]= -862265664;
assign addr[31659]= -720088517;
assign addr[31660]= -574258580;
assign addr[31661]= -425515602;
assign addr[31662]= -274614114;
assign addr[31663]= -122319591;
assign addr[31664]= 30595422;
assign addr[31665]= 183355234;
assign addr[31666]= 335184940;
assign addr[31667]= 485314355;
assign addr[31668]= 632981917;
assign addr[31669]= 777438554;
assign addr[31670]= 917951481;
assign addr[31671]= 1053807919;
assign addr[31672]= 1184318708;
assign addr[31673]= 1308821808;
assign addr[31674]= 1426685652;
assign addr[31675]= 1537312353;
assign addr[31676]= 1640140734;
assign addr[31677]= 1734649179;
assign addr[31678]= 1820358275;
assign addr[31679]= 1896833245;
assign addr[31680]= 1963686155;
assign addr[31681]= 2020577882;
assign addr[31682]= 2067219829;
assign addr[31683]= 2103375398;
assign addr[31684]= 2128861181;
assign addr[31685]= 2143547897;
assign addr[31686]= 2147361045;
assign addr[31687]= 2140281282;
assign addr[31688]= 2122344521;
assign addr[31689]= 2093641749;
assign addr[31690]= 2054318569;
assign addr[31691]= 2004574453;
assign addr[31692]= 1944661739;
assign addr[31693]= 1874884346;
assign addr[31694]= 1795596234;
assign addr[31695]= 1707199606;
assign addr[31696]= 1610142873;
assign addr[31697]= 1504918373;
assign addr[31698]= 1392059879;
assign addr[31699]= 1272139887;
assign addr[31700]= 1145766716;
assign addr[31701]= 1013581418;
assign addr[31702]= 876254528;
assign addr[31703]= 734482665;
assign addr[31704]= 588984994;
assign addr[31705]= 440499581;
assign addr[31706]= 289779648;
assign addr[31707]= 137589750;
assign addr[31708]= -15298099;
assign addr[31709]= -168108346;
assign addr[31710]= -320065829;
assign addr[31711]= -470399716;
assign addr[31712]= -618347408;
assign addr[31713]= -763158411;
assign addr[31714]= -904098143;
assign addr[31715]= -1040451659;
assign addr[31716]= -1171527280;
assign addr[31717]= -1296660098;
assign addr[31718]= -1415215352;
assign addr[31719]= -1526591649;
assign addr[31720]= -1630224009;
assign addr[31721]= -1725586737;
assign addr[31722]= -1812196087;
assign addr[31723]= -1889612716;
assign addr[31724]= -1957443913;
assign addr[31725]= -2015345591;
assign addr[31726]= -2063024031;
assign addr[31727]= -2100237377;
assign addr[31728]= -2126796855;
assign addr[31729]= -2142567738;
assign addr[31730]= -2147470025;
assign addr[31731]= -2141478848;
assign addr[31732]= -2124624598;
assign addr[31733]= -2096992772;
assign addr[31734]= -2058723538;
assign addr[31735]= -2010011024;
assign addr[31736]= -1951102334;
assign addr[31737]= -1882296293;
assign addr[31738]= -1803941934;
assign addr[31739]= -1716436725;
assign addr[31740]= -1620224553;
assign addr[31741]= -1515793473;
assign addr[31742]= -1403673233;
assign addr[31743]= -1284432584;
assign addr[31744]= -1158676398;
assign addr[31745]= -1027042599;
assign addr[31746]= -890198924;
assign addr[31747]= -748839539;
assign addr[31748]= -603681519;
assign addr[31749]= -455461206;
assign addr[31750]= -304930476;
assign addr[31751]= -152852926;
assign addr[31752]= 0;
assign addr[31753]= 152852926;
assign addr[31754]= 304930476;
assign addr[31755]= 455461206;
assign addr[31756]= 603681519;
assign addr[31757]= 748839539;
assign addr[31758]= 890198924;
assign addr[31759]= 1027042599;
assign addr[31760]= 1158676398;
assign addr[31761]= 1284432584;
assign addr[31762]= 1403673233;
assign addr[31763]= 1515793473;
assign addr[31764]= 1620224553;
assign addr[31765]= 1716436725;
assign addr[31766]= 1803941934;
assign addr[31767]= 1882296293;
assign addr[31768]= 1951102334;
assign addr[31769]= 2010011024;
assign addr[31770]= 2058723538;
assign addr[31771]= 2096992772;
assign addr[31772]= 2124624598;
assign addr[31773]= 2141478848;
assign addr[31774]= 2147470025;
assign addr[31775]= 2142567738;
assign addr[31776]= 2126796855;
assign addr[31777]= 2100237377;
assign addr[31778]= 2063024031;
assign addr[31779]= 2015345591;
assign addr[31780]= 1957443913;
assign addr[31781]= 1889612716;
assign addr[31782]= 1812196087;
assign addr[31783]= 1725586737;
assign addr[31784]= 1630224009;
assign addr[31785]= 1526591649;
assign addr[31786]= 1415215352;
assign addr[31787]= 1296660098;
assign addr[31788]= 1171527280;
assign addr[31789]= 1040451659;
assign addr[31790]= 904098143;
assign addr[31791]= 763158411;
assign addr[31792]= 618347408;
assign addr[31793]= 470399716;
assign addr[31794]= 320065829;
assign addr[31795]= 168108346;
assign addr[31796]= 15298099;
assign addr[31797]= -137589750;
assign addr[31798]= -289779648;
assign addr[31799]= -440499581;
assign addr[31800]= -588984994;
assign addr[31801]= -734482665;
assign addr[31802]= -876254528;
assign addr[31803]= -1013581418;
assign addr[31804]= -1145766716;
assign addr[31805]= -1272139887;
assign addr[31806]= -1392059879;
assign addr[31807]= -1504918373;
assign addr[31808]= -1610142873;
assign addr[31809]= -1707199606;
assign addr[31810]= -1795596234;
assign addr[31811]= -1874884346;
assign addr[31812]= -1944661739;
assign addr[31813]= -2004574453;
assign addr[31814]= -2054318569;
assign addr[31815]= -2093641749;
assign addr[31816]= -2122344521;
assign addr[31817]= -2140281282;
assign addr[31818]= -2147361045;
assign addr[31819]= -2143547897;
assign addr[31820]= -2128861181;
assign addr[31821]= -2103375398;
assign addr[31822]= -2067219829;
assign addr[31823]= -2020577882;
assign addr[31824]= -1963686155;
assign addr[31825]= -1896833245;
assign addr[31826]= -1820358275;
assign addr[31827]= -1734649179;
assign addr[31828]= -1640140734;
assign addr[31829]= -1537312353;
assign addr[31830]= -1426685652;
assign addr[31831]= -1308821808;
assign addr[31832]= -1184318708;
assign addr[31833]= -1053807919;
assign addr[31834]= -917951481;
assign addr[31835]= -777438554;
assign addr[31836]= -632981917;
assign addr[31837]= -485314355;
assign addr[31838]= -335184940;
assign addr[31839]= -183355234;
assign addr[31840]= -30595422;
assign addr[31841]= 122319591;
assign addr[31842]= 274614114;
assign addr[31843]= 425515602;
assign addr[31844]= 574258580;
assign addr[31845]= 720088517;
assign addr[31846]= 862265664;
assign addr[31847]= 1000068799;
assign addr[31848]= 1132798888;
assign addr[31849]= 1259782632;
assign addr[31850]= 1380375881;
assign addr[31851]= 1493966902;
assign addr[31852]= 1599979481;
assign addr[31853]= 1697875851;
assign addr[31854]= 1787159411;
assign addr[31855]= 1867377253;
assign addr[31856]= 1938122457;
assign addr[31857]= 1999036154;
assign addr[31858]= 2049809346;
assign addr[31859]= 2090184478;
assign addr[31860]= 2119956737;
assign addr[31861]= 2138975100;
assign addr[31862]= 2147143090;
assign addr[31863]= 2144419275;
assign addr[31864]= 2130817471;
assign addr[31865]= 2106406677;
assign addr[31866]= 2071310720;
assign addr[31867]= 2025707632;
assign addr[31868]= 1969828744;
assign addr[31869]= 1903957513;
assign addr[31870]= 1828428082;
assign addr[31871]= 1743623590;
assign addr[31872]= 1649974225;
assign addr[31873]= 1547955041;
assign addr[31874]= 1438083551;
assign addr[31875]= 1320917099;
assign addr[31876]= 1197050035;
assign addr[31877]= 1067110699;
assign addr[31878]= 931758235;
assign addr[31879]= 791679244;
assign addr[31880]= 647584304;
assign addr[31881]= 500204365;
assign addr[31882]= 350287041;
assign addr[31883]= 198592817;
assign addr[31884]= 45891193;
assign addr[31885]= -107043224;
assign addr[31886]= -259434643;
assign addr[31887]= -410510029;
assign addr[31888]= -559503022;
assign addr[31889]= -705657826;
assign addr[31890]= -848233042;
assign addr[31891]= -986505429;
assign addr[31892]= -1119773573;
assign addr[31893]= -1247361445;
assign addr[31894]= -1368621831;
assign addr[31895]= -1482939614;
assign addr[31896]= -1589734894;
assign addr[31897]= -1688465931;
assign addr[31898]= -1778631892;
assign addr[31899]= -1859775393;
assign addr[31900]= -1931484818;
assign addr[31901]= -1993396407;
assign addr[31902]= -2045196100;
assign addr[31903]= -2086621133;
assign addr[31904]= -2117461370;
assign addr[31905]= -2137560369;
assign addr[31906]= -2146816171;
assign addr[31907]= -2145181827;
assign addr[31908]= -2132665626;
assign addr[31909]= -2109331059;
assign addr[31910]= -2075296495;
assign addr[31911]= -2030734582;
assign addr[31912]= -1975871368;
assign addr[31913]= -1910985158;
assign addr[31914]= -1836405100;
assign addr[31915]= -1752509516;
assign addr[31916]= -1659723983;
assign addr[31917]= -1558519173;
assign addr[31918]= -1449408469;
assign addr[31919]= -1332945355;
assign addr[31920]= -1209720613;
assign addr[31921]= -1080359326;
assign addr[31922]= -945517704;
assign addr[31923]= -805879757;
assign addr[31924]= -662153826;
assign addr[31925]= -515068990;
assign addr[31926]= -365371365;
assign addr[31927]= -213820322;
assign addr[31928]= -61184634;
assign addr[31929]= 91761426;
assign addr[31930]= 244242007;
assign addr[31931]= 395483624;
assign addr[31932]= 544719071;
assign addr[31933]= 691191324;
assign addr[31934]= 834157373;
assign addr[31935]= 972891995;
assign addr[31936]= 1106691431;
assign addr[31937]= 1234876957;
assign addr[31938]= 1356798326;
assign addr[31939]= 1471837070;
assign addr[31940]= 1579409630;
assign addr[31941]= 1678970324;
assign addr[31942]= 1770014111;
assign addr[31943]= 1852079154;
assign addr[31944]= 1924749160;
assign addr[31945]= 1987655498;
assign addr[31946]= 2040479063;
assign addr[31947]= 2082951896;
assign addr[31948]= 2114858546;
assign addr[31949]= 2136037160;
assign addr[31950]= 2146380306;
assign addr[31951]= 2145835515;
assign addr[31952]= 2134405552;
assign addr[31953]= 2112148396;
assign addr[31954]= 2079176953;
assign addr[31955]= 2035658475;
assign addr[31956]= 1981813720;
assign addr[31957]= 1917915825;
assign addr[31958]= 1844288924;
assign addr[31959]= 1761306505;
assign addr[31960]= 1669389513;
assign addr[31961]= 1569004214;
assign addr[31962]= 1460659832;
assign addr[31963]= 1344905966;
assign addr[31964]= 1222329801;
assign addr[31965]= 1093553126;
assign addr[31966]= 959229189;
assign addr[31967]= 820039373;
assign addr[31968]= 676689746;
assign addr[31969]= 529907477;
assign addr[31970]= 380437148;
assign addr[31971]= 229036977;
assign addr[31972]= 76474970;
assign addr[31973]= -76474970;
assign addr[31974]= -229036977;
assign addr[31975]= -380437148;
assign addr[31976]= -529907477;
assign addr[31977]= -676689746;
assign addr[31978]= -820039373;
assign addr[31979]= -959229189;
assign addr[31980]= -1093553126;
assign addr[31981]= -1222329801;
assign addr[31982]= -1344905966;
assign addr[31983]= -1460659832;
assign addr[31984]= -1569004214;
assign addr[31985]= -1669389513;
assign addr[31986]= -1761306505;
assign addr[31987]= -1844288924;
assign addr[31988]= -1917915825;
assign addr[31989]= -1981813720;
assign addr[31990]= -2035658475;
assign addr[31991]= -2079176953;
assign addr[31992]= -2112148396;
assign addr[31993]= -2134405552;
assign addr[31994]= -2145835515;
assign addr[31995]= -2146380306;
assign addr[31996]= -2136037160;
assign addr[31997]= -2114858546;
assign addr[31998]= -2082951896;
assign addr[31999]= -2040479063;
assign addr[32000]= -1987655498;
assign addr[32001]= -1924749160;
assign addr[32002]= -1852079154;
assign addr[32003]= -1770014111;
assign addr[32004]= -1678970324;
assign addr[32005]= -1579409630;
assign addr[32006]= -1471837070;
assign addr[32007]= -1356798326;
assign addr[32008]= -1234876957;
assign addr[32009]= -1106691431;
assign addr[32010]= -972891995;
assign addr[32011]= -834157373;
assign addr[32012]= -691191324;
assign addr[32013]= -544719071;
assign addr[32014]= -395483624;
assign addr[32015]= -244242007;
assign addr[32016]= -91761426;
assign addr[32017]= 61184634;
assign addr[32018]= 213820322;
assign addr[32019]= 365371365;
assign addr[32020]= 515068990;
assign addr[32021]= 662153826;
assign addr[32022]= 805879757;
assign addr[32023]= 945517704;
assign addr[32024]= 1080359326;
assign addr[32025]= 1209720613;
assign addr[32026]= 1332945355;
assign addr[32027]= 1449408469;
assign addr[32028]= 1558519173;
assign addr[32029]= 1659723983;
assign addr[32030]= 1752509516;
assign addr[32031]= 1836405100;
assign addr[32032]= 1910985158;
assign addr[32033]= 1975871368;
assign addr[32034]= 2030734582;
assign addr[32035]= 2075296495;
assign addr[32036]= 2109331059;
assign addr[32037]= 2132665626;
assign addr[32038]= 2145181827;
assign addr[32039]= 2146816171;
assign addr[32040]= 2137560369;
assign addr[32041]= 2117461370;
assign addr[32042]= 2086621133;
assign addr[32043]= 2045196100;
assign addr[32044]= 1993396407;
assign addr[32045]= 1931484818;
assign addr[32046]= 1859775393;
assign addr[32047]= 1778631892;
assign addr[32048]= 1688465931;
assign addr[32049]= 1589734894;
assign addr[32050]= 1482939614;
assign addr[32051]= 1368621831;
assign addr[32052]= 1247361445;
assign addr[32053]= 1119773573;
assign addr[32054]= 986505429;
assign addr[32055]= 848233042;
assign addr[32056]= 705657826;
assign addr[32057]= 559503022;
assign addr[32058]= 410510029;
assign addr[32059]= 259434643;
assign addr[32060]= 107043224;
assign addr[32061]= -45891193;
assign addr[32062]= -198592817;
assign addr[32063]= -350287041;
assign addr[32064]= -500204365;
assign addr[32065]= -647584304;
assign addr[32066]= -791679244;
assign addr[32067]= -931758235;
assign addr[32068]= -1067110699;
assign addr[32069]= -1197050035;
assign addr[32070]= -1320917099;
assign addr[32071]= -1438083551;
assign addr[32072]= -1547955041;
assign addr[32073]= -1649974225;
assign addr[32074]= -1743623590;
assign addr[32075]= -1828428082;
assign addr[32076]= -1903957513;
assign addr[32077]= -1969828744;
assign addr[32078]= -2025707632;
assign addr[32079]= -2071310720;
assign addr[32080]= -2106406677;
assign addr[32081]= -2130817471;
assign addr[32082]= -2144419275;
assign addr[32083]= -2147143090;
assign addr[32084]= -2138975100;
assign addr[32085]= -2119956737;
assign addr[32086]= -2090184478;
assign addr[32087]= -2049809346;
assign addr[32088]= -1999036154;
assign addr[32089]= -1938122457;
assign addr[32090]= -1867377253;
assign addr[32091]= -1787159411;
assign addr[32092]= -1697875851;
assign addr[32093]= -1599979481;
assign addr[32094]= -1493966902;
assign addr[32095]= -1380375881;
assign addr[32096]= -1259782632;
assign addr[32097]= -1132798888;
assign addr[32098]= -1000068799;
assign addr[32099]= -862265664;
assign addr[32100]= -720088517;
assign addr[32101]= -574258580;
assign addr[32102]= -425515602;
assign addr[32103]= -274614114;
assign addr[32104]= -122319591;
assign addr[32105]= 30595422;
assign addr[32106]= 183355234;
assign addr[32107]= 335184940;
assign addr[32108]= 485314355;
assign addr[32109]= 632981917;
assign addr[32110]= 777438554;
assign addr[32111]= 917951481;
assign addr[32112]= 1053807919;
assign addr[32113]= 1184318708;
assign addr[32114]= 1308821808;
assign addr[32115]= 1426685652;
assign addr[32116]= 1537312353;
assign addr[32117]= 1640140734;
assign addr[32118]= 1734649179;
assign addr[32119]= 1820358275;
assign addr[32120]= 1896833245;
assign addr[32121]= 1963686155;
assign addr[32122]= 2020577882;
assign addr[32123]= 2067219829;
assign addr[32124]= 2103375398;
assign addr[32125]= 2128861181;
assign addr[32126]= 2143547897;
assign addr[32127]= 2147361045;
assign addr[32128]= 2140281282;
assign addr[32129]= 2122344521;
assign addr[32130]= 2093641749;
assign addr[32131]= 2054318569;
assign addr[32132]= 2004574453;
assign addr[32133]= 1944661739;
assign addr[32134]= 1874884346;
assign addr[32135]= 1795596234;
assign addr[32136]= 1707199606;
assign addr[32137]= 1610142873;
assign addr[32138]= 1504918373;
assign addr[32139]= 1392059879;
assign addr[32140]= 1272139887;
assign addr[32141]= 1145766716;
assign addr[32142]= 1013581418;
assign addr[32143]= 876254528;
assign addr[32144]= 734482665;
assign addr[32145]= 588984994;
assign addr[32146]= 440499581;
assign addr[32147]= 289779648;
assign addr[32148]= 137589750;
assign addr[32149]= -15298099;
assign addr[32150]= -168108346;
assign addr[32151]= -320065829;
assign addr[32152]= -470399716;
assign addr[32153]= -618347408;
assign addr[32154]= -763158411;
assign addr[32155]= -904098143;
assign addr[32156]= -1040451659;
assign addr[32157]= -1171527280;
assign addr[32158]= -1296660098;
assign addr[32159]= -1415215352;
assign addr[32160]= -1526591649;
assign addr[32161]= -1630224009;
assign addr[32162]= -1725586737;
assign addr[32163]= -1812196087;
assign addr[32164]= -1889612716;
assign addr[32165]= -1957443913;
assign addr[32166]= -2015345591;
assign addr[32167]= -2063024031;
assign addr[32168]= -2100237377;
assign addr[32169]= -2126796855;
assign addr[32170]= -2142567738;
assign addr[32171]= -2147470025;
assign addr[32172]= -2141478848;
assign addr[32173]= -2124624598;
assign addr[32174]= -2096992772;
assign addr[32175]= -2058723538;
assign addr[32176]= -2010011024;
assign addr[32177]= -1951102334;
assign addr[32178]= -1882296293;
assign addr[32179]= -1803941934;
assign addr[32180]= -1716436725;
assign addr[32181]= -1620224553;
assign addr[32182]= -1515793473;
assign addr[32183]= -1403673233;
assign addr[32184]= -1284432584;
assign addr[32185]= -1158676398;
assign addr[32186]= -1027042599;
assign addr[32187]= -890198924;
assign addr[32188]= -748839539;
assign addr[32189]= -603681519;
assign addr[32190]= -455461206;
assign addr[32191]= -304930476;
assign addr[32192]= -152852926;
assign addr[32193]= 0;
assign addr[32194]= 152852926;
assign addr[32195]= 304930476;
assign addr[32196]= 455461206;
assign addr[32197]= 603681519;
assign addr[32198]= 748839539;
assign addr[32199]= 890198924;
assign addr[32200]= 1027042599;
assign addr[32201]= 1158676398;
assign addr[32202]= 1284432584;
assign addr[32203]= 1403673233;
assign addr[32204]= 1515793473;
assign addr[32205]= 1620224553;
assign addr[32206]= 1716436725;
assign addr[32207]= 1803941934;
assign addr[32208]= 1882296293;
assign addr[32209]= 1951102334;
assign addr[32210]= 2010011024;
assign addr[32211]= 2058723538;
assign addr[32212]= 2096992772;
assign addr[32213]= 2124624598;
assign addr[32214]= 2141478848;
assign addr[32215]= 2147470025;
assign addr[32216]= 2142567738;
assign addr[32217]= 2126796855;
assign addr[32218]= 2100237377;
assign addr[32219]= 2063024031;
assign addr[32220]= 2015345591;
assign addr[32221]= 1957443913;
assign addr[32222]= 1889612716;
assign addr[32223]= 1812196087;
assign addr[32224]= 1725586737;
assign addr[32225]= 1630224009;
assign addr[32226]= 1526591649;
assign addr[32227]= 1415215352;
assign addr[32228]= 1296660098;
assign addr[32229]= 1171527280;
assign addr[32230]= 1040451659;
assign addr[32231]= 904098143;
assign addr[32232]= 763158411;
assign addr[32233]= 618347408;
assign addr[32234]= 470399716;
assign addr[32235]= 320065829;
assign addr[32236]= 168108346;
assign addr[32237]= 15298099;
assign addr[32238]= -137589750;
assign addr[32239]= -289779648;
assign addr[32240]= -440499581;
assign addr[32241]= -588984994;
assign addr[32242]= -734482665;
assign addr[32243]= -876254528;
assign addr[32244]= -1013581418;
assign addr[32245]= -1145766716;
assign addr[32246]= -1272139887;
assign addr[32247]= -1392059879;
assign addr[32248]= -1504918373;
assign addr[32249]= -1610142873;
assign addr[32250]= -1707199606;
assign addr[32251]= -1795596234;
assign addr[32252]= -1874884346;
assign addr[32253]= -1944661739;
assign addr[32254]= -2004574453;
assign addr[32255]= -2054318569;
assign addr[32256]= -2093641749;
assign addr[32257]= -2122344521;
assign addr[32258]= -2140281282;
assign addr[32259]= -2147361045;
assign addr[32260]= -2143547897;
assign addr[32261]= -2128861181;
assign addr[32262]= -2103375398;
assign addr[32263]= -2067219829;
assign addr[32264]= -2020577882;
assign addr[32265]= -1963686155;
assign addr[32266]= -1896833245;
assign addr[32267]= -1820358275;
assign addr[32268]= -1734649179;
assign addr[32269]= -1640140734;
assign addr[32270]= -1537312353;
assign addr[32271]= -1426685652;
assign addr[32272]= -1308821808;
assign addr[32273]= -1184318708;
assign addr[32274]= -1053807919;
assign addr[32275]= -917951481;
assign addr[32276]= -777438554;
assign addr[32277]= -632981917;
assign addr[32278]= -485314355;
assign addr[32279]= -335184940;
assign addr[32280]= -183355234;
assign addr[32281]= -30595422;
assign addr[32282]= 122319591;
assign addr[32283]= 274614114;
assign addr[32284]= 425515602;
assign addr[32285]= 574258580;
assign addr[32286]= 720088517;
assign addr[32287]= 862265664;
assign addr[32288]= 1000068799;
assign addr[32289]= 1132798888;
assign addr[32290]= 1259782632;
assign addr[32291]= 1380375881;
assign addr[32292]= 1493966902;
assign addr[32293]= 1599979481;
assign addr[32294]= 1697875851;
assign addr[32295]= 1787159411;
assign addr[32296]= 1867377253;
assign addr[32297]= 1938122457;
assign addr[32298]= 1999036154;
assign addr[32299]= 2049809346;
assign addr[32300]= 2090184478;
assign addr[32301]= 2119956737;
assign addr[32302]= 2138975100;
assign addr[32303]= 2147143090;
assign addr[32304]= 2144419275;
assign addr[32305]= 2130817471;
assign addr[32306]= 2106406677;
assign addr[32307]= 2071310720;
assign addr[32308]= 2025707632;
assign addr[32309]= 1969828744;
assign addr[32310]= 1903957513;
assign addr[32311]= 1828428082;
assign addr[32312]= 1743623590;
assign addr[32313]= 1649974225;
assign addr[32314]= 1547955041;
assign addr[32315]= 1438083551;
assign addr[32316]= 1320917099;
assign addr[32317]= 1197050035;
assign addr[32318]= 1067110699;
assign addr[32319]= 931758235;
assign addr[32320]= 791679244;
assign addr[32321]= 647584304;
assign addr[32322]= 500204365;
assign addr[32323]= 350287041;
assign addr[32324]= 198592817;
assign addr[32325]= 45891193;
assign addr[32326]= -107043224;
assign addr[32327]= -259434643;
assign addr[32328]= -410510029;
assign addr[32329]= -559503022;
assign addr[32330]= -705657826;
assign addr[32331]= -848233042;
assign addr[32332]= -986505429;
assign addr[32333]= -1119773573;
assign addr[32334]= -1247361445;
assign addr[32335]= -1368621831;
assign addr[32336]= -1482939614;
assign addr[32337]= -1589734894;
assign addr[32338]= -1688465931;
assign addr[32339]= -1778631892;
assign addr[32340]= -1859775393;
assign addr[32341]= -1931484818;
assign addr[32342]= -1993396407;
assign addr[32343]= -2045196100;
assign addr[32344]= -2086621133;
assign addr[32345]= -2117461370;
assign addr[32346]= -2137560369;
assign addr[32347]= -2146816171;
assign addr[32348]= -2145181827;
assign addr[32349]= -2132665626;
assign addr[32350]= -2109331059;
assign addr[32351]= -2075296495;
assign addr[32352]= -2030734582;
assign addr[32353]= -1975871368;
assign addr[32354]= -1910985158;
assign addr[32355]= -1836405100;
assign addr[32356]= -1752509516;
assign addr[32357]= -1659723983;
assign addr[32358]= -1558519173;
assign addr[32359]= -1449408469;
assign addr[32360]= -1332945355;
assign addr[32361]= -1209720613;
assign addr[32362]= -1080359326;
assign addr[32363]= -945517704;
assign addr[32364]= -805879757;
assign addr[32365]= -662153826;
assign addr[32366]= -515068990;
assign addr[32367]= -365371365;
assign addr[32368]= -213820322;
assign addr[32369]= -61184634;
assign addr[32370]= 91761426;
assign addr[32371]= 244242007;
assign addr[32372]= 395483624;
assign addr[32373]= 544719071;
assign addr[32374]= 691191324;
assign addr[32375]= 834157373;
assign addr[32376]= 972891995;
assign addr[32377]= 1106691431;
assign addr[32378]= 1234876957;
assign addr[32379]= 1356798326;
assign addr[32380]= 1471837070;
assign addr[32381]= 1579409630;
assign addr[32382]= 1678970324;
assign addr[32383]= 1770014111;
assign addr[32384]= 1852079154;
assign addr[32385]= 1924749160;
assign addr[32386]= 1987655498;
assign addr[32387]= 2040479063;
assign addr[32388]= 2082951896;
assign addr[32389]= 2114858546;
assign addr[32390]= 2136037160;
assign addr[32391]= 2146380306;
assign addr[32392]= 2145835515;
assign addr[32393]= 2134405552;
assign addr[32394]= 2112148396;
assign addr[32395]= 2079176953;
assign addr[32396]= 2035658475;
assign addr[32397]= 1981813720;
assign addr[32398]= 1917915825;
assign addr[32399]= 1844288924;
assign addr[32400]= 1761306505;
assign addr[32401]= 1669389513;
assign addr[32402]= 1569004214;
assign addr[32403]= 1460659832;
assign addr[32404]= 1344905966;
assign addr[32405]= 1222329801;
assign addr[32406]= 1093553126;
assign addr[32407]= 959229189;
assign addr[32408]= 820039373;
assign addr[32409]= 676689746;
assign addr[32410]= 529907477;
assign addr[32411]= 380437148;
assign addr[32412]= 229036977;
assign addr[32413]= 76474970;
assign addr[32414]= -76474970;
assign addr[32415]= -229036977;
assign addr[32416]= -380437148;
assign addr[32417]= -529907477;
assign addr[32418]= -676689746;
assign addr[32419]= -820039373;
assign addr[32420]= -959229189;
assign addr[32421]= -1093553126;
assign addr[32422]= -1222329801;
assign addr[32423]= -1344905966;
assign addr[32424]= -1460659832;
assign addr[32425]= -1569004214;
assign addr[32426]= -1669389513;
assign addr[32427]= -1761306505;
assign addr[32428]= -1844288924;
assign addr[32429]= -1917915825;
assign addr[32430]= -1981813720;
assign addr[32431]= -2035658475;
assign addr[32432]= -2079176953;
assign addr[32433]= -2112148396;
assign addr[32434]= -2134405552;
assign addr[32435]= -2145835515;
assign addr[32436]= -2146380306;
assign addr[32437]= -2136037160;
assign addr[32438]= -2114858546;
assign addr[32439]= -2082951896;
assign addr[32440]= -2040479063;
assign addr[32441]= -1987655498;
assign addr[32442]= -1924749160;
assign addr[32443]= -1852079154;
assign addr[32444]= -1770014111;
assign addr[32445]= -1678970324;
assign addr[32446]= -1579409630;
assign addr[32447]= -1471837070;
assign addr[32448]= -1356798326;
assign addr[32449]= -1234876957;
assign addr[32450]= -1106691431;
assign addr[32451]= -972891995;
assign addr[32452]= -834157373;
assign addr[32453]= -691191324;
assign addr[32454]= -544719071;
assign addr[32455]= -395483624;
assign addr[32456]= -244242007;
assign addr[32457]= -91761426;
assign addr[32458]= 61184634;
assign addr[32459]= 213820322;
assign addr[32460]= 365371365;
assign addr[32461]= 515068990;
assign addr[32462]= 662153826;
assign addr[32463]= 805879757;
assign addr[32464]= 945517704;
assign addr[32465]= 1080359326;
assign addr[32466]= 1209720613;
assign addr[32467]= 1332945355;
assign addr[32468]= 1449408469;
assign addr[32469]= 1558519173;
assign addr[32470]= 1659723983;
assign addr[32471]= 1752509516;
assign addr[32472]= 1836405100;
assign addr[32473]= 1910985158;
assign addr[32474]= 1975871368;
assign addr[32475]= 2030734582;
assign addr[32476]= 2075296495;
assign addr[32477]= 2109331059;
assign addr[32478]= 2132665626;
assign addr[32479]= 2145181827;
assign addr[32480]= 2146816171;
assign addr[32481]= 2137560369;
assign addr[32482]= 2117461370;
assign addr[32483]= 2086621133;
assign addr[32484]= 2045196100;
assign addr[32485]= 1993396407;
assign addr[32486]= 1931484818;
assign addr[32487]= 1859775393;
assign addr[32488]= 1778631892;
assign addr[32489]= 1688465931;
assign addr[32490]= 1589734894;
assign addr[32491]= 1482939614;
assign addr[32492]= 1368621831;
assign addr[32493]= 1247361445;
assign addr[32494]= 1119773573;
assign addr[32495]= 986505429;
assign addr[32496]= 848233042;
assign addr[32497]= 705657826;
assign addr[32498]= 559503022;
assign addr[32499]= 410510029;
assign addr[32500]= 259434643;
assign addr[32501]= 107043224;
assign addr[32502]= -45891193;
assign addr[32503]= -198592817;
assign addr[32504]= -350287041;
assign addr[32505]= -500204365;
assign addr[32506]= -647584304;
assign addr[32507]= -791679244;
assign addr[32508]= -931758235;
assign addr[32509]= -1067110699;
assign addr[32510]= -1197050035;
assign addr[32511]= -1320917099;
assign addr[32512]= -1438083551;
assign addr[32513]= -1547955041;
assign addr[32514]= -1649974225;
assign addr[32515]= -1743623590;
assign addr[32516]= -1828428082;
assign addr[32517]= -1903957513;
assign addr[32518]= -1969828744;
assign addr[32519]= -2025707632;
assign addr[32520]= -2071310720;
assign addr[32521]= -2106406677;
assign addr[32522]= -2130817471;
assign addr[32523]= -2144419275;
assign addr[32524]= -2147143090;
assign addr[32525]= -2138975100;
assign addr[32526]= -2119956737;
assign addr[32527]= -2090184478;
assign addr[32528]= -2049809346;
assign addr[32529]= -1999036154;
assign addr[32530]= -1938122457;
assign addr[32531]= -1867377253;
assign addr[32532]= -1787159411;
assign addr[32533]= -1697875851;
assign addr[32534]= -1599979481;
assign addr[32535]= -1493966902;
assign addr[32536]= -1380375881;
assign addr[32537]= -1259782632;
assign addr[32538]= -1132798888;
assign addr[32539]= -1000068799;
assign addr[32540]= -862265664;
assign addr[32541]= -720088517;
assign addr[32542]= -574258580;
assign addr[32543]= -425515602;
assign addr[32544]= -274614114;
assign addr[32545]= -122319591;
assign addr[32546]= 30595422;
assign addr[32547]= 183355234;
assign addr[32548]= 335184940;
assign addr[32549]= 485314355;
assign addr[32550]= 632981917;
assign addr[32551]= 777438554;
assign addr[32552]= 917951481;
assign addr[32553]= 1053807919;
assign addr[32554]= 1184318708;
assign addr[32555]= 1308821808;
assign addr[32556]= 1426685652;
assign addr[32557]= 1537312353;
assign addr[32558]= 1640140734;
assign addr[32559]= 1734649179;
assign addr[32560]= 1820358275;
assign addr[32561]= 1896833245;
assign addr[32562]= 1963686155;
assign addr[32563]= 2020577882;
assign addr[32564]= 2067219829;
assign addr[32565]= 2103375398;
assign addr[32566]= 2128861181;
assign addr[32567]= 2143547897;
assign addr[32568]= 2147361045;
assign addr[32569]= 2140281282;
assign addr[32570]= 2122344521;
assign addr[32571]= 2093641749;
assign addr[32572]= 2054318569;
assign addr[32573]= 2004574453;
assign addr[32574]= 1944661739;
assign addr[32575]= 1874884346;
assign addr[32576]= 1795596234;
assign addr[32577]= 1707199606;
assign addr[32578]= 1610142873;
assign addr[32579]= 1504918373;
assign addr[32580]= 1392059879;
assign addr[32581]= 1272139887;
assign addr[32582]= 1145766716;
assign addr[32583]= 1013581418;
assign addr[32584]= 876254528;
assign addr[32585]= 734482665;
assign addr[32586]= 588984994;
assign addr[32587]= 440499581;
assign addr[32588]= 289779648;
assign addr[32589]= 137589750;
assign addr[32590]= -15298099;
assign addr[32591]= -168108346;
assign addr[32592]= -320065829;
assign addr[32593]= -470399716;
assign addr[32594]= -618347408;
assign addr[32595]= -763158411;
assign addr[32596]= -904098143;
assign addr[32597]= -1040451659;
assign addr[32598]= -1171527280;
assign addr[32599]= -1296660098;
assign addr[32600]= -1415215352;
assign addr[32601]= -1526591649;
assign addr[32602]= -1630224009;
assign addr[32603]= -1725586737;
assign addr[32604]= -1812196087;
assign addr[32605]= -1889612716;
assign addr[32606]= -1957443913;
assign addr[32607]= -2015345591;
assign addr[32608]= -2063024031;
assign addr[32609]= -2100237377;
assign addr[32610]= -2126796855;
assign addr[32611]= -2142567738;
assign addr[32612]= -2147470025;
assign addr[32613]= -2141478848;
assign addr[32614]= -2124624598;
assign addr[32615]= -2096992772;
assign addr[32616]= -2058723538;
assign addr[32617]= -2010011024;
assign addr[32618]= -1951102334;
assign addr[32619]= -1882296293;
assign addr[32620]= -1803941934;
assign addr[32621]= -1716436725;
assign addr[32622]= -1620224553;
assign addr[32623]= -1515793473;
assign addr[32624]= -1403673233;
assign addr[32625]= -1284432584;
assign addr[32626]= -1158676398;
assign addr[32627]= -1027042599;
assign addr[32628]= -890198924;
assign addr[32629]= -748839539;
assign addr[32630]= -603681519;
assign addr[32631]= -455461206;
assign addr[32632]= -304930476;
assign addr[32633]= -152852926;
assign addr[32634]= 0;
assign addr[32635]= 152852926;
assign addr[32636]= 304930476;
assign addr[32637]= 455461206;
assign addr[32638]= 603681519;
assign addr[32639]= 748839539;
assign addr[32640]= 890198924;
assign addr[32641]= 1027042599;
assign addr[32642]= 1158676398;
assign addr[32643]= 1284432584;
assign addr[32644]= 1403673233;
assign addr[32645]= 1515793473;
assign addr[32646]= 1620224553;
assign addr[32647]= 1716436725;
assign addr[32648]= 1803941934;
assign addr[32649]= 1882296293;
assign addr[32650]= 1951102334;
assign addr[32651]= 2010011024;
assign addr[32652]= 2058723538;
assign addr[32653]= 2096992772;
assign addr[32654]= 2124624598;
assign addr[32655]= 2141478848;
assign addr[32656]= 2147470025;
assign addr[32657]= 2142567738;
assign addr[32658]= 2126796855;
assign addr[32659]= 2100237377;
assign addr[32660]= 2063024031;
assign addr[32661]= 2015345591;
assign addr[32662]= 1957443913;
assign addr[32663]= 1889612716;
assign addr[32664]= 1812196087;
assign addr[32665]= 1725586737;
assign addr[32666]= 1630224009;
assign addr[32667]= 1526591649;
assign addr[32668]= 1415215352;
assign addr[32669]= 1296660098;
assign addr[32670]= 1171527280;
assign addr[32671]= 1040451659;
assign addr[32672]= 904098143;
assign addr[32673]= 763158411;
assign addr[32674]= 618347408;
assign addr[32675]= 470399716;
assign addr[32676]= 320065829;
assign addr[32677]= 168108346;
assign addr[32678]= 15298099;
assign addr[32679]= -137589750;
assign addr[32680]= -289779648;
assign addr[32681]= -440499581;
assign addr[32682]= -588984994;
assign addr[32683]= -734482665;
assign addr[32684]= -876254528;
assign addr[32685]= -1013581418;
assign addr[32686]= -1145766716;
assign addr[32687]= -1272139887;
assign addr[32688]= -1392059879;
assign addr[32689]= -1504918373;
assign addr[32690]= -1610142873;
assign addr[32691]= -1707199606;
assign addr[32692]= -1795596234;
assign addr[32693]= -1874884346;
assign addr[32694]= -1944661739;
assign addr[32695]= -2004574453;
assign addr[32696]= -2054318569;
assign addr[32697]= -2093641749;
assign addr[32698]= -2122344521;
assign addr[32699]= -2140281282;
assign addr[32700]= -2147361045;
assign addr[32701]= -2143547897;
assign addr[32702]= -2128861181;
assign addr[32703]= -2103375398;
assign addr[32704]= -2067219829;
assign addr[32705]= -2020577882;
assign addr[32706]= -1963686155;
assign addr[32707]= -1896833245;
assign addr[32708]= -1820358275;
assign addr[32709]= -1734649179;
assign addr[32710]= -1640140734;
assign addr[32711]= -1537312353;
assign addr[32712]= -1426685652;
assign addr[32713]= -1308821808;
assign addr[32714]= -1184318708;
assign addr[32715]= -1053807919;
assign addr[32716]= -917951481;
assign addr[32717]= -777438554;
assign addr[32718]= -632981917;
assign addr[32719]= -485314355;
assign addr[32720]= -335184940;
assign addr[32721]= -183355234;
assign addr[32722]= -30595422;
assign addr[32723]= 122319591;
assign addr[32724]= 274614114;
assign addr[32725]= 425515602;
assign addr[32726]= 574258580;
assign addr[32727]= 720088517;
assign addr[32728]= 862265664;
assign addr[32729]= 1000068799;
assign addr[32730]= 1132798888;
assign addr[32731]= 1259782632;
assign addr[32732]= 1380375881;
assign addr[32733]= 1493966902;
assign addr[32734]= 1599979481;
assign addr[32735]= 1697875851;
assign addr[32736]= 1787159411;
assign addr[32737]= 1867377253;
assign addr[32738]= 1938122457;
assign addr[32739]= 1999036154;
assign addr[32740]= 2049809346;
assign addr[32741]= 2090184478;
assign addr[32742]= 2119956737;
assign addr[32743]= 2138975100;
assign addr[32744]= 2147143090;
assign addr[32745]= 2144419275;
assign addr[32746]= 2130817471;
assign addr[32747]= 2106406677;
assign addr[32748]= 2071310720;
assign addr[32749]= 2025707632;
assign addr[32750]= 1969828744;
assign addr[32751]= 1903957513;
assign addr[32752]= 1828428082;
assign addr[32753]= 1743623590;
assign addr[32754]= 1649974225;
assign addr[32755]= 1547955041;
assign addr[32756]= 1438083551;
assign addr[32757]= 1320917099;
assign addr[32758]= 1197050035;
assign addr[32759]= 1067110699;
assign addr[32760]= 931758235;
assign addr[32761]= 791679244;
assign addr[32762]= 647584304;
assign addr[32763]= 500204365;
assign addr[32764]= 350287041;
assign addr[32765]= 198592817;
assign addr[32766]= 45891193;
assign addr[32767]= -107043224;
assign addr[32768]= -259434643;
assign addr[32769]= -410510029;
assign addr[32770]= -559503022;
assign addr[32771]= -705657826;
assign addr[32772]= -848233042;
assign addr[32773]= -986505429;
assign addr[32774]= -1119773573;
assign addr[32775]= -1247361445;
assign addr[32776]= -1368621831;
assign addr[32777]= -1482939614;
assign addr[32778]= -1589734894;
assign addr[32779]= -1688465931;
assign addr[32780]= -1778631892;
assign addr[32781]= -1859775393;
assign addr[32782]= -1931484818;
assign addr[32783]= -1993396407;
assign addr[32784]= -2045196100;
assign addr[32785]= -2086621133;
assign addr[32786]= -2117461370;
assign addr[32787]= -2137560369;
assign addr[32788]= -2146816171;
assign addr[32789]= -2145181827;
assign addr[32790]= -2132665626;
assign addr[32791]= -2109331059;
assign addr[32792]= -2075296495;
assign addr[32793]= -2030734582;
assign addr[32794]= -1975871368;
assign addr[32795]= -1910985158;
assign addr[32796]= -1836405100;
assign addr[32797]= -1752509516;
assign addr[32798]= -1659723983;
assign addr[32799]= -1558519173;
assign addr[32800]= -1449408469;
assign addr[32801]= -1332945355;
assign addr[32802]= -1209720613;
assign addr[32803]= -1080359326;
assign addr[32804]= -945517704;
assign addr[32805]= -805879757;
assign addr[32806]= -662153826;
assign addr[32807]= -515068990;
assign addr[32808]= -365371365;
assign addr[32809]= -213820322;
assign addr[32810]= -61184634;
assign addr[32811]= 91761426;
assign addr[32812]= 244242007;
assign addr[32813]= 395483624;
assign addr[32814]= 544719071;
assign addr[32815]= 691191324;
assign addr[32816]= 834157373;
assign addr[32817]= 972891995;
assign addr[32818]= 1106691431;
assign addr[32819]= 1234876957;
assign addr[32820]= 1356798326;
assign addr[32821]= 1471837070;
assign addr[32822]= 1579409630;
assign addr[32823]= 1678970324;
assign addr[32824]= 1770014111;
assign addr[32825]= 1852079154;
assign addr[32826]= 1924749160;
assign addr[32827]= 1987655498;
assign addr[32828]= 2040479063;
assign addr[32829]= 2082951896;
assign addr[32830]= 2114858546;
assign addr[32831]= 2136037160;
assign addr[32832]= 2146380306;
assign addr[32833]= 2145835515;
assign addr[32834]= 2134405552;
assign addr[32835]= 2112148396;
assign addr[32836]= 2079176953;
assign addr[32837]= 2035658475;
assign addr[32838]= 1981813720;
assign addr[32839]= 1917915825;
assign addr[32840]= 1844288924;
assign addr[32841]= 1761306505;
assign addr[32842]= 1669389513;
assign addr[32843]= 1569004214;
assign addr[32844]= 1460659832;
assign addr[32845]= 1344905966;
assign addr[32846]= 1222329801;
assign addr[32847]= 1093553126;
assign addr[32848]= 959229189;
assign addr[32849]= 820039373;
assign addr[32850]= 676689746;
assign addr[32851]= 529907477;
assign addr[32852]= 380437148;
assign addr[32853]= 229036977;
assign addr[32854]= 76474970;
assign addr[32855]= -76474970;
assign addr[32856]= -229036977;
assign addr[32857]= -380437148;
assign addr[32858]= -529907477;
assign addr[32859]= -676689746;
assign addr[32860]= -820039373;
assign addr[32861]= -959229189;
assign addr[32862]= -1093553126;
assign addr[32863]= -1222329801;
assign addr[32864]= -1344905966;
assign addr[32865]= -1460659832;
assign addr[32866]= -1569004214;
assign addr[32867]= -1669389513;
assign addr[32868]= -1761306505;
assign addr[32869]= -1844288924;
assign addr[32870]= -1917915825;
assign addr[32871]= -1981813720;
assign addr[32872]= -2035658475;
assign addr[32873]= -2079176953;
assign addr[32874]= -2112148396;
assign addr[32875]= -2134405552;
assign addr[32876]= -2145835515;
assign addr[32877]= -2146380306;
assign addr[32878]= -2136037160;
assign addr[32879]= -2114858546;
assign addr[32880]= -2082951896;
assign addr[32881]= -2040479063;
assign addr[32882]= -1987655498;
assign addr[32883]= -1924749160;
assign addr[32884]= -1852079154;
assign addr[32885]= -1770014111;
assign addr[32886]= -1678970324;
assign addr[32887]= -1579409630;
assign addr[32888]= -1471837070;
assign addr[32889]= -1356798326;
assign addr[32890]= -1234876957;
assign addr[32891]= -1106691431;
assign addr[32892]= -972891995;
assign addr[32893]= -834157373;
assign addr[32894]= -691191324;
assign addr[32895]= -544719071;
assign addr[32896]= -395483624;
assign addr[32897]= -244242007;
assign addr[32898]= -91761426;
assign addr[32899]= 61184634;
assign addr[32900]= 213820322;
assign addr[32901]= 365371365;
assign addr[32902]= 515068990;
assign addr[32903]= 662153826;
assign addr[32904]= 805879757;
assign addr[32905]= 945517704;
assign addr[32906]= 1080359326;
assign addr[32907]= 1209720613;
assign addr[32908]= 1332945355;
assign addr[32909]= 1449408469;
assign addr[32910]= 1558519173;
assign addr[32911]= 1659723983;
assign addr[32912]= 1752509516;
assign addr[32913]= 1836405100;
assign addr[32914]= 1910985158;
assign addr[32915]= 1975871368;
assign addr[32916]= 2030734582;
assign addr[32917]= 2075296495;
assign addr[32918]= 2109331059;
assign addr[32919]= 2132665626;
assign addr[32920]= 2145181827;
assign addr[32921]= 2146816171;
assign addr[32922]= 2137560369;
assign addr[32923]= 2117461370;
assign addr[32924]= 2086621133;
assign addr[32925]= 2045196100;
assign addr[32926]= 1993396407;
assign addr[32927]= 1931484818;
assign addr[32928]= 1859775393;
assign addr[32929]= 1778631892;
assign addr[32930]= 1688465931;
assign addr[32931]= 1589734894;
assign addr[32932]= 1482939614;
assign addr[32933]= 1368621831;
assign addr[32934]= 1247361445;
assign addr[32935]= 1119773573;
assign addr[32936]= 986505429;
assign addr[32937]= 848233042;
assign addr[32938]= 705657826;
assign addr[32939]= 559503022;
assign addr[32940]= 410510029;
assign addr[32941]= 259434643;
assign addr[32942]= 107043224;
assign addr[32943]= -45891193;
assign addr[32944]= -198592817;
assign addr[32945]= -350287041;
assign addr[32946]= -500204365;
assign addr[32947]= -647584304;
assign addr[32948]= -791679244;
assign addr[32949]= -931758235;
assign addr[32950]= -1067110699;
assign addr[32951]= -1197050035;
assign addr[32952]= -1320917099;
assign addr[32953]= -1438083551;
assign addr[32954]= -1547955041;
assign addr[32955]= -1649974225;
assign addr[32956]= -1743623590;
assign addr[32957]= -1828428082;
assign addr[32958]= -1903957513;
assign addr[32959]= -1969828744;
assign addr[32960]= -2025707632;
assign addr[32961]= -2071310720;
assign addr[32962]= -2106406677;
assign addr[32963]= -2130817471;
assign addr[32964]= -2144419275;
assign addr[32965]= -2147143090;
assign addr[32966]= -2138975100;
assign addr[32967]= -2119956737;
assign addr[32968]= -2090184478;
assign addr[32969]= -2049809346;
assign addr[32970]= -1999036154;
assign addr[32971]= -1938122457;
assign addr[32972]= -1867377253;
assign addr[32973]= -1787159411;
assign addr[32974]= -1697875851;
assign addr[32975]= -1599979481;
assign addr[32976]= -1493966902;
assign addr[32977]= -1380375881;
assign addr[32978]= -1259782632;
assign addr[32979]= -1132798888;
assign addr[32980]= -1000068799;
assign addr[32981]= -862265664;
assign addr[32982]= -720088517;
assign addr[32983]= -574258580;
assign addr[32984]= -425515602;
assign addr[32985]= -274614114;
assign addr[32986]= -122319591;
assign addr[32987]= 30595422;
assign addr[32988]= 183355234;
assign addr[32989]= 335184940;
assign addr[32990]= 485314355;
assign addr[32991]= 632981917;
assign addr[32992]= 777438554;
assign addr[32993]= 917951481;
assign addr[32994]= 1053807919;
assign addr[32995]= 1184318708;
assign addr[32996]= 1308821808;
assign addr[32997]= 1426685652;
assign addr[32998]= 1537312353;
assign addr[32999]= 1640140734;
assign addr[33000]= 1734649179;
assign addr[33001]= 1820358275;
assign addr[33002]= 1896833245;
assign addr[33003]= 1963686155;
assign addr[33004]= 2020577882;
assign addr[33005]= 2067219829;
assign addr[33006]= 2103375398;
assign addr[33007]= 2128861181;
assign addr[33008]= 2143547897;
assign addr[33009]= 2147361045;
assign addr[33010]= 2140281282;
assign addr[33011]= 2122344521;
assign addr[33012]= 2093641749;
assign addr[33013]= 2054318569;
assign addr[33014]= 2004574453;
assign addr[33015]= 1944661739;
assign addr[33016]= 1874884346;
assign addr[33017]= 1795596234;
assign addr[33018]= 1707199606;
assign addr[33019]= 1610142873;
assign addr[33020]= 1504918373;
assign addr[33021]= 1392059879;
assign addr[33022]= 1272139887;
assign addr[33023]= 1145766716;
assign addr[33024]= 1013581418;
assign addr[33025]= 876254528;
assign addr[33026]= 734482665;
assign addr[33027]= 588984994;
assign addr[33028]= 440499581;
assign addr[33029]= 289779648;
assign addr[33030]= 137589750;
assign addr[33031]= -15298099;
assign addr[33032]= -168108346;
assign addr[33033]= -320065829;
assign addr[33034]= -470399716;
assign addr[33035]= -618347408;
assign addr[33036]= -763158411;
assign addr[33037]= -904098143;
assign addr[33038]= -1040451659;
assign addr[33039]= -1171527280;
assign addr[33040]= -1296660098;
assign addr[33041]= -1415215352;
assign addr[33042]= -1526591649;
assign addr[33043]= -1630224009;
assign addr[33044]= -1725586737;
assign addr[33045]= -1812196087;
assign addr[33046]= -1889612716;
assign addr[33047]= -1957443913;
assign addr[33048]= -2015345591;
assign addr[33049]= -2063024031;
assign addr[33050]= -2100237377;
assign addr[33051]= -2126796855;
assign addr[33052]= -2142567738;
assign addr[33053]= -2147470025;
assign addr[33054]= -2141478848;
assign addr[33055]= -2124624598;
assign addr[33056]= -2096992772;
assign addr[33057]= -2058723538;
assign addr[33058]= -2010011024;
assign addr[33059]= -1951102334;
assign addr[33060]= -1882296293;
assign addr[33061]= -1803941934;
assign addr[33062]= -1716436725;
assign addr[33063]= -1620224553;
assign addr[33064]= -1515793473;
assign addr[33065]= -1403673233;
assign addr[33066]= -1284432584;
assign addr[33067]= -1158676398;
assign addr[33068]= -1027042599;
assign addr[33069]= -890198924;
assign addr[33070]= -748839539;
assign addr[33071]= -603681519;
assign addr[33072]= -455461206;
assign addr[33073]= -304930476;
assign addr[33074]= -152852926;
assign addr[33075]= 0;
assign addr[33076]= 152852926;
assign addr[33077]= 304930476;
assign addr[33078]= 455461206;
assign addr[33079]= 603681519;
assign addr[33080]= 748839539;
assign addr[33081]= 890198924;
assign addr[33082]= 1027042599;
assign addr[33083]= 1158676398;
assign addr[33084]= 1284432584;
assign addr[33085]= 1403673233;
assign addr[33086]= 1515793473;
assign addr[33087]= 1620224553;
assign addr[33088]= 1716436725;
assign addr[33089]= 1803941934;
assign addr[33090]= 1882296293;
assign addr[33091]= 1951102334;
assign addr[33092]= 2010011024;
assign addr[33093]= 2058723538;
assign addr[33094]= 2096992772;
assign addr[33095]= 2124624598;
assign addr[33096]= 2141478848;
assign addr[33097]= 2147470025;
assign addr[33098]= 2142567738;
assign addr[33099]= 2126796855;
assign addr[33100]= 2100237377;
assign addr[33101]= 2063024031;
assign addr[33102]= 2015345591;
assign addr[33103]= 1957443913;
assign addr[33104]= 1889612716;
assign addr[33105]= 1812196087;
assign addr[33106]= 1725586737;
assign addr[33107]= 1630224009;
assign addr[33108]= 1526591649;
assign addr[33109]= 1415215352;
assign addr[33110]= 1296660098;
assign addr[33111]= 1171527280;
assign addr[33112]= 1040451659;
assign addr[33113]= 904098143;
assign addr[33114]= 763158411;
assign addr[33115]= 618347408;
assign addr[33116]= 470399716;
assign addr[33117]= 320065829;
assign addr[33118]= 168108346;
assign addr[33119]= 15298099;
assign addr[33120]= -137589750;
assign addr[33121]= -289779648;
assign addr[33122]= -440499581;
assign addr[33123]= -588984994;
assign addr[33124]= -734482665;
assign addr[33125]= -876254528;
assign addr[33126]= -1013581418;
assign addr[33127]= -1145766716;
assign addr[33128]= -1272139887;
assign addr[33129]= -1392059879;
assign addr[33130]= -1504918373;
assign addr[33131]= -1610142873;
assign addr[33132]= -1707199606;
assign addr[33133]= -1795596234;
assign addr[33134]= -1874884346;
assign addr[33135]= -1944661739;
assign addr[33136]= -2004574453;
assign addr[33137]= -2054318569;
assign addr[33138]= -2093641749;
assign addr[33139]= -2122344521;
assign addr[33140]= -2140281282;
assign addr[33141]= -2147361045;
assign addr[33142]= -2143547897;
assign addr[33143]= -2128861181;
assign addr[33144]= -2103375398;
assign addr[33145]= -2067219829;
assign addr[33146]= -2020577882;
assign addr[33147]= -1963686155;
assign addr[33148]= -1896833245;
assign addr[33149]= -1820358275;
assign addr[33150]= -1734649179;
assign addr[33151]= -1640140734;
assign addr[33152]= -1537312353;
assign addr[33153]= -1426685652;
assign addr[33154]= -1308821808;
assign addr[33155]= -1184318708;
assign addr[33156]= -1053807919;
assign addr[33157]= -917951481;
assign addr[33158]= -777438554;
assign addr[33159]= -632981917;
assign addr[33160]= -485314355;
assign addr[33161]= -335184940;
assign addr[33162]= -183355234;
assign addr[33163]= -30595422;
assign addr[33164]= 122319591;
assign addr[33165]= 274614114;
assign addr[33166]= 425515602;
assign addr[33167]= 574258580;
assign addr[33168]= 720088517;
assign addr[33169]= 862265664;
assign addr[33170]= 1000068799;
assign addr[33171]= 1132798888;
assign addr[33172]= 1259782632;
assign addr[33173]= 1380375881;
assign addr[33174]= 1493966902;
assign addr[33175]= 1599979481;
assign addr[33176]= 1697875851;
assign addr[33177]= 1787159411;
assign addr[33178]= 1867377253;
assign addr[33179]= 1938122457;
assign addr[33180]= 1999036154;
assign addr[33181]= 2049809346;
assign addr[33182]= 2090184478;
assign addr[33183]= 2119956737;
assign addr[33184]= 2138975100;
assign addr[33185]= 2147143090;
assign addr[33186]= 2144419275;
assign addr[33187]= 2130817471;
assign addr[33188]= 2106406677;
assign addr[33189]= 2071310720;
assign addr[33190]= 2025707632;
assign addr[33191]= 1969828744;
assign addr[33192]= 1903957513;
assign addr[33193]= 1828428082;
assign addr[33194]= 1743623590;
assign addr[33195]= 1649974225;
assign addr[33196]= 1547955041;
assign addr[33197]= 1438083551;
assign addr[33198]= 1320917099;
assign addr[33199]= 1197050035;
assign addr[33200]= 1067110699;
assign addr[33201]= 931758235;
assign addr[33202]= 791679244;
assign addr[33203]= 647584304;
assign addr[33204]= 500204365;
assign addr[33205]= 350287041;
assign addr[33206]= 198592817;
assign addr[33207]= 45891193;
assign addr[33208]= -107043224;
assign addr[33209]= -259434643;
assign addr[33210]= -410510029;
assign addr[33211]= -559503022;
assign addr[33212]= -705657826;
assign addr[33213]= -848233042;
assign addr[33214]= -986505429;
assign addr[33215]= -1119773573;
assign addr[33216]= -1247361445;
assign addr[33217]= -1368621831;
assign addr[33218]= -1482939614;
assign addr[33219]= -1589734894;
assign addr[33220]= -1688465931;
assign addr[33221]= -1778631892;
assign addr[33222]= -1859775393;
assign addr[33223]= -1931484818;
assign addr[33224]= -1993396407;
assign addr[33225]= -2045196100;
assign addr[33226]= -2086621133;
assign addr[33227]= -2117461370;
assign addr[33228]= -2137560369;
assign addr[33229]= -2146816171;
assign addr[33230]= -2145181827;
assign addr[33231]= -2132665626;
assign addr[33232]= -2109331059;
assign addr[33233]= -2075296495;
assign addr[33234]= -2030734582;
assign addr[33235]= -1975871368;
assign addr[33236]= -1910985158;
assign addr[33237]= -1836405100;
assign addr[33238]= -1752509516;
assign addr[33239]= -1659723983;
assign addr[33240]= -1558519173;
assign addr[33241]= -1449408469;
assign addr[33242]= -1332945355;
assign addr[33243]= -1209720613;
assign addr[33244]= -1080359326;
assign addr[33245]= -945517704;
assign addr[33246]= -805879757;
assign addr[33247]= -662153826;
assign addr[33248]= -515068990;
assign addr[33249]= -365371365;
assign addr[33250]= -213820322;
assign addr[33251]= -61184634;
assign addr[33252]= 91761426;
assign addr[33253]= 244242007;
assign addr[33254]= 395483624;
assign addr[33255]= 544719071;
assign addr[33256]= 691191324;
assign addr[33257]= 834157373;
assign addr[33258]= 972891995;
assign addr[33259]= 1106691431;
assign addr[33260]= 1234876957;
assign addr[33261]= 1356798326;
assign addr[33262]= 1471837070;
assign addr[33263]= 1579409630;
assign addr[33264]= 1678970324;
assign addr[33265]= 1770014111;
assign addr[33266]= 1852079154;
assign addr[33267]= 1924749160;
assign addr[33268]= 1987655498;
assign addr[33269]= 2040479063;
assign addr[33270]= 2082951896;
assign addr[33271]= 2114858546;
assign addr[33272]= 2136037160;
assign addr[33273]= 2146380306;
assign addr[33274]= 2145835515;
assign addr[33275]= 2134405552;
assign addr[33276]= 2112148396;
assign addr[33277]= 2079176953;
assign addr[33278]= 2035658475;
assign addr[33279]= 1981813720;
assign addr[33280]= 1917915825;
assign addr[33281]= 1844288924;
assign addr[33282]= 1761306505;
assign addr[33283]= 1669389513;
assign addr[33284]= 1569004214;
assign addr[33285]= 1460659832;
assign addr[33286]= 1344905966;
assign addr[33287]= 1222329801;
assign addr[33288]= 1093553126;
assign addr[33289]= 959229189;
assign addr[33290]= 820039373;
assign addr[33291]= 676689746;
assign addr[33292]= 529907477;
assign addr[33293]= 380437148;
assign addr[33294]= 229036977;
assign addr[33295]= 76474970;
assign addr[33296]= -76474970;
assign addr[33297]= -229036977;
assign addr[33298]= -380437148;
assign addr[33299]= -529907477;
assign addr[33300]= -676689746;
assign addr[33301]= -820039373;
assign addr[33302]= -959229189;
assign addr[33303]= -1093553126;
assign addr[33304]= -1222329801;
assign addr[33305]= -1344905966;
assign addr[33306]= -1460659832;
assign addr[33307]= -1569004214;
assign addr[33308]= -1669389513;
assign addr[33309]= -1761306505;
assign addr[33310]= -1844288924;
assign addr[33311]= -1917915825;
assign addr[33312]= -1981813720;
assign addr[33313]= -2035658475;
assign addr[33314]= -2079176953;
assign addr[33315]= -2112148396;
assign addr[33316]= -2134405552;
assign addr[33317]= -2145835515;
assign addr[33318]= -2146380306;
assign addr[33319]= -2136037160;
assign addr[33320]= -2114858546;
assign addr[33321]= -2082951896;
assign addr[33322]= -2040479063;
assign addr[33323]= -1987655498;
assign addr[33324]= -1924749160;
assign addr[33325]= -1852079154;
assign addr[33326]= -1770014111;
assign addr[33327]= -1678970324;
assign addr[33328]= -1579409630;
assign addr[33329]= -1471837070;
assign addr[33330]= -1356798326;
assign addr[33331]= -1234876957;
assign addr[33332]= -1106691431;
assign addr[33333]= -972891995;
assign addr[33334]= -834157373;
assign addr[33335]= -691191324;
assign addr[33336]= -544719071;
assign addr[33337]= -395483624;
assign addr[33338]= -244242007;
assign addr[33339]= -91761426;
assign addr[33340]= 61184634;
assign addr[33341]= 213820322;
assign addr[33342]= 365371365;
assign addr[33343]= 515068990;
assign addr[33344]= 662153826;
assign addr[33345]= 805879757;
assign addr[33346]= 945517704;
assign addr[33347]= 1080359326;
assign addr[33348]= 1209720613;
assign addr[33349]= 1332945355;
assign addr[33350]= 1449408469;
assign addr[33351]= 1558519173;
assign addr[33352]= 1659723983;
assign addr[33353]= 1752509516;
assign addr[33354]= 1836405100;
assign addr[33355]= 1910985158;
assign addr[33356]= 1975871368;
assign addr[33357]= 2030734582;
assign addr[33358]= 2075296495;
assign addr[33359]= 2109331059;
assign addr[33360]= 2132665626;
assign addr[33361]= 2145181827;
assign addr[33362]= 2146816171;
assign addr[33363]= 2137560369;
assign addr[33364]= 2117461370;
assign addr[33365]= 2086621133;
assign addr[33366]= 2045196100;
assign addr[33367]= 1993396407;
assign addr[33368]= 1931484818;
assign addr[33369]= 1859775393;
assign addr[33370]= 1778631892;
assign addr[33371]= 1688465931;
assign addr[33372]= 1589734894;
assign addr[33373]= 1482939614;
assign addr[33374]= 1368621831;
assign addr[33375]= 1247361445;
assign addr[33376]= 1119773573;
assign addr[33377]= 986505429;
assign addr[33378]= 848233042;
assign addr[33379]= 705657826;
assign addr[33380]= 559503022;
assign addr[33381]= 410510029;
assign addr[33382]= 259434643;
assign addr[33383]= 107043224;
assign addr[33384]= -45891193;
assign addr[33385]= -198592817;
assign addr[33386]= -350287041;
assign addr[33387]= -500204365;
assign addr[33388]= -647584304;
assign addr[33389]= -791679244;
assign addr[33390]= -931758235;
assign addr[33391]= -1067110699;
assign addr[33392]= -1197050035;
assign addr[33393]= -1320917099;
assign addr[33394]= -1438083551;
assign addr[33395]= -1547955041;
assign addr[33396]= -1649974225;
assign addr[33397]= -1743623590;
assign addr[33398]= -1828428082;
assign addr[33399]= -1903957513;
assign addr[33400]= -1969828744;
assign addr[33401]= -2025707632;
assign addr[33402]= -2071310720;
assign addr[33403]= -2106406677;
assign addr[33404]= -2130817471;
assign addr[33405]= -2144419275;
assign addr[33406]= -2147143090;
assign addr[33407]= -2138975100;
assign addr[33408]= -2119956737;
assign addr[33409]= -2090184478;
assign addr[33410]= -2049809346;
assign addr[33411]= -1999036154;
assign addr[33412]= -1938122457;
assign addr[33413]= -1867377253;
assign addr[33414]= -1787159411;
assign addr[33415]= -1697875851;
assign addr[33416]= -1599979481;
assign addr[33417]= -1493966902;
assign addr[33418]= -1380375881;
assign addr[33419]= -1259782632;
assign addr[33420]= -1132798888;
assign addr[33421]= -1000068799;
assign addr[33422]= -862265664;
assign addr[33423]= -720088517;
assign addr[33424]= -574258580;
assign addr[33425]= -425515602;
assign addr[33426]= -274614114;
assign addr[33427]= -122319591;
assign addr[33428]= 30595422;
assign addr[33429]= 183355234;
assign addr[33430]= 335184940;
assign addr[33431]= 485314355;
assign addr[33432]= 632981917;
assign addr[33433]= 777438554;
assign addr[33434]= 917951481;
assign addr[33435]= 1053807919;
assign addr[33436]= 1184318708;
assign addr[33437]= 1308821808;
assign addr[33438]= 1426685652;
assign addr[33439]= 1537312353;
assign addr[33440]= 1640140734;
assign addr[33441]= 1734649179;
assign addr[33442]= 1820358275;
assign addr[33443]= 1896833245;
assign addr[33444]= 1963686155;
assign addr[33445]= 2020577882;
assign addr[33446]= 2067219829;
assign addr[33447]= 2103375398;
assign addr[33448]= 2128861181;
assign addr[33449]= 2143547897;
assign addr[33450]= 2147361045;
assign addr[33451]= 2140281282;
assign addr[33452]= 2122344521;
assign addr[33453]= 2093641749;
assign addr[33454]= 2054318569;
assign addr[33455]= 2004574453;
assign addr[33456]= 1944661739;
assign addr[33457]= 1874884346;
assign addr[33458]= 1795596234;
assign addr[33459]= 1707199606;
assign addr[33460]= 1610142873;
assign addr[33461]= 1504918373;
assign addr[33462]= 1392059879;
assign addr[33463]= 1272139887;
assign addr[33464]= 1145766716;
assign addr[33465]= 1013581418;
assign addr[33466]= 876254528;
assign addr[33467]= 734482665;
assign addr[33468]= 588984994;
assign addr[33469]= 440499581;
assign addr[33470]= 289779648;
assign addr[33471]= 137589750;
assign addr[33472]= -15298099;
assign addr[33473]= -168108346;
assign addr[33474]= -320065829;
assign addr[33475]= -470399716;
assign addr[33476]= -618347408;
assign addr[33477]= -763158411;
assign addr[33478]= -904098143;
assign addr[33479]= -1040451659;
assign addr[33480]= -1171527280;
assign addr[33481]= -1296660098;
assign addr[33482]= -1415215352;
assign addr[33483]= -1526591649;
assign addr[33484]= -1630224009;
assign addr[33485]= -1725586737;
assign addr[33486]= -1812196087;
assign addr[33487]= -1889612716;
assign addr[33488]= -1957443913;
assign addr[33489]= -2015345591;
assign addr[33490]= -2063024031;
assign addr[33491]= -2100237377;
assign addr[33492]= -2126796855;
assign addr[33493]= -2142567738;
assign addr[33494]= -2147470025;
assign addr[33495]= -2141478848;
assign addr[33496]= -2124624598;
assign addr[33497]= -2096992772;
assign addr[33498]= -2058723538;
assign addr[33499]= -2010011024;
assign addr[33500]= -1951102334;
assign addr[33501]= -1882296293;
assign addr[33502]= -1803941934;
assign addr[33503]= -1716436725;
assign addr[33504]= -1620224553;
assign addr[33505]= -1515793473;
assign addr[33506]= -1403673233;
assign addr[33507]= -1284432584;
assign addr[33508]= -1158676398;
assign addr[33509]= -1027042599;
assign addr[33510]= -890198924;
assign addr[33511]= -748839539;
assign addr[33512]= -603681519;
assign addr[33513]= -455461206;
assign addr[33514]= -304930476;
assign addr[33515]= -152852926;
assign addr[33516]= 0;
assign addr[33517]= 152852926;
assign addr[33518]= 304930476;
assign addr[33519]= 455461206;
assign addr[33520]= 603681519;
assign addr[33521]= 748839539;
assign addr[33522]= 890198924;
assign addr[33523]= 1027042599;
assign addr[33524]= 1158676398;
assign addr[33525]= 1284432584;
assign addr[33526]= 1403673233;
assign addr[33527]= 1515793473;
assign addr[33528]= 1620224553;
assign addr[33529]= 1716436725;
assign addr[33530]= 1803941934;
assign addr[33531]= 1882296293;
assign addr[33532]= 1951102334;
assign addr[33533]= 2010011024;
assign addr[33534]= 2058723538;
assign addr[33535]= 2096992772;
assign addr[33536]= 2124624598;
assign addr[33537]= 2141478848;
assign addr[33538]= 2147470025;
assign addr[33539]= 2142567738;
assign addr[33540]= 2126796855;
assign addr[33541]= 2100237377;
assign addr[33542]= 2063024031;
assign addr[33543]= 2015345591;
assign addr[33544]= 1957443913;
assign addr[33545]= 1889612716;
assign addr[33546]= 1812196087;
assign addr[33547]= 1725586737;
assign addr[33548]= 1630224009;
assign addr[33549]= 1526591649;
assign addr[33550]= 1415215352;
assign addr[33551]= 1296660098;
assign addr[33552]= 1171527280;
assign addr[33553]= 1040451659;
assign addr[33554]= 904098143;
assign addr[33555]= 763158411;
assign addr[33556]= 618347408;
assign addr[33557]= 470399716;
assign addr[33558]= 320065829;
assign addr[33559]= 168108346;
assign addr[33560]= 15298099;
assign addr[33561]= -137589750;
assign addr[33562]= -289779648;
assign addr[33563]= -440499581;
assign addr[33564]= -588984994;
assign addr[33565]= -734482665;
assign addr[33566]= -876254528;
assign addr[33567]= -1013581418;
assign addr[33568]= -1145766716;
assign addr[33569]= -1272139887;
assign addr[33570]= -1392059879;
assign addr[33571]= -1504918373;
assign addr[33572]= -1610142873;
assign addr[33573]= -1707199606;
assign addr[33574]= -1795596234;
assign addr[33575]= -1874884346;
assign addr[33576]= -1944661739;
assign addr[33577]= -2004574453;
assign addr[33578]= -2054318569;
assign addr[33579]= -2093641749;
assign addr[33580]= -2122344521;
assign addr[33581]= -2140281282;
assign addr[33582]= -2147361045;
assign addr[33583]= -2143547897;
assign addr[33584]= -2128861181;
assign addr[33585]= -2103375398;
assign addr[33586]= -2067219829;
assign addr[33587]= -2020577882;
assign addr[33588]= -1963686155;
assign addr[33589]= -1896833245;
assign addr[33590]= -1820358275;
assign addr[33591]= -1734649179;
assign addr[33592]= -1640140734;
assign addr[33593]= -1537312353;
assign addr[33594]= -1426685652;
assign addr[33595]= -1308821808;
assign addr[33596]= -1184318708;
assign addr[33597]= -1053807919;
assign addr[33598]= -917951481;
assign addr[33599]= -777438554;
assign addr[33600]= -632981917;
assign addr[33601]= -485314355;
assign addr[33602]= -335184940;
assign addr[33603]= -183355234;
assign addr[33604]= -30595422;
assign addr[33605]= 122319591;
assign addr[33606]= 274614114;
assign addr[33607]= 425515602;
assign addr[33608]= 574258580;
assign addr[33609]= 720088517;
assign addr[33610]= 862265664;
assign addr[33611]= 1000068799;
assign addr[33612]= 1132798888;
assign addr[33613]= 1259782632;
assign addr[33614]= 1380375881;
assign addr[33615]= 1493966902;
assign addr[33616]= 1599979481;
assign addr[33617]= 1697875851;
assign addr[33618]= 1787159411;
assign addr[33619]= 1867377253;
assign addr[33620]= 1938122457;
assign addr[33621]= 1999036154;
assign addr[33622]= 2049809346;
assign addr[33623]= 2090184478;
assign addr[33624]= 2119956737;
assign addr[33625]= 2138975100;
assign addr[33626]= 2147143090;
assign addr[33627]= 2144419275;
assign addr[33628]= 2130817471;
assign addr[33629]= 2106406677;
assign addr[33630]= 2071310720;
assign addr[33631]= 2025707632;
assign addr[33632]= 1969828744;
assign addr[33633]= 1903957513;
assign addr[33634]= 1828428082;
assign addr[33635]= 1743623590;
assign addr[33636]= 1649974225;
assign addr[33637]= 1547955041;
assign addr[33638]= 1438083551;
assign addr[33639]= 1320917099;
assign addr[33640]= 1197050035;
assign addr[33641]= 1067110699;
assign addr[33642]= 931758235;
assign addr[33643]= 791679244;
assign addr[33644]= 647584304;
assign addr[33645]= 500204365;
assign addr[33646]= 350287041;
assign addr[33647]= 198592817;
assign addr[33648]= 45891193;
assign addr[33649]= -107043224;
assign addr[33650]= -259434643;
assign addr[33651]= -410510029;
assign addr[33652]= -559503022;
assign addr[33653]= -705657826;
assign addr[33654]= -848233042;
assign addr[33655]= -986505429;
assign addr[33656]= -1119773573;
assign addr[33657]= -1247361445;
assign addr[33658]= -1368621831;
assign addr[33659]= -1482939614;
assign addr[33660]= -1589734894;
assign addr[33661]= -1688465931;
assign addr[33662]= -1778631892;
assign addr[33663]= -1859775393;
assign addr[33664]= -1931484818;
assign addr[33665]= -1993396407;
assign addr[33666]= -2045196100;
assign addr[33667]= -2086621133;
assign addr[33668]= -2117461370;
assign addr[33669]= -2137560369;
assign addr[33670]= -2146816171;
assign addr[33671]= -2145181827;
assign addr[33672]= -2132665626;
assign addr[33673]= -2109331059;
assign addr[33674]= -2075296495;
assign addr[33675]= -2030734582;
assign addr[33676]= -1975871368;
assign addr[33677]= -1910985158;
assign addr[33678]= -1836405100;
assign addr[33679]= -1752509516;
assign addr[33680]= -1659723983;
assign addr[33681]= -1558519173;
assign addr[33682]= -1449408469;
assign addr[33683]= -1332945355;
assign addr[33684]= -1209720613;
assign addr[33685]= -1080359326;
assign addr[33686]= -945517704;
assign addr[33687]= -805879757;
assign addr[33688]= -662153826;
assign addr[33689]= -515068990;
assign addr[33690]= -365371365;
assign addr[33691]= -213820322;
assign addr[33692]= -61184634;
assign addr[33693]= 91761426;
assign addr[33694]= 244242007;
assign addr[33695]= 395483624;
assign addr[33696]= 544719071;
assign addr[33697]= 691191324;
assign addr[33698]= 834157373;
assign addr[33699]= 972891995;
assign addr[33700]= 1106691431;
assign addr[33701]= 1234876957;
assign addr[33702]= 1356798326;
assign addr[33703]= 1471837070;
assign addr[33704]= 1579409630;
assign addr[33705]= 1678970324;
assign addr[33706]= 1770014111;
assign addr[33707]= 1852079154;
assign addr[33708]= 1924749160;
assign addr[33709]= 1987655498;
assign addr[33710]= 2040479063;
assign addr[33711]= 2082951896;
assign addr[33712]= 2114858546;
assign addr[33713]= 2136037160;
assign addr[33714]= 2146380306;
assign addr[33715]= 2145835515;
assign addr[33716]= 2134405552;
assign addr[33717]= 2112148396;
assign addr[33718]= 2079176953;
assign addr[33719]= 2035658475;
assign addr[33720]= 1981813720;
assign addr[33721]= 1917915825;
assign addr[33722]= 1844288924;
assign addr[33723]= 1761306505;
assign addr[33724]= 1669389513;
assign addr[33725]= 1569004214;
assign addr[33726]= 1460659832;
assign addr[33727]= 1344905966;
assign addr[33728]= 1222329801;
assign addr[33729]= 1093553126;
assign addr[33730]= 959229189;
assign addr[33731]= 820039373;
assign addr[33732]= 676689746;
assign addr[33733]= 529907477;
assign addr[33734]= 380437148;
assign addr[33735]= 229036977;
assign addr[33736]= 76474970;
assign addr[33737]= -76474970;
assign addr[33738]= -229036977;
assign addr[33739]= -380437148;
assign addr[33740]= -529907477;
assign addr[33741]= -676689746;
assign addr[33742]= -820039373;
assign addr[33743]= -959229189;
assign addr[33744]= -1093553126;
assign addr[33745]= -1222329801;
assign addr[33746]= -1344905966;
assign addr[33747]= -1460659832;
assign addr[33748]= -1569004214;
assign addr[33749]= -1669389513;
assign addr[33750]= -1761306505;
assign addr[33751]= -1844288924;
assign addr[33752]= -1917915825;
assign addr[33753]= -1981813720;
assign addr[33754]= -2035658475;
assign addr[33755]= -2079176953;
assign addr[33756]= -2112148396;
assign addr[33757]= -2134405552;
assign addr[33758]= -2145835515;
assign addr[33759]= -2146380306;
assign addr[33760]= -2136037160;
assign addr[33761]= -2114858546;
assign addr[33762]= -2082951896;
assign addr[33763]= -2040479063;
assign addr[33764]= -1987655498;
assign addr[33765]= -1924749160;
assign addr[33766]= -1852079154;
assign addr[33767]= -1770014111;
assign addr[33768]= -1678970324;
assign addr[33769]= -1579409630;
assign addr[33770]= -1471837070;
assign addr[33771]= -1356798326;
assign addr[33772]= -1234876957;
assign addr[33773]= -1106691431;
assign addr[33774]= -972891995;
assign addr[33775]= -834157373;
assign addr[33776]= -691191324;
assign addr[33777]= -544719071;
assign addr[33778]= -395483624;
assign addr[33779]= -244242007;
assign addr[33780]= -91761426;
assign addr[33781]= 61184634;
assign addr[33782]= 213820322;
assign addr[33783]= 365371365;
assign addr[33784]= 515068990;
assign addr[33785]= 662153826;
assign addr[33786]= 805879757;
assign addr[33787]= 945517704;
assign addr[33788]= 1080359326;
assign addr[33789]= 1209720613;
assign addr[33790]= 1332945355;
assign addr[33791]= 1449408469;
assign addr[33792]= 1558519173;
assign addr[33793]= 1659723983;
assign addr[33794]= 1752509516;
assign addr[33795]= 1836405100;
assign addr[33796]= 1910985158;
assign addr[33797]= 1975871368;
assign addr[33798]= 2030734582;
assign addr[33799]= 2075296495;
assign addr[33800]= 2109331059;
assign addr[33801]= 2132665626;
assign addr[33802]= 2145181827;
assign addr[33803]= 2146816171;
assign addr[33804]= 2137560369;
assign addr[33805]= 2117461370;
assign addr[33806]= 2086621133;
assign addr[33807]= 2045196100;
assign addr[33808]= 1993396407;
assign addr[33809]= 1931484818;
assign addr[33810]= 1859775393;
assign addr[33811]= 1778631892;
assign addr[33812]= 1688465931;
assign addr[33813]= 1589734894;
assign addr[33814]= 1482939614;
assign addr[33815]= 1368621831;
assign addr[33816]= 1247361445;
assign addr[33817]= 1119773573;
assign addr[33818]= 986505429;
assign addr[33819]= 848233042;
assign addr[33820]= 705657826;
assign addr[33821]= 559503022;
assign addr[33822]= 410510029;
assign addr[33823]= 259434643;
assign addr[33824]= 107043224;
assign addr[33825]= -45891193;
assign addr[33826]= -198592817;
assign addr[33827]= -350287041;
assign addr[33828]= -500204365;
assign addr[33829]= -647584304;
assign addr[33830]= -791679244;
assign addr[33831]= -931758235;
assign addr[33832]= -1067110699;
assign addr[33833]= -1197050035;
assign addr[33834]= -1320917099;
assign addr[33835]= -1438083551;
assign addr[33836]= -1547955041;
assign addr[33837]= -1649974225;
assign addr[33838]= -1743623590;
assign addr[33839]= -1828428082;
assign addr[33840]= -1903957513;
assign addr[33841]= -1969828744;
assign addr[33842]= -2025707632;
assign addr[33843]= -2071310720;
assign addr[33844]= -2106406677;
assign addr[33845]= -2130817471;
assign addr[33846]= -2144419275;
assign addr[33847]= -2147143090;
assign addr[33848]= -2138975100;
assign addr[33849]= -2119956737;
assign addr[33850]= -2090184478;
assign addr[33851]= -2049809346;
assign addr[33852]= -1999036154;
assign addr[33853]= -1938122457;
assign addr[33854]= -1867377253;
assign addr[33855]= -1787159411;
assign addr[33856]= -1697875851;
assign addr[33857]= -1599979481;
assign addr[33858]= -1493966902;
assign addr[33859]= -1380375881;
assign addr[33860]= -1259782632;
assign addr[33861]= -1132798888;
assign addr[33862]= -1000068799;
assign addr[33863]= -862265664;
assign addr[33864]= -720088517;
assign addr[33865]= -574258580;
assign addr[33866]= -425515602;
assign addr[33867]= -274614114;
assign addr[33868]= -122319591;
assign addr[33869]= 30595422;
assign addr[33870]= 183355234;
assign addr[33871]= 335184940;
assign addr[33872]= 485314355;
assign addr[33873]= 632981917;
assign addr[33874]= 777438554;
assign addr[33875]= 917951481;
assign addr[33876]= 1053807919;
assign addr[33877]= 1184318708;
assign addr[33878]= 1308821808;
assign addr[33879]= 1426685652;
assign addr[33880]= 1537312353;
assign addr[33881]= 1640140734;
assign addr[33882]= 1734649179;
assign addr[33883]= 1820358275;
assign addr[33884]= 1896833245;
assign addr[33885]= 1963686155;
assign addr[33886]= 2020577882;
assign addr[33887]= 2067219829;
assign addr[33888]= 2103375398;
assign addr[33889]= 2128861181;
assign addr[33890]= 2143547897;
assign addr[33891]= 2147361045;
assign addr[33892]= 2140281282;
assign addr[33893]= 2122344521;
assign addr[33894]= 2093641749;
assign addr[33895]= 2054318569;
assign addr[33896]= 2004574453;
assign addr[33897]= 1944661739;
assign addr[33898]= 1874884346;
assign addr[33899]= 1795596234;
assign addr[33900]= 1707199606;
assign addr[33901]= 1610142873;
assign addr[33902]= 1504918373;
assign addr[33903]= 1392059879;
assign addr[33904]= 1272139887;
assign addr[33905]= 1145766716;
assign addr[33906]= 1013581418;
assign addr[33907]= 876254528;
assign addr[33908]= 734482665;
assign addr[33909]= 588984994;
assign addr[33910]= 440499581;
assign addr[33911]= 289779648;
assign addr[33912]= 137589750;
assign addr[33913]= -15298099;
assign addr[33914]= -168108346;
assign addr[33915]= -320065829;
assign addr[33916]= -470399716;
assign addr[33917]= -618347408;
assign addr[33918]= -763158411;
assign addr[33919]= -904098143;
assign addr[33920]= -1040451659;
assign addr[33921]= -1171527280;
assign addr[33922]= -1296660098;
assign addr[33923]= -1415215352;
assign addr[33924]= -1526591649;
assign addr[33925]= -1630224009;
assign addr[33926]= -1725586737;
assign addr[33927]= -1812196087;
assign addr[33928]= -1889612716;
assign addr[33929]= -1957443913;
assign addr[33930]= -2015345591;
assign addr[33931]= -2063024031;
assign addr[33932]= -2100237377;
assign addr[33933]= -2126796855;
assign addr[33934]= -2142567738;
assign addr[33935]= -2147470025;
assign addr[33936]= -2141478848;
assign addr[33937]= -2124624598;
assign addr[33938]= -2096992772;
assign addr[33939]= -2058723538;
assign addr[33940]= -2010011024;
assign addr[33941]= -1951102334;
assign addr[33942]= -1882296293;
assign addr[33943]= -1803941934;
assign addr[33944]= -1716436725;
assign addr[33945]= -1620224553;
assign addr[33946]= -1515793473;
assign addr[33947]= -1403673233;
assign addr[33948]= -1284432584;
assign addr[33949]= -1158676398;
assign addr[33950]= -1027042599;
assign addr[33951]= -890198924;
assign addr[33952]= -748839539;
assign addr[33953]= -603681519;
assign addr[33954]= -455461206;
assign addr[33955]= -304930476;
assign addr[33956]= -152852926;
assign addr[33957]= 0;
assign addr[33958]= 152852926;
assign addr[33959]= 304930476;
assign addr[33960]= 455461206;
assign addr[33961]= 603681519;
assign addr[33962]= 748839539;
assign addr[33963]= 890198924;
assign addr[33964]= 1027042599;
assign addr[33965]= 1158676398;
assign addr[33966]= 1284432584;
assign addr[33967]= 1403673233;
assign addr[33968]= 1515793473;
assign addr[33969]= 1620224553;
assign addr[33970]= 1716436725;
assign addr[33971]= 1803941934;
assign addr[33972]= 1882296293;
assign addr[33973]= 1951102334;
assign addr[33974]= 2010011024;
assign addr[33975]= 2058723538;
assign addr[33976]= 2096992772;
assign addr[33977]= 2124624598;
assign addr[33978]= 2141478848;
assign addr[33979]= 2147470025;
assign addr[33980]= 2142567738;
assign addr[33981]= 2126796855;
assign addr[33982]= 2100237377;
assign addr[33983]= 2063024031;
assign addr[33984]= 2015345591;
assign addr[33985]= 1957443913;
assign addr[33986]= 1889612716;
assign addr[33987]= 1812196087;
assign addr[33988]= 1725586737;
assign addr[33989]= 1630224009;
assign addr[33990]= 1526591649;
assign addr[33991]= 1415215352;
assign addr[33992]= 1296660098;
assign addr[33993]= 1171527280;
assign addr[33994]= 1040451659;
assign addr[33995]= 904098143;
assign addr[33996]= 763158411;
assign addr[33997]= 618347408;
assign addr[33998]= 470399716;
assign addr[33999]= 320065829;
assign addr[34000]= 168108346;
assign addr[34001]= 15298099;
assign addr[34002]= -137589750;
assign addr[34003]= -289779648;
assign addr[34004]= -440499581;
assign addr[34005]= -588984994;
assign addr[34006]= -734482665;
assign addr[34007]= -876254528;
assign addr[34008]= -1013581418;
assign addr[34009]= -1145766716;
assign addr[34010]= -1272139887;
assign addr[34011]= -1392059879;
assign addr[34012]= -1504918373;
assign addr[34013]= -1610142873;
assign addr[34014]= -1707199606;
assign addr[34015]= -1795596234;
assign addr[34016]= -1874884346;
assign addr[34017]= -1944661739;
assign addr[34018]= -2004574453;
assign addr[34019]= -2054318569;
assign addr[34020]= -2093641749;
assign addr[34021]= -2122344521;
assign addr[34022]= -2140281282;
assign addr[34023]= -2147361045;
assign addr[34024]= -2143547897;
assign addr[34025]= -2128861181;
assign addr[34026]= -2103375398;
assign addr[34027]= -2067219829;
assign addr[34028]= -2020577882;
assign addr[34029]= -1963686155;
assign addr[34030]= -1896833245;
assign addr[34031]= -1820358275;
assign addr[34032]= -1734649179;
assign addr[34033]= -1640140734;
assign addr[34034]= -1537312353;
assign addr[34035]= -1426685652;
assign addr[34036]= -1308821808;
assign addr[34037]= -1184318708;
assign addr[34038]= -1053807919;
assign addr[34039]= -917951481;
assign addr[34040]= -777438554;
assign addr[34041]= -632981917;
assign addr[34042]= -485314355;
assign addr[34043]= -335184940;
assign addr[34044]= -183355234;
assign addr[34045]= -30595422;
assign addr[34046]= 122319591;
assign addr[34047]= 274614114;
assign addr[34048]= 425515602;
assign addr[34049]= 574258580;
assign addr[34050]= 720088517;
assign addr[34051]= 862265664;
assign addr[34052]= 1000068799;
assign addr[34053]= 1132798888;
assign addr[34054]= 1259782632;
assign addr[34055]= 1380375881;
assign addr[34056]= 1493966902;
assign addr[34057]= 1599979481;
assign addr[34058]= 1697875851;
assign addr[34059]= 1787159411;
assign addr[34060]= 1867377253;
assign addr[34061]= 1938122457;
assign addr[34062]= 1999036154;
assign addr[34063]= 2049809346;
assign addr[34064]= 2090184478;
assign addr[34065]= 2119956737;
assign addr[34066]= 2138975100;
assign addr[34067]= 2147143090;
assign addr[34068]= 2144419275;
assign addr[34069]= 2130817471;
assign addr[34070]= 2106406677;
assign addr[34071]= 2071310720;
assign addr[34072]= 2025707632;
assign addr[34073]= 1969828744;
assign addr[34074]= 1903957513;
assign addr[34075]= 1828428082;
assign addr[34076]= 1743623590;
assign addr[34077]= 1649974225;
assign addr[34078]= 1547955041;
assign addr[34079]= 1438083551;
assign addr[34080]= 1320917099;
assign addr[34081]= 1197050035;
assign addr[34082]= 1067110699;
assign addr[34083]= 931758235;
assign addr[34084]= 791679244;
assign addr[34085]= 647584304;
assign addr[34086]= 500204365;
assign addr[34087]= 350287041;
assign addr[34088]= 198592817;
assign addr[34089]= 45891193;
assign addr[34090]= -107043224;
assign addr[34091]= -259434643;
assign addr[34092]= -410510029;
assign addr[34093]= -559503022;
assign addr[34094]= -705657826;
assign addr[34095]= -848233042;
assign addr[34096]= -986505429;
assign addr[34097]= -1119773573;
assign addr[34098]= -1247361445;
assign addr[34099]= -1368621831;
assign addr[34100]= -1482939614;
assign addr[34101]= -1589734894;
assign addr[34102]= -1688465931;
assign addr[34103]= -1778631892;
assign addr[34104]= -1859775393;
assign addr[34105]= -1931484818;
assign addr[34106]= -1993396407;
assign addr[34107]= -2045196100;
assign addr[34108]= -2086621133;
assign addr[34109]= -2117461370;
assign addr[34110]= -2137560369;
assign addr[34111]= -2146816171;
assign addr[34112]= -2145181827;
assign addr[34113]= -2132665626;
assign addr[34114]= -2109331059;
assign addr[34115]= -2075296495;
assign addr[34116]= -2030734582;
assign addr[34117]= -1975871368;
assign addr[34118]= -1910985158;
assign addr[34119]= -1836405100;
assign addr[34120]= -1752509516;
assign addr[34121]= -1659723983;
assign addr[34122]= -1558519173;
assign addr[34123]= -1449408469;
assign addr[34124]= -1332945355;
assign addr[34125]= -1209720613;
assign addr[34126]= -1080359326;
assign addr[34127]= -945517704;
assign addr[34128]= -805879757;
assign addr[34129]= -662153826;
assign addr[34130]= -515068990;
assign addr[34131]= -365371365;
assign addr[34132]= -213820322;
assign addr[34133]= -61184634;
assign addr[34134]= 91761426;
assign addr[34135]= 244242007;
assign addr[34136]= 395483624;
assign addr[34137]= 544719071;
assign addr[34138]= 691191324;
assign addr[34139]= 834157373;
assign addr[34140]= 972891995;
assign addr[34141]= 1106691431;
assign addr[34142]= 1234876957;
assign addr[34143]= 1356798326;
assign addr[34144]= 1471837070;
assign addr[34145]= 1579409630;
assign addr[34146]= 1678970324;
assign addr[34147]= 1770014111;
assign addr[34148]= 1852079154;
assign addr[34149]= 1924749160;
assign addr[34150]= 1987655498;
assign addr[34151]= 2040479063;
assign addr[34152]= 2082951896;
assign addr[34153]= 2114858546;
assign addr[34154]= 2136037160;
assign addr[34155]= 2146380306;
assign addr[34156]= 2145835515;
assign addr[34157]= 2134405552;
assign addr[34158]= 2112148396;
assign addr[34159]= 2079176953;
assign addr[34160]= 2035658475;
assign addr[34161]= 1981813720;
assign addr[34162]= 1917915825;
assign addr[34163]= 1844288924;
assign addr[34164]= 1761306505;
assign addr[34165]= 1669389513;
assign addr[34166]= 1569004214;
assign addr[34167]= 1460659832;
assign addr[34168]= 1344905966;
assign addr[34169]= 1222329801;
assign addr[34170]= 1093553126;
assign addr[34171]= 959229189;
assign addr[34172]= 820039373;
assign addr[34173]= 676689746;
assign addr[34174]= 529907477;
assign addr[34175]= 380437148;
assign addr[34176]= 229036977;
assign addr[34177]= 76474970;
assign addr[34178]= -76474970;
assign addr[34179]= -229036977;
assign addr[34180]= -380437148;
assign addr[34181]= -529907477;
assign addr[34182]= -676689746;
assign addr[34183]= -820039373;
assign addr[34184]= -959229189;
assign addr[34185]= -1093553126;
assign addr[34186]= -1222329801;
assign addr[34187]= -1344905966;
assign addr[34188]= -1460659832;
assign addr[34189]= -1569004214;
assign addr[34190]= -1669389513;
assign addr[34191]= -1761306505;
assign addr[34192]= -1844288924;
assign addr[34193]= -1917915825;
assign addr[34194]= -1981813720;
assign addr[34195]= -2035658475;
assign addr[34196]= -2079176953;
assign addr[34197]= -2112148396;
assign addr[34198]= -2134405552;
assign addr[34199]= -2145835515;
assign addr[34200]= -2146380306;
assign addr[34201]= -2136037160;
assign addr[34202]= -2114858546;
assign addr[34203]= -2082951896;
assign addr[34204]= -2040479063;
assign addr[34205]= -1987655498;
assign addr[34206]= -1924749160;
assign addr[34207]= -1852079154;
assign addr[34208]= -1770014111;
assign addr[34209]= -1678970324;
assign addr[34210]= -1579409630;
assign addr[34211]= -1471837070;
assign addr[34212]= -1356798326;
assign addr[34213]= -1234876957;
assign addr[34214]= -1106691431;
assign addr[34215]= -972891995;
assign addr[34216]= -834157373;
assign addr[34217]= -691191324;
assign addr[34218]= -544719071;
assign addr[34219]= -395483624;
assign addr[34220]= -244242007;
assign addr[34221]= -91761426;
assign addr[34222]= 61184634;
assign addr[34223]= 213820322;
assign addr[34224]= 365371365;
assign addr[34225]= 515068990;
assign addr[34226]= 662153826;
assign addr[34227]= 805879757;
assign addr[34228]= 945517704;
assign addr[34229]= 1080359326;
assign addr[34230]= 1209720613;
assign addr[34231]= 1332945355;
assign addr[34232]= 1449408469;
assign addr[34233]= 1558519173;
assign addr[34234]= 1659723983;
assign addr[34235]= 1752509516;
assign addr[34236]= 1836405100;
assign addr[34237]= 1910985158;
assign addr[34238]= 1975871368;
assign addr[34239]= 2030734582;
assign addr[34240]= 2075296495;
assign addr[34241]= 2109331059;
assign addr[34242]= 2132665626;
assign addr[34243]= 2145181827;
assign addr[34244]= 2146816171;
assign addr[34245]= 2137560369;
assign addr[34246]= 2117461370;
assign addr[34247]= 2086621133;
assign addr[34248]= 2045196100;
assign addr[34249]= 1993396407;
assign addr[34250]= 1931484818;
assign addr[34251]= 1859775393;
assign addr[34252]= 1778631892;
assign addr[34253]= 1688465931;
assign addr[34254]= 1589734894;
assign addr[34255]= 1482939614;
assign addr[34256]= 1368621831;
assign addr[34257]= 1247361445;
assign addr[34258]= 1119773573;
assign addr[34259]= 986505429;
assign addr[34260]= 848233042;
assign addr[34261]= 705657826;
assign addr[34262]= 559503022;
assign addr[34263]= 410510029;
assign addr[34264]= 259434643;
assign addr[34265]= 107043224;
assign addr[34266]= -45891193;
assign addr[34267]= -198592817;
assign addr[34268]= -350287041;
assign addr[34269]= -500204365;
assign addr[34270]= -647584304;
assign addr[34271]= -791679244;
assign addr[34272]= -931758235;
assign addr[34273]= -1067110699;
assign addr[34274]= -1197050035;
assign addr[34275]= -1320917099;
assign addr[34276]= -1438083551;
assign addr[34277]= -1547955041;
assign addr[34278]= -1649974225;
assign addr[34279]= -1743623590;
assign addr[34280]= -1828428082;
assign addr[34281]= -1903957513;
assign addr[34282]= -1969828744;
assign addr[34283]= -2025707632;
assign addr[34284]= -2071310720;
assign addr[34285]= -2106406677;
assign addr[34286]= -2130817471;
assign addr[34287]= -2144419275;
assign addr[34288]= -2147143090;
assign addr[34289]= -2138975100;
assign addr[34290]= -2119956737;
assign addr[34291]= -2090184478;
assign addr[34292]= -2049809346;
assign addr[34293]= -1999036154;
assign addr[34294]= -1938122457;
assign addr[34295]= -1867377253;
assign addr[34296]= -1787159411;
assign addr[34297]= -1697875851;
assign addr[34298]= -1599979481;
assign addr[34299]= -1493966902;
assign addr[34300]= -1380375881;
assign addr[34301]= -1259782632;
assign addr[34302]= -1132798888;
assign addr[34303]= -1000068799;
assign addr[34304]= -862265664;
assign addr[34305]= -720088517;
assign addr[34306]= -574258580;
assign addr[34307]= -425515602;
assign addr[34308]= -274614114;
assign addr[34309]= -122319591;
assign addr[34310]= 30595422;
assign addr[34311]= 183355234;
assign addr[34312]= 335184940;
assign addr[34313]= 485314355;
assign addr[34314]= 632981917;
assign addr[34315]= 777438554;
assign addr[34316]= 917951481;
assign addr[34317]= 1053807919;
assign addr[34318]= 1184318708;
assign addr[34319]= 1308821808;
assign addr[34320]= 1426685652;
assign addr[34321]= 1537312353;
assign addr[34322]= 1640140734;
assign addr[34323]= 1734649179;
assign addr[34324]= 1820358275;
assign addr[34325]= 1896833245;
assign addr[34326]= 1963686155;
assign addr[34327]= 2020577882;
assign addr[34328]= 2067219829;
assign addr[34329]= 2103375398;
assign addr[34330]= 2128861181;
assign addr[34331]= 2143547897;
assign addr[34332]= 2147361045;
assign addr[34333]= 2140281282;
assign addr[34334]= 2122344521;
assign addr[34335]= 2093641749;
assign addr[34336]= 2054318569;
assign addr[34337]= 2004574453;
assign addr[34338]= 1944661739;
assign addr[34339]= 1874884346;
assign addr[34340]= 1795596234;
assign addr[34341]= 1707199606;
assign addr[34342]= 1610142873;
assign addr[34343]= 1504918373;
assign addr[34344]= 1392059879;
assign addr[34345]= 1272139887;
assign addr[34346]= 1145766716;
assign addr[34347]= 1013581418;
assign addr[34348]= 876254528;
assign addr[34349]= 734482665;
assign addr[34350]= 588984994;
assign addr[34351]= 440499581;
assign addr[34352]= 289779648;
assign addr[34353]= 137589750;
assign addr[34354]= -15298099;
assign addr[34355]= -168108346;
assign addr[34356]= -320065829;
assign addr[34357]= -470399716;
assign addr[34358]= -618347408;
assign addr[34359]= -763158411;
assign addr[34360]= -904098143;
assign addr[34361]= -1040451659;
assign addr[34362]= -1171527280;
assign addr[34363]= -1296660098;
assign addr[34364]= -1415215352;
assign addr[34365]= -1526591649;
assign addr[34366]= -1630224009;
assign addr[34367]= -1725586737;
assign addr[34368]= -1812196087;
assign addr[34369]= -1889612716;
assign addr[34370]= -1957443913;
assign addr[34371]= -2015345591;
assign addr[34372]= -2063024031;
assign addr[34373]= -2100237377;
assign addr[34374]= -2126796855;
assign addr[34375]= -2142567738;
assign addr[34376]= -2147470025;
assign addr[34377]= -2141478848;
assign addr[34378]= -2124624598;
assign addr[34379]= -2096992772;
assign addr[34380]= -2058723538;
assign addr[34381]= -2010011024;
assign addr[34382]= -1951102334;
assign addr[34383]= -1882296293;
assign addr[34384]= -1803941934;
assign addr[34385]= -1716436725;
assign addr[34386]= -1620224553;
assign addr[34387]= -1515793473;
assign addr[34388]= -1403673233;
assign addr[34389]= -1284432584;
assign addr[34390]= -1158676398;
assign addr[34391]= -1027042599;
assign addr[34392]= -890198924;
assign addr[34393]= -748839539;
assign addr[34394]= -603681519;
assign addr[34395]= -455461206;
assign addr[34396]= -304930476;
assign addr[34397]= -152852926;
assign addr[34398]= 0;
assign addr[34399]= 152852926;
assign addr[34400]= 304930476;
assign addr[34401]= 455461206;
assign addr[34402]= 603681519;
assign addr[34403]= 748839539;
assign addr[34404]= 890198924;
assign addr[34405]= 1027042599;
assign addr[34406]= 1158676398;
assign addr[34407]= 1284432584;
assign addr[34408]= 1403673233;
assign addr[34409]= 1515793473;
assign addr[34410]= 1620224553;
assign addr[34411]= 1716436725;
assign addr[34412]= 1803941934;
assign addr[34413]= 1882296293;
assign addr[34414]= 1951102334;
assign addr[34415]= 2010011024;
assign addr[34416]= 2058723538;
assign addr[34417]= 2096992772;
assign addr[34418]= 2124624598;
assign addr[34419]= 2141478848;
assign addr[34420]= 2147470025;
assign addr[34421]= 2142567738;
assign addr[34422]= 2126796855;
assign addr[34423]= 2100237377;
assign addr[34424]= 2063024031;
assign addr[34425]= 2015345591;
assign addr[34426]= 1957443913;
assign addr[34427]= 1889612716;
assign addr[34428]= 1812196087;
assign addr[34429]= 1725586737;
assign addr[34430]= 1630224009;
assign addr[34431]= 1526591649;
assign addr[34432]= 1415215352;
assign addr[34433]= 1296660098;
assign addr[34434]= 1171527280;
assign addr[34435]= 1040451659;
assign addr[34436]= 904098143;
assign addr[34437]= 763158411;
assign addr[34438]= 618347408;
assign addr[34439]= 470399716;
assign addr[34440]= 320065829;
assign addr[34441]= 168108346;
assign addr[34442]= 15298099;
assign addr[34443]= -137589750;
assign addr[34444]= -289779648;
assign addr[34445]= -440499581;
assign addr[34446]= -588984994;
assign addr[34447]= -734482665;
assign addr[34448]= -876254528;
assign addr[34449]= -1013581418;
assign addr[34450]= -1145766716;
assign addr[34451]= -1272139887;
assign addr[34452]= -1392059879;
assign addr[34453]= -1504918373;
assign addr[34454]= -1610142873;
assign addr[34455]= -1707199606;
assign addr[34456]= -1795596234;
assign addr[34457]= -1874884346;
assign addr[34458]= -1944661739;
assign addr[34459]= -2004574453;
assign addr[34460]= -2054318569;
assign addr[34461]= -2093641749;
assign addr[34462]= -2122344521;
assign addr[34463]= -2140281282;
assign addr[34464]= -2147361045;
assign addr[34465]= -2143547897;
assign addr[34466]= -2128861181;
assign addr[34467]= -2103375398;
assign addr[34468]= -2067219829;
assign addr[34469]= -2020577882;
assign addr[34470]= -1963686155;
assign addr[34471]= -1896833245;
assign addr[34472]= -1820358275;
assign addr[34473]= -1734649179;
assign addr[34474]= -1640140734;
assign addr[34475]= -1537312353;
assign addr[34476]= -1426685652;
assign addr[34477]= -1308821808;
assign addr[34478]= -1184318708;
assign addr[34479]= -1053807919;
assign addr[34480]= -917951481;
assign addr[34481]= -777438554;
assign addr[34482]= -632981917;
assign addr[34483]= -485314355;
assign addr[34484]= -335184940;
assign addr[34485]= -183355234;
assign addr[34486]= -30595422;
assign addr[34487]= 122319591;
assign addr[34488]= 274614114;
assign addr[34489]= 425515602;
assign addr[34490]= 574258580;
assign addr[34491]= 720088517;
assign addr[34492]= 862265664;
assign addr[34493]= 1000068799;
assign addr[34494]= 1132798888;
assign addr[34495]= 1259782632;
assign addr[34496]= 1380375881;
assign addr[34497]= 1493966902;
assign addr[34498]= 1599979481;
assign addr[34499]= 1697875851;
assign addr[34500]= 1787159411;
assign addr[34501]= 1867377253;
assign addr[34502]= 1938122457;
assign addr[34503]= 1999036154;
assign addr[34504]= 2049809346;
assign addr[34505]= 2090184478;
assign addr[34506]= 2119956737;
assign addr[34507]= 2138975100;
assign addr[34508]= 2147143090;
assign addr[34509]= 2144419275;
assign addr[34510]= 2130817471;
assign addr[34511]= 2106406677;
assign addr[34512]= 2071310720;
assign addr[34513]= 2025707632;
assign addr[34514]= 1969828744;
assign addr[34515]= 1903957513;
assign addr[34516]= 1828428082;
assign addr[34517]= 1743623590;
assign addr[34518]= 1649974225;
assign addr[34519]= 1547955041;
assign addr[34520]= 1438083551;
assign addr[34521]= 1320917099;
assign addr[34522]= 1197050035;
assign addr[34523]= 1067110699;
assign addr[34524]= 931758235;
assign addr[34525]= 791679244;
assign addr[34526]= 647584304;
assign addr[34527]= 500204365;
assign addr[34528]= 350287041;
assign addr[34529]= 198592817;
assign addr[34530]= 45891193;
assign addr[34531]= -107043224;
assign addr[34532]= -259434643;
assign addr[34533]= -410510029;
assign addr[34534]= -559503022;
assign addr[34535]= -705657826;
assign addr[34536]= -848233042;
assign addr[34537]= -986505429;
assign addr[34538]= -1119773573;
assign addr[34539]= -1247361445;
assign addr[34540]= -1368621831;
assign addr[34541]= -1482939614;
assign addr[34542]= -1589734894;
assign addr[34543]= -1688465931;
assign addr[34544]= -1778631892;
assign addr[34545]= -1859775393;
assign addr[34546]= -1931484818;
assign addr[34547]= -1993396407;
assign addr[34548]= -2045196100;
assign addr[34549]= -2086621133;
assign addr[34550]= -2117461370;
assign addr[34551]= -2137560369;
assign addr[34552]= -2146816171;
assign addr[34553]= -2145181827;
assign addr[34554]= -2132665626;
assign addr[34555]= -2109331059;
assign addr[34556]= -2075296495;
assign addr[34557]= -2030734582;
assign addr[34558]= -1975871368;
assign addr[34559]= -1910985158;
assign addr[34560]= -1836405100;
assign addr[34561]= -1752509516;
assign addr[34562]= -1659723983;
assign addr[34563]= -1558519173;
assign addr[34564]= -1449408469;
assign addr[34565]= -1332945355;
assign addr[34566]= -1209720613;
assign addr[34567]= -1080359326;
assign addr[34568]= -945517704;
assign addr[34569]= -805879757;
assign addr[34570]= -662153826;
assign addr[34571]= -515068990;
assign addr[34572]= -365371365;
assign addr[34573]= -213820322;
assign addr[34574]= -61184634;
assign addr[34575]= 91761426;
assign addr[34576]= 244242007;
assign addr[34577]= 395483624;
assign addr[34578]= 544719071;
assign addr[34579]= 691191324;
assign addr[34580]= 834157373;
assign addr[34581]= 972891995;
assign addr[34582]= 1106691431;
assign addr[34583]= 1234876957;
assign addr[34584]= 1356798326;
assign addr[34585]= 1471837070;
assign addr[34586]= 1579409630;
assign addr[34587]= 1678970324;
assign addr[34588]= 1770014111;
assign addr[34589]= 1852079154;
assign addr[34590]= 1924749160;
assign addr[34591]= 1987655498;
assign addr[34592]= 2040479063;
assign addr[34593]= 2082951896;
assign addr[34594]= 2114858546;
assign addr[34595]= 2136037160;
assign addr[34596]= 2146380306;
assign addr[34597]= 2145835515;
assign addr[34598]= 2134405552;
assign addr[34599]= 2112148396;
assign addr[34600]= 2079176953;
assign addr[34601]= 2035658475;
assign addr[34602]= 1981813720;
assign addr[34603]= 1917915825;
assign addr[34604]= 1844288924;
assign addr[34605]= 1761306505;
assign addr[34606]= 1669389513;
assign addr[34607]= 1569004214;
assign addr[34608]= 1460659832;
assign addr[34609]= 1344905966;
assign addr[34610]= 1222329801;
assign addr[34611]= 1093553126;
assign addr[34612]= 959229189;
assign addr[34613]= 820039373;
assign addr[34614]= 676689746;
assign addr[34615]= 529907477;
assign addr[34616]= 380437148;
assign addr[34617]= 229036977;
assign addr[34618]= 76474970;
assign addr[34619]= -76474970;
assign addr[34620]= -229036977;
assign addr[34621]= -380437148;
assign addr[34622]= -529907477;
assign addr[34623]= -676689746;
assign addr[34624]= -820039373;
assign addr[34625]= -959229189;
assign addr[34626]= -1093553126;
assign addr[34627]= -1222329801;
assign addr[34628]= -1344905966;
assign addr[34629]= -1460659832;
assign addr[34630]= -1569004214;
assign addr[34631]= -1669389513;
assign addr[34632]= -1761306505;
assign addr[34633]= -1844288924;
assign addr[34634]= -1917915825;
assign addr[34635]= -1981813720;
assign addr[34636]= -2035658475;
assign addr[34637]= -2079176953;
assign addr[34638]= -2112148396;
assign addr[34639]= -2134405552;
assign addr[34640]= -2145835515;
assign addr[34641]= -2146380306;
assign addr[34642]= -2136037160;
assign addr[34643]= -2114858546;
assign addr[34644]= -2082951896;
assign addr[34645]= -2040479063;
assign addr[34646]= -1987655498;
assign addr[34647]= -1924749160;
assign addr[34648]= -1852079154;
assign addr[34649]= -1770014111;
assign addr[34650]= -1678970324;
assign addr[34651]= -1579409630;
assign addr[34652]= -1471837070;
assign addr[34653]= -1356798326;
assign addr[34654]= -1234876957;
assign addr[34655]= -1106691431;
assign addr[34656]= -972891995;
assign addr[34657]= -834157373;
assign addr[34658]= -691191324;
assign addr[34659]= -544719071;
assign addr[34660]= -395483624;
assign addr[34661]= -244242007;
assign addr[34662]= -91761426;
assign addr[34663]= 61184634;
assign addr[34664]= 213820322;
assign addr[34665]= 365371365;
assign addr[34666]= 515068990;
assign addr[34667]= 662153826;
assign addr[34668]= 805879757;
assign addr[34669]= 945517704;
assign addr[34670]= 1080359326;
assign addr[34671]= 1209720613;
assign addr[34672]= 1332945355;
assign addr[34673]= 1449408469;
assign addr[34674]= 1558519173;
assign addr[34675]= 1659723983;
assign addr[34676]= 1752509516;
assign addr[34677]= 1836405100;
assign addr[34678]= 1910985158;
assign addr[34679]= 1975871368;
assign addr[34680]= 2030734582;
assign addr[34681]= 2075296495;
assign addr[34682]= 2109331059;
assign addr[34683]= 2132665626;
assign addr[34684]= 2145181827;
assign addr[34685]= 2146816171;
assign addr[34686]= 2137560369;
assign addr[34687]= 2117461370;
assign addr[34688]= 2086621133;
assign addr[34689]= 2045196100;
assign addr[34690]= 1993396407;
assign addr[34691]= 1931484818;
assign addr[34692]= 1859775393;
assign addr[34693]= 1778631892;
assign addr[34694]= 1688465931;
assign addr[34695]= 1589734894;
assign addr[34696]= 1482939614;
assign addr[34697]= 1368621831;
assign addr[34698]= 1247361445;
assign addr[34699]= 1119773573;
assign addr[34700]= 986505429;
assign addr[34701]= 848233042;
assign addr[34702]= 705657826;
assign addr[34703]= 559503022;
assign addr[34704]= 410510029;
assign addr[34705]= 259434643;
assign addr[34706]= 107043224;
assign addr[34707]= -45891193;
assign addr[34708]= -198592817;
assign addr[34709]= -350287041;
assign addr[34710]= -500204365;
assign addr[34711]= -647584304;
assign addr[34712]= -791679244;
assign addr[34713]= -931758235;
assign addr[34714]= -1067110699;
assign addr[34715]= -1197050035;
assign addr[34716]= -1320917099;
assign addr[34717]= -1438083551;
assign addr[34718]= -1547955041;
assign addr[34719]= -1649974225;
assign addr[34720]= -1743623590;
assign addr[34721]= -1828428082;
assign addr[34722]= -1903957513;
assign addr[34723]= -1969828744;
assign addr[34724]= -2025707632;
assign addr[34725]= -2071310720;
assign addr[34726]= -2106406677;
assign addr[34727]= -2130817471;
assign addr[34728]= -2144419275;
assign addr[34729]= -2147143090;
assign addr[34730]= -2138975100;
assign addr[34731]= -2119956737;
assign addr[34732]= -2090184478;
assign addr[34733]= -2049809346;
assign addr[34734]= -1999036154;
assign addr[34735]= -1938122457;
assign addr[34736]= -1867377253;
assign addr[34737]= -1787159411;
assign addr[34738]= -1697875851;
assign addr[34739]= -1599979481;
assign addr[34740]= -1493966902;
assign addr[34741]= -1380375881;
assign addr[34742]= -1259782632;
assign addr[34743]= -1132798888;
assign addr[34744]= -1000068799;
assign addr[34745]= -862265664;
assign addr[34746]= -720088517;
assign addr[34747]= -574258580;
assign addr[34748]= -425515602;
assign addr[34749]= -274614114;
assign addr[34750]= -122319591;
assign addr[34751]= 30595422;
assign addr[34752]= 183355234;
assign addr[34753]= 335184940;
assign addr[34754]= 485314355;
assign addr[34755]= 632981917;
assign addr[34756]= 777438554;
assign addr[34757]= 917951481;
assign addr[34758]= 1053807919;
assign addr[34759]= 1184318708;
assign addr[34760]= 1308821808;
assign addr[34761]= 1426685652;
assign addr[34762]= 1537312353;
assign addr[34763]= 1640140734;
assign addr[34764]= 1734649179;
assign addr[34765]= 1820358275;
assign addr[34766]= 1896833245;
assign addr[34767]= 1963686155;
assign addr[34768]= 2020577882;
assign addr[34769]= 2067219829;
assign addr[34770]= 2103375398;
assign addr[34771]= 2128861181;
assign addr[34772]= 2143547897;
assign addr[34773]= 2147361045;
assign addr[34774]= 2140281282;
assign addr[34775]= 2122344521;
assign addr[34776]= 2093641749;
assign addr[34777]= 2054318569;
assign addr[34778]= 2004574453;
assign addr[34779]= 1944661739;
assign addr[34780]= 1874884346;
assign addr[34781]= 1795596234;
assign addr[34782]= 1707199606;
assign addr[34783]= 1610142873;
assign addr[34784]= 1504918373;
assign addr[34785]= 1392059879;
assign addr[34786]= 1272139887;
assign addr[34787]= 1145766716;
assign addr[34788]= 1013581418;
assign addr[34789]= 876254528;
assign addr[34790]= 734482665;
assign addr[34791]= 588984994;
assign addr[34792]= 440499581;
assign addr[34793]= 289779648;
assign addr[34794]= 137589750;
assign addr[34795]= -15298099;
assign addr[34796]= -168108346;
assign addr[34797]= -320065829;
assign addr[34798]= -470399716;
assign addr[34799]= -618347408;
assign addr[34800]= -763158411;
assign addr[34801]= -904098143;
assign addr[34802]= -1040451659;
assign addr[34803]= -1171527280;
assign addr[34804]= -1296660098;
assign addr[34805]= -1415215352;
assign addr[34806]= -1526591649;
assign addr[34807]= -1630224009;
assign addr[34808]= -1725586737;
assign addr[34809]= -1812196087;
assign addr[34810]= -1889612716;
assign addr[34811]= -1957443913;
assign addr[34812]= -2015345591;
assign addr[34813]= -2063024031;
assign addr[34814]= -2100237377;
assign addr[34815]= -2126796855;
assign addr[34816]= -2142567738;
assign addr[34817]= -2147470025;
assign addr[34818]= -2141478848;
assign addr[34819]= -2124624598;
assign addr[34820]= -2096992772;
assign addr[34821]= -2058723538;
assign addr[34822]= -2010011024;
assign addr[34823]= -1951102334;
assign addr[34824]= -1882296293;
assign addr[34825]= -1803941934;
assign addr[34826]= -1716436725;
assign addr[34827]= -1620224553;
assign addr[34828]= -1515793473;
assign addr[34829]= -1403673233;
assign addr[34830]= -1284432584;
assign addr[34831]= -1158676398;
assign addr[34832]= -1027042599;
assign addr[34833]= -890198924;
assign addr[34834]= -748839539;
assign addr[34835]= -603681519;
assign addr[34836]= -455461206;
assign addr[34837]= -304930476;
assign addr[34838]= -152852926;
assign addr[34839]= 0;
assign addr[34840]= 152852926;
assign addr[34841]= 304930476;
assign addr[34842]= 455461206;
assign addr[34843]= 603681519;
assign addr[34844]= 748839539;
assign addr[34845]= 890198924;
assign addr[34846]= 1027042599;
assign addr[34847]= 1158676398;
assign addr[34848]= 1284432584;
assign addr[34849]= 1403673233;
assign addr[34850]= 1515793473;
assign addr[34851]= 1620224553;
assign addr[34852]= 1716436725;
assign addr[34853]= 1803941934;
assign addr[34854]= 1882296293;
assign addr[34855]= 1951102334;
assign addr[34856]= 2010011024;
assign addr[34857]= 2058723538;
assign addr[34858]= 2096992772;
assign addr[34859]= 2124624598;
assign addr[34860]= 2141478848;
assign addr[34861]= 2147470025;
assign addr[34862]= 2142567738;
assign addr[34863]= 2126796855;
assign addr[34864]= 2100237377;
assign addr[34865]= 2063024031;
assign addr[34866]= 2015345591;
assign addr[34867]= 1957443913;
assign addr[34868]= 1889612716;
assign addr[34869]= 1812196087;
assign addr[34870]= 1725586737;
assign addr[34871]= 1630224009;
assign addr[34872]= 1526591649;
assign addr[34873]= 1415215352;
assign addr[34874]= 1296660098;
assign addr[34875]= 1171527280;
assign addr[34876]= 1040451659;
assign addr[34877]= 904098143;
assign addr[34878]= 763158411;
assign addr[34879]= 618347408;
assign addr[34880]= 470399716;
assign addr[34881]= 320065829;
assign addr[34882]= 168108346;
assign addr[34883]= 15298099;
assign addr[34884]= -137589750;
assign addr[34885]= -289779648;
assign addr[34886]= -440499581;
assign addr[34887]= -588984994;
assign addr[34888]= -734482665;
assign addr[34889]= -876254528;
assign addr[34890]= -1013581418;
assign addr[34891]= -1145766716;
assign addr[34892]= -1272139887;
assign addr[34893]= -1392059879;
assign addr[34894]= -1504918373;
assign addr[34895]= -1610142873;
assign addr[34896]= -1707199606;
assign addr[34897]= -1795596234;
assign addr[34898]= -1874884346;
assign addr[34899]= -1944661739;
assign addr[34900]= -2004574453;
assign addr[34901]= -2054318569;
assign addr[34902]= -2093641749;
assign addr[34903]= -2122344521;
assign addr[34904]= -2140281282;
assign addr[34905]= -2147361045;
assign addr[34906]= -2143547897;
assign addr[34907]= -2128861181;
assign addr[34908]= -2103375398;
assign addr[34909]= -2067219829;
assign addr[34910]= -2020577882;
assign addr[34911]= -1963686155;
assign addr[34912]= -1896833245;
assign addr[34913]= -1820358275;
assign addr[34914]= -1734649179;
assign addr[34915]= -1640140734;
assign addr[34916]= -1537312353;
assign addr[34917]= -1426685652;
assign addr[34918]= -1308821808;
assign addr[34919]= -1184318708;
assign addr[34920]= -1053807919;
assign addr[34921]= -917951481;
assign addr[34922]= -777438554;
assign addr[34923]= -632981917;
assign addr[34924]= -485314355;
assign addr[34925]= -335184940;
assign addr[34926]= -183355234;
assign addr[34927]= -30595422;
assign addr[34928]= 122319591;
assign addr[34929]= 274614114;
assign addr[34930]= 425515602;
assign addr[34931]= 574258580;
assign addr[34932]= 720088517;
assign addr[34933]= 862265664;
assign addr[34934]= 1000068799;
assign addr[34935]= 1132798888;
assign addr[34936]= 1259782632;
assign addr[34937]= 1380375881;
assign addr[34938]= 1493966902;
assign addr[34939]= 1599979481;
assign addr[34940]= 1697875851;
assign addr[34941]= 1787159411;
assign addr[34942]= 1867377253;
assign addr[34943]= 1938122457;
assign addr[34944]= 1999036154;
assign addr[34945]= 2049809346;
assign addr[34946]= 2090184478;
assign addr[34947]= 2119956737;
assign addr[34948]= 2138975100;
assign addr[34949]= 2147143090;
assign addr[34950]= 2144419275;
assign addr[34951]= 2130817471;
assign addr[34952]= 2106406677;
assign addr[34953]= 2071310720;
assign addr[34954]= 2025707632;
assign addr[34955]= 1969828744;
assign addr[34956]= 1903957513;
assign addr[34957]= 1828428082;
assign addr[34958]= 1743623590;
assign addr[34959]= 1649974225;
assign addr[34960]= 1547955041;
assign addr[34961]= 1438083551;
assign addr[34962]= 1320917099;
assign addr[34963]= 1197050035;
assign addr[34964]= 1067110699;
assign addr[34965]= 931758235;
assign addr[34966]= 791679244;
assign addr[34967]= 647584304;
assign addr[34968]= 500204365;
assign addr[34969]= 350287041;
assign addr[34970]= 198592817;
assign addr[34971]= 45891193;
assign addr[34972]= -107043224;
assign addr[34973]= -259434643;
assign addr[34974]= -410510029;
assign addr[34975]= -559503022;
assign addr[34976]= -705657826;
assign addr[34977]= -848233042;
assign addr[34978]= -986505429;
assign addr[34979]= -1119773573;
assign addr[34980]= -1247361445;
assign addr[34981]= -1368621831;
assign addr[34982]= -1482939614;
assign addr[34983]= -1589734894;
assign addr[34984]= -1688465931;
assign addr[34985]= -1778631892;
assign addr[34986]= -1859775393;
assign addr[34987]= -1931484818;
assign addr[34988]= -1993396407;
assign addr[34989]= -2045196100;
assign addr[34990]= -2086621133;
assign addr[34991]= -2117461370;
assign addr[34992]= -2137560369;
assign addr[34993]= -2146816171;
assign addr[34994]= -2145181827;
assign addr[34995]= -2132665626;
assign addr[34996]= -2109331059;
assign addr[34997]= -2075296495;
assign addr[34998]= -2030734582;
assign addr[34999]= -1975871368;
assign addr[35000]= -1910985158;
assign addr[35001]= -1836405100;
assign addr[35002]= -1752509516;
assign addr[35003]= -1659723983;
assign addr[35004]= -1558519173;
assign addr[35005]= -1449408469;
assign addr[35006]= -1332945355;
assign addr[35007]= -1209720613;
assign addr[35008]= -1080359326;
assign addr[35009]= -945517704;
assign addr[35010]= -805879757;
assign addr[35011]= -662153826;
assign addr[35012]= -515068990;
assign addr[35013]= -365371365;
assign addr[35014]= -213820322;
assign addr[35015]= -61184634;
assign addr[35016]= 91761426;
assign addr[35017]= 244242007;
assign addr[35018]= 395483624;
assign addr[35019]= 544719071;
assign addr[35020]= 691191324;
assign addr[35021]= 834157373;
assign addr[35022]= 972891995;
assign addr[35023]= 1106691431;
assign addr[35024]= 1234876957;
assign addr[35025]= 1356798326;
assign addr[35026]= 1471837070;
assign addr[35027]= 1579409630;
assign addr[35028]= 1678970324;
assign addr[35029]= 1770014111;
assign addr[35030]= 1852079154;
assign addr[35031]= 1924749160;
assign addr[35032]= 1987655498;
assign addr[35033]= 2040479063;
assign addr[35034]= 2082951896;
assign addr[35035]= 2114858546;
assign addr[35036]= 2136037160;
assign addr[35037]= 2146380306;
assign addr[35038]= 2145835515;
assign addr[35039]= 2134405552;
assign addr[35040]= 2112148396;
assign addr[35041]= 2079176953;
assign addr[35042]= 2035658475;
assign addr[35043]= 1981813720;
assign addr[35044]= 1917915825;
assign addr[35045]= 1844288924;
assign addr[35046]= 1761306505;
assign addr[35047]= 1669389513;
assign addr[35048]= 1569004214;
assign addr[35049]= 1460659832;
assign addr[35050]= 1344905966;
assign addr[35051]= 1222329801;
assign addr[35052]= 1093553126;
assign addr[35053]= 959229189;
assign addr[35054]= 820039373;
assign addr[35055]= 676689746;
assign addr[35056]= 529907477;
assign addr[35057]= 380437148;
assign addr[35058]= 229036977;
assign addr[35059]= 76474970;
assign addr[35060]= -76474970;
assign addr[35061]= -229036977;
assign addr[35062]= -380437148;
assign addr[35063]= -529907477;
assign addr[35064]= -676689746;
assign addr[35065]= -820039373;
assign addr[35066]= -959229189;
assign addr[35067]= -1093553126;
assign addr[35068]= -1222329801;
assign addr[35069]= -1344905966;
assign addr[35070]= -1460659832;
assign addr[35071]= -1569004214;
assign addr[35072]= -1669389513;
assign addr[35073]= -1761306505;
assign addr[35074]= -1844288924;
assign addr[35075]= -1917915825;
assign addr[35076]= -1981813720;
assign addr[35077]= -2035658475;
assign addr[35078]= -2079176953;
assign addr[35079]= -2112148396;
assign addr[35080]= -2134405552;
assign addr[35081]= -2145835515;
assign addr[35082]= -2146380306;
assign addr[35083]= -2136037160;
assign addr[35084]= -2114858546;
assign addr[35085]= -2082951896;
assign addr[35086]= -2040479063;
assign addr[35087]= -1987655498;
assign addr[35088]= -1924749160;
assign addr[35089]= -1852079154;
assign addr[35090]= -1770014111;
assign addr[35091]= -1678970324;
assign addr[35092]= -1579409630;
assign addr[35093]= -1471837070;
assign addr[35094]= -1356798326;
assign addr[35095]= -1234876957;
assign addr[35096]= -1106691431;
assign addr[35097]= -972891995;
assign addr[35098]= -834157373;
assign addr[35099]= -691191324;
assign addr[35100]= -544719071;
assign addr[35101]= -395483624;
assign addr[35102]= -244242007;
assign addr[35103]= -91761426;
assign addr[35104]= 61184634;
assign addr[35105]= 213820322;
assign addr[35106]= 365371365;
assign addr[35107]= 515068990;
assign addr[35108]= 662153826;
assign addr[35109]= 805879757;
assign addr[35110]= 945517704;
assign addr[35111]= 1080359326;
assign addr[35112]= 1209720613;
assign addr[35113]= 1332945355;
assign addr[35114]= 1449408469;
assign addr[35115]= 1558519173;
assign addr[35116]= 1659723983;
assign addr[35117]= 1752509516;
assign addr[35118]= 1836405100;
assign addr[35119]= 1910985158;
assign addr[35120]= 1975871368;
assign addr[35121]= 2030734582;
assign addr[35122]= 2075296495;
assign addr[35123]= 2109331059;
assign addr[35124]= 2132665626;
assign addr[35125]= 2145181827;
assign addr[35126]= 2146816171;
assign addr[35127]= 2137560369;
assign addr[35128]= 2117461370;
assign addr[35129]= 2086621133;
assign addr[35130]= 2045196100;
assign addr[35131]= 1993396407;
assign addr[35132]= 1931484818;
assign addr[35133]= 1859775393;
assign addr[35134]= 1778631892;
assign addr[35135]= 1688465931;
assign addr[35136]= 1589734894;
assign addr[35137]= 1482939614;
assign addr[35138]= 1368621831;
assign addr[35139]= 1247361445;
assign addr[35140]= 1119773573;
assign addr[35141]= 986505429;
assign addr[35142]= 848233042;
assign addr[35143]= 705657826;
assign addr[35144]= 559503022;
assign addr[35145]= 410510029;
assign addr[35146]= 259434643;
assign addr[35147]= 107043224;
assign addr[35148]= -45891193;
assign addr[35149]= -198592817;
assign addr[35150]= -350287041;
assign addr[35151]= -500204365;
assign addr[35152]= -647584304;
assign addr[35153]= -791679244;
assign addr[35154]= -931758235;
assign addr[35155]= -1067110699;
assign addr[35156]= -1197050035;
assign addr[35157]= -1320917099;
assign addr[35158]= -1438083551;
assign addr[35159]= -1547955041;
assign addr[35160]= -1649974225;
assign addr[35161]= -1743623590;
assign addr[35162]= -1828428082;
assign addr[35163]= -1903957513;
assign addr[35164]= -1969828744;
assign addr[35165]= -2025707632;
assign addr[35166]= -2071310720;
assign addr[35167]= -2106406677;
assign addr[35168]= -2130817471;
assign addr[35169]= -2144419275;
assign addr[35170]= -2147143090;
assign addr[35171]= -2138975100;
assign addr[35172]= -2119956737;
assign addr[35173]= -2090184478;
assign addr[35174]= -2049809346;
assign addr[35175]= -1999036154;
assign addr[35176]= -1938122457;
assign addr[35177]= -1867377253;
assign addr[35178]= -1787159411;
assign addr[35179]= -1697875851;
assign addr[35180]= -1599979481;
assign addr[35181]= -1493966902;
assign addr[35182]= -1380375881;
assign addr[35183]= -1259782632;
assign addr[35184]= -1132798888;
assign addr[35185]= -1000068799;
assign addr[35186]= -862265664;
assign addr[35187]= -720088517;
assign addr[35188]= -574258580;
assign addr[35189]= -425515602;
assign addr[35190]= -274614114;
assign addr[35191]= -122319591;
assign addr[35192]= 30595422;
assign addr[35193]= 183355234;
assign addr[35194]= 335184940;
assign addr[35195]= 485314355;
assign addr[35196]= 632981917;
assign addr[35197]= 777438554;
assign addr[35198]= 917951481;
assign addr[35199]= 1053807919;
assign addr[35200]= 1184318708;
assign addr[35201]= 1308821808;
assign addr[35202]= 1426685652;
assign addr[35203]= 1537312353;
assign addr[35204]= 1640140734;
assign addr[35205]= 1734649179;
assign addr[35206]= 1820358275;
assign addr[35207]= 1896833245;
assign addr[35208]= 1963686155;
assign addr[35209]= 2020577882;
assign addr[35210]= 2067219829;
assign addr[35211]= 2103375398;
assign addr[35212]= 2128861181;
assign addr[35213]= 2143547897;
assign addr[35214]= 2147361045;
assign addr[35215]= 2140281282;
assign addr[35216]= 2122344521;
assign addr[35217]= 2093641749;
assign addr[35218]= 2054318569;
assign addr[35219]= 2004574453;
assign addr[35220]= 1944661739;
assign addr[35221]= 1874884346;
assign addr[35222]= 1795596234;
assign addr[35223]= 1707199606;
assign addr[35224]= 1610142873;
assign addr[35225]= 1504918373;
assign addr[35226]= 1392059879;
assign addr[35227]= 1272139887;
assign addr[35228]= 1145766716;
assign addr[35229]= 1013581418;
assign addr[35230]= 876254528;
assign addr[35231]= 734482665;
assign addr[35232]= 588984994;
assign addr[35233]= 440499581;
assign addr[35234]= 289779648;
assign addr[35235]= 137589750;
assign addr[35236]= -15298099;
assign addr[35237]= -168108346;
assign addr[35238]= -320065829;
assign addr[35239]= -470399716;
assign addr[35240]= -618347408;
assign addr[35241]= -763158411;
assign addr[35242]= -904098143;
assign addr[35243]= -1040451659;
assign addr[35244]= -1171527280;
assign addr[35245]= -1296660098;
assign addr[35246]= -1415215352;
assign addr[35247]= -1526591649;
assign addr[35248]= -1630224009;
assign addr[35249]= -1725586737;
assign addr[35250]= -1812196087;
assign addr[35251]= -1889612716;
assign addr[35252]= -1957443913;
assign addr[35253]= -2015345591;
assign addr[35254]= -2063024031;
assign addr[35255]= -2100237377;
assign addr[35256]= -2126796855;
assign addr[35257]= -2142567738;
assign addr[35258]= -2147470025;
assign addr[35259]= -2141478848;
assign addr[35260]= -2124624598;
assign addr[35261]= -2096992772;
assign addr[35262]= -2058723538;
assign addr[35263]= -2010011024;
assign addr[35264]= -1951102334;
assign addr[35265]= -1882296293;
assign addr[35266]= -1803941934;
assign addr[35267]= -1716436725;
assign addr[35268]= -1620224553;
assign addr[35269]= -1515793473;
assign addr[35270]= -1403673233;
assign addr[35271]= -1284432584;
assign addr[35272]= -1158676398;
assign addr[35273]= -1027042599;
assign addr[35274]= -890198924;
assign addr[35275]= -748839539;
assign addr[35276]= -603681519;
assign addr[35277]= -455461206;
assign addr[35278]= -304930476;
assign addr[35279]= -152852926;
assign addr[35280]= 0;
assign addr[35281]= 152852926;
assign addr[35282]= 304930476;
assign addr[35283]= 455461206;
assign addr[35284]= 603681519;
assign addr[35285]= 748839539;
assign addr[35286]= 890198924;
assign addr[35287]= 1027042599;
assign addr[35288]= 1158676398;
assign addr[35289]= 1284432584;
assign addr[35290]= 1403673233;
assign addr[35291]= 1515793473;
assign addr[35292]= 1620224553;
assign addr[35293]= 1716436725;
assign addr[35294]= 1803941934;
assign addr[35295]= 1882296293;
assign addr[35296]= 1951102334;
assign addr[35297]= 2010011024;
assign addr[35298]= 2058723538;
assign addr[35299]= 2096992772;
assign addr[35300]= 2124624598;
assign addr[35301]= 2141478848;
assign addr[35302]= 2147470025;
assign addr[35303]= 2142567738;
assign addr[35304]= 2126796855;
assign addr[35305]= 2100237377;
assign addr[35306]= 2063024031;
assign addr[35307]= 2015345591;
assign addr[35308]= 1957443913;
assign addr[35309]= 1889612716;
assign addr[35310]= 1812196087;
assign addr[35311]= 1725586737;
assign addr[35312]= 1630224009;
assign addr[35313]= 1526591649;
assign addr[35314]= 1415215352;
assign addr[35315]= 1296660098;
assign addr[35316]= 1171527280;
assign addr[35317]= 1040451659;
assign addr[35318]= 904098143;
assign addr[35319]= 763158411;
assign addr[35320]= 618347408;
assign addr[35321]= 470399716;
assign addr[35322]= 320065829;
assign addr[35323]= 168108346;
assign addr[35324]= 15298099;
assign addr[35325]= -137589750;
assign addr[35326]= -289779648;
assign addr[35327]= -440499581;
assign addr[35328]= -588984994;
assign addr[35329]= -734482665;
assign addr[35330]= -876254528;
assign addr[35331]= -1013581418;
assign addr[35332]= -1145766716;
assign addr[35333]= -1272139887;
assign addr[35334]= -1392059879;
assign addr[35335]= -1504918373;
assign addr[35336]= -1610142873;
assign addr[35337]= -1707199606;
assign addr[35338]= -1795596234;
assign addr[35339]= -1874884346;
assign addr[35340]= -1944661739;
assign addr[35341]= -2004574453;
assign addr[35342]= -2054318569;
assign addr[35343]= -2093641749;
assign addr[35344]= -2122344521;
assign addr[35345]= -2140281282;
assign addr[35346]= -2147361045;
assign addr[35347]= -2143547897;
assign addr[35348]= -2128861181;
assign addr[35349]= -2103375398;
assign addr[35350]= -2067219829;
assign addr[35351]= -2020577882;
assign addr[35352]= -1963686155;
assign addr[35353]= -1896833245;
assign addr[35354]= -1820358275;
assign addr[35355]= -1734649179;
assign addr[35356]= -1640140734;
assign addr[35357]= -1537312353;
assign addr[35358]= -1426685652;
assign addr[35359]= -1308821808;
assign addr[35360]= -1184318708;
assign addr[35361]= -1053807919;
assign addr[35362]= -917951481;
assign addr[35363]= -777438554;
assign addr[35364]= -632981917;
assign addr[35365]= -485314355;
assign addr[35366]= -335184940;
assign addr[35367]= -183355234;
assign addr[35368]= -30595422;
assign addr[35369]= 122319591;
assign addr[35370]= 274614114;
assign addr[35371]= 425515602;
assign addr[35372]= 574258580;
assign addr[35373]= 720088517;
assign addr[35374]= 862265664;
assign addr[35375]= 1000068799;
assign addr[35376]= 1132798888;
assign addr[35377]= 1259782632;
assign addr[35378]= 1380375881;
assign addr[35379]= 1493966902;
assign addr[35380]= 1599979481;
assign addr[35381]= 1697875851;
assign addr[35382]= 1787159411;
assign addr[35383]= 1867377253;
assign addr[35384]= 1938122457;
assign addr[35385]= 1999036154;
assign addr[35386]= 2049809346;
assign addr[35387]= 2090184478;
assign addr[35388]= 2119956737;
assign addr[35389]= 2138975100;
assign addr[35390]= 2147143090;
assign addr[35391]= 2144419275;
assign addr[35392]= 2130817471;
assign addr[35393]= 2106406677;
assign addr[35394]= 2071310720;
assign addr[35395]= 2025707632;
assign addr[35396]= 1969828744;
assign addr[35397]= 1903957513;
assign addr[35398]= 1828428082;
assign addr[35399]= 1743623590;
assign addr[35400]= 1649974225;
assign addr[35401]= 1547955041;
assign addr[35402]= 1438083551;
assign addr[35403]= 1320917099;
assign addr[35404]= 1197050035;
assign addr[35405]= 1067110699;
assign addr[35406]= 931758235;
assign addr[35407]= 791679244;
assign addr[35408]= 647584304;
assign addr[35409]= 500204365;
assign addr[35410]= 350287041;
assign addr[35411]= 198592817;
assign addr[35412]= 45891193;
assign addr[35413]= -107043224;
assign addr[35414]= -259434643;
assign addr[35415]= -410510029;
assign addr[35416]= -559503022;
assign addr[35417]= -705657826;
assign addr[35418]= -848233042;
assign addr[35419]= -986505429;
assign addr[35420]= -1119773573;
assign addr[35421]= -1247361445;
assign addr[35422]= -1368621831;
assign addr[35423]= -1482939614;
assign addr[35424]= -1589734894;
assign addr[35425]= -1688465931;
assign addr[35426]= -1778631892;
assign addr[35427]= -1859775393;
assign addr[35428]= -1931484818;
assign addr[35429]= -1993396407;
assign addr[35430]= -2045196100;
assign addr[35431]= -2086621133;
assign addr[35432]= -2117461370;
assign addr[35433]= -2137560369;
assign addr[35434]= -2146816171;
assign addr[35435]= -2145181827;
assign addr[35436]= -2132665626;
assign addr[35437]= -2109331059;
assign addr[35438]= -2075296495;
assign addr[35439]= -2030734582;
assign addr[35440]= -1975871368;
assign addr[35441]= -1910985158;
assign addr[35442]= -1836405100;
assign addr[35443]= -1752509516;
assign addr[35444]= -1659723983;
assign addr[35445]= -1558519173;
assign addr[35446]= -1449408469;
assign addr[35447]= -1332945355;
assign addr[35448]= -1209720613;
assign addr[35449]= -1080359326;
assign addr[35450]= -945517704;
assign addr[35451]= -805879757;
assign addr[35452]= -662153826;
assign addr[35453]= -515068990;
assign addr[35454]= -365371365;
assign addr[35455]= -213820322;
assign addr[35456]= -61184634;
assign addr[35457]= 91761426;
assign addr[35458]= 244242007;
assign addr[35459]= 395483624;
assign addr[35460]= 544719071;
assign addr[35461]= 691191324;
assign addr[35462]= 834157373;
assign addr[35463]= 972891995;
assign addr[35464]= 1106691431;
assign addr[35465]= 1234876957;
assign addr[35466]= 1356798326;
assign addr[35467]= 1471837070;
assign addr[35468]= 1579409630;
assign addr[35469]= 1678970324;
assign addr[35470]= 1770014111;
assign addr[35471]= 1852079154;
assign addr[35472]= 1924749160;
assign addr[35473]= 1987655498;
assign addr[35474]= 2040479063;
assign addr[35475]= 2082951896;
assign addr[35476]= 2114858546;
assign addr[35477]= 2136037160;
assign addr[35478]= 2146380306;
assign addr[35479]= 2145835515;
assign addr[35480]= 2134405552;
assign addr[35481]= 2112148396;
assign addr[35482]= 2079176953;
assign addr[35483]= 2035658475;
assign addr[35484]= 1981813720;
assign addr[35485]= 1917915825;
assign addr[35486]= 1844288924;
assign addr[35487]= 1761306505;
assign addr[35488]= 1669389513;
assign addr[35489]= 1569004214;
assign addr[35490]= 1460659832;
assign addr[35491]= 1344905966;
assign addr[35492]= 1222329801;
assign addr[35493]= 1093553126;
assign addr[35494]= 959229189;
assign addr[35495]= 820039373;
assign addr[35496]= 676689746;
assign addr[35497]= 529907477;
assign addr[35498]= 380437148;
assign addr[35499]= 229036977;
assign addr[35500]= 76474970;
assign addr[35501]= -76474970;
assign addr[35502]= -229036977;
assign addr[35503]= -380437148;
assign addr[35504]= -529907477;
assign addr[35505]= -676689746;
assign addr[35506]= -820039373;
assign addr[35507]= -959229189;
assign addr[35508]= -1093553126;
assign addr[35509]= -1222329801;
assign addr[35510]= -1344905966;
assign addr[35511]= -1460659832;
assign addr[35512]= -1569004214;
assign addr[35513]= -1669389513;
assign addr[35514]= -1761306505;
assign addr[35515]= -1844288924;
assign addr[35516]= -1917915825;
assign addr[35517]= -1981813720;
assign addr[35518]= -2035658475;
assign addr[35519]= -2079176953;
assign addr[35520]= -2112148396;
assign addr[35521]= -2134405552;
assign addr[35522]= -2145835515;
assign addr[35523]= -2146380306;
assign addr[35524]= -2136037160;
assign addr[35525]= -2114858546;
assign addr[35526]= -2082951896;
assign addr[35527]= -2040479063;
assign addr[35528]= -1987655498;
assign addr[35529]= -1924749160;
assign addr[35530]= -1852079154;
assign addr[35531]= -1770014111;
assign addr[35532]= -1678970324;
assign addr[35533]= -1579409630;
assign addr[35534]= -1471837070;
assign addr[35535]= -1356798326;
assign addr[35536]= -1234876957;
assign addr[35537]= -1106691431;
assign addr[35538]= -972891995;
assign addr[35539]= -834157373;
assign addr[35540]= -691191324;
assign addr[35541]= -544719071;
assign addr[35542]= -395483624;
assign addr[35543]= -244242007;
assign addr[35544]= -91761426;
assign addr[35545]= 61184634;
assign addr[35546]= 213820322;
assign addr[35547]= 365371365;
assign addr[35548]= 515068990;
assign addr[35549]= 662153826;
assign addr[35550]= 805879757;
assign addr[35551]= 945517704;
assign addr[35552]= 1080359326;
assign addr[35553]= 1209720613;
assign addr[35554]= 1332945355;
assign addr[35555]= 1449408469;
assign addr[35556]= 1558519173;
assign addr[35557]= 1659723983;
assign addr[35558]= 1752509516;
assign addr[35559]= 1836405100;
assign addr[35560]= 1910985158;
assign addr[35561]= 1975871368;
assign addr[35562]= 2030734582;
assign addr[35563]= 2075296495;
assign addr[35564]= 2109331059;
assign addr[35565]= 2132665626;
assign addr[35566]= 2145181827;
assign addr[35567]= 2146816171;
assign addr[35568]= 2137560369;
assign addr[35569]= 2117461370;
assign addr[35570]= 2086621133;
assign addr[35571]= 2045196100;
assign addr[35572]= 1993396407;
assign addr[35573]= 1931484818;
assign addr[35574]= 1859775393;
assign addr[35575]= 1778631892;
assign addr[35576]= 1688465931;
assign addr[35577]= 1589734894;
assign addr[35578]= 1482939614;
assign addr[35579]= 1368621831;
assign addr[35580]= 1247361445;
assign addr[35581]= 1119773573;
assign addr[35582]= 986505429;
assign addr[35583]= 848233042;
assign addr[35584]= 705657826;
assign addr[35585]= 559503022;
assign addr[35586]= 410510029;
assign addr[35587]= 259434643;
assign addr[35588]= 107043224;
assign addr[35589]= -45891193;
assign addr[35590]= -198592817;
assign addr[35591]= -350287041;
assign addr[35592]= -500204365;
assign addr[35593]= -647584304;
assign addr[35594]= -791679244;
assign addr[35595]= -931758235;
assign addr[35596]= -1067110699;
assign addr[35597]= -1197050035;
assign addr[35598]= -1320917099;
assign addr[35599]= -1438083551;
assign addr[35600]= -1547955041;
assign addr[35601]= -1649974225;
assign addr[35602]= -1743623590;
assign addr[35603]= -1828428082;
assign addr[35604]= -1903957513;
assign addr[35605]= -1969828744;
assign addr[35606]= -2025707632;
assign addr[35607]= -2071310720;
assign addr[35608]= -2106406677;
assign addr[35609]= -2130817471;
assign addr[35610]= -2144419275;
assign addr[35611]= -2147143090;
assign addr[35612]= -2138975100;
assign addr[35613]= -2119956737;
assign addr[35614]= -2090184478;
assign addr[35615]= -2049809346;
assign addr[35616]= -1999036154;
assign addr[35617]= -1938122457;
assign addr[35618]= -1867377253;
assign addr[35619]= -1787159411;
assign addr[35620]= -1697875851;
assign addr[35621]= -1599979481;
assign addr[35622]= -1493966902;
assign addr[35623]= -1380375881;
assign addr[35624]= -1259782632;
assign addr[35625]= -1132798888;
assign addr[35626]= -1000068799;
assign addr[35627]= -862265664;
assign addr[35628]= -720088517;
assign addr[35629]= -574258580;
assign addr[35630]= -425515602;
assign addr[35631]= -274614114;
assign addr[35632]= -122319591;
assign addr[35633]= 30595422;
assign addr[35634]= 183355234;
assign addr[35635]= 335184940;
assign addr[35636]= 485314355;
assign addr[35637]= 632981917;
assign addr[35638]= 777438554;
assign addr[35639]= 917951481;
assign addr[35640]= 1053807919;
assign addr[35641]= 1184318708;
assign addr[35642]= 1308821808;
assign addr[35643]= 1426685652;
assign addr[35644]= 1537312353;
assign addr[35645]= 1640140734;
assign addr[35646]= 1734649179;
assign addr[35647]= 1820358275;
assign addr[35648]= 1896833245;
assign addr[35649]= 1963686155;
assign addr[35650]= 2020577882;
assign addr[35651]= 2067219829;
assign addr[35652]= 2103375398;
assign addr[35653]= 2128861181;
assign addr[35654]= 2143547897;
assign addr[35655]= 2147361045;
assign addr[35656]= 2140281282;
assign addr[35657]= 2122344521;
assign addr[35658]= 2093641749;
assign addr[35659]= 2054318569;
assign addr[35660]= 2004574453;
assign addr[35661]= 1944661739;
assign addr[35662]= 1874884346;
assign addr[35663]= 1795596234;
assign addr[35664]= 1707199606;
assign addr[35665]= 1610142873;
assign addr[35666]= 1504918373;
assign addr[35667]= 1392059879;
assign addr[35668]= 1272139887;
assign addr[35669]= 1145766716;
assign addr[35670]= 1013581418;
assign addr[35671]= 876254528;
assign addr[35672]= 734482665;
assign addr[35673]= 588984994;
assign addr[35674]= 440499581;
assign addr[35675]= 289779648;
assign addr[35676]= 137589750;
assign addr[35677]= -15298099;
assign addr[35678]= -168108346;
assign addr[35679]= -320065829;
assign addr[35680]= -470399716;
assign addr[35681]= -618347408;
assign addr[35682]= -763158411;
assign addr[35683]= -904098143;
assign addr[35684]= -1040451659;
assign addr[35685]= -1171527280;
assign addr[35686]= -1296660098;
assign addr[35687]= -1415215352;
assign addr[35688]= -1526591649;
assign addr[35689]= -1630224009;
assign addr[35690]= -1725586737;
assign addr[35691]= -1812196087;
assign addr[35692]= -1889612716;
assign addr[35693]= -1957443913;
assign addr[35694]= -2015345591;
assign addr[35695]= -2063024031;
assign addr[35696]= -2100237377;
assign addr[35697]= -2126796855;
assign addr[35698]= -2142567738;
assign addr[35699]= -2147470025;
assign addr[35700]= -2141478848;
assign addr[35701]= -2124624598;
assign addr[35702]= -2096992772;
assign addr[35703]= -2058723538;
assign addr[35704]= -2010011024;
assign addr[35705]= -1951102334;
assign addr[35706]= -1882296293;
assign addr[35707]= -1803941934;
assign addr[35708]= -1716436725;
assign addr[35709]= -1620224553;
assign addr[35710]= -1515793473;
assign addr[35711]= -1403673233;
assign addr[35712]= -1284432584;
assign addr[35713]= -1158676398;
assign addr[35714]= -1027042599;
assign addr[35715]= -890198924;
assign addr[35716]= -748839539;
assign addr[35717]= -603681519;
assign addr[35718]= -455461206;
assign addr[35719]= -304930476;
assign addr[35720]= -152852926;
assign addr[35721]= 0;
assign addr[35722]= 152852926;
assign addr[35723]= 304930476;
assign addr[35724]= 455461206;
assign addr[35725]= 603681519;
assign addr[35726]= 748839539;
assign addr[35727]= 890198924;
assign addr[35728]= 1027042599;
assign addr[35729]= 1158676398;
assign addr[35730]= 1284432584;
assign addr[35731]= 1403673233;
assign addr[35732]= 1515793473;
assign addr[35733]= 1620224553;
assign addr[35734]= 1716436725;
assign addr[35735]= 1803941934;
assign addr[35736]= 1882296293;
assign addr[35737]= 1951102334;
assign addr[35738]= 2010011024;
assign addr[35739]= 2058723538;
assign addr[35740]= 2096992772;
assign addr[35741]= 2124624598;
assign addr[35742]= 2141478848;
assign addr[35743]= 2147470025;
assign addr[35744]= 2142567738;
assign addr[35745]= 2126796855;
assign addr[35746]= 2100237377;
assign addr[35747]= 2063024031;
assign addr[35748]= 2015345591;
assign addr[35749]= 1957443913;
assign addr[35750]= 1889612716;
assign addr[35751]= 1812196087;
assign addr[35752]= 1725586737;
assign addr[35753]= 1630224009;
assign addr[35754]= 1526591649;
assign addr[35755]= 1415215352;
assign addr[35756]= 1296660098;
assign addr[35757]= 1171527280;
assign addr[35758]= 1040451659;
assign addr[35759]= 904098143;
assign addr[35760]= 763158411;
assign addr[35761]= 618347408;
assign addr[35762]= 470399716;
assign addr[35763]= 320065829;
assign addr[35764]= 168108346;
assign addr[35765]= 15298099;
assign addr[35766]= -137589750;
assign addr[35767]= -289779648;
assign addr[35768]= -440499581;
assign addr[35769]= -588984994;
assign addr[35770]= -734482665;
assign addr[35771]= -876254528;
assign addr[35772]= -1013581418;
assign addr[35773]= -1145766716;
assign addr[35774]= -1272139887;
assign addr[35775]= -1392059879;
assign addr[35776]= -1504918373;
assign addr[35777]= -1610142873;
assign addr[35778]= -1707199606;
assign addr[35779]= -1795596234;
assign addr[35780]= -1874884346;
assign addr[35781]= -1944661739;
assign addr[35782]= -2004574453;
assign addr[35783]= -2054318569;
assign addr[35784]= -2093641749;
assign addr[35785]= -2122344521;
assign addr[35786]= -2140281282;
assign addr[35787]= -2147361045;
assign addr[35788]= -2143547897;
assign addr[35789]= -2128861181;
assign addr[35790]= -2103375398;
assign addr[35791]= -2067219829;
assign addr[35792]= -2020577882;
assign addr[35793]= -1963686155;
assign addr[35794]= -1896833245;
assign addr[35795]= -1820358275;
assign addr[35796]= -1734649179;
assign addr[35797]= -1640140734;
assign addr[35798]= -1537312353;
assign addr[35799]= -1426685652;
assign addr[35800]= -1308821808;
assign addr[35801]= -1184318708;
assign addr[35802]= -1053807919;
assign addr[35803]= -917951481;
assign addr[35804]= -777438554;
assign addr[35805]= -632981917;
assign addr[35806]= -485314355;
assign addr[35807]= -335184940;
assign addr[35808]= -183355234;
assign addr[35809]= -30595422;
assign addr[35810]= 122319591;
assign addr[35811]= 274614114;
assign addr[35812]= 425515602;
assign addr[35813]= 574258580;
assign addr[35814]= 720088517;
assign addr[35815]= 862265664;
assign addr[35816]= 1000068799;
assign addr[35817]= 1132798888;
assign addr[35818]= 1259782632;
assign addr[35819]= 1380375881;
assign addr[35820]= 1493966902;
assign addr[35821]= 1599979481;
assign addr[35822]= 1697875851;
assign addr[35823]= 1787159411;
assign addr[35824]= 1867377253;
assign addr[35825]= 1938122457;
assign addr[35826]= 1999036154;
assign addr[35827]= 2049809346;
assign addr[35828]= 2090184478;
assign addr[35829]= 2119956737;
assign addr[35830]= 2138975100;
assign addr[35831]= 2147143090;
assign addr[35832]= 2144419275;
assign addr[35833]= 2130817471;
assign addr[35834]= 2106406677;
assign addr[35835]= 2071310720;
assign addr[35836]= 2025707632;
assign addr[35837]= 1969828744;
assign addr[35838]= 1903957513;
assign addr[35839]= 1828428082;
assign addr[35840]= 1743623590;
assign addr[35841]= 1649974225;
assign addr[35842]= 1547955041;
assign addr[35843]= 1438083551;
assign addr[35844]= 1320917099;
assign addr[35845]= 1197050035;
assign addr[35846]= 1067110699;
assign addr[35847]= 931758235;
assign addr[35848]= 791679244;
assign addr[35849]= 647584304;
assign addr[35850]= 500204365;
assign addr[35851]= 350287041;
assign addr[35852]= 198592817;
assign addr[35853]= 45891193;
assign addr[35854]= -107043224;
assign addr[35855]= -259434643;
assign addr[35856]= -410510029;
assign addr[35857]= -559503022;
assign addr[35858]= -705657826;
assign addr[35859]= -848233042;
assign addr[35860]= -986505429;
assign addr[35861]= -1119773573;
assign addr[35862]= -1247361445;
assign addr[35863]= -1368621831;
assign addr[35864]= -1482939614;
assign addr[35865]= -1589734894;
assign addr[35866]= -1688465931;
assign addr[35867]= -1778631892;
assign addr[35868]= -1859775393;
assign addr[35869]= -1931484818;
assign addr[35870]= -1993396407;
assign addr[35871]= -2045196100;
assign addr[35872]= -2086621133;
assign addr[35873]= -2117461370;
assign addr[35874]= -2137560369;
assign addr[35875]= -2146816171;
assign addr[35876]= -2145181827;
assign addr[35877]= -2132665626;
assign addr[35878]= -2109331059;
assign addr[35879]= -2075296495;
assign addr[35880]= -2030734582;
assign addr[35881]= -1975871368;
assign addr[35882]= -1910985158;
assign addr[35883]= -1836405100;
assign addr[35884]= -1752509516;
assign addr[35885]= -1659723983;
assign addr[35886]= -1558519173;
assign addr[35887]= -1449408469;
assign addr[35888]= -1332945355;
assign addr[35889]= -1209720613;
assign addr[35890]= -1080359326;
assign addr[35891]= -945517704;
assign addr[35892]= -805879757;
assign addr[35893]= -662153826;
assign addr[35894]= -515068990;
assign addr[35895]= -365371365;
assign addr[35896]= -213820322;
assign addr[35897]= -61184634;
assign addr[35898]= 91761426;
assign addr[35899]= 244242007;
assign addr[35900]= 395483624;
assign addr[35901]= 544719071;
assign addr[35902]= 691191324;
assign addr[35903]= 834157373;
assign addr[35904]= 972891995;
assign addr[35905]= 1106691431;
assign addr[35906]= 1234876957;
assign addr[35907]= 1356798326;
assign addr[35908]= 1471837070;
assign addr[35909]= 1579409630;
assign addr[35910]= 1678970324;
assign addr[35911]= 1770014111;
assign addr[35912]= 1852079154;
assign addr[35913]= 1924749160;
assign addr[35914]= 1987655498;
assign addr[35915]= 2040479063;
assign addr[35916]= 2082951896;
assign addr[35917]= 2114858546;
assign addr[35918]= 2136037160;
assign addr[35919]= 2146380306;
assign addr[35920]= 2145835515;
assign addr[35921]= 2134405552;
assign addr[35922]= 2112148396;
assign addr[35923]= 2079176953;
assign addr[35924]= 2035658475;
assign addr[35925]= 1981813720;
assign addr[35926]= 1917915825;
assign addr[35927]= 1844288924;
assign addr[35928]= 1761306505;
assign addr[35929]= 1669389513;
assign addr[35930]= 1569004214;
assign addr[35931]= 1460659832;
assign addr[35932]= 1344905966;
assign addr[35933]= 1222329801;
assign addr[35934]= 1093553126;
assign addr[35935]= 959229189;
assign addr[35936]= 820039373;
assign addr[35937]= 676689746;
assign addr[35938]= 529907477;
assign addr[35939]= 380437148;
assign addr[35940]= 229036977;
assign addr[35941]= 76474970;
assign addr[35942]= -76474970;
assign addr[35943]= -229036977;
assign addr[35944]= -380437148;
assign addr[35945]= -529907477;
assign addr[35946]= -676689746;
assign addr[35947]= -820039373;
assign addr[35948]= -959229189;
assign addr[35949]= -1093553126;
assign addr[35950]= -1222329801;
assign addr[35951]= -1344905966;
assign addr[35952]= -1460659832;
assign addr[35953]= -1569004214;
assign addr[35954]= -1669389513;
assign addr[35955]= -1761306505;
assign addr[35956]= -1844288924;
assign addr[35957]= -1917915825;
assign addr[35958]= -1981813720;
assign addr[35959]= -2035658475;
assign addr[35960]= -2079176953;
assign addr[35961]= -2112148396;
assign addr[35962]= -2134405552;
assign addr[35963]= -2145835515;
assign addr[35964]= -2146380306;
assign addr[35965]= -2136037160;
assign addr[35966]= -2114858546;
assign addr[35967]= -2082951896;
assign addr[35968]= -2040479063;
assign addr[35969]= -1987655498;
assign addr[35970]= -1924749160;
assign addr[35971]= -1852079154;
assign addr[35972]= -1770014111;
assign addr[35973]= -1678970324;
assign addr[35974]= -1579409630;
assign addr[35975]= -1471837070;
assign addr[35976]= -1356798326;
assign addr[35977]= -1234876957;
assign addr[35978]= -1106691431;
assign addr[35979]= -972891995;
assign addr[35980]= -834157373;
assign addr[35981]= -691191324;
assign addr[35982]= -544719071;
assign addr[35983]= -395483624;
assign addr[35984]= -244242007;
assign addr[35985]= -91761426;
assign addr[35986]= 61184634;
assign addr[35987]= 213820322;
assign addr[35988]= 365371365;
assign addr[35989]= 515068990;
assign addr[35990]= 662153826;
assign addr[35991]= 805879757;
assign addr[35992]= 945517704;
assign addr[35993]= 1080359326;
assign addr[35994]= 1209720613;
assign addr[35995]= 1332945355;
assign addr[35996]= 1449408469;
assign addr[35997]= 1558519173;
assign addr[35998]= 1659723983;
assign addr[35999]= 1752509516;
assign addr[36000]= 1836405100;
assign addr[36001]= 1910985158;
assign addr[36002]= 1975871368;
assign addr[36003]= 2030734582;
assign addr[36004]= 2075296495;
assign addr[36005]= 2109331059;
assign addr[36006]= 2132665626;
assign addr[36007]= 2145181827;
assign addr[36008]= 2146816171;
assign addr[36009]= 2137560369;
assign addr[36010]= 2117461370;
assign addr[36011]= 2086621133;
assign addr[36012]= 2045196100;
assign addr[36013]= 1993396407;
assign addr[36014]= 1931484818;
assign addr[36015]= 1859775393;
assign addr[36016]= 1778631892;
assign addr[36017]= 1688465931;
assign addr[36018]= 1589734894;
assign addr[36019]= 1482939614;
assign addr[36020]= 1368621831;
assign addr[36021]= 1247361445;
assign addr[36022]= 1119773573;
assign addr[36023]= 986505429;
assign addr[36024]= 848233042;
assign addr[36025]= 705657826;
assign addr[36026]= 559503022;
assign addr[36027]= 410510029;
assign addr[36028]= 259434643;
assign addr[36029]= 107043224;
assign addr[36030]= -45891193;
assign addr[36031]= -198592817;
assign addr[36032]= -350287041;
assign addr[36033]= -500204365;
assign addr[36034]= -647584304;
assign addr[36035]= -791679244;
assign addr[36036]= -931758235;
assign addr[36037]= -1067110699;
assign addr[36038]= -1197050035;
assign addr[36039]= -1320917099;
assign addr[36040]= -1438083551;
assign addr[36041]= -1547955041;
assign addr[36042]= -1649974225;
assign addr[36043]= -1743623590;
assign addr[36044]= -1828428082;
assign addr[36045]= -1903957513;
assign addr[36046]= -1969828744;
assign addr[36047]= -2025707632;
assign addr[36048]= -2071310720;
assign addr[36049]= -2106406677;
assign addr[36050]= -2130817471;
assign addr[36051]= -2144419275;
assign addr[36052]= -2147143090;
assign addr[36053]= -2138975100;
assign addr[36054]= -2119956737;
assign addr[36055]= -2090184478;
assign addr[36056]= -2049809346;
assign addr[36057]= -1999036154;
assign addr[36058]= -1938122457;
assign addr[36059]= -1867377253;
assign addr[36060]= -1787159411;
assign addr[36061]= -1697875851;
assign addr[36062]= -1599979481;
assign addr[36063]= -1493966902;
assign addr[36064]= -1380375881;
assign addr[36065]= -1259782632;
assign addr[36066]= -1132798888;
assign addr[36067]= -1000068799;
assign addr[36068]= -862265664;
assign addr[36069]= -720088517;
assign addr[36070]= -574258580;
assign addr[36071]= -425515602;
assign addr[36072]= -274614114;
assign addr[36073]= -122319591;
assign addr[36074]= 30595422;
assign addr[36075]= 183355234;
assign addr[36076]= 335184940;
assign addr[36077]= 485314355;
assign addr[36078]= 632981917;
assign addr[36079]= 777438554;
assign addr[36080]= 917951481;
assign addr[36081]= 1053807919;
assign addr[36082]= 1184318708;
assign addr[36083]= 1308821808;
assign addr[36084]= 1426685652;
assign addr[36085]= 1537312353;
assign addr[36086]= 1640140734;
assign addr[36087]= 1734649179;
assign addr[36088]= 1820358275;
assign addr[36089]= 1896833245;
assign addr[36090]= 1963686155;
assign addr[36091]= 2020577882;
assign addr[36092]= 2067219829;
assign addr[36093]= 2103375398;
assign addr[36094]= 2128861181;
assign addr[36095]= 2143547897;
assign addr[36096]= 2147361045;
assign addr[36097]= 2140281282;
assign addr[36098]= 2122344521;
assign addr[36099]= 2093641749;
assign addr[36100]= 2054318569;
assign addr[36101]= 2004574453;
assign addr[36102]= 1944661739;
assign addr[36103]= 1874884346;
assign addr[36104]= 1795596234;
assign addr[36105]= 1707199606;
assign addr[36106]= 1610142873;
assign addr[36107]= 1504918373;
assign addr[36108]= 1392059879;
assign addr[36109]= 1272139887;
assign addr[36110]= 1145766716;
assign addr[36111]= 1013581418;
assign addr[36112]= 876254528;
assign addr[36113]= 734482665;
assign addr[36114]= 588984994;
assign addr[36115]= 440499581;
assign addr[36116]= 289779648;
assign addr[36117]= 137589750;
assign addr[36118]= -15298099;
assign addr[36119]= -168108346;
assign addr[36120]= -320065829;
assign addr[36121]= -470399716;
assign addr[36122]= -618347408;
assign addr[36123]= -763158411;
assign addr[36124]= -904098143;
assign addr[36125]= -1040451659;
assign addr[36126]= -1171527280;
assign addr[36127]= -1296660098;
assign addr[36128]= -1415215352;
assign addr[36129]= -1526591649;
assign addr[36130]= -1630224009;
assign addr[36131]= -1725586737;
assign addr[36132]= -1812196087;
assign addr[36133]= -1889612716;
assign addr[36134]= -1957443913;
assign addr[36135]= -2015345591;
assign addr[36136]= -2063024031;
assign addr[36137]= -2100237377;
assign addr[36138]= -2126796855;
assign addr[36139]= -2142567738;
assign addr[36140]= -2147470025;
assign addr[36141]= -2141478848;
assign addr[36142]= -2124624598;
assign addr[36143]= -2096992772;
assign addr[36144]= -2058723538;
assign addr[36145]= -2010011024;
assign addr[36146]= -1951102334;
assign addr[36147]= -1882296293;
assign addr[36148]= -1803941934;
assign addr[36149]= -1716436725;
assign addr[36150]= -1620224553;
assign addr[36151]= -1515793473;
assign addr[36152]= -1403673233;
assign addr[36153]= -1284432584;
assign addr[36154]= -1158676398;
assign addr[36155]= -1027042599;
assign addr[36156]= -890198924;
assign addr[36157]= -748839539;
assign addr[36158]= -603681519;
assign addr[36159]= -455461206;
assign addr[36160]= -304930476;
assign addr[36161]= -152852926;
assign addr[36162]= 0;
assign addr[36163]= 152852926;
assign addr[36164]= 304930476;
assign addr[36165]= 455461206;
assign addr[36166]= 603681519;
assign addr[36167]= 748839539;
assign addr[36168]= 890198924;
assign addr[36169]= 1027042599;
assign addr[36170]= 1158676398;
assign addr[36171]= 1284432584;
assign addr[36172]= 1403673233;
assign addr[36173]= 1515793473;
assign addr[36174]= 1620224553;
assign addr[36175]= 1716436725;
assign addr[36176]= 1803941934;
assign addr[36177]= 1882296293;
assign addr[36178]= 1951102334;
assign addr[36179]= 2010011024;
assign addr[36180]= 2058723538;
assign addr[36181]= 2096992772;
assign addr[36182]= 2124624598;
assign addr[36183]= 2141478848;
assign addr[36184]= 2147470025;
assign addr[36185]= 2142567738;
assign addr[36186]= 2126796855;
assign addr[36187]= 2100237377;
assign addr[36188]= 2063024031;
assign addr[36189]= 2015345591;
assign addr[36190]= 1957443913;
assign addr[36191]= 1889612716;
assign addr[36192]= 1812196087;
assign addr[36193]= 1725586737;
assign addr[36194]= 1630224009;
assign addr[36195]= 1526591649;
assign addr[36196]= 1415215352;
assign addr[36197]= 1296660098;
assign addr[36198]= 1171527280;
assign addr[36199]= 1040451659;
assign addr[36200]= 904098143;
assign addr[36201]= 763158411;
assign addr[36202]= 618347408;
assign addr[36203]= 470399716;
assign addr[36204]= 320065829;
assign addr[36205]= 168108346;
assign addr[36206]= 15298099;
assign addr[36207]= -137589750;
assign addr[36208]= -289779648;
assign addr[36209]= -440499581;
assign addr[36210]= -588984994;
assign addr[36211]= -734482665;
assign addr[36212]= -876254528;
assign addr[36213]= -1013581418;
assign addr[36214]= -1145766716;
assign addr[36215]= -1272139887;
assign addr[36216]= -1392059879;
assign addr[36217]= -1504918373;
assign addr[36218]= -1610142873;
assign addr[36219]= -1707199606;
assign addr[36220]= -1795596234;
assign addr[36221]= -1874884346;
assign addr[36222]= -1944661739;
assign addr[36223]= -2004574453;
assign addr[36224]= -2054318569;
assign addr[36225]= -2093641749;
assign addr[36226]= -2122344521;
assign addr[36227]= -2140281282;
assign addr[36228]= -2147361045;
assign addr[36229]= -2143547897;
assign addr[36230]= -2128861181;
assign addr[36231]= -2103375398;
assign addr[36232]= -2067219829;
assign addr[36233]= -2020577882;
assign addr[36234]= -1963686155;
assign addr[36235]= -1896833245;
assign addr[36236]= -1820358275;
assign addr[36237]= -1734649179;
assign addr[36238]= -1640140734;
assign addr[36239]= -1537312353;
assign addr[36240]= -1426685652;
assign addr[36241]= -1308821808;
assign addr[36242]= -1184318708;
assign addr[36243]= -1053807919;
assign addr[36244]= -917951481;
assign addr[36245]= -777438554;
assign addr[36246]= -632981917;
assign addr[36247]= -485314355;
assign addr[36248]= -335184940;
assign addr[36249]= -183355234;
assign addr[36250]= -30595422;
assign addr[36251]= 122319591;
assign addr[36252]= 274614114;
assign addr[36253]= 425515602;
assign addr[36254]= 574258580;
assign addr[36255]= 720088517;
assign addr[36256]= 862265664;
assign addr[36257]= 1000068799;
assign addr[36258]= 1132798888;
assign addr[36259]= 1259782632;
assign addr[36260]= 1380375881;
assign addr[36261]= 1493966902;
assign addr[36262]= 1599979481;
assign addr[36263]= 1697875851;
assign addr[36264]= 1787159411;
assign addr[36265]= 1867377253;
assign addr[36266]= 1938122457;
assign addr[36267]= 1999036154;
assign addr[36268]= 2049809346;
assign addr[36269]= 2090184478;
assign addr[36270]= 2119956737;
assign addr[36271]= 2138975100;
assign addr[36272]= 2147143090;
assign addr[36273]= 2144419275;
assign addr[36274]= 2130817471;
assign addr[36275]= 2106406677;
assign addr[36276]= 2071310720;
assign addr[36277]= 2025707632;
assign addr[36278]= 1969828744;
assign addr[36279]= 1903957513;
assign addr[36280]= 1828428082;
assign addr[36281]= 1743623590;
assign addr[36282]= 1649974225;
assign addr[36283]= 1547955041;
assign addr[36284]= 1438083551;
assign addr[36285]= 1320917099;
assign addr[36286]= 1197050035;
assign addr[36287]= 1067110699;
assign addr[36288]= 931758235;
assign addr[36289]= 791679244;
assign addr[36290]= 647584304;
assign addr[36291]= 500204365;
assign addr[36292]= 350287041;
assign addr[36293]= 198592817;
assign addr[36294]= 45891193;
assign addr[36295]= -107043224;
assign addr[36296]= -259434643;
assign addr[36297]= -410510029;
assign addr[36298]= -559503022;
assign addr[36299]= -705657826;
assign addr[36300]= -848233042;
assign addr[36301]= -986505429;
assign addr[36302]= -1119773573;
assign addr[36303]= -1247361445;
assign addr[36304]= -1368621831;
assign addr[36305]= -1482939614;
assign addr[36306]= -1589734894;
assign addr[36307]= -1688465931;
assign addr[36308]= -1778631892;
assign addr[36309]= -1859775393;
assign addr[36310]= -1931484818;
assign addr[36311]= -1993396407;
assign addr[36312]= -2045196100;
assign addr[36313]= -2086621133;
assign addr[36314]= -2117461370;
assign addr[36315]= -2137560369;
assign addr[36316]= -2146816171;
assign addr[36317]= -2145181827;
assign addr[36318]= -2132665626;
assign addr[36319]= -2109331059;
assign addr[36320]= -2075296495;
assign addr[36321]= -2030734582;
assign addr[36322]= -1975871368;
assign addr[36323]= -1910985158;
assign addr[36324]= -1836405100;
assign addr[36325]= -1752509516;
assign addr[36326]= -1659723983;
assign addr[36327]= -1558519173;
assign addr[36328]= -1449408469;
assign addr[36329]= -1332945355;
assign addr[36330]= -1209720613;
assign addr[36331]= -1080359326;
assign addr[36332]= -945517704;
assign addr[36333]= -805879757;
assign addr[36334]= -662153826;
assign addr[36335]= -515068990;
assign addr[36336]= -365371365;
assign addr[36337]= -213820322;
assign addr[36338]= -61184634;
assign addr[36339]= 91761426;
assign addr[36340]= 244242007;
assign addr[36341]= 395483624;
assign addr[36342]= 544719071;
assign addr[36343]= 691191324;
assign addr[36344]= 834157373;
assign addr[36345]= 972891995;
assign addr[36346]= 1106691431;
assign addr[36347]= 1234876957;
assign addr[36348]= 1356798326;
assign addr[36349]= 1471837070;
assign addr[36350]= 1579409630;
assign addr[36351]= 1678970324;
assign addr[36352]= 1770014111;
assign addr[36353]= 1852079154;
assign addr[36354]= 1924749160;
assign addr[36355]= 1987655498;
assign addr[36356]= 2040479063;
assign addr[36357]= 2082951896;
assign addr[36358]= 2114858546;
assign addr[36359]= 2136037160;
assign addr[36360]= 2146380306;
assign addr[36361]= 2145835515;
assign addr[36362]= 2134405552;
assign addr[36363]= 2112148396;
assign addr[36364]= 2079176953;
assign addr[36365]= 2035658475;
assign addr[36366]= 1981813720;
assign addr[36367]= 1917915825;
assign addr[36368]= 1844288924;
assign addr[36369]= 1761306505;
assign addr[36370]= 1669389513;
assign addr[36371]= 1569004214;
assign addr[36372]= 1460659832;
assign addr[36373]= 1344905966;
assign addr[36374]= 1222329801;
assign addr[36375]= 1093553126;
assign addr[36376]= 959229189;
assign addr[36377]= 820039373;
assign addr[36378]= 676689746;
assign addr[36379]= 529907477;
assign addr[36380]= 380437148;
assign addr[36381]= 229036977;
assign addr[36382]= 76474970;
assign addr[36383]= -76474970;
assign addr[36384]= -229036977;
assign addr[36385]= -380437148;
assign addr[36386]= -529907477;
assign addr[36387]= -676689746;
assign addr[36388]= -820039373;
assign addr[36389]= -959229189;
assign addr[36390]= -1093553126;
assign addr[36391]= -1222329801;
assign addr[36392]= -1344905966;
assign addr[36393]= -1460659832;
assign addr[36394]= -1569004214;
assign addr[36395]= -1669389513;
assign addr[36396]= -1761306505;
assign addr[36397]= -1844288924;
assign addr[36398]= -1917915825;
assign addr[36399]= -1981813720;
assign addr[36400]= -2035658475;
assign addr[36401]= -2079176953;
assign addr[36402]= -2112148396;
assign addr[36403]= -2134405552;
assign addr[36404]= -2145835515;
assign addr[36405]= -2146380306;
assign addr[36406]= -2136037160;
assign addr[36407]= -2114858546;
assign addr[36408]= -2082951896;
assign addr[36409]= -2040479063;
assign addr[36410]= -1987655498;
assign addr[36411]= -1924749160;
assign addr[36412]= -1852079154;
assign addr[36413]= -1770014111;
assign addr[36414]= -1678970324;
assign addr[36415]= -1579409630;
assign addr[36416]= -1471837070;
assign addr[36417]= -1356798326;
assign addr[36418]= -1234876957;
assign addr[36419]= -1106691431;
assign addr[36420]= -972891995;
assign addr[36421]= -834157373;
assign addr[36422]= -691191324;
assign addr[36423]= -544719071;
assign addr[36424]= -395483624;
assign addr[36425]= -244242007;
assign addr[36426]= -91761426;
assign addr[36427]= 61184634;
assign addr[36428]= 213820322;
assign addr[36429]= 365371365;
assign addr[36430]= 515068990;
assign addr[36431]= 662153826;
assign addr[36432]= 805879757;
assign addr[36433]= 945517704;
assign addr[36434]= 1080359326;
assign addr[36435]= 1209720613;
assign addr[36436]= 1332945355;
assign addr[36437]= 1449408469;
assign addr[36438]= 1558519173;
assign addr[36439]= 1659723983;
assign addr[36440]= 1752509516;
assign addr[36441]= 1836405100;
assign addr[36442]= 1910985158;
assign addr[36443]= 1975871368;
assign addr[36444]= 2030734582;
assign addr[36445]= 2075296495;
assign addr[36446]= 2109331059;
assign addr[36447]= 2132665626;
assign addr[36448]= 2145181827;
assign addr[36449]= 2146816171;
assign addr[36450]= 2137560369;
assign addr[36451]= 2117461370;
assign addr[36452]= 2086621133;
assign addr[36453]= 2045196100;
assign addr[36454]= 1993396407;
assign addr[36455]= 1931484818;
assign addr[36456]= 1859775393;
assign addr[36457]= 1778631892;
assign addr[36458]= 1688465931;
assign addr[36459]= 1589734894;
assign addr[36460]= 1482939614;
assign addr[36461]= 1368621831;
assign addr[36462]= 1247361445;
assign addr[36463]= 1119773573;
assign addr[36464]= 986505429;
assign addr[36465]= 848233042;
assign addr[36466]= 705657826;
assign addr[36467]= 559503022;
assign addr[36468]= 410510029;
assign addr[36469]= 259434643;
assign addr[36470]= 107043224;
assign addr[36471]= -45891193;
assign addr[36472]= -198592817;
assign addr[36473]= -350287041;
assign addr[36474]= -500204365;
assign addr[36475]= -647584304;
assign addr[36476]= -791679244;
assign addr[36477]= -931758235;
assign addr[36478]= -1067110699;
assign addr[36479]= -1197050035;
assign addr[36480]= -1320917099;
assign addr[36481]= -1438083551;
assign addr[36482]= -1547955041;
assign addr[36483]= -1649974225;
assign addr[36484]= -1743623590;
assign addr[36485]= -1828428082;
assign addr[36486]= -1903957513;
assign addr[36487]= -1969828744;
assign addr[36488]= -2025707632;
assign addr[36489]= -2071310720;
assign addr[36490]= -2106406677;
assign addr[36491]= -2130817471;
assign addr[36492]= -2144419275;
assign addr[36493]= -2147143090;
assign addr[36494]= -2138975100;
assign addr[36495]= -2119956737;
assign addr[36496]= -2090184478;
assign addr[36497]= -2049809346;
assign addr[36498]= -1999036154;
assign addr[36499]= -1938122457;
assign addr[36500]= -1867377253;
assign addr[36501]= -1787159411;
assign addr[36502]= -1697875851;
assign addr[36503]= -1599979481;
assign addr[36504]= -1493966902;
assign addr[36505]= -1380375881;
assign addr[36506]= -1259782632;
assign addr[36507]= -1132798888;
assign addr[36508]= -1000068799;
assign addr[36509]= -862265664;
assign addr[36510]= -720088517;
assign addr[36511]= -574258580;
assign addr[36512]= -425515602;
assign addr[36513]= -274614114;
assign addr[36514]= -122319591;
assign addr[36515]= 30595422;
assign addr[36516]= 183355234;
assign addr[36517]= 335184940;
assign addr[36518]= 485314355;
assign addr[36519]= 632981917;
assign addr[36520]= 777438554;
assign addr[36521]= 917951481;
assign addr[36522]= 1053807919;
assign addr[36523]= 1184318708;
assign addr[36524]= 1308821808;
assign addr[36525]= 1426685652;
assign addr[36526]= 1537312353;
assign addr[36527]= 1640140734;
assign addr[36528]= 1734649179;
assign addr[36529]= 1820358275;
assign addr[36530]= 1896833245;
assign addr[36531]= 1963686155;
assign addr[36532]= 2020577882;
assign addr[36533]= 2067219829;
assign addr[36534]= 2103375398;
assign addr[36535]= 2128861181;
assign addr[36536]= 2143547897;
assign addr[36537]= 2147361045;
assign addr[36538]= 2140281282;
assign addr[36539]= 2122344521;
assign addr[36540]= 2093641749;
assign addr[36541]= 2054318569;
assign addr[36542]= 2004574453;
assign addr[36543]= 1944661739;
assign addr[36544]= 1874884346;
assign addr[36545]= 1795596234;
assign addr[36546]= 1707199606;
assign addr[36547]= 1610142873;
assign addr[36548]= 1504918373;
assign addr[36549]= 1392059879;
assign addr[36550]= 1272139887;
assign addr[36551]= 1145766716;
assign addr[36552]= 1013581418;
assign addr[36553]= 876254528;
assign addr[36554]= 734482665;
assign addr[36555]= 588984994;
assign addr[36556]= 440499581;
assign addr[36557]= 289779648;
assign addr[36558]= 137589750;
assign addr[36559]= -15298099;
assign addr[36560]= -168108346;
assign addr[36561]= -320065829;
assign addr[36562]= -470399716;
assign addr[36563]= -618347408;
assign addr[36564]= -763158411;
assign addr[36565]= -904098143;
assign addr[36566]= -1040451659;
assign addr[36567]= -1171527280;
assign addr[36568]= -1296660098;
assign addr[36569]= -1415215352;
assign addr[36570]= -1526591649;
assign addr[36571]= -1630224009;
assign addr[36572]= -1725586737;
assign addr[36573]= -1812196087;
assign addr[36574]= -1889612716;
assign addr[36575]= -1957443913;
assign addr[36576]= -2015345591;
assign addr[36577]= -2063024031;
assign addr[36578]= -2100237377;
assign addr[36579]= -2126796855;
assign addr[36580]= -2142567738;
assign addr[36581]= -2147470025;
assign addr[36582]= -2141478848;
assign addr[36583]= -2124624598;
assign addr[36584]= -2096992772;
assign addr[36585]= -2058723538;
assign addr[36586]= -2010011024;
assign addr[36587]= -1951102334;
assign addr[36588]= -1882296293;
assign addr[36589]= -1803941934;
assign addr[36590]= -1716436725;
assign addr[36591]= -1620224553;
assign addr[36592]= -1515793473;
assign addr[36593]= -1403673233;
assign addr[36594]= -1284432584;
assign addr[36595]= -1158676398;
assign addr[36596]= -1027042599;
assign addr[36597]= -890198924;
assign addr[36598]= -748839539;
assign addr[36599]= -603681519;
assign addr[36600]= -455461206;
assign addr[36601]= -304930476;
assign addr[36602]= -152852926;
assign addr[36603]= 0;
assign addr[36604]= 152852926;
assign addr[36605]= 304930476;
assign addr[36606]= 455461206;
assign addr[36607]= 603681519;
assign addr[36608]= 748839539;
assign addr[36609]= 890198924;
assign addr[36610]= 1027042599;
assign addr[36611]= 1158676398;
assign addr[36612]= 1284432584;
assign addr[36613]= 1403673233;
assign addr[36614]= 1515793473;
assign addr[36615]= 1620224553;
assign addr[36616]= 1716436725;
assign addr[36617]= 1803941934;
assign addr[36618]= 1882296293;
assign addr[36619]= 1951102334;
assign addr[36620]= 2010011024;
assign addr[36621]= 2058723538;
assign addr[36622]= 2096992772;
assign addr[36623]= 2124624598;
assign addr[36624]= 2141478848;
assign addr[36625]= 2147470025;
assign addr[36626]= 2142567738;
assign addr[36627]= 2126796855;
assign addr[36628]= 2100237377;
assign addr[36629]= 2063024031;
assign addr[36630]= 2015345591;
assign addr[36631]= 1957443913;
assign addr[36632]= 1889612716;
assign addr[36633]= 1812196087;
assign addr[36634]= 1725586737;
assign addr[36635]= 1630224009;
assign addr[36636]= 1526591649;
assign addr[36637]= 1415215352;
assign addr[36638]= 1296660098;
assign addr[36639]= 1171527280;
assign addr[36640]= 1040451659;
assign addr[36641]= 904098143;
assign addr[36642]= 763158411;
assign addr[36643]= 618347408;
assign addr[36644]= 470399716;
assign addr[36645]= 320065829;
assign addr[36646]= 168108346;
assign addr[36647]= 15298099;
assign addr[36648]= -137589750;
assign addr[36649]= -289779648;
assign addr[36650]= -440499581;
assign addr[36651]= -588984994;
assign addr[36652]= -734482665;
assign addr[36653]= -876254528;
assign addr[36654]= -1013581418;
assign addr[36655]= -1145766716;
assign addr[36656]= -1272139887;
assign addr[36657]= -1392059879;
assign addr[36658]= -1504918373;
assign addr[36659]= -1610142873;
assign addr[36660]= -1707199606;
assign addr[36661]= -1795596234;
assign addr[36662]= -1874884346;
assign addr[36663]= -1944661739;
assign addr[36664]= -2004574453;
assign addr[36665]= -2054318569;
assign addr[36666]= -2093641749;
assign addr[36667]= -2122344521;
assign addr[36668]= -2140281282;
assign addr[36669]= -2147361045;
assign addr[36670]= -2143547897;
assign addr[36671]= -2128861181;
assign addr[36672]= -2103375398;
assign addr[36673]= -2067219829;
assign addr[36674]= -2020577882;
assign addr[36675]= -1963686155;
assign addr[36676]= -1896833245;
assign addr[36677]= -1820358275;
assign addr[36678]= -1734649179;
assign addr[36679]= -1640140734;
assign addr[36680]= -1537312353;
assign addr[36681]= -1426685652;
assign addr[36682]= -1308821808;
assign addr[36683]= -1184318708;
assign addr[36684]= -1053807919;
assign addr[36685]= -917951481;
assign addr[36686]= -777438554;
assign addr[36687]= -632981917;
assign addr[36688]= -485314355;
assign addr[36689]= -335184940;
assign addr[36690]= -183355234;
assign addr[36691]= -30595422;
assign addr[36692]= 122319591;
assign addr[36693]= 274614114;
assign addr[36694]= 425515602;
assign addr[36695]= 574258580;
assign addr[36696]= 720088517;
assign addr[36697]= 862265664;
assign addr[36698]= 1000068799;
assign addr[36699]= 1132798888;
assign addr[36700]= 1259782632;
assign addr[36701]= 1380375881;
assign addr[36702]= 1493966902;
assign addr[36703]= 1599979481;
assign addr[36704]= 1697875851;
assign addr[36705]= 1787159411;
assign addr[36706]= 1867377253;
assign addr[36707]= 1938122457;
assign addr[36708]= 1999036154;
assign addr[36709]= 2049809346;
assign addr[36710]= 2090184478;
assign addr[36711]= 2119956737;
assign addr[36712]= 2138975100;
assign addr[36713]= 2147143090;
assign addr[36714]= 2144419275;
assign addr[36715]= 2130817471;
assign addr[36716]= 2106406677;
assign addr[36717]= 2071310720;
assign addr[36718]= 2025707632;
assign addr[36719]= 1969828744;
assign addr[36720]= 1903957513;
assign addr[36721]= 1828428082;
assign addr[36722]= 1743623590;
assign addr[36723]= 1649974225;
assign addr[36724]= 1547955041;
assign addr[36725]= 1438083551;
assign addr[36726]= 1320917099;
assign addr[36727]= 1197050035;
assign addr[36728]= 1067110699;
assign addr[36729]= 931758235;
assign addr[36730]= 791679244;
assign addr[36731]= 647584304;
assign addr[36732]= 500204365;
assign addr[36733]= 350287041;
assign addr[36734]= 198592817;
assign addr[36735]= 45891193;
assign addr[36736]= -107043224;
assign addr[36737]= -259434643;
assign addr[36738]= -410510029;
assign addr[36739]= -559503022;
assign addr[36740]= -705657826;
assign addr[36741]= -848233042;
assign addr[36742]= -986505429;
assign addr[36743]= -1119773573;
assign addr[36744]= -1247361445;
assign addr[36745]= -1368621831;
assign addr[36746]= -1482939614;
assign addr[36747]= -1589734894;
assign addr[36748]= -1688465931;
assign addr[36749]= -1778631892;
assign addr[36750]= -1859775393;
assign addr[36751]= -1931484818;
assign addr[36752]= -1993396407;
assign addr[36753]= -2045196100;
assign addr[36754]= -2086621133;
assign addr[36755]= -2117461370;
assign addr[36756]= -2137560369;
assign addr[36757]= -2146816171;
assign addr[36758]= -2145181827;
assign addr[36759]= -2132665626;
assign addr[36760]= -2109331059;
assign addr[36761]= -2075296495;
assign addr[36762]= -2030734582;
assign addr[36763]= -1975871368;
assign addr[36764]= -1910985158;
assign addr[36765]= -1836405100;
assign addr[36766]= -1752509516;
assign addr[36767]= -1659723983;
assign addr[36768]= -1558519173;
assign addr[36769]= -1449408469;
assign addr[36770]= -1332945355;
assign addr[36771]= -1209720613;
assign addr[36772]= -1080359326;
assign addr[36773]= -945517704;
assign addr[36774]= -805879757;
assign addr[36775]= -662153826;
assign addr[36776]= -515068990;
assign addr[36777]= -365371365;
assign addr[36778]= -213820322;
assign addr[36779]= -61184634;
assign addr[36780]= 91761426;
assign addr[36781]= 244242007;
assign addr[36782]= 395483624;
assign addr[36783]= 544719071;
assign addr[36784]= 691191324;
assign addr[36785]= 834157373;
assign addr[36786]= 972891995;
assign addr[36787]= 1106691431;
assign addr[36788]= 1234876957;
assign addr[36789]= 1356798326;
assign addr[36790]= 1471837070;
assign addr[36791]= 1579409630;
assign addr[36792]= 1678970324;
assign addr[36793]= 1770014111;
assign addr[36794]= 1852079154;
assign addr[36795]= 1924749160;
assign addr[36796]= 1987655498;
assign addr[36797]= 2040479063;
assign addr[36798]= 2082951896;
assign addr[36799]= 2114858546;
assign addr[36800]= 2136037160;
assign addr[36801]= 2146380306;
assign addr[36802]= 2145835515;
assign addr[36803]= 2134405552;
assign addr[36804]= 2112148396;
assign addr[36805]= 2079176953;
assign addr[36806]= 2035658475;
assign addr[36807]= 1981813720;
assign addr[36808]= 1917915825;
assign addr[36809]= 1844288924;
assign addr[36810]= 1761306505;
assign addr[36811]= 1669389513;
assign addr[36812]= 1569004214;
assign addr[36813]= 1460659832;
assign addr[36814]= 1344905966;
assign addr[36815]= 1222329801;
assign addr[36816]= 1093553126;
assign addr[36817]= 959229189;
assign addr[36818]= 820039373;
assign addr[36819]= 676689746;
assign addr[36820]= 529907477;
assign addr[36821]= 380437148;
assign addr[36822]= 229036977;
assign addr[36823]= 76474970;
assign addr[36824]= -76474970;
assign addr[36825]= -229036977;
assign addr[36826]= -380437148;
assign addr[36827]= -529907477;
assign addr[36828]= -676689746;
assign addr[36829]= -820039373;
assign addr[36830]= -959229189;
assign addr[36831]= -1093553126;
assign addr[36832]= -1222329801;
assign addr[36833]= -1344905966;
assign addr[36834]= -1460659832;
assign addr[36835]= -1569004214;
assign addr[36836]= -1669389513;
assign addr[36837]= -1761306505;
assign addr[36838]= -1844288924;
assign addr[36839]= -1917915825;
assign addr[36840]= -1981813720;
assign addr[36841]= -2035658475;
assign addr[36842]= -2079176953;
assign addr[36843]= -2112148396;
assign addr[36844]= -2134405552;
assign addr[36845]= -2145835515;
assign addr[36846]= -2146380306;
assign addr[36847]= -2136037160;
assign addr[36848]= -2114858546;
assign addr[36849]= -2082951896;
assign addr[36850]= -2040479063;
assign addr[36851]= -1987655498;
assign addr[36852]= -1924749160;
assign addr[36853]= -1852079154;
assign addr[36854]= -1770014111;
assign addr[36855]= -1678970324;
assign addr[36856]= -1579409630;
assign addr[36857]= -1471837070;
assign addr[36858]= -1356798326;
assign addr[36859]= -1234876957;
assign addr[36860]= -1106691431;
assign addr[36861]= -972891995;
assign addr[36862]= -834157373;
assign addr[36863]= -691191324;
assign addr[36864]= -544719071;
assign addr[36865]= -395483624;
assign addr[36866]= -244242007;
assign addr[36867]= -91761426;
assign addr[36868]= 61184634;
assign addr[36869]= 213820322;
assign addr[36870]= 365371365;
assign addr[36871]= 515068990;
assign addr[36872]= 662153826;
assign addr[36873]= 805879757;
assign addr[36874]= 945517704;
assign addr[36875]= 1080359326;
assign addr[36876]= 1209720613;
assign addr[36877]= 1332945355;
assign addr[36878]= 1449408469;
assign addr[36879]= 1558519173;
assign addr[36880]= 1659723983;
assign addr[36881]= 1752509516;
assign addr[36882]= 1836405100;
assign addr[36883]= 1910985158;
assign addr[36884]= 1975871368;
assign addr[36885]= 2030734582;
assign addr[36886]= 2075296495;
assign addr[36887]= 2109331059;
assign addr[36888]= 2132665626;
assign addr[36889]= 2145181827;
assign addr[36890]= 2146816171;
assign addr[36891]= 2137560369;
assign addr[36892]= 2117461370;
assign addr[36893]= 2086621133;
assign addr[36894]= 2045196100;
assign addr[36895]= 1993396407;
assign addr[36896]= 1931484818;
assign addr[36897]= 1859775393;
assign addr[36898]= 1778631892;
assign addr[36899]= 1688465931;
assign addr[36900]= 1589734894;
assign addr[36901]= 1482939614;
assign addr[36902]= 1368621831;
assign addr[36903]= 1247361445;
assign addr[36904]= 1119773573;
assign addr[36905]= 986505429;
assign addr[36906]= 848233042;
assign addr[36907]= 705657826;
assign addr[36908]= 559503022;
assign addr[36909]= 410510029;
assign addr[36910]= 259434643;
assign addr[36911]= 107043224;
assign addr[36912]= -45891193;
assign addr[36913]= -198592817;
assign addr[36914]= -350287041;
assign addr[36915]= -500204365;
assign addr[36916]= -647584304;
assign addr[36917]= -791679244;
assign addr[36918]= -931758235;
assign addr[36919]= -1067110699;
assign addr[36920]= -1197050035;
assign addr[36921]= -1320917099;
assign addr[36922]= -1438083551;
assign addr[36923]= -1547955041;
assign addr[36924]= -1649974225;
assign addr[36925]= -1743623590;
assign addr[36926]= -1828428082;
assign addr[36927]= -1903957513;
assign addr[36928]= -1969828744;
assign addr[36929]= -2025707632;
assign addr[36930]= -2071310720;
assign addr[36931]= -2106406677;
assign addr[36932]= -2130817471;
assign addr[36933]= -2144419275;
assign addr[36934]= -2147143090;
assign addr[36935]= -2138975100;
assign addr[36936]= -2119956737;
assign addr[36937]= -2090184478;
assign addr[36938]= -2049809346;
assign addr[36939]= -1999036154;
assign addr[36940]= -1938122457;
assign addr[36941]= -1867377253;
assign addr[36942]= -1787159411;
assign addr[36943]= -1697875851;
assign addr[36944]= -1599979481;
assign addr[36945]= -1493966902;
assign addr[36946]= -1380375881;
assign addr[36947]= -1259782632;
assign addr[36948]= -1132798888;
assign addr[36949]= -1000068799;
assign addr[36950]= -862265664;
assign addr[36951]= -720088517;
assign addr[36952]= -574258580;
assign addr[36953]= -425515602;
assign addr[36954]= -274614114;
assign addr[36955]= -122319591;
assign addr[36956]= 30595422;
assign addr[36957]= 183355234;
assign addr[36958]= 335184940;
assign addr[36959]= 485314355;
assign addr[36960]= 632981917;
assign addr[36961]= 777438554;
assign addr[36962]= 917951481;
assign addr[36963]= 1053807919;
assign addr[36964]= 1184318708;
assign addr[36965]= 1308821808;
assign addr[36966]= 1426685652;
assign addr[36967]= 1537312353;
assign addr[36968]= 1640140734;
assign addr[36969]= 1734649179;
assign addr[36970]= 1820358275;
assign addr[36971]= 1896833245;
assign addr[36972]= 1963686155;
assign addr[36973]= 2020577882;
assign addr[36974]= 2067219829;
assign addr[36975]= 2103375398;
assign addr[36976]= 2128861181;
assign addr[36977]= 2143547897;
assign addr[36978]= 2147361045;
assign addr[36979]= 2140281282;
assign addr[36980]= 2122344521;
assign addr[36981]= 2093641749;
assign addr[36982]= 2054318569;
assign addr[36983]= 2004574453;
assign addr[36984]= 1944661739;
assign addr[36985]= 1874884346;
assign addr[36986]= 1795596234;
assign addr[36987]= 1707199606;
assign addr[36988]= 1610142873;
assign addr[36989]= 1504918373;
assign addr[36990]= 1392059879;
assign addr[36991]= 1272139887;
assign addr[36992]= 1145766716;
assign addr[36993]= 1013581418;
assign addr[36994]= 876254528;
assign addr[36995]= 734482665;
assign addr[36996]= 588984994;
assign addr[36997]= 440499581;
assign addr[36998]= 289779648;
assign addr[36999]= 137589750;
assign addr[37000]= -15298099;
assign addr[37001]= -168108346;
assign addr[37002]= -320065829;
assign addr[37003]= -470399716;
assign addr[37004]= -618347408;
assign addr[37005]= -763158411;
assign addr[37006]= -904098143;
assign addr[37007]= -1040451659;
assign addr[37008]= -1171527280;
assign addr[37009]= -1296660098;
assign addr[37010]= -1415215352;
assign addr[37011]= -1526591649;
assign addr[37012]= -1630224009;
assign addr[37013]= -1725586737;
assign addr[37014]= -1812196087;
assign addr[37015]= -1889612716;
assign addr[37016]= -1957443913;
assign addr[37017]= -2015345591;
assign addr[37018]= -2063024031;
assign addr[37019]= -2100237377;
assign addr[37020]= -2126796855;
assign addr[37021]= -2142567738;
assign addr[37022]= -2147470025;
assign addr[37023]= -2141478848;
assign addr[37024]= -2124624598;
assign addr[37025]= -2096992772;
assign addr[37026]= -2058723538;
assign addr[37027]= -2010011024;
assign addr[37028]= -1951102334;
assign addr[37029]= -1882296293;
assign addr[37030]= -1803941934;
assign addr[37031]= -1716436725;
assign addr[37032]= -1620224553;
assign addr[37033]= -1515793473;
assign addr[37034]= -1403673233;
assign addr[37035]= -1284432584;
assign addr[37036]= -1158676398;
assign addr[37037]= -1027042599;
assign addr[37038]= -890198924;
assign addr[37039]= -748839539;
assign addr[37040]= -603681519;
assign addr[37041]= -455461206;
assign addr[37042]= -304930476;
assign addr[37043]= -152852926;
assign addr[37044]= 0;
assign addr[37045]= 152852926;
assign addr[37046]= 304930476;
assign addr[37047]= 455461206;
assign addr[37048]= 603681519;
assign addr[37049]= 748839539;
assign addr[37050]= 890198924;
assign addr[37051]= 1027042599;
assign addr[37052]= 1158676398;
assign addr[37053]= 1284432584;
assign addr[37054]= 1403673233;
assign addr[37055]= 1515793473;
assign addr[37056]= 1620224553;
assign addr[37057]= 1716436725;
assign addr[37058]= 1803941934;
assign addr[37059]= 1882296293;
assign addr[37060]= 1951102334;
assign addr[37061]= 2010011024;
assign addr[37062]= 2058723538;
assign addr[37063]= 2096992772;
assign addr[37064]= 2124624598;
assign addr[37065]= 2141478848;
assign addr[37066]= 2147470025;
assign addr[37067]= 2142567738;
assign addr[37068]= 2126796855;
assign addr[37069]= 2100237377;
assign addr[37070]= 2063024031;
assign addr[37071]= 2015345591;
assign addr[37072]= 1957443913;
assign addr[37073]= 1889612716;
assign addr[37074]= 1812196087;
assign addr[37075]= 1725586737;
assign addr[37076]= 1630224009;
assign addr[37077]= 1526591649;
assign addr[37078]= 1415215352;
assign addr[37079]= 1296660098;
assign addr[37080]= 1171527280;
assign addr[37081]= 1040451659;
assign addr[37082]= 904098143;
assign addr[37083]= 763158411;
assign addr[37084]= 618347408;
assign addr[37085]= 470399716;
assign addr[37086]= 320065829;
assign addr[37087]= 168108346;
assign addr[37088]= 15298099;
assign addr[37089]= -137589750;
assign addr[37090]= -289779648;
assign addr[37091]= -440499581;
assign addr[37092]= -588984994;
assign addr[37093]= -734482665;
assign addr[37094]= -876254528;
assign addr[37095]= -1013581418;
assign addr[37096]= -1145766716;
assign addr[37097]= -1272139887;
assign addr[37098]= -1392059879;
assign addr[37099]= -1504918373;
assign addr[37100]= -1610142873;
assign addr[37101]= -1707199606;
assign addr[37102]= -1795596234;
assign addr[37103]= -1874884346;
assign addr[37104]= -1944661739;
assign addr[37105]= -2004574453;
assign addr[37106]= -2054318569;
assign addr[37107]= -2093641749;
assign addr[37108]= -2122344521;
assign addr[37109]= -2140281282;
assign addr[37110]= -2147361045;
assign addr[37111]= -2143547897;
assign addr[37112]= -2128861181;
assign addr[37113]= -2103375398;
assign addr[37114]= -2067219829;
assign addr[37115]= -2020577882;
assign addr[37116]= -1963686155;
assign addr[37117]= -1896833245;
assign addr[37118]= -1820358275;
assign addr[37119]= -1734649179;
assign addr[37120]= -1640140734;
assign addr[37121]= -1537312353;
assign addr[37122]= -1426685652;
assign addr[37123]= -1308821808;
assign addr[37124]= -1184318708;
assign addr[37125]= -1053807919;
assign addr[37126]= -917951481;
assign addr[37127]= -777438554;
assign addr[37128]= -632981917;
assign addr[37129]= -485314355;
assign addr[37130]= -335184940;
assign addr[37131]= -183355234;
assign addr[37132]= -30595422;
assign addr[37133]= 122319591;
assign addr[37134]= 274614114;
assign addr[37135]= 425515602;
assign addr[37136]= 574258580;
assign addr[37137]= 720088517;
assign addr[37138]= 862265664;
assign addr[37139]= 1000068799;
assign addr[37140]= 1132798888;
assign addr[37141]= 1259782632;
assign addr[37142]= 1380375881;
assign addr[37143]= 1493966902;
assign addr[37144]= 1599979481;
assign addr[37145]= 1697875851;
assign addr[37146]= 1787159411;
assign addr[37147]= 1867377253;
assign addr[37148]= 1938122457;
assign addr[37149]= 1999036154;
assign addr[37150]= 2049809346;
assign addr[37151]= 2090184478;
assign addr[37152]= 2119956737;
assign addr[37153]= 2138975100;
assign addr[37154]= 2147143090;
assign addr[37155]= 2144419275;
assign addr[37156]= 2130817471;
assign addr[37157]= 2106406677;
assign addr[37158]= 2071310720;
assign addr[37159]= 2025707632;
assign addr[37160]= 1969828744;
assign addr[37161]= 1903957513;
assign addr[37162]= 1828428082;
assign addr[37163]= 1743623590;
assign addr[37164]= 1649974225;
assign addr[37165]= 1547955041;
assign addr[37166]= 1438083551;
assign addr[37167]= 1320917099;
assign addr[37168]= 1197050035;
assign addr[37169]= 1067110699;
assign addr[37170]= 931758235;
assign addr[37171]= 791679244;
assign addr[37172]= 647584304;
assign addr[37173]= 500204365;
assign addr[37174]= 350287041;
assign addr[37175]= 198592817;
assign addr[37176]= 45891193;
assign addr[37177]= -107043224;
assign addr[37178]= -259434643;
assign addr[37179]= -410510029;
assign addr[37180]= -559503022;
assign addr[37181]= -705657826;
assign addr[37182]= -848233042;
assign addr[37183]= -986505429;
assign addr[37184]= -1119773573;
assign addr[37185]= -1247361445;
assign addr[37186]= -1368621831;
assign addr[37187]= -1482939614;
assign addr[37188]= -1589734894;
assign addr[37189]= -1688465931;
assign addr[37190]= -1778631892;
assign addr[37191]= -1859775393;
assign addr[37192]= -1931484818;
assign addr[37193]= -1993396407;
assign addr[37194]= -2045196100;
assign addr[37195]= -2086621133;
assign addr[37196]= -2117461370;
assign addr[37197]= -2137560369;
assign addr[37198]= -2146816171;
assign addr[37199]= -2145181827;
assign addr[37200]= -2132665626;
assign addr[37201]= -2109331059;
assign addr[37202]= -2075296495;
assign addr[37203]= -2030734582;
assign addr[37204]= -1975871368;
assign addr[37205]= -1910985158;
assign addr[37206]= -1836405100;
assign addr[37207]= -1752509516;
assign addr[37208]= -1659723983;
assign addr[37209]= -1558519173;
assign addr[37210]= -1449408469;
assign addr[37211]= -1332945355;
assign addr[37212]= -1209720613;
assign addr[37213]= -1080359326;
assign addr[37214]= -945517704;
assign addr[37215]= -805879757;
assign addr[37216]= -662153826;
assign addr[37217]= -515068990;
assign addr[37218]= -365371365;
assign addr[37219]= -213820322;
assign addr[37220]= -61184634;
assign addr[37221]= 91761426;
assign addr[37222]= 244242007;
assign addr[37223]= 395483624;
assign addr[37224]= 544719071;
assign addr[37225]= 691191324;
assign addr[37226]= 834157373;
assign addr[37227]= 972891995;
assign addr[37228]= 1106691431;
assign addr[37229]= 1234876957;
assign addr[37230]= 1356798326;
assign addr[37231]= 1471837070;
assign addr[37232]= 1579409630;
assign addr[37233]= 1678970324;
assign addr[37234]= 1770014111;
assign addr[37235]= 1852079154;
assign addr[37236]= 1924749160;
assign addr[37237]= 1987655498;
assign addr[37238]= 2040479063;
assign addr[37239]= 2082951896;
assign addr[37240]= 2114858546;
assign addr[37241]= 2136037160;
assign addr[37242]= 2146380306;
assign addr[37243]= 2145835515;
assign addr[37244]= 2134405552;
assign addr[37245]= 2112148396;
assign addr[37246]= 2079176953;
assign addr[37247]= 2035658475;
assign addr[37248]= 1981813720;
assign addr[37249]= 1917915825;
assign addr[37250]= 1844288924;
assign addr[37251]= 1761306505;
assign addr[37252]= 1669389513;
assign addr[37253]= 1569004214;
assign addr[37254]= 1460659832;
assign addr[37255]= 1344905966;
assign addr[37256]= 1222329801;
assign addr[37257]= 1093553126;
assign addr[37258]= 959229189;
assign addr[37259]= 820039373;
assign addr[37260]= 676689746;
assign addr[37261]= 529907477;
assign addr[37262]= 380437148;
assign addr[37263]= 229036977;
assign addr[37264]= 76474970;
assign addr[37265]= -76474970;
assign addr[37266]= -229036977;
assign addr[37267]= -380437148;
assign addr[37268]= -529907477;
assign addr[37269]= -676689746;
assign addr[37270]= -820039373;
assign addr[37271]= -959229189;
assign addr[37272]= -1093553126;
assign addr[37273]= -1222329801;
assign addr[37274]= -1344905966;
assign addr[37275]= -1460659832;
assign addr[37276]= -1569004214;
assign addr[37277]= -1669389513;
assign addr[37278]= -1761306505;
assign addr[37279]= -1844288924;
assign addr[37280]= -1917915825;
assign addr[37281]= -1981813720;
assign addr[37282]= -2035658475;
assign addr[37283]= -2079176953;
assign addr[37284]= -2112148396;
assign addr[37285]= -2134405552;
assign addr[37286]= -2145835515;
assign addr[37287]= -2146380306;
assign addr[37288]= -2136037160;
assign addr[37289]= -2114858546;
assign addr[37290]= -2082951896;
assign addr[37291]= -2040479063;
assign addr[37292]= -1987655498;
assign addr[37293]= -1924749160;
assign addr[37294]= -1852079154;
assign addr[37295]= -1770014111;
assign addr[37296]= -1678970324;
assign addr[37297]= -1579409630;
assign addr[37298]= -1471837070;
assign addr[37299]= -1356798326;
assign addr[37300]= -1234876957;
assign addr[37301]= -1106691431;
assign addr[37302]= -972891995;
assign addr[37303]= -834157373;
assign addr[37304]= -691191324;
assign addr[37305]= -544719071;
assign addr[37306]= -395483624;
assign addr[37307]= -244242007;
assign addr[37308]= -91761426;
assign addr[37309]= 61184634;
assign addr[37310]= 213820322;
assign addr[37311]= 365371365;
assign addr[37312]= 515068990;
assign addr[37313]= 662153826;
assign addr[37314]= 805879757;
assign addr[37315]= 945517704;
assign addr[37316]= 1080359326;
assign addr[37317]= 1209720613;
assign addr[37318]= 1332945355;
assign addr[37319]= 1449408469;
assign addr[37320]= 1558519173;
assign addr[37321]= 1659723983;
assign addr[37322]= 1752509516;
assign addr[37323]= 1836405100;
assign addr[37324]= 1910985158;
assign addr[37325]= 1975871368;
assign addr[37326]= 2030734582;
assign addr[37327]= 2075296495;
assign addr[37328]= 2109331059;
assign addr[37329]= 2132665626;
assign addr[37330]= 2145181827;
assign addr[37331]= 2146816171;
assign addr[37332]= 2137560369;
assign addr[37333]= 2117461370;
assign addr[37334]= 2086621133;
assign addr[37335]= 2045196100;
assign addr[37336]= 1993396407;
assign addr[37337]= 1931484818;
assign addr[37338]= 1859775393;
assign addr[37339]= 1778631892;
assign addr[37340]= 1688465931;
assign addr[37341]= 1589734894;
assign addr[37342]= 1482939614;
assign addr[37343]= 1368621831;
assign addr[37344]= 1247361445;
assign addr[37345]= 1119773573;
assign addr[37346]= 986505429;
assign addr[37347]= 848233042;
assign addr[37348]= 705657826;
assign addr[37349]= 559503022;
assign addr[37350]= 410510029;
assign addr[37351]= 259434643;
assign addr[37352]= 107043224;
assign addr[37353]= -45891193;
assign addr[37354]= -198592817;
assign addr[37355]= -350287041;
assign addr[37356]= -500204365;
assign addr[37357]= -647584304;
assign addr[37358]= -791679244;
assign addr[37359]= -931758235;
assign addr[37360]= -1067110699;
assign addr[37361]= -1197050035;
assign addr[37362]= -1320917099;
assign addr[37363]= -1438083551;
assign addr[37364]= -1547955041;
assign addr[37365]= -1649974225;
assign addr[37366]= -1743623590;
assign addr[37367]= -1828428082;
assign addr[37368]= -1903957513;
assign addr[37369]= -1969828744;
assign addr[37370]= -2025707632;
assign addr[37371]= -2071310720;
assign addr[37372]= -2106406677;
assign addr[37373]= -2130817471;
assign addr[37374]= -2144419275;
assign addr[37375]= -2147143090;
assign addr[37376]= -2138975100;
assign addr[37377]= -2119956737;
assign addr[37378]= -2090184478;
assign addr[37379]= -2049809346;
assign addr[37380]= -1999036154;
assign addr[37381]= -1938122457;
assign addr[37382]= -1867377253;
assign addr[37383]= -1787159411;
assign addr[37384]= -1697875851;
assign addr[37385]= -1599979481;
assign addr[37386]= -1493966902;
assign addr[37387]= -1380375881;
assign addr[37388]= -1259782632;
assign addr[37389]= -1132798888;
assign addr[37390]= -1000068799;
assign addr[37391]= -862265664;
assign addr[37392]= -720088517;
assign addr[37393]= -574258580;
assign addr[37394]= -425515602;
assign addr[37395]= -274614114;
assign addr[37396]= -122319591;
assign addr[37397]= 30595422;
assign addr[37398]= 183355234;
assign addr[37399]= 335184940;
assign addr[37400]= 485314355;
assign addr[37401]= 632981917;
assign addr[37402]= 777438554;
assign addr[37403]= 917951481;
assign addr[37404]= 1053807919;
assign addr[37405]= 1184318708;
assign addr[37406]= 1308821808;
assign addr[37407]= 1426685652;
assign addr[37408]= 1537312353;
assign addr[37409]= 1640140734;
assign addr[37410]= 1734649179;
assign addr[37411]= 1820358275;
assign addr[37412]= 1896833245;
assign addr[37413]= 1963686155;
assign addr[37414]= 2020577882;
assign addr[37415]= 2067219829;
assign addr[37416]= 2103375398;
assign addr[37417]= 2128861181;
assign addr[37418]= 2143547897;
assign addr[37419]= 2147361045;
assign addr[37420]= 2140281282;
assign addr[37421]= 2122344521;
assign addr[37422]= 2093641749;
assign addr[37423]= 2054318569;
assign addr[37424]= 2004574453;
assign addr[37425]= 1944661739;
assign addr[37426]= 1874884346;
assign addr[37427]= 1795596234;
assign addr[37428]= 1707199606;
assign addr[37429]= 1610142873;
assign addr[37430]= 1504918373;
assign addr[37431]= 1392059879;
assign addr[37432]= 1272139887;
assign addr[37433]= 1145766716;
assign addr[37434]= 1013581418;
assign addr[37435]= 876254528;
assign addr[37436]= 734482665;
assign addr[37437]= 588984994;
assign addr[37438]= 440499581;
assign addr[37439]= 289779648;
assign addr[37440]= 137589750;
assign addr[37441]= -15298099;
assign addr[37442]= -168108346;
assign addr[37443]= -320065829;
assign addr[37444]= -470399716;
assign addr[37445]= -618347408;
assign addr[37446]= -763158411;
assign addr[37447]= -904098143;
assign addr[37448]= -1040451659;
assign addr[37449]= -1171527280;
assign addr[37450]= -1296660098;
assign addr[37451]= -1415215352;
assign addr[37452]= -1526591649;
assign addr[37453]= -1630224009;
assign addr[37454]= -1725586737;
assign addr[37455]= -1812196087;
assign addr[37456]= -1889612716;
assign addr[37457]= -1957443913;
assign addr[37458]= -2015345591;
assign addr[37459]= -2063024031;
assign addr[37460]= -2100237377;
assign addr[37461]= -2126796855;
assign addr[37462]= -2142567738;
assign addr[37463]= -2147470025;
assign addr[37464]= -2141478848;
assign addr[37465]= -2124624598;
assign addr[37466]= -2096992772;
assign addr[37467]= -2058723538;
assign addr[37468]= -2010011024;
assign addr[37469]= -1951102334;
assign addr[37470]= -1882296293;
assign addr[37471]= -1803941934;
assign addr[37472]= -1716436725;
assign addr[37473]= -1620224553;
assign addr[37474]= -1515793473;
assign addr[37475]= -1403673233;
assign addr[37476]= -1284432584;
assign addr[37477]= -1158676398;
assign addr[37478]= -1027042599;
assign addr[37479]= -890198924;
assign addr[37480]= -748839539;
assign addr[37481]= -603681519;
assign addr[37482]= -455461206;
assign addr[37483]= -304930476;
assign addr[37484]= -152852926;
assign addr[37485]= 0;
assign addr[37486]= 152852926;
assign addr[37487]= 304930476;
assign addr[37488]= 455461206;
assign addr[37489]= 603681519;
assign addr[37490]= 748839539;
assign addr[37491]= 890198924;
assign addr[37492]= 1027042599;
assign addr[37493]= 1158676398;
assign addr[37494]= 1284432584;
assign addr[37495]= 1403673233;
assign addr[37496]= 1515793473;
assign addr[37497]= 1620224553;
assign addr[37498]= 1716436725;
assign addr[37499]= 1803941934;
assign addr[37500]= 1882296293;
assign addr[37501]= 1951102334;
assign addr[37502]= 2010011024;
assign addr[37503]= 2058723538;
assign addr[37504]= 2096992772;
assign addr[37505]= 2124624598;
assign addr[37506]= 2141478848;
assign addr[37507]= 2147470025;
assign addr[37508]= 2142567738;
assign addr[37509]= 2126796855;
assign addr[37510]= 2100237377;
assign addr[37511]= 2063024031;
assign addr[37512]= 2015345591;
assign addr[37513]= 1957443913;
assign addr[37514]= 1889612716;
assign addr[37515]= 1812196087;
assign addr[37516]= 1725586737;
assign addr[37517]= 1630224009;
assign addr[37518]= 1526591649;
assign addr[37519]= 1415215352;
assign addr[37520]= 1296660098;
assign addr[37521]= 1171527280;
assign addr[37522]= 1040451659;
assign addr[37523]= 904098143;
assign addr[37524]= 763158411;
assign addr[37525]= 618347408;
assign addr[37526]= 470399716;
assign addr[37527]= 320065829;
assign addr[37528]= 168108346;
assign addr[37529]= 15298099;
assign addr[37530]= -137589750;
assign addr[37531]= -289779648;
assign addr[37532]= -440499581;
assign addr[37533]= -588984994;
assign addr[37534]= -734482665;
assign addr[37535]= -876254528;
assign addr[37536]= -1013581418;
assign addr[37537]= -1145766716;
assign addr[37538]= -1272139887;
assign addr[37539]= -1392059879;
assign addr[37540]= -1504918373;
assign addr[37541]= -1610142873;
assign addr[37542]= -1707199606;
assign addr[37543]= -1795596234;
assign addr[37544]= -1874884346;
assign addr[37545]= -1944661739;
assign addr[37546]= -2004574453;
assign addr[37547]= -2054318569;
assign addr[37548]= -2093641749;
assign addr[37549]= -2122344521;
assign addr[37550]= -2140281282;
assign addr[37551]= -2147361045;
assign addr[37552]= -2143547897;
assign addr[37553]= -2128861181;
assign addr[37554]= -2103375398;
assign addr[37555]= -2067219829;
assign addr[37556]= -2020577882;
assign addr[37557]= -1963686155;
assign addr[37558]= -1896833245;
assign addr[37559]= -1820358275;
assign addr[37560]= -1734649179;
assign addr[37561]= -1640140734;
assign addr[37562]= -1537312353;
assign addr[37563]= -1426685652;
assign addr[37564]= -1308821808;
assign addr[37565]= -1184318708;
assign addr[37566]= -1053807919;
assign addr[37567]= -917951481;
assign addr[37568]= -777438554;
assign addr[37569]= -632981917;
assign addr[37570]= -485314355;
assign addr[37571]= -335184940;
assign addr[37572]= -183355234;
assign addr[37573]= -30595422;
assign addr[37574]= 122319591;
assign addr[37575]= 274614114;
assign addr[37576]= 425515602;
assign addr[37577]= 574258580;
assign addr[37578]= 720088517;
assign addr[37579]= 862265664;
assign addr[37580]= 1000068799;
assign addr[37581]= 1132798888;
assign addr[37582]= 1259782632;
assign addr[37583]= 1380375881;
assign addr[37584]= 1493966902;
assign addr[37585]= 1599979481;
assign addr[37586]= 1697875851;
assign addr[37587]= 1787159411;
assign addr[37588]= 1867377253;
assign addr[37589]= 1938122457;
assign addr[37590]= 1999036154;
assign addr[37591]= 2049809346;
assign addr[37592]= 2090184478;
assign addr[37593]= 2119956737;
assign addr[37594]= 2138975100;
assign addr[37595]= 2147143090;
assign addr[37596]= 2144419275;
assign addr[37597]= 2130817471;
assign addr[37598]= 2106406677;
assign addr[37599]= 2071310720;
assign addr[37600]= 2025707632;
assign addr[37601]= 1969828744;
assign addr[37602]= 1903957513;
assign addr[37603]= 1828428082;
assign addr[37604]= 1743623590;
assign addr[37605]= 1649974225;
assign addr[37606]= 1547955041;
assign addr[37607]= 1438083551;
assign addr[37608]= 1320917099;
assign addr[37609]= 1197050035;
assign addr[37610]= 1067110699;
assign addr[37611]= 931758235;
assign addr[37612]= 791679244;
assign addr[37613]= 647584304;
assign addr[37614]= 500204365;
assign addr[37615]= 350287041;
assign addr[37616]= 198592817;
assign addr[37617]= 45891193;
assign addr[37618]= -107043224;
assign addr[37619]= -259434643;
assign addr[37620]= -410510029;
assign addr[37621]= -559503022;
assign addr[37622]= -705657826;
assign addr[37623]= -848233042;
assign addr[37624]= -986505429;
assign addr[37625]= -1119773573;
assign addr[37626]= -1247361445;
assign addr[37627]= -1368621831;
assign addr[37628]= -1482939614;
assign addr[37629]= -1589734894;
assign addr[37630]= -1688465931;
assign addr[37631]= -1778631892;
assign addr[37632]= -1859775393;
assign addr[37633]= -1931484818;
assign addr[37634]= -1993396407;
assign addr[37635]= -2045196100;
assign addr[37636]= -2086621133;
assign addr[37637]= -2117461370;
assign addr[37638]= -2137560369;
assign addr[37639]= -2146816171;
assign addr[37640]= -2145181827;
assign addr[37641]= -2132665626;
assign addr[37642]= -2109331059;
assign addr[37643]= -2075296495;
assign addr[37644]= -2030734582;
assign addr[37645]= -1975871368;
assign addr[37646]= -1910985158;
assign addr[37647]= -1836405100;
assign addr[37648]= -1752509516;
assign addr[37649]= -1659723983;
assign addr[37650]= -1558519173;
assign addr[37651]= -1449408469;
assign addr[37652]= -1332945355;
assign addr[37653]= -1209720613;
assign addr[37654]= -1080359326;
assign addr[37655]= -945517704;
assign addr[37656]= -805879757;
assign addr[37657]= -662153826;
assign addr[37658]= -515068990;
assign addr[37659]= -365371365;
assign addr[37660]= -213820322;
assign addr[37661]= -61184634;
assign addr[37662]= 91761426;
assign addr[37663]= 244242007;
assign addr[37664]= 395483624;
assign addr[37665]= 544719071;
assign addr[37666]= 691191324;
assign addr[37667]= 834157373;
assign addr[37668]= 972891995;
assign addr[37669]= 1106691431;
assign addr[37670]= 1234876957;
assign addr[37671]= 1356798326;
assign addr[37672]= 1471837070;
assign addr[37673]= 1579409630;
assign addr[37674]= 1678970324;
assign addr[37675]= 1770014111;
assign addr[37676]= 1852079154;
assign addr[37677]= 1924749160;
assign addr[37678]= 1987655498;
assign addr[37679]= 2040479063;
assign addr[37680]= 2082951896;
assign addr[37681]= 2114858546;
assign addr[37682]= 2136037160;
assign addr[37683]= 2146380306;
assign addr[37684]= 2145835515;
assign addr[37685]= 2134405552;
assign addr[37686]= 2112148396;
assign addr[37687]= 2079176953;
assign addr[37688]= 2035658475;
assign addr[37689]= 1981813720;
assign addr[37690]= 1917915825;
assign addr[37691]= 1844288924;
assign addr[37692]= 1761306505;
assign addr[37693]= 1669389513;
assign addr[37694]= 1569004214;
assign addr[37695]= 1460659832;
assign addr[37696]= 1344905966;
assign addr[37697]= 1222329801;
assign addr[37698]= 1093553126;
assign addr[37699]= 959229189;
assign addr[37700]= 820039373;
assign addr[37701]= 676689746;
assign addr[37702]= 529907477;
assign addr[37703]= 380437148;
assign addr[37704]= 229036977;
assign addr[37705]= 76474970;
assign addr[37706]= -76474970;
assign addr[37707]= -229036977;
assign addr[37708]= -380437148;
assign addr[37709]= -529907477;
assign addr[37710]= -676689746;
assign addr[37711]= -820039373;
assign addr[37712]= -959229189;
assign addr[37713]= -1093553126;
assign addr[37714]= -1222329801;
assign addr[37715]= -1344905966;
assign addr[37716]= -1460659832;
assign addr[37717]= -1569004214;
assign addr[37718]= -1669389513;
assign addr[37719]= -1761306505;
assign addr[37720]= -1844288924;
assign addr[37721]= -1917915825;
assign addr[37722]= -1981813720;
assign addr[37723]= -2035658475;
assign addr[37724]= -2079176953;
assign addr[37725]= -2112148396;
assign addr[37726]= -2134405552;
assign addr[37727]= -2145835515;
assign addr[37728]= -2146380306;
assign addr[37729]= -2136037160;
assign addr[37730]= -2114858546;
assign addr[37731]= -2082951896;
assign addr[37732]= -2040479063;
assign addr[37733]= -1987655498;
assign addr[37734]= -1924749160;
assign addr[37735]= -1852079154;
assign addr[37736]= -1770014111;
assign addr[37737]= -1678970324;
assign addr[37738]= -1579409630;
assign addr[37739]= -1471837070;
assign addr[37740]= -1356798326;
assign addr[37741]= -1234876957;
assign addr[37742]= -1106691431;
assign addr[37743]= -972891995;
assign addr[37744]= -834157373;
assign addr[37745]= -691191324;
assign addr[37746]= -544719071;
assign addr[37747]= -395483624;
assign addr[37748]= -244242007;
assign addr[37749]= -91761426;
assign addr[37750]= 61184634;
assign addr[37751]= 213820322;
assign addr[37752]= 365371365;
assign addr[37753]= 515068990;
assign addr[37754]= 662153826;
assign addr[37755]= 805879757;
assign addr[37756]= 945517704;
assign addr[37757]= 1080359326;
assign addr[37758]= 1209720613;
assign addr[37759]= 1332945355;
assign addr[37760]= 1449408469;
assign addr[37761]= 1558519173;
assign addr[37762]= 1659723983;
assign addr[37763]= 1752509516;
assign addr[37764]= 1836405100;
assign addr[37765]= 1910985158;
assign addr[37766]= 1975871368;
assign addr[37767]= 2030734582;
assign addr[37768]= 2075296495;
assign addr[37769]= 2109331059;
assign addr[37770]= 2132665626;
assign addr[37771]= 2145181827;
assign addr[37772]= 2146816171;
assign addr[37773]= 2137560369;
assign addr[37774]= 2117461370;
assign addr[37775]= 2086621133;
assign addr[37776]= 2045196100;
assign addr[37777]= 1993396407;
assign addr[37778]= 1931484818;
assign addr[37779]= 1859775393;
assign addr[37780]= 1778631892;
assign addr[37781]= 1688465931;
assign addr[37782]= 1589734894;
assign addr[37783]= 1482939614;
assign addr[37784]= 1368621831;
assign addr[37785]= 1247361445;
assign addr[37786]= 1119773573;
assign addr[37787]= 986505429;
assign addr[37788]= 848233042;
assign addr[37789]= 705657826;
assign addr[37790]= 559503022;
assign addr[37791]= 410510029;
assign addr[37792]= 259434643;
assign addr[37793]= 107043224;
assign addr[37794]= -45891193;
assign addr[37795]= -198592817;
assign addr[37796]= -350287041;
assign addr[37797]= -500204365;
assign addr[37798]= -647584304;
assign addr[37799]= -791679244;
assign addr[37800]= -931758235;
assign addr[37801]= -1067110699;
assign addr[37802]= -1197050035;
assign addr[37803]= -1320917099;
assign addr[37804]= -1438083551;
assign addr[37805]= -1547955041;
assign addr[37806]= -1649974225;
assign addr[37807]= -1743623590;
assign addr[37808]= -1828428082;
assign addr[37809]= -1903957513;
assign addr[37810]= -1969828744;
assign addr[37811]= -2025707632;
assign addr[37812]= -2071310720;
assign addr[37813]= -2106406677;
assign addr[37814]= -2130817471;
assign addr[37815]= -2144419275;
assign addr[37816]= -2147143090;
assign addr[37817]= -2138975100;
assign addr[37818]= -2119956737;
assign addr[37819]= -2090184478;
assign addr[37820]= -2049809346;
assign addr[37821]= -1999036154;
assign addr[37822]= -1938122457;
assign addr[37823]= -1867377253;
assign addr[37824]= -1787159411;
assign addr[37825]= -1697875851;
assign addr[37826]= -1599979481;
assign addr[37827]= -1493966902;
assign addr[37828]= -1380375881;
assign addr[37829]= -1259782632;
assign addr[37830]= -1132798888;
assign addr[37831]= -1000068799;
assign addr[37832]= -862265664;
assign addr[37833]= -720088517;
assign addr[37834]= -574258580;
assign addr[37835]= -425515602;
assign addr[37836]= -274614114;
assign addr[37837]= -122319591;
assign addr[37838]= 30595422;
assign addr[37839]= 183355234;
assign addr[37840]= 335184940;
assign addr[37841]= 485314355;
assign addr[37842]= 632981917;
assign addr[37843]= 777438554;
assign addr[37844]= 917951481;
assign addr[37845]= 1053807919;
assign addr[37846]= 1184318708;
assign addr[37847]= 1308821808;
assign addr[37848]= 1426685652;
assign addr[37849]= 1537312353;
assign addr[37850]= 1640140734;
assign addr[37851]= 1734649179;
assign addr[37852]= 1820358275;
assign addr[37853]= 1896833245;
assign addr[37854]= 1963686155;
assign addr[37855]= 2020577882;
assign addr[37856]= 2067219829;
assign addr[37857]= 2103375398;
assign addr[37858]= 2128861181;
assign addr[37859]= 2143547897;
assign addr[37860]= 2147361045;
assign addr[37861]= 2140281282;
assign addr[37862]= 2122344521;
assign addr[37863]= 2093641749;
assign addr[37864]= 2054318569;
assign addr[37865]= 2004574453;
assign addr[37866]= 1944661739;
assign addr[37867]= 1874884346;
assign addr[37868]= 1795596234;
assign addr[37869]= 1707199606;
assign addr[37870]= 1610142873;
assign addr[37871]= 1504918373;
assign addr[37872]= 1392059879;
assign addr[37873]= 1272139887;
assign addr[37874]= 1145766716;
assign addr[37875]= 1013581418;
assign addr[37876]= 876254528;
assign addr[37877]= 734482665;
assign addr[37878]= 588984994;
assign addr[37879]= 440499581;
assign addr[37880]= 289779648;
assign addr[37881]= 137589750;
assign addr[37882]= -15298099;
assign addr[37883]= -168108346;
assign addr[37884]= -320065829;
assign addr[37885]= -470399716;
assign addr[37886]= -618347408;
assign addr[37887]= -763158411;
assign addr[37888]= -904098143;
assign addr[37889]= -1040451659;
assign addr[37890]= -1171527280;
assign addr[37891]= -1296660098;
assign addr[37892]= -1415215352;
assign addr[37893]= -1526591649;
assign addr[37894]= -1630224009;
assign addr[37895]= -1725586737;
assign addr[37896]= -1812196087;
assign addr[37897]= -1889612716;
assign addr[37898]= -1957443913;
assign addr[37899]= -2015345591;
assign addr[37900]= -2063024031;
assign addr[37901]= -2100237377;
assign addr[37902]= -2126796855;
assign addr[37903]= -2142567738;
assign addr[37904]= -2147470025;
assign addr[37905]= -2141478848;
assign addr[37906]= -2124624598;
assign addr[37907]= -2096992772;
assign addr[37908]= -2058723538;
assign addr[37909]= -2010011024;
assign addr[37910]= -1951102334;
assign addr[37911]= -1882296293;
assign addr[37912]= -1803941934;
assign addr[37913]= -1716436725;
assign addr[37914]= -1620224553;
assign addr[37915]= -1515793473;
assign addr[37916]= -1403673233;
assign addr[37917]= -1284432584;
assign addr[37918]= -1158676398;
assign addr[37919]= -1027042599;
assign addr[37920]= -890198924;
assign addr[37921]= -748839539;
assign addr[37922]= -603681519;
assign addr[37923]= -455461206;
assign addr[37924]= -304930476;
assign addr[37925]= -152852926;
assign addr[37926]= 0;
assign addr[37927]= 152852926;
assign addr[37928]= 304930476;
assign addr[37929]= 455461206;
assign addr[37930]= 603681519;
assign addr[37931]= 748839539;
assign addr[37932]= 890198924;
assign addr[37933]= 1027042599;
assign addr[37934]= 1158676398;
assign addr[37935]= 1284432584;
assign addr[37936]= 1403673233;
assign addr[37937]= 1515793473;
assign addr[37938]= 1620224553;
assign addr[37939]= 1716436725;
assign addr[37940]= 1803941934;
assign addr[37941]= 1882296293;
assign addr[37942]= 1951102334;
assign addr[37943]= 2010011024;
assign addr[37944]= 2058723538;
assign addr[37945]= 2096992772;
assign addr[37946]= 2124624598;
assign addr[37947]= 2141478848;
assign addr[37948]= 2147470025;
assign addr[37949]= 2142567738;
assign addr[37950]= 2126796855;
assign addr[37951]= 2100237377;
assign addr[37952]= 2063024031;
assign addr[37953]= 2015345591;
assign addr[37954]= 1957443913;
assign addr[37955]= 1889612716;
assign addr[37956]= 1812196087;
assign addr[37957]= 1725586737;
assign addr[37958]= 1630224009;
assign addr[37959]= 1526591649;
assign addr[37960]= 1415215352;
assign addr[37961]= 1296660098;
assign addr[37962]= 1171527280;
assign addr[37963]= 1040451659;
assign addr[37964]= 904098143;
assign addr[37965]= 763158411;
assign addr[37966]= 618347408;
assign addr[37967]= 470399716;
assign addr[37968]= 320065829;
assign addr[37969]= 168108346;
assign addr[37970]= 15298099;
assign addr[37971]= -137589750;
assign addr[37972]= -289779648;
assign addr[37973]= -440499581;
assign addr[37974]= -588984994;
assign addr[37975]= -734482665;
assign addr[37976]= -876254528;
assign addr[37977]= -1013581418;
assign addr[37978]= -1145766716;
assign addr[37979]= -1272139887;
assign addr[37980]= -1392059879;
assign addr[37981]= -1504918373;
assign addr[37982]= -1610142873;
assign addr[37983]= -1707199606;
assign addr[37984]= -1795596234;
assign addr[37985]= -1874884346;
assign addr[37986]= -1944661739;
assign addr[37987]= -2004574453;
assign addr[37988]= -2054318569;
assign addr[37989]= -2093641749;
assign addr[37990]= -2122344521;
assign addr[37991]= -2140281282;
assign addr[37992]= -2147361045;
assign addr[37993]= -2143547897;
assign addr[37994]= -2128861181;
assign addr[37995]= -2103375398;
assign addr[37996]= -2067219829;
assign addr[37997]= -2020577882;
assign addr[37998]= -1963686155;
assign addr[37999]= -1896833245;
assign addr[38000]= -1820358275;
assign addr[38001]= -1734649179;
assign addr[38002]= -1640140734;
assign addr[38003]= -1537312353;
assign addr[38004]= -1426685652;
assign addr[38005]= -1308821808;
assign addr[38006]= -1184318708;
assign addr[38007]= -1053807919;
assign addr[38008]= -917951481;
assign addr[38009]= -777438554;
assign addr[38010]= -632981917;
assign addr[38011]= -485314355;
assign addr[38012]= -335184940;
assign addr[38013]= -183355234;
assign addr[38014]= -30595422;
assign addr[38015]= 122319591;
assign addr[38016]= 274614114;
assign addr[38017]= 425515602;
assign addr[38018]= 574258580;
assign addr[38019]= 720088517;
assign addr[38020]= 862265664;
assign addr[38021]= 1000068799;
assign addr[38022]= 1132798888;
assign addr[38023]= 1259782632;
assign addr[38024]= 1380375881;
assign addr[38025]= 1493966902;
assign addr[38026]= 1599979481;
assign addr[38027]= 1697875851;
assign addr[38028]= 1787159411;
assign addr[38029]= 1867377253;
assign addr[38030]= 1938122457;
assign addr[38031]= 1999036154;
assign addr[38032]= 2049809346;
assign addr[38033]= 2090184478;
assign addr[38034]= 2119956737;
assign addr[38035]= 2138975100;
assign addr[38036]= 2147143090;
assign addr[38037]= 2144419275;
assign addr[38038]= 2130817471;
assign addr[38039]= 2106406677;
assign addr[38040]= 2071310720;
assign addr[38041]= 2025707632;
assign addr[38042]= 1969828744;
assign addr[38043]= 1903957513;
assign addr[38044]= 1828428082;
assign addr[38045]= 1743623590;
assign addr[38046]= 1649974225;
assign addr[38047]= 1547955041;
assign addr[38048]= 1438083551;
assign addr[38049]= 1320917099;
assign addr[38050]= 1197050035;
assign addr[38051]= 1067110699;
assign addr[38052]= 931758235;
assign addr[38053]= 791679244;
assign addr[38054]= 647584304;
assign addr[38055]= 500204365;
assign addr[38056]= 350287041;
assign addr[38057]= 198592817;
assign addr[38058]= 45891193;
assign addr[38059]= -107043224;
assign addr[38060]= -259434643;
assign addr[38061]= -410510029;
assign addr[38062]= -559503022;
assign addr[38063]= -705657826;
assign addr[38064]= -848233042;
assign addr[38065]= -986505429;
assign addr[38066]= -1119773573;
assign addr[38067]= -1247361445;
assign addr[38068]= -1368621831;
assign addr[38069]= -1482939614;
assign addr[38070]= -1589734894;
assign addr[38071]= -1688465931;
assign addr[38072]= -1778631892;
assign addr[38073]= -1859775393;
assign addr[38074]= -1931484818;
assign addr[38075]= -1993396407;
assign addr[38076]= -2045196100;
assign addr[38077]= -2086621133;
assign addr[38078]= -2117461370;
assign addr[38079]= -2137560369;
assign addr[38080]= -2146816171;
assign addr[38081]= -2145181827;
assign addr[38082]= -2132665626;
assign addr[38083]= -2109331059;
assign addr[38084]= -2075296495;
assign addr[38085]= -2030734582;
assign addr[38086]= -1975871368;
assign addr[38087]= -1910985158;
assign addr[38088]= -1836405100;
assign addr[38089]= -1752509516;
assign addr[38090]= -1659723983;
assign addr[38091]= -1558519173;
assign addr[38092]= -1449408469;
assign addr[38093]= -1332945355;
assign addr[38094]= -1209720613;
assign addr[38095]= -1080359326;
assign addr[38096]= -945517704;
assign addr[38097]= -805879757;
assign addr[38098]= -662153826;
assign addr[38099]= -515068990;
assign addr[38100]= -365371365;
assign addr[38101]= -213820322;
assign addr[38102]= -61184634;
assign addr[38103]= 91761426;
assign addr[38104]= 244242007;
assign addr[38105]= 395483624;
assign addr[38106]= 544719071;
assign addr[38107]= 691191324;
assign addr[38108]= 834157373;
assign addr[38109]= 972891995;
assign addr[38110]= 1106691431;
assign addr[38111]= 1234876957;
assign addr[38112]= 1356798326;
assign addr[38113]= 1471837070;
assign addr[38114]= 1579409630;
assign addr[38115]= 1678970324;
assign addr[38116]= 1770014111;
assign addr[38117]= 1852079154;
assign addr[38118]= 1924749160;
assign addr[38119]= 1987655498;
assign addr[38120]= 2040479063;
assign addr[38121]= 2082951896;
assign addr[38122]= 2114858546;
assign addr[38123]= 2136037160;
assign addr[38124]= 2146380306;
assign addr[38125]= 2145835515;
assign addr[38126]= 2134405552;
assign addr[38127]= 2112148396;
assign addr[38128]= 2079176953;
assign addr[38129]= 2035658475;
assign addr[38130]= 1981813720;
assign addr[38131]= 1917915825;
assign addr[38132]= 1844288924;
assign addr[38133]= 1761306505;
assign addr[38134]= 1669389513;
assign addr[38135]= 1569004214;
assign addr[38136]= 1460659832;
assign addr[38137]= 1344905966;
assign addr[38138]= 1222329801;
assign addr[38139]= 1093553126;
assign addr[38140]= 959229189;
assign addr[38141]= 820039373;
assign addr[38142]= 676689746;
assign addr[38143]= 529907477;
assign addr[38144]= 380437148;
assign addr[38145]= 229036977;
assign addr[38146]= 76474970;
assign addr[38147]= -76474970;
assign addr[38148]= -229036977;
assign addr[38149]= -380437148;
assign addr[38150]= -529907477;
assign addr[38151]= -676689746;
assign addr[38152]= -820039373;
assign addr[38153]= -959229189;
assign addr[38154]= -1093553126;
assign addr[38155]= -1222329801;
assign addr[38156]= -1344905966;
assign addr[38157]= -1460659832;
assign addr[38158]= -1569004214;
assign addr[38159]= -1669389513;
assign addr[38160]= -1761306505;
assign addr[38161]= -1844288924;
assign addr[38162]= -1917915825;
assign addr[38163]= -1981813720;
assign addr[38164]= -2035658475;
assign addr[38165]= -2079176953;
assign addr[38166]= -2112148396;
assign addr[38167]= -2134405552;
assign addr[38168]= -2145835515;
assign addr[38169]= -2146380306;
assign addr[38170]= -2136037160;
assign addr[38171]= -2114858546;
assign addr[38172]= -2082951896;
assign addr[38173]= -2040479063;
assign addr[38174]= -1987655498;
assign addr[38175]= -1924749160;
assign addr[38176]= -1852079154;
assign addr[38177]= -1770014111;
assign addr[38178]= -1678970324;
assign addr[38179]= -1579409630;
assign addr[38180]= -1471837070;
assign addr[38181]= -1356798326;
assign addr[38182]= -1234876957;
assign addr[38183]= -1106691431;
assign addr[38184]= -972891995;
assign addr[38185]= -834157373;
assign addr[38186]= -691191324;
assign addr[38187]= -544719071;
assign addr[38188]= -395483624;
assign addr[38189]= -244242007;
assign addr[38190]= -91761426;
assign addr[38191]= 61184634;
assign addr[38192]= 213820322;
assign addr[38193]= 365371365;
assign addr[38194]= 515068990;
assign addr[38195]= 662153826;
assign addr[38196]= 805879757;
assign addr[38197]= 945517704;
assign addr[38198]= 1080359326;
assign addr[38199]= 1209720613;
assign addr[38200]= 1332945355;
assign addr[38201]= 1449408469;
assign addr[38202]= 1558519173;
assign addr[38203]= 1659723983;
assign addr[38204]= 1752509516;
assign addr[38205]= 1836405100;
assign addr[38206]= 1910985158;
assign addr[38207]= 1975871368;
assign addr[38208]= 2030734582;
assign addr[38209]= 2075296495;
assign addr[38210]= 2109331059;
assign addr[38211]= 2132665626;
assign addr[38212]= 2145181827;
assign addr[38213]= 2146816171;
assign addr[38214]= 2137560369;
assign addr[38215]= 2117461370;
assign addr[38216]= 2086621133;
assign addr[38217]= 2045196100;
assign addr[38218]= 1993396407;
assign addr[38219]= 1931484818;
assign addr[38220]= 1859775393;
assign addr[38221]= 1778631892;
assign addr[38222]= 1688465931;
assign addr[38223]= 1589734894;
assign addr[38224]= 1482939614;
assign addr[38225]= 1368621831;
assign addr[38226]= 1247361445;
assign addr[38227]= 1119773573;
assign addr[38228]= 986505429;
assign addr[38229]= 848233042;
assign addr[38230]= 705657826;
assign addr[38231]= 559503022;
assign addr[38232]= 410510029;
assign addr[38233]= 259434643;
assign addr[38234]= 107043224;
assign addr[38235]= -45891193;
assign addr[38236]= -198592817;
assign addr[38237]= -350287041;
assign addr[38238]= -500204365;
assign addr[38239]= -647584304;
assign addr[38240]= -791679244;
assign addr[38241]= -931758235;
assign addr[38242]= -1067110699;
assign addr[38243]= -1197050035;
assign addr[38244]= -1320917099;
assign addr[38245]= -1438083551;
assign addr[38246]= -1547955041;
assign addr[38247]= -1649974225;
assign addr[38248]= -1743623590;
assign addr[38249]= -1828428082;
assign addr[38250]= -1903957513;
assign addr[38251]= -1969828744;
assign addr[38252]= -2025707632;
assign addr[38253]= -2071310720;
assign addr[38254]= -2106406677;
assign addr[38255]= -2130817471;
assign addr[38256]= -2144419275;
assign addr[38257]= -2147143090;
assign addr[38258]= -2138975100;
assign addr[38259]= -2119956737;
assign addr[38260]= -2090184478;
assign addr[38261]= -2049809346;
assign addr[38262]= -1999036154;
assign addr[38263]= -1938122457;
assign addr[38264]= -1867377253;
assign addr[38265]= -1787159411;
assign addr[38266]= -1697875851;
assign addr[38267]= -1599979481;
assign addr[38268]= -1493966902;
assign addr[38269]= -1380375881;
assign addr[38270]= -1259782632;
assign addr[38271]= -1132798888;
assign addr[38272]= -1000068799;
assign addr[38273]= -862265664;
assign addr[38274]= -720088517;
assign addr[38275]= -574258580;
assign addr[38276]= -425515602;
assign addr[38277]= -274614114;
assign addr[38278]= -122319591;
assign addr[38279]= 30595422;
assign addr[38280]= 183355234;
assign addr[38281]= 335184940;
assign addr[38282]= 485314355;
assign addr[38283]= 632981917;
assign addr[38284]= 777438554;
assign addr[38285]= 917951481;
assign addr[38286]= 1053807919;
assign addr[38287]= 1184318708;
assign addr[38288]= 1308821808;
assign addr[38289]= 1426685652;
assign addr[38290]= 1537312353;
assign addr[38291]= 1640140734;
assign addr[38292]= 1734649179;
assign addr[38293]= 1820358275;
assign addr[38294]= 1896833245;
assign addr[38295]= 1963686155;
assign addr[38296]= 2020577882;
assign addr[38297]= 2067219829;
assign addr[38298]= 2103375398;
assign addr[38299]= 2128861181;
assign addr[38300]= 2143547897;
assign addr[38301]= 2147361045;
assign addr[38302]= 2140281282;
assign addr[38303]= 2122344521;
assign addr[38304]= 2093641749;
assign addr[38305]= 2054318569;
assign addr[38306]= 2004574453;
assign addr[38307]= 1944661739;
assign addr[38308]= 1874884346;
assign addr[38309]= 1795596234;
assign addr[38310]= 1707199606;
assign addr[38311]= 1610142873;
assign addr[38312]= 1504918373;
assign addr[38313]= 1392059879;
assign addr[38314]= 1272139887;
assign addr[38315]= 1145766716;
assign addr[38316]= 1013581418;
assign addr[38317]= 876254528;
assign addr[38318]= 734482665;
assign addr[38319]= 588984994;
assign addr[38320]= 440499581;
assign addr[38321]= 289779648;
assign addr[38322]= 137589750;
assign addr[38323]= -15298099;
assign addr[38324]= -168108346;
assign addr[38325]= -320065829;
assign addr[38326]= -470399716;
assign addr[38327]= -618347408;
assign addr[38328]= -763158411;
assign addr[38329]= -904098143;
assign addr[38330]= -1040451659;
assign addr[38331]= -1171527280;
assign addr[38332]= -1296660098;
assign addr[38333]= -1415215352;
assign addr[38334]= -1526591649;
assign addr[38335]= -1630224009;
assign addr[38336]= -1725586737;
assign addr[38337]= -1812196087;
assign addr[38338]= -1889612716;
assign addr[38339]= -1957443913;
assign addr[38340]= -2015345591;
assign addr[38341]= -2063024031;
assign addr[38342]= -2100237377;
assign addr[38343]= -2126796855;
assign addr[38344]= -2142567738;
assign addr[38345]= -2147470025;
assign addr[38346]= -2141478848;
assign addr[38347]= -2124624598;
assign addr[38348]= -2096992772;
assign addr[38349]= -2058723538;
assign addr[38350]= -2010011024;
assign addr[38351]= -1951102334;
assign addr[38352]= -1882296293;
assign addr[38353]= -1803941934;
assign addr[38354]= -1716436725;
assign addr[38355]= -1620224553;
assign addr[38356]= -1515793473;
assign addr[38357]= -1403673233;
assign addr[38358]= -1284432584;
assign addr[38359]= -1158676398;
assign addr[38360]= -1027042599;
assign addr[38361]= -890198924;
assign addr[38362]= -748839539;
assign addr[38363]= -603681519;
assign addr[38364]= -455461206;
assign addr[38365]= -304930476;
assign addr[38366]= -152852926;
assign addr[38367]= 0;
assign addr[38368]= 152852926;
assign addr[38369]= 304930476;
assign addr[38370]= 455461206;
assign addr[38371]= 603681519;
assign addr[38372]= 748839539;
assign addr[38373]= 890198924;
assign addr[38374]= 1027042599;
assign addr[38375]= 1158676398;
assign addr[38376]= 1284432584;
assign addr[38377]= 1403673233;
assign addr[38378]= 1515793473;
assign addr[38379]= 1620224553;
assign addr[38380]= 1716436725;
assign addr[38381]= 1803941934;
assign addr[38382]= 1882296293;
assign addr[38383]= 1951102334;
assign addr[38384]= 2010011024;
assign addr[38385]= 2058723538;
assign addr[38386]= 2096992772;
assign addr[38387]= 2124624598;
assign addr[38388]= 2141478848;
assign addr[38389]= 2147470025;
assign addr[38390]= 2142567738;
assign addr[38391]= 2126796855;
assign addr[38392]= 2100237377;
assign addr[38393]= 2063024031;
assign addr[38394]= 2015345591;
assign addr[38395]= 1957443913;
assign addr[38396]= 1889612716;
assign addr[38397]= 1812196087;
assign addr[38398]= 1725586737;
assign addr[38399]= 1630224009;
assign addr[38400]= 1526591649;
assign addr[38401]= 1415215352;
assign addr[38402]= 1296660098;
assign addr[38403]= 1171527280;
assign addr[38404]= 1040451659;
assign addr[38405]= 904098143;
assign addr[38406]= 763158411;
assign addr[38407]= 618347408;
assign addr[38408]= 470399716;
assign addr[38409]= 320065829;
assign addr[38410]= 168108346;
assign addr[38411]= 15298099;
assign addr[38412]= -137589750;
assign addr[38413]= -289779648;
assign addr[38414]= -440499581;
assign addr[38415]= -588984994;
assign addr[38416]= -734482665;
assign addr[38417]= -876254528;
assign addr[38418]= -1013581418;
assign addr[38419]= -1145766716;
assign addr[38420]= -1272139887;
assign addr[38421]= -1392059879;
assign addr[38422]= -1504918373;
assign addr[38423]= -1610142873;
assign addr[38424]= -1707199606;
assign addr[38425]= -1795596234;
assign addr[38426]= -1874884346;
assign addr[38427]= -1944661739;
assign addr[38428]= -2004574453;
assign addr[38429]= -2054318569;
assign addr[38430]= -2093641749;
assign addr[38431]= -2122344521;
assign addr[38432]= -2140281282;
assign addr[38433]= -2147361045;
assign addr[38434]= -2143547897;
assign addr[38435]= -2128861181;
assign addr[38436]= -2103375398;
assign addr[38437]= -2067219829;
assign addr[38438]= -2020577882;
assign addr[38439]= -1963686155;
assign addr[38440]= -1896833245;
assign addr[38441]= -1820358275;
assign addr[38442]= -1734649179;
assign addr[38443]= -1640140734;
assign addr[38444]= -1537312353;
assign addr[38445]= -1426685652;
assign addr[38446]= -1308821808;
assign addr[38447]= -1184318708;
assign addr[38448]= -1053807919;
assign addr[38449]= -917951481;
assign addr[38450]= -777438554;
assign addr[38451]= -632981917;
assign addr[38452]= -485314355;
assign addr[38453]= -335184940;
assign addr[38454]= -183355234;
assign addr[38455]= -30595422;
assign addr[38456]= 122319591;
assign addr[38457]= 274614114;
assign addr[38458]= 425515602;
assign addr[38459]= 574258580;
assign addr[38460]= 720088517;
assign addr[38461]= 862265664;
assign addr[38462]= 1000068799;
assign addr[38463]= 1132798888;
assign addr[38464]= 1259782632;
assign addr[38465]= 1380375881;
assign addr[38466]= 1493966902;
assign addr[38467]= 1599979481;
assign addr[38468]= 1697875851;
assign addr[38469]= 1787159411;
assign addr[38470]= 1867377253;
assign addr[38471]= 1938122457;
assign addr[38472]= 1999036154;
assign addr[38473]= 2049809346;
assign addr[38474]= 2090184478;
assign addr[38475]= 2119956737;
assign addr[38476]= 2138975100;
assign addr[38477]= 2147143090;
assign addr[38478]= 2144419275;
assign addr[38479]= 2130817471;
assign addr[38480]= 2106406677;
assign addr[38481]= 2071310720;
assign addr[38482]= 2025707632;
assign addr[38483]= 1969828744;
assign addr[38484]= 1903957513;
assign addr[38485]= 1828428082;
assign addr[38486]= 1743623590;
assign addr[38487]= 1649974225;
assign addr[38488]= 1547955041;
assign addr[38489]= 1438083551;
assign addr[38490]= 1320917099;
assign addr[38491]= 1197050035;
assign addr[38492]= 1067110699;
assign addr[38493]= 931758235;
assign addr[38494]= 791679244;
assign addr[38495]= 647584304;
assign addr[38496]= 500204365;
assign addr[38497]= 350287041;
assign addr[38498]= 198592817;
assign addr[38499]= 45891193;
assign addr[38500]= -107043224;
assign addr[38501]= -259434643;
assign addr[38502]= -410510029;
assign addr[38503]= -559503022;
assign addr[38504]= -705657826;
assign addr[38505]= -848233042;
assign addr[38506]= -986505429;
assign addr[38507]= -1119773573;
assign addr[38508]= -1247361445;
assign addr[38509]= -1368621831;
assign addr[38510]= -1482939614;
assign addr[38511]= -1589734894;
assign addr[38512]= -1688465931;
assign addr[38513]= -1778631892;
assign addr[38514]= -1859775393;
assign addr[38515]= -1931484818;
assign addr[38516]= -1993396407;
assign addr[38517]= -2045196100;
assign addr[38518]= -2086621133;
assign addr[38519]= -2117461370;
assign addr[38520]= -2137560369;
assign addr[38521]= -2146816171;
assign addr[38522]= -2145181827;
assign addr[38523]= -2132665626;
assign addr[38524]= -2109331059;
assign addr[38525]= -2075296495;
assign addr[38526]= -2030734582;
assign addr[38527]= -1975871368;
assign addr[38528]= -1910985158;
assign addr[38529]= -1836405100;
assign addr[38530]= -1752509516;
assign addr[38531]= -1659723983;
assign addr[38532]= -1558519173;
assign addr[38533]= -1449408469;
assign addr[38534]= -1332945355;
assign addr[38535]= -1209720613;
assign addr[38536]= -1080359326;
assign addr[38537]= -945517704;
assign addr[38538]= -805879757;
assign addr[38539]= -662153826;
assign addr[38540]= -515068990;
assign addr[38541]= -365371365;
assign addr[38542]= -213820322;
assign addr[38543]= -61184634;
assign addr[38544]= 91761426;
assign addr[38545]= 244242007;
assign addr[38546]= 395483624;
assign addr[38547]= 544719071;
assign addr[38548]= 691191324;
assign addr[38549]= 834157373;
assign addr[38550]= 972891995;
assign addr[38551]= 1106691431;
assign addr[38552]= 1234876957;
assign addr[38553]= 1356798326;
assign addr[38554]= 1471837070;
assign addr[38555]= 1579409630;
assign addr[38556]= 1678970324;
assign addr[38557]= 1770014111;
assign addr[38558]= 1852079154;
assign addr[38559]= 1924749160;
assign addr[38560]= 1987655498;
assign addr[38561]= 2040479063;
assign addr[38562]= 2082951896;
assign addr[38563]= 2114858546;
assign addr[38564]= 2136037160;
assign addr[38565]= 2146380306;
assign addr[38566]= 2145835515;
assign addr[38567]= 2134405552;
assign addr[38568]= 2112148396;
assign addr[38569]= 2079176953;
assign addr[38570]= 2035658475;
assign addr[38571]= 1981813720;
assign addr[38572]= 1917915825;
assign addr[38573]= 1844288924;
assign addr[38574]= 1761306505;
assign addr[38575]= 1669389513;
assign addr[38576]= 1569004214;
assign addr[38577]= 1460659832;
assign addr[38578]= 1344905966;
assign addr[38579]= 1222329801;
assign addr[38580]= 1093553126;
assign addr[38581]= 959229189;
assign addr[38582]= 820039373;
assign addr[38583]= 676689746;
assign addr[38584]= 529907477;
assign addr[38585]= 380437148;
assign addr[38586]= 229036977;
assign addr[38587]= 76474970;
assign addr[38588]= -76474970;
assign addr[38589]= -229036977;
assign addr[38590]= -380437148;
assign addr[38591]= -529907477;
assign addr[38592]= -676689746;
assign addr[38593]= -820039373;
assign addr[38594]= -959229189;
assign addr[38595]= -1093553126;
assign addr[38596]= -1222329801;
assign addr[38597]= -1344905966;
assign addr[38598]= -1460659832;
assign addr[38599]= -1569004214;
assign addr[38600]= -1669389513;
assign addr[38601]= -1761306505;
assign addr[38602]= -1844288924;
assign addr[38603]= -1917915825;
assign addr[38604]= -1981813720;
assign addr[38605]= -2035658475;
assign addr[38606]= -2079176953;
assign addr[38607]= -2112148396;
assign addr[38608]= -2134405552;
assign addr[38609]= -2145835515;
assign addr[38610]= -2146380306;
assign addr[38611]= -2136037160;
assign addr[38612]= -2114858546;
assign addr[38613]= -2082951896;
assign addr[38614]= -2040479063;
assign addr[38615]= -1987655498;
assign addr[38616]= -1924749160;
assign addr[38617]= -1852079154;
assign addr[38618]= -1770014111;
assign addr[38619]= -1678970324;
assign addr[38620]= -1579409630;
assign addr[38621]= -1471837070;
assign addr[38622]= -1356798326;
assign addr[38623]= -1234876957;
assign addr[38624]= -1106691431;
assign addr[38625]= -972891995;
assign addr[38626]= -834157373;
assign addr[38627]= -691191324;
assign addr[38628]= -544719071;
assign addr[38629]= -395483624;
assign addr[38630]= -244242007;
assign addr[38631]= -91761426;
assign addr[38632]= 61184634;
assign addr[38633]= 213820322;
assign addr[38634]= 365371365;
assign addr[38635]= 515068990;
assign addr[38636]= 662153826;
assign addr[38637]= 805879757;
assign addr[38638]= 945517704;
assign addr[38639]= 1080359326;
assign addr[38640]= 1209720613;
assign addr[38641]= 1332945355;
assign addr[38642]= 1449408469;
assign addr[38643]= 1558519173;
assign addr[38644]= 1659723983;
assign addr[38645]= 1752509516;
assign addr[38646]= 1836405100;
assign addr[38647]= 1910985158;
assign addr[38648]= 1975871368;
assign addr[38649]= 2030734582;
assign addr[38650]= 2075296495;
assign addr[38651]= 2109331059;
assign addr[38652]= 2132665626;
assign addr[38653]= 2145181827;
assign addr[38654]= 2146816171;
assign addr[38655]= 2137560369;
assign addr[38656]= 2117461370;
assign addr[38657]= 2086621133;
assign addr[38658]= 2045196100;
assign addr[38659]= 1993396407;
assign addr[38660]= 1931484818;
assign addr[38661]= 1859775393;
assign addr[38662]= 1778631892;
assign addr[38663]= 1688465931;
assign addr[38664]= 1589734894;
assign addr[38665]= 1482939614;
assign addr[38666]= 1368621831;
assign addr[38667]= 1247361445;
assign addr[38668]= 1119773573;
assign addr[38669]= 986505429;
assign addr[38670]= 848233042;
assign addr[38671]= 705657826;
assign addr[38672]= 559503022;
assign addr[38673]= 410510029;
assign addr[38674]= 259434643;
assign addr[38675]= 107043224;
assign addr[38676]= -45891193;
assign addr[38677]= -198592817;
assign addr[38678]= -350287041;
assign addr[38679]= -500204365;
assign addr[38680]= -647584304;
assign addr[38681]= -791679244;
assign addr[38682]= -931758235;
assign addr[38683]= -1067110699;
assign addr[38684]= -1197050035;
assign addr[38685]= -1320917099;
assign addr[38686]= -1438083551;
assign addr[38687]= -1547955041;
assign addr[38688]= -1649974225;
assign addr[38689]= -1743623590;
assign addr[38690]= -1828428082;
assign addr[38691]= -1903957513;
assign addr[38692]= -1969828744;
assign addr[38693]= -2025707632;
assign addr[38694]= -2071310720;
assign addr[38695]= -2106406677;
assign addr[38696]= -2130817471;
assign addr[38697]= -2144419275;
assign addr[38698]= -2147143090;
assign addr[38699]= -2138975100;
assign addr[38700]= -2119956737;
assign addr[38701]= -2090184478;
assign addr[38702]= -2049809346;
assign addr[38703]= -1999036154;
assign addr[38704]= -1938122457;
assign addr[38705]= -1867377253;
assign addr[38706]= -1787159411;
assign addr[38707]= -1697875851;
assign addr[38708]= -1599979481;
assign addr[38709]= -1493966902;
assign addr[38710]= -1380375881;
assign addr[38711]= -1259782632;
assign addr[38712]= -1132798888;
assign addr[38713]= -1000068799;
assign addr[38714]= -862265664;
assign addr[38715]= -720088517;
assign addr[38716]= -574258580;
assign addr[38717]= -425515602;
assign addr[38718]= -274614114;
assign addr[38719]= -122319591;
assign addr[38720]= 30595422;
assign addr[38721]= 183355234;
assign addr[38722]= 335184940;
assign addr[38723]= 485314355;
assign addr[38724]= 632981917;
assign addr[38725]= 777438554;
assign addr[38726]= 917951481;
assign addr[38727]= 1053807919;
assign addr[38728]= 1184318708;
assign addr[38729]= 1308821808;
assign addr[38730]= 1426685652;
assign addr[38731]= 1537312353;
assign addr[38732]= 1640140734;
assign addr[38733]= 1734649179;
assign addr[38734]= 1820358275;
assign addr[38735]= 1896833245;
assign addr[38736]= 1963686155;
assign addr[38737]= 2020577882;
assign addr[38738]= 2067219829;
assign addr[38739]= 2103375398;
assign addr[38740]= 2128861181;
assign addr[38741]= 2143547897;
assign addr[38742]= 2147361045;
assign addr[38743]= 2140281282;
assign addr[38744]= 2122344521;
assign addr[38745]= 2093641749;
assign addr[38746]= 2054318569;
assign addr[38747]= 2004574453;
assign addr[38748]= 1944661739;
assign addr[38749]= 1874884346;
assign addr[38750]= 1795596234;
assign addr[38751]= 1707199606;
assign addr[38752]= 1610142873;
assign addr[38753]= 1504918373;
assign addr[38754]= 1392059879;
assign addr[38755]= 1272139887;
assign addr[38756]= 1145766716;
assign addr[38757]= 1013581418;
assign addr[38758]= 876254528;
assign addr[38759]= 734482665;
assign addr[38760]= 588984994;
assign addr[38761]= 440499581;
assign addr[38762]= 289779648;
assign addr[38763]= 137589750;
assign addr[38764]= -15298099;
assign addr[38765]= -168108346;
assign addr[38766]= -320065829;
assign addr[38767]= -470399716;
assign addr[38768]= -618347408;
assign addr[38769]= -763158411;
assign addr[38770]= -904098143;
assign addr[38771]= -1040451659;
assign addr[38772]= -1171527280;
assign addr[38773]= -1296660098;
assign addr[38774]= -1415215352;
assign addr[38775]= -1526591649;
assign addr[38776]= -1630224009;
assign addr[38777]= -1725586737;
assign addr[38778]= -1812196087;
assign addr[38779]= -1889612716;
assign addr[38780]= -1957443913;
assign addr[38781]= -2015345591;
assign addr[38782]= -2063024031;
assign addr[38783]= -2100237377;
assign addr[38784]= -2126796855;
assign addr[38785]= -2142567738;
assign addr[38786]= -2147470025;
assign addr[38787]= -2141478848;
assign addr[38788]= -2124624598;
assign addr[38789]= -2096992772;
assign addr[38790]= -2058723538;
assign addr[38791]= -2010011024;
assign addr[38792]= -1951102334;
assign addr[38793]= -1882296293;
assign addr[38794]= -1803941934;
assign addr[38795]= -1716436725;
assign addr[38796]= -1620224553;
assign addr[38797]= -1515793473;
assign addr[38798]= -1403673233;
assign addr[38799]= -1284432584;
assign addr[38800]= -1158676398;
assign addr[38801]= -1027042599;
assign addr[38802]= -890198924;
assign addr[38803]= -748839539;
assign addr[38804]= -603681519;
assign addr[38805]= -455461206;
assign addr[38806]= -304930476;
assign addr[38807]= -152852926;
assign addr[38808]= 0;
assign addr[38809]= 152852926;
assign addr[38810]= 304930476;
assign addr[38811]= 455461206;
assign addr[38812]= 603681519;
assign addr[38813]= 748839539;
assign addr[38814]= 890198924;
assign addr[38815]= 1027042599;
assign addr[38816]= 1158676398;
assign addr[38817]= 1284432584;
assign addr[38818]= 1403673233;
assign addr[38819]= 1515793473;
assign addr[38820]= 1620224553;
assign addr[38821]= 1716436725;
assign addr[38822]= 1803941934;
assign addr[38823]= 1882296293;
assign addr[38824]= 1951102334;
assign addr[38825]= 2010011024;
assign addr[38826]= 2058723538;
assign addr[38827]= 2096992772;
assign addr[38828]= 2124624598;
assign addr[38829]= 2141478848;
assign addr[38830]= 2147470025;
assign addr[38831]= 2142567738;
assign addr[38832]= 2126796855;
assign addr[38833]= 2100237377;
assign addr[38834]= 2063024031;
assign addr[38835]= 2015345591;
assign addr[38836]= 1957443913;
assign addr[38837]= 1889612716;
assign addr[38838]= 1812196087;
assign addr[38839]= 1725586737;
assign addr[38840]= 1630224009;
assign addr[38841]= 1526591649;
assign addr[38842]= 1415215352;
assign addr[38843]= 1296660098;
assign addr[38844]= 1171527280;
assign addr[38845]= 1040451659;
assign addr[38846]= 904098143;
assign addr[38847]= 763158411;
assign addr[38848]= 618347408;
assign addr[38849]= 470399716;
assign addr[38850]= 320065829;
assign addr[38851]= 168108346;
assign addr[38852]= 15298099;
assign addr[38853]= -137589750;
assign addr[38854]= -289779648;
assign addr[38855]= -440499581;
assign addr[38856]= -588984994;
assign addr[38857]= -734482665;
assign addr[38858]= -876254528;
assign addr[38859]= -1013581418;
assign addr[38860]= -1145766716;
assign addr[38861]= -1272139887;
assign addr[38862]= -1392059879;
assign addr[38863]= -1504918373;
assign addr[38864]= -1610142873;
assign addr[38865]= -1707199606;
assign addr[38866]= -1795596234;
assign addr[38867]= -1874884346;
assign addr[38868]= -1944661739;
assign addr[38869]= -2004574453;
assign addr[38870]= -2054318569;
assign addr[38871]= -2093641749;
assign addr[38872]= -2122344521;
assign addr[38873]= -2140281282;
assign addr[38874]= -2147361045;
assign addr[38875]= -2143547897;
assign addr[38876]= -2128861181;
assign addr[38877]= -2103375398;
assign addr[38878]= -2067219829;
assign addr[38879]= -2020577882;
assign addr[38880]= -1963686155;
assign addr[38881]= -1896833245;
assign addr[38882]= -1820358275;
assign addr[38883]= -1734649179;
assign addr[38884]= -1640140734;
assign addr[38885]= -1537312353;
assign addr[38886]= -1426685652;
assign addr[38887]= -1308821808;
assign addr[38888]= -1184318708;
assign addr[38889]= -1053807919;
assign addr[38890]= -917951481;
assign addr[38891]= -777438554;
assign addr[38892]= -632981917;
assign addr[38893]= -485314355;
assign addr[38894]= -335184940;
assign addr[38895]= -183355234;
assign addr[38896]= -30595422;
assign addr[38897]= 122319591;
assign addr[38898]= 274614114;
assign addr[38899]= 425515602;
assign addr[38900]= 574258580;
assign addr[38901]= 720088517;
assign addr[38902]= 862265664;
assign addr[38903]= 1000068799;
assign addr[38904]= 1132798888;
assign addr[38905]= 1259782632;
assign addr[38906]= 1380375881;
assign addr[38907]= 1493966902;
assign addr[38908]= 1599979481;
assign addr[38909]= 1697875851;
assign addr[38910]= 1787159411;
assign addr[38911]= 1867377253;
assign addr[38912]= 1938122457;
assign addr[38913]= 1999036154;
assign addr[38914]= 2049809346;
assign addr[38915]= 2090184478;
assign addr[38916]= 2119956737;
assign addr[38917]= 2138975100;
assign addr[38918]= 2147143090;
assign addr[38919]= 2144419275;
assign addr[38920]= 2130817471;
assign addr[38921]= 2106406677;
assign addr[38922]= 2071310720;
assign addr[38923]= 2025707632;
assign addr[38924]= 1969828744;
assign addr[38925]= 1903957513;
assign addr[38926]= 1828428082;
assign addr[38927]= 1743623590;
assign addr[38928]= 1649974225;
assign addr[38929]= 1547955041;
assign addr[38930]= 1438083551;
assign addr[38931]= 1320917099;
assign addr[38932]= 1197050035;
assign addr[38933]= 1067110699;
assign addr[38934]= 931758235;
assign addr[38935]= 791679244;
assign addr[38936]= 647584304;
assign addr[38937]= 500204365;
assign addr[38938]= 350287041;
assign addr[38939]= 198592817;
assign addr[38940]= 45891193;
assign addr[38941]= -107043224;
assign addr[38942]= -259434643;
assign addr[38943]= -410510029;
assign addr[38944]= -559503022;
assign addr[38945]= -705657826;
assign addr[38946]= -848233042;
assign addr[38947]= -986505429;
assign addr[38948]= -1119773573;
assign addr[38949]= -1247361445;
assign addr[38950]= -1368621831;
assign addr[38951]= -1482939614;
assign addr[38952]= -1589734894;
assign addr[38953]= -1688465931;
assign addr[38954]= -1778631892;
assign addr[38955]= -1859775393;
assign addr[38956]= -1931484818;
assign addr[38957]= -1993396407;
assign addr[38958]= -2045196100;
assign addr[38959]= -2086621133;
assign addr[38960]= -2117461370;
assign addr[38961]= -2137560369;
assign addr[38962]= -2146816171;
assign addr[38963]= -2145181827;
assign addr[38964]= -2132665626;
assign addr[38965]= -2109331059;
assign addr[38966]= -2075296495;
assign addr[38967]= -2030734582;
assign addr[38968]= -1975871368;
assign addr[38969]= -1910985158;
assign addr[38970]= -1836405100;
assign addr[38971]= -1752509516;
assign addr[38972]= -1659723983;
assign addr[38973]= -1558519173;
assign addr[38974]= -1449408469;
assign addr[38975]= -1332945355;
assign addr[38976]= -1209720613;
assign addr[38977]= -1080359326;
assign addr[38978]= -945517704;
assign addr[38979]= -805879757;
assign addr[38980]= -662153826;
assign addr[38981]= -515068990;
assign addr[38982]= -365371365;
assign addr[38983]= -213820322;
assign addr[38984]= -61184634;
assign addr[38985]= 91761426;
assign addr[38986]= 244242007;
assign addr[38987]= 395483624;
assign addr[38988]= 544719071;
assign addr[38989]= 691191324;
assign addr[38990]= 834157373;
assign addr[38991]= 972891995;
assign addr[38992]= 1106691431;
assign addr[38993]= 1234876957;
assign addr[38994]= 1356798326;
assign addr[38995]= 1471837070;
assign addr[38996]= 1579409630;
assign addr[38997]= 1678970324;
assign addr[38998]= 1770014111;
assign addr[38999]= 1852079154;
assign addr[39000]= 1924749160;
assign addr[39001]= 1987655498;
assign addr[39002]= 2040479063;
assign addr[39003]= 2082951896;
assign addr[39004]= 2114858546;
assign addr[39005]= 2136037160;
assign addr[39006]= 2146380306;
assign addr[39007]= 2145835515;
assign addr[39008]= 2134405552;
assign addr[39009]= 2112148396;
assign addr[39010]= 2079176953;
assign addr[39011]= 2035658475;
assign addr[39012]= 1981813720;
assign addr[39013]= 1917915825;
assign addr[39014]= 1844288924;
assign addr[39015]= 1761306505;
assign addr[39016]= 1669389513;
assign addr[39017]= 1569004214;
assign addr[39018]= 1460659832;
assign addr[39019]= 1344905966;
assign addr[39020]= 1222329801;
assign addr[39021]= 1093553126;
assign addr[39022]= 959229189;
assign addr[39023]= 820039373;
assign addr[39024]= 676689746;
assign addr[39025]= 529907477;
assign addr[39026]= 380437148;
assign addr[39027]= 229036977;
assign addr[39028]= 76474970;
assign addr[39029]= -76474970;
assign addr[39030]= -229036977;
assign addr[39031]= -380437148;
assign addr[39032]= -529907477;
assign addr[39033]= -676689746;
assign addr[39034]= -820039373;
assign addr[39035]= -959229189;
assign addr[39036]= -1093553126;
assign addr[39037]= -1222329801;
assign addr[39038]= -1344905966;
assign addr[39039]= -1460659832;
assign addr[39040]= -1569004214;
assign addr[39041]= -1669389513;
assign addr[39042]= -1761306505;
assign addr[39043]= -1844288924;
assign addr[39044]= -1917915825;
assign addr[39045]= -1981813720;
assign addr[39046]= -2035658475;
assign addr[39047]= -2079176953;
assign addr[39048]= -2112148396;
assign addr[39049]= -2134405552;
assign addr[39050]= -2145835515;
assign addr[39051]= -2146380306;
assign addr[39052]= -2136037160;
assign addr[39053]= -2114858546;
assign addr[39054]= -2082951896;
assign addr[39055]= -2040479063;
assign addr[39056]= -1987655498;
assign addr[39057]= -1924749160;
assign addr[39058]= -1852079154;
assign addr[39059]= -1770014111;
assign addr[39060]= -1678970324;
assign addr[39061]= -1579409630;
assign addr[39062]= -1471837070;
assign addr[39063]= -1356798326;
assign addr[39064]= -1234876957;
assign addr[39065]= -1106691431;
assign addr[39066]= -972891995;
assign addr[39067]= -834157373;
assign addr[39068]= -691191324;
assign addr[39069]= -544719071;
assign addr[39070]= -395483624;
assign addr[39071]= -244242007;
assign addr[39072]= -91761426;
assign addr[39073]= 61184634;
assign addr[39074]= 213820322;
assign addr[39075]= 365371365;
assign addr[39076]= 515068990;
assign addr[39077]= 662153826;
assign addr[39078]= 805879757;
assign addr[39079]= 945517704;
assign addr[39080]= 1080359326;
assign addr[39081]= 1209720613;
assign addr[39082]= 1332945355;
assign addr[39083]= 1449408469;
assign addr[39084]= 1558519173;
assign addr[39085]= 1659723983;
assign addr[39086]= 1752509516;
assign addr[39087]= 1836405100;
assign addr[39088]= 1910985158;
assign addr[39089]= 1975871368;
assign addr[39090]= 2030734582;
assign addr[39091]= 2075296495;
assign addr[39092]= 2109331059;
assign addr[39093]= 2132665626;
assign addr[39094]= 2145181827;
assign addr[39095]= 2146816171;
assign addr[39096]= 2137560369;
assign addr[39097]= 2117461370;
assign addr[39098]= 2086621133;
assign addr[39099]= 2045196100;
assign addr[39100]= 1993396407;
assign addr[39101]= 1931484818;
assign addr[39102]= 1859775393;
assign addr[39103]= 1778631892;
assign addr[39104]= 1688465931;
assign addr[39105]= 1589734894;
assign addr[39106]= 1482939614;
assign addr[39107]= 1368621831;
assign addr[39108]= 1247361445;
assign addr[39109]= 1119773573;
assign addr[39110]= 986505429;
assign addr[39111]= 848233042;
assign addr[39112]= 705657826;
assign addr[39113]= 559503022;
assign addr[39114]= 410510029;
assign addr[39115]= 259434643;
assign addr[39116]= 107043224;
assign addr[39117]= -45891193;
assign addr[39118]= -198592817;
assign addr[39119]= -350287041;
assign addr[39120]= -500204365;
assign addr[39121]= -647584304;
assign addr[39122]= -791679244;
assign addr[39123]= -931758235;
assign addr[39124]= -1067110699;
assign addr[39125]= -1197050035;
assign addr[39126]= -1320917099;
assign addr[39127]= -1438083551;
assign addr[39128]= -1547955041;
assign addr[39129]= -1649974225;
assign addr[39130]= -1743623590;
assign addr[39131]= -1828428082;
assign addr[39132]= -1903957513;
assign addr[39133]= -1969828744;
assign addr[39134]= -2025707632;
assign addr[39135]= -2071310720;
assign addr[39136]= -2106406677;
assign addr[39137]= -2130817471;
assign addr[39138]= -2144419275;
assign addr[39139]= -2147143090;
assign addr[39140]= -2138975100;
assign addr[39141]= -2119956737;
assign addr[39142]= -2090184478;
assign addr[39143]= -2049809346;
assign addr[39144]= -1999036154;
assign addr[39145]= -1938122457;
assign addr[39146]= -1867377253;
assign addr[39147]= -1787159411;
assign addr[39148]= -1697875851;
assign addr[39149]= -1599979481;
assign addr[39150]= -1493966902;
assign addr[39151]= -1380375881;
assign addr[39152]= -1259782632;
assign addr[39153]= -1132798888;
assign addr[39154]= -1000068799;
assign addr[39155]= -862265664;
assign addr[39156]= -720088517;
assign addr[39157]= -574258580;
assign addr[39158]= -425515602;
assign addr[39159]= -274614114;
assign addr[39160]= -122319591;
assign addr[39161]= 30595422;
assign addr[39162]= 183355234;
assign addr[39163]= 335184940;
assign addr[39164]= 485314355;
assign addr[39165]= 632981917;
assign addr[39166]= 777438554;
assign addr[39167]= 917951481;
assign addr[39168]= 1053807919;
assign addr[39169]= 1184318708;
assign addr[39170]= 1308821808;
assign addr[39171]= 1426685652;
assign addr[39172]= 1537312353;
assign addr[39173]= 1640140734;
assign addr[39174]= 1734649179;
assign addr[39175]= 1820358275;
assign addr[39176]= 1896833245;
assign addr[39177]= 1963686155;
assign addr[39178]= 2020577882;
assign addr[39179]= 2067219829;
assign addr[39180]= 2103375398;
assign addr[39181]= 2128861181;
assign addr[39182]= 2143547897;
assign addr[39183]= 2147361045;
assign addr[39184]= 2140281282;
assign addr[39185]= 2122344521;
assign addr[39186]= 2093641749;
assign addr[39187]= 2054318569;
assign addr[39188]= 2004574453;
assign addr[39189]= 1944661739;
assign addr[39190]= 1874884346;
assign addr[39191]= 1795596234;
assign addr[39192]= 1707199606;
assign addr[39193]= 1610142873;
assign addr[39194]= 1504918373;
assign addr[39195]= 1392059879;
assign addr[39196]= 1272139887;
assign addr[39197]= 1145766716;
assign addr[39198]= 1013581418;
assign addr[39199]= 876254528;
assign addr[39200]= 734482665;
assign addr[39201]= 588984994;
assign addr[39202]= 440499581;
assign addr[39203]= 289779648;
assign addr[39204]= 137589750;
assign addr[39205]= -15298099;
assign addr[39206]= -168108346;
assign addr[39207]= -320065829;
assign addr[39208]= -470399716;
assign addr[39209]= -618347408;
assign addr[39210]= -763158411;
assign addr[39211]= -904098143;
assign addr[39212]= -1040451659;
assign addr[39213]= -1171527280;
assign addr[39214]= -1296660098;
assign addr[39215]= -1415215352;
assign addr[39216]= -1526591649;
assign addr[39217]= -1630224009;
assign addr[39218]= -1725586737;
assign addr[39219]= -1812196087;
assign addr[39220]= -1889612716;
assign addr[39221]= -1957443913;
assign addr[39222]= -2015345591;
assign addr[39223]= -2063024031;
assign addr[39224]= -2100237377;
assign addr[39225]= -2126796855;
assign addr[39226]= -2142567738;
assign addr[39227]= -2147470025;
assign addr[39228]= -2141478848;
assign addr[39229]= -2124624598;
assign addr[39230]= -2096992772;
assign addr[39231]= -2058723538;
assign addr[39232]= -2010011024;
assign addr[39233]= -1951102334;
assign addr[39234]= -1882296293;
assign addr[39235]= -1803941934;
assign addr[39236]= -1716436725;
assign addr[39237]= -1620224553;
assign addr[39238]= -1515793473;
assign addr[39239]= -1403673233;
assign addr[39240]= -1284432584;
assign addr[39241]= -1158676398;
assign addr[39242]= -1027042599;
assign addr[39243]= -890198924;
assign addr[39244]= -748839539;
assign addr[39245]= -603681519;
assign addr[39246]= -455461206;
assign addr[39247]= -304930476;
assign addr[39248]= -152852926;
assign addr[39249]= 0;
assign addr[39250]= 152852926;
assign addr[39251]= 304930476;
assign addr[39252]= 455461206;
assign addr[39253]= 603681519;
assign addr[39254]= 748839539;
assign addr[39255]= 890198924;
assign addr[39256]= 1027042599;
assign addr[39257]= 1158676398;
assign addr[39258]= 1284432584;
assign addr[39259]= 1403673233;
assign addr[39260]= 1515793473;
assign addr[39261]= 1620224553;
assign addr[39262]= 1716436725;
assign addr[39263]= 1803941934;
assign addr[39264]= 1882296293;
assign addr[39265]= 1951102334;
assign addr[39266]= 2010011024;
assign addr[39267]= 2058723538;
assign addr[39268]= 2096992772;
assign addr[39269]= 2124624598;
assign addr[39270]= 2141478848;
assign addr[39271]= 2147470025;
assign addr[39272]= 2142567738;
assign addr[39273]= 2126796855;
assign addr[39274]= 2100237377;
assign addr[39275]= 2063024031;
assign addr[39276]= 2015345591;
assign addr[39277]= 1957443913;
assign addr[39278]= 1889612716;
assign addr[39279]= 1812196087;
assign addr[39280]= 1725586737;
assign addr[39281]= 1630224009;
assign addr[39282]= 1526591649;
assign addr[39283]= 1415215352;
assign addr[39284]= 1296660098;
assign addr[39285]= 1171527280;
assign addr[39286]= 1040451659;
assign addr[39287]= 904098143;
assign addr[39288]= 763158411;
assign addr[39289]= 618347408;
assign addr[39290]= 470399716;
assign addr[39291]= 320065829;
assign addr[39292]= 168108346;
assign addr[39293]= 15298099;
assign addr[39294]= -137589750;
assign addr[39295]= -289779648;
assign addr[39296]= -440499581;
assign addr[39297]= -588984994;
assign addr[39298]= -734482665;
assign addr[39299]= -876254528;
assign addr[39300]= -1013581418;
assign addr[39301]= -1145766716;
assign addr[39302]= -1272139887;
assign addr[39303]= -1392059879;
assign addr[39304]= -1504918373;
assign addr[39305]= -1610142873;
assign addr[39306]= -1707199606;
assign addr[39307]= -1795596234;
assign addr[39308]= -1874884346;
assign addr[39309]= -1944661739;
assign addr[39310]= -2004574453;
assign addr[39311]= -2054318569;
assign addr[39312]= -2093641749;
assign addr[39313]= -2122344521;
assign addr[39314]= -2140281282;
assign addr[39315]= -2147361045;
assign addr[39316]= -2143547897;
assign addr[39317]= -2128861181;
assign addr[39318]= -2103375398;
assign addr[39319]= -2067219829;
assign addr[39320]= -2020577882;
assign addr[39321]= -1963686155;
assign addr[39322]= -1896833245;
assign addr[39323]= -1820358275;
assign addr[39324]= -1734649179;
assign addr[39325]= -1640140734;
assign addr[39326]= -1537312353;
assign addr[39327]= -1426685652;
assign addr[39328]= -1308821808;
assign addr[39329]= -1184318708;
assign addr[39330]= -1053807919;
assign addr[39331]= -917951481;
assign addr[39332]= -777438554;
assign addr[39333]= -632981917;
assign addr[39334]= -485314355;
assign addr[39335]= -335184940;
assign addr[39336]= -183355234;
assign addr[39337]= -30595422;
assign addr[39338]= 122319591;
assign addr[39339]= 274614114;
assign addr[39340]= 425515602;
assign addr[39341]= 574258580;
assign addr[39342]= 720088517;
assign addr[39343]= 862265664;
assign addr[39344]= 1000068799;
assign addr[39345]= 1132798888;
assign addr[39346]= 1259782632;
assign addr[39347]= 1380375881;
assign addr[39348]= 1493966902;
assign addr[39349]= 1599979481;
assign addr[39350]= 1697875851;
assign addr[39351]= 1787159411;
assign addr[39352]= 1867377253;
assign addr[39353]= 1938122457;
assign addr[39354]= 1999036154;
assign addr[39355]= 2049809346;
assign addr[39356]= 2090184478;
assign addr[39357]= 2119956737;
assign addr[39358]= 2138975100;
assign addr[39359]= 2147143090;
assign addr[39360]= 2144419275;
assign addr[39361]= 2130817471;
assign addr[39362]= 2106406677;
assign addr[39363]= 2071310720;
assign addr[39364]= 2025707632;
assign addr[39365]= 1969828744;
assign addr[39366]= 1903957513;
assign addr[39367]= 1828428082;
assign addr[39368]= 1743623590;
assign addr[39369]= 1649974225;
assign addr[39370]= 1547955041;
assign addr[39371]= 1438083551;
assign addr[39372]= 1320917099;
assign addr[39373]= 1197050035;
assign addr[39374]= 1067110699;
assign addr[39375]= 931758235;
assign addr[39376]= 791679244;
assign addr[39377]= 647584304;
assign addr[39378]= 500204365;
assign addr[39379]= 350287041;
assign addr[39380]= 198592817;
assign addr[39381]= 45891193;
assign addr[39382]= -107043224;
assign addr[39383]= -259434643;
assign addr[39384]= -410510029;
assign addr[39385]= -559503022;
assign addr[39386]= -705657826;
assign addr[39387]= -848233042;
assign addr[39388]= -986505429;
assign addr[39389]= -1119773573;
assign addr[39390]= -1247361445;
assign addr[39391]= -1368621831;
assign addr[39392]= -1482939614;
assign addr[39393]= -1589734894;
assign addr[39394]= -1688465931;
assign addr[39395]= -1778631892;
assign addr[39396]= -1859775393;
assign addr[39397]= -1931484818;
assign addr[39398]= -1993396407;
assign addr[39399]= -2045196100;
assign addr[39400]= -2086621133;
assign addr[39401]= -2117461370;
assign addr[39402]= -2137560369;
assign addr[39403]= -2146816171;
assign addr[39404]= -2145181827;
assign addr[39405]= -2132665626;
assign addr[39406]= -2109331059;
assign addr[39407]= -2075296495;
assign addr[39408]= -2030734582;
assign addr[39409]= -1975871368;
assign addr[39410]= -1910985158;
assign addr[39411]= -1836405100;
assign addr[39412]= -1752509516;
assign addr[39413]= -1659723983;
assign addr[39414]= -1558519173;
assign addr[39415]= -1449408469;
assign addr[39416]= -1332945355;
assign addr[39417]= -1209720613;
assign addr[39418]= -1080359326;
assign addr[39419]= -945517704;
assign addr[39420]= -805879757;
assign addr[39421]= -662153826;
assign addr[39422]= -515068990;
assign addr[39423]= -365371365;
assign addr[39424]= -213820322;
assign addr[39425]= -61184634;
assign addr[39426]= 91761426;
assign addr[39427]= 244242007;
assign addr[39428]= 395483624;
assign addr[39429]= 544719071;
assign addr[39430]= 691191324;
assign addr[39431]= 834157373;
assign addr[39432]= 972891995;
assign addr[39433]= 1106691431;
assign addr[39434]= 1234876957;
assign addr[39435]= 1356798326;
assign addr[39436]= 1471837070;
assign addr[39437]= 1579409630;
assign addr[39438]= 1678970324;
assign addr[39439]= 1770014111;
assign addr[39440]= 1852079154;
assign addr[39441]= 1924749160;
assign addr[39442]= 1987655498;
assign addr[39443]= 2040479063;
assign addr[39444]= 2082951896;
assign addr[39445]= 2114858546;
assign addr[39446]= 2136037160;
assign addr[39447]= 2146380306;
assign addr[39448]= 2145835515;
assign addr[39449]= 2134405552;
assign addr[39450]= 2112148396;
assign addr[39451]= 2079176953;
assign addr[39452]= 2035658475;
assign addr[39453]= 1981813720;
assign addr[39454]= 1917915825;
assign addr[39455]= 1844288924;
assign addr[39456]= 1761306505;
assign addr[39457]= 1669389513;
assign addr[39458]= 1569004214;
assign addr[39459]= 1460659832;
assign addr[39460]= 1344905966;
assign addr[39461]= 1222329801;
assign addr[39462]= 1093553126;
assign addr[39463]= 959229189;
assign addr[39464]= 820039373;
assign addr[39465]= 676689746;
assign addr[39466]= 529907477;
assign addr[39467]= 380437148;
assign addr[39468]= 229036977;
assign addr[39469]= 76474970;
assign addr[39470]= -76474970;
assign addr[39471]= -229036977;
assign addr[39472]= -380437148;
assign addr[39473]= -529907477;
assign addr[39474]= -676689746;
assign addr[39475]= -820039373;
assign addr[39476]= -959229189;
assign addr[39477]= -1093553126;
assign addr[39478]= -1222329801;
assign addr[39479]= -1344905966;
assign addr[39480]= -1460659832;
assign addr[39481]= -1569004214;
assign addr[39482]= -1669389513;
assign addr[39483]= -1761306505;
assign addr[39484]= -1844288924;
assign addr[39485]= -1917915825;
assign addr[39486]= -1981813720;
assign addr[39487]= -2035658475;
assign addr[39488]= -2079176953;
assign addr[39489]= -2112148396;
assign addr[39490]= -2134405552;
assign addr[39491]= -2145835515;
assign addr[39492]= -2146380306;
assign addr[39493]= -2136037160;
assign addr[39494]= -2114858546;
assign addr[39495]= -2082951896;
assign addr[39496]= -2040479063;
assign addr[39497]= -1987655498;
assign addr[39498]= -1924749160;
assign addr[39499]= -1852079154;
assign addr[39500]= -1770014111;
assign addr[39501]= -1678970324;
assign addr[39502]= -1579409630;
assign addr[39503]= -1471837070;
assign addr[39504]= -1356798326;
assign addr[39505]= -1234876957;
assign addr[39506]= -1106691431;
assign addr[39507]= -972891995;
assign addr[39508]= -834157373;
assign addr[39509]= -691191324;
assign addr[39510]= -544719071;
assign addr[39511]= -395483624;
assign addr[39512]= -244242007;
assign addr[39513]= -91761426;
assign addr[39514]= 61184634;
assign addr[39515]= 213820322;
assign addr[39516]= 365371365;
assign addr[39517]= 515068990;
assign addr[39518]= 662153826;
assign addr[39519]= 805879757;
assign addr[39520]= 945517704;
assign addr[39521]= 1080359326;
assign addr[39522]= 1209720613;
assign addr[39523]= 1332945355;
assign addr[39524]= 1449408469;
assign addr[39525]= 1558519173;
assign addr[39526]= 1659723983;
assign addr[39527]= 1752509516;
assign addr[39528]= 1836405100;
assign addr[39529]= 1910985158;
assign addr[39530]= 1975871368;
assign addr[39531]= 2030734582;
assign addr[39532]= 2075296495;
assign addr[39533]= 2109331059;
assign addr[39534]= 2132665626;
assign addr[39535]= 2145181827;
assign addr[39536]= 2146816171;
assign addr[39537]= 2137560369;
assign addr[39538]= 2117461370;
assign addr[39539]= 2086621133;
assign addr[39540]= 2045196100;
assign addr[39541]= 1993396407;
assign addr[39542]= 1931484818;
assign addr[39543]= 1859775393;
assign addr[39544]= 1778631892;
assign addr[39545]= 1688465931;
assign addr[39546]= 1589734894;
assign addr[39547]= 1482939614;
assign addr[39548]= 1368621831;
assign addr[39549]= 1247361445;
assign addr[39550]= 1119773573;
assign addr[39551]= 986505429;
assign addr[39552]= 848233042;
assign addr[39553]= 705657826;
assign addr[39554]= 559503022;
assign addr[39555]= 410510029;
assign addr[39556]= 259434643;
assign addr[39557]= 107043224;
assign addr[39558]= -45891193;
assign addr[39559]= -198592817;
assign addr[39560]= -350287041;
assign addr[39561]= -500204365;
assign addr[39562]= -647584304;
assign addr[39563]= -791679244;
assign addr[39564]= -931758235;
assign addr[39565]= -1067110699;
assign addr[39566]= -1197050035;
assign addr[39567]= -1320917099;
assign addr[39568]= -1438083551;
assign addr[39569]= -1547955041;
assign addr[39570]= -1649974225;
assign addr[39571]= -1743623590;
assign addr[39572]= -1828428082;
assign addr[39573]= -1903957513;
assign addr[39574]= -1969828744;
assign addr[39575]= -2025707632;
assign addr[39576]= -2071310720;
assign addr[39577]= -2106406677;
assign addr[39578]= -2130817471;
assign addr[39579]= -2144419275;
assign addr[39580]= -2147143090;
assign addr[39581]= -2138975100;
assign addr[39582]= -2119956737;
assign addr[39583]= -2090184478;
assign addr[39584]= -2049809346;
assign addr[39585]= -1999036154;
assign addr[39586]= -1938122457;
assign addr[39587]= -1867377253;
assign addr[39588]= -1787159411;
assign addr[39589]= -1697875851;
assign addr[39590]= -1599979481;
assign addr[39591]= -1493966902;
assign addr[39592]= -1380375881;
assign addr[39593]= -1259782632;
assign addr[39594]= -1132798888;
assign addr[39595]= -1000068799;
assign addr[39596]= -862265664;
assign addr[39597]= -720088517;
assign addr[39598]= -574258580;
assign addr[39599]= -425515602;
assign addr[39600]= -274614114;
assign addr[39601]= -122319591;
assign addr[39602]= 30595422;
assign addr[39603]= 183355234;
assign addr[39604]= 335184940;
assign addr[39605]= 485314355;
assign addr[39606]= 632981917;
assign addr[39607]= 777438554;
assign addr[39608]= 917951481;
assign addr[39609]= 1053807919;
assign addr[39610]= 1184318708;
assign addr[39611]= 1308821808;
assign addr[39612]= 1426685652;
assign addr[39613]= 1537312353;
assign addr[39614]= 1640140734;
assign addr[39615]= 1734649179;
assign addr[39616]= 1820358275;
assign addr[39617]= 1896833245;
assign addr[39618]= 1963686155;
assign addr[39619]= 2020577882;
assign addr[39620]= 2067219829;
assign addr[39621]= 2103375398;
assign addr[39622]= 2128861181;
assign addr[39623]= 2143547897;
assign addr[39624]= 2147361045;
assign addr[39625]= 2140281282;
assign addr[39626]= 2122344521;
assign addr[39627]= 2093641749;
assign addr[39628]= 2054318569;
assign addr[39629]= 2004574453;
assign addr[39630]= 1944661739;
assign addr[39631]= 1874884346;
assign addr[39632]= 1795596234;
assign addr[39633]= 1707199606;
assign addr[39634]= 1610142873;
assign addr[39635]= 1504918373;
assign addr[39636]= 1392059879;
assign addr[39637]= 1272139887;
assign addr[39638]= 1145766716;
assign addr[39639]= 1013581418;
assign addr[39640]= 876254528;
assign addr[39641]= 734482665;
assign addr[39642]= 588984994;
assign addr[39643]= 440499581;
assign addr[39644]= 289779648;
assign addr[39645]= 137589750;
assign addr[39646]= -15298099;
assign addr[39647]= -168108346;
assign addr[39648]= -320065829;
assign addr[39649]= -470399716;
assign addr[39650]= -618347408;
assign addr[39651]= -763158411;
assign addr[39652]= -904098143;
assign addr[39653]= -1040451659;
assign addr[39654]= -1171527280;
assign addr[39655]= -1296660098;
assign addr[39656]= -1415215352;
assign addr[39657]= -1526591649;
assign addr[39658]= -1630224009;
assign addr[39659]= -1725586737;
assign addr[39660]= -1812196087;
assign addr[39661]= -1889612716;
assign addr[39662]= -1957443913;
assign addr[39663]= -2015345591;
assign addr[39664]= -2063024031;
assign addr[39665]= -2100237377;
assign addr[39666]= -2126796855;
assign addr[39667]= -2142567738;
assign addr[39668]= -2147470025;
assign addr[39669]= -2141478848;
assign addr[39670]= -2124624598;
assign addr[39671]= -2096992772;
assign addr[39672]= -2058723538;
assign addr[39673]= -2010011024;
assign addr[39674]= -1951102334;
assign addr[39675]= -1882296293;
assign addr[39676]= -1803941934;
assign addr[39677]= -1716436725;
assign addr[39678]= -1620224553;
assign addr[39679]= -1515793473;
assign addr[39680]= -1403673233;
assign addr[39681]= -1284432584;
assign addr[39682]= -1158676398;
assign addr[39683]= -1027042599;
assign addr[39684]= -890198924;
assign addr[39685]= -748839539;
assign addr[39686]= -603681519;
assign addr[39687]= -455461206;
assign addr[39688]= -304930476;
assign addr[39689]= -152852926;
assign addr[39690]= 0;
assign addr[39691]= 152852926;
assign addr[39692]= 304930476;
assign addr[39693]= 455461206;
assign addr[39694]= 603681519;
assign addr[39695]= 748839539;
assign addr[39696]= 890198924;
assign addr[39697]= 1027042599;
assign addr[39698]= 1158676398;
assign addr[39699]= 1284432584;
assign addr[39700]= 1403673233;
assign addr[39701]= 1515793473;
assign addr[39702]= 1620224553;
assign addr[39703]= 1716436725;
assign addr[39704]= 1803941934;
assign addr[39705]= 1882296293;
assign addr[39706]= 1951102334;
assign addr[39707]= 2010011024;
assign addr[39708]= 2058723538;
assign addr[39709]= 2096992772;
assign addr[39710]= 2124624598;
assign addr[39711]= 2141478848;
assign addr[39712]= 2147470025;
assign addr[39713]= 2142567738;
assign addr[39714]= 2126796855;
assign addr[39715]= 2100237377;
assign addr[39716]= 2063024031;
assign addr[39717]= 2015345591;
assign addr[39718]= 1957443913;
assign addr[39719]= 1889612716;
assign addr[39720]= 1812196087;
assign addr[39721]= 1725586737;
assign addr[39722]= 1630224009;
assign addr[39723]= 1526591649;
assign addr[39724]= 1415215352;
assign addr[39725]= 1296660098;
assign addr[39726]= 1171527280;
assign addr[39727]= 1040451659;
assign addr[39728]= 904098143;
assign addr[39729]= 763158411;
assign addr[39730]= 618347408;
assign addr[39731]= 470399716;
assign addr[39732]= 320065829;
assign addr[39733]= 168108346;
assign addr[39734]= 15298099;
assign addr[39735]= -137589750;
assign addr[39736]= -289779648;
assign addr[39737]= -440499581;
assign addr[39738]= -588984994;
assign addr[39739]= -734482665;
assign addr[39740]= -876254528;
assign addr[39741]= -1013581418;
assign addr[39742]= -1145766716;
assign addr[39743]= -1272139887;
assign addr[39744]= -1392059879;
assign addr[39745]= -1504918373;
assign addr[39746]= -1610142873;
assign addr[39747]= -1707199606;
assign addr[39748]= -1795596234;
assign addr[39749]= -1874884346;
assign addr[39750]= -1944661739;
assign addr[39751]= -2004574453;
assign addr[39752]= -2054318569;
assign addr[39753]= -2093641749;
assign addr[39754]= -2122344521;
assign addr[39755]= -2140281282;
assign addr[39756]= -2147361045;
assign addr[39757]= -2143547897;
assign addr[39758]= -2128861181;
assign addr[39759]= -2103375398;
assign addr[39760]= -2067219829;
assign addr[39761]= -2020577882;
assign addr[39762]= -1963686155;
assign addr[39763]= -1896833245;
assign addr[39764]= -1820358275;
assign addr[39765]= -1734649179;
assign addr[39766]= -1640140734;
assign addr[39767]= -1537312353;
assign addr[39768]= -1426685652;
assign addr[39769]= -1308821808;
assign addr[39770]= -1184318708;
assign addr[39771]= -1053807919;
assign addr[39772]= -917951481;
assign addr[39773]= -777438554;
assign addr[39774]= -632981917;
assign addr[39775]= -485314355;
assign addr[39776]= -335184940;
assign addr[39777]= -183355234;
assign addr[39778]= -30595422;
assign addr[39779]= 122319591;
assign addr[39780]= 274614114;
assign addr[39781]= 425515602;
assign addr[39782]= 574258580;
assign addr[39783]= 720088517;
assign addr[39784]= 862265664;
assign addr[39785]= 1000068799;
assign addr[39786]= 1132798888;
assign addr[39787]= 1259782632;
assign addr[39788]= 1380375881;
assign addr[39789]= 1493966902;
assign addr[39790]= 1599979481;
assign addr[39791]= 1697875851;
assign addr[39792]= 1787159411;
assign addr[39793]= 1867377253;
assign addr[39794]= 1938122457;
assign addr[39795]= 1999036154;
assign addr[39796]= 2049809346;
assign addr[39797]= 2090184478;
assign addr[39798]= 2119956737;
assign addr[39799]= 2138975100;
assign addr[39800]= 2147143090;
assign addr[39801]= 2144419275;
assign addr[39802]= 2130817471;
assign addr[39803]= 2106406677;
assign addr[39804]= 2071310720;
assign addr[39805]= 2025707632;
assign addr[39806]= 1969828744;
assign addr[39807]= 1903957513;
assign addr[39808]= 1828428082;
assign addr[39809]= 1743623590;
assign addr[39810]= 1649974225;
assign addr[39811]= 1547955041;
assign addr[39812]= 1438083551;
assign addr[39813]= 1320917099;
assign addr[39814]= 1197050035;
assign addr[39815]= 1067110699;
assign addr[39816]= 931758235;
assign addr[39817]= 791679244;
assign addr[39818]= 647584304;
assign addr[39819]= 500204365;
assign addr[39820]= 350287041;
assign addr[39821]= 198592817;
assign addr[39822]= 45891193;
assign addr[39823]= -107043224;
assign addr[39824]= -259434643;
assign addr[39825]= -410510029;
assign addr[39826]= -559503022;
assign addr[39827]= -705657826;
assign addr[39828]= -848233042;
assign addr[39829]= -986505429;
assign addr[39830]= -1119773573;
assign addr[39831]= -1247361445;
assign addr[39832]= -1368621831;
assign addr[39833]= -1482939614;
assign addr[39834]= -1589734894;
assign addr[39835]= -1688465931;
assign addr[39836]= -1778631892;
assign addr[39837]= -1859775393;
assign addr[39838]= -1931484818;
assign addr[39839]= -1993396407;
assign addr[39840]= -2045196100;
assign addr[39841]= -2086621133;
assign addr[39842]= -2117461370;
assign addr[39843]= -2137560369;
assign addr[39844]= -2146816171;
assign addr[39845]= -2145181827;
assign addr[39846]= -2132665626;
assign addr[39847]= -2109331059;
assign addr[39848]= -2075296495;
assign addr[39849]= -2030734582;
assign addr[39850]= -1975871368;
assign addr[39851]= -1910985158;
assign addr[39852]= -1836405100;
assign addr[39853]= -1752509516;
assign addr[39854]= -1659723983;
assign addr[39855]= -1558519173;
assign addr[39856]= -1449408469;
assign addr[39857]= -1332945355;
assign addr[39858]= -1209720613;
assign addr[39859]= -1080359326;
assign addr[39860]= -945517704;
assign addr[39861]= -805879757;
assign addr[39862]= -662153826;
assign addr[39863]= -515068990;
assign addr[39864]= -365371365;
assign addr[39865]= -213820322;
assign addr[39866]= -61184634;
assign addr[39867]= 91761426;
assign addr[39868]= 244242007;
assign addr[39869]= 395483624;
assign addr[39870]= 544719071;
assign addr[39871]= 691191324;
assign addr[39872]= 834157373;
assign addr[39873]= 972891995;
assign addr[39874]= 1106691431;
assign addr[39875]= 1234876957;
assign addr[39876]= 1356798326;
assign addr[39877]= 1471837070;
assign addr[39878]= 1579409630;
assign addr[39879]= 1678970324;
assign addr[39880]= 1770014111;
assign addr[39881]= 1852079154;
assign addr[39882]= 1924749160;
assign addr[39883]= 1987655498;
assign addr[39884]= 2040479063;
assign addr[39885]= 2082951896;
assign addr[39886]= 2114858546;
assign addr[39887]= 2136037160;
assign addr[39888]= 2146380306;
assign addr[39889]= 2145835515;
assign addr[39890]= 2134405552;
assign addr[39891]= 2112148396;
assign addr[39892]= 2079176953;
assign addr[39893]= 2035658475;
assign addr[39894]= 1981813720;
assign addr[39895]= 1917915825;
assign addr[39896]= 1844288924;
assign addr[39897]= 1761306505;
assign addr[39898]= 1669389513;
assign addr[39899]= 1569004214;
assign addr[39900]= 1460659832;
assign addr[39901]= 1344905966;
assign addr[39902]= 1222329801;
assign addr[39903]= 1093553126;
assign addr[39904]= 959229189;
assign addr[39905]= 820039373;
assign addr[39906]= 676689746;
assign addr[39907]= 529907477;
assign addr[39908]= 380437148;
assign addr[39909]= 229036977;
assign addr[39910]= 76474970;
assign addr[39911]= -76474970;
assign addr[39912]= -229036977;
assign addr[39913]= -380437148;
assign addr[39914]= -529907477;
assign addr[39915]= -676689746;
assign addr[39916]= -820039373;
assign addr[39917]= -959229189;
assign addr[39918]= -1093553126;
assign addr[39919]= -1222329801;
assign addr[39920]= -1344905966;
assign addr[39921]= -1460659832;
assign addr[39922]= -1569004214;
assign addr[39923]= -1669389513;
assign addr[39924]= -1761306505;
assign addr[39925]= -1844288924;
assign addr[39926]= -1917915825;
assign addr[39927]= -1981813720;
assign addr[39928]= -2035658475;
assign addr[39929]= -2079176953;
assign addr[39930]= -2112148396;
assign addr[39931]= -2134405552;
assign addr[39932]= -2145835515;
assign addr[39933]= -2146380306;
assign addr[39934]= -2136037160;
assign addr[39935]= -2114858546;
assign addr[39936]= -2082951896;
assign addr[39937]= -2040479063;
assign addr[39938]= -1987655498;
assign addr[39939]= -1924749160;
assign addr[39940]= -1852079154;
assign addr[39941]= -1770014111;
assign addr[39942]= -1678970324;
assign addr[39943]= -1579409630;
assign addr[39944]= -1471837070;
assign addr[39945]= -1356798326;
assign addr[39946]= -1234876957;
assign addr[39947]= -1106691431;
assign addr[39948]= -972891995;
assign addr[39949]= -834157373;
assign addr[39950]= -691191324;
assign addr[39951]= -544719071;
assign addr[39952]= -395483624;
assign addr[39953]= -244242007;
assign addr[39954]= -91761426;
assign addr[39955]= 61184634;
assign addr[39956]= 213820322;
assign addr[39957]= 365371365;
assign addr[39958]= 515068990;
assign addr[39959]= 662153826;
assign addr[39960]= 805879757;
assign addr[39961]= 945517704;
assign addr[39962]= 1080359326;
assign addr[39963]= 1209720613;
assign addr[39964]= 1332945355;
assign addr[39965]= 1449408469;
assign addr[39966]= 1558519173;
assign addr[39967]= 1659723983;
assign addr[39968]= 1752509516;
assign addr[39969]= 1836405100;
assign addr[39970]= 1910985158;
assign addr[39971]= 1975871368;
assign addr[39972]= 2030734582;
assign addr[39973]= 2075296495;
assign addr[39974]= 2109331059;
assign addr[39975]= 2132665626;
assign addr[39976]= 2145181827;
assign addr[39977]= 2146816171;
assign addr[39978]= 2137560369;
assign addr[39979]= 2117461370;
assign addr[39980]= 2086621133;
assign addr[39981]= 2045196100;
assign addr[39982]= 1993396407;
assign addr[39983]= 1931484818;
assign addr[39984]= 1859775393;
assign addr[39985]= 1778631892;
assign addr[39986]= 1688465931;
assign addr[39987]= 1589734894;
assign addr[39988]= 1482939614;
assign addr[39989]= 1368621831;
assign addr[39990]= 1247361445;
assign addr[39991]= 1119773573;
assign addr[39992]= 986505429;
assign addr[39993]= 848233042;
assign addr[39994]= 705657826;
assign addr[39995]= 559503022;
assign addr[39996]= 410510029;
assign addr[39997]= 259434643;
assign addr[39998]= 107043224;
assign addr[39999]= -45891193;
assign addr[40000]= -198592817;
assign addr[40001]= -350287041;
assign addr[40002]= -500204365;
assign addr[40003]= -647584304;
assign addr[40004]= -791679244;
assign addr[40005]= -931758235;
assign addr[40006]= -1067110699;
assign addr[40007]= -1197050035;
assign addr[40008]= -1320917099;
assign addr[40009]= -1438083551;
assign addr[40010]= -1547955041;
assign addr[40011]= -1649974225;
assign addr[40012]= -1743623590;
assign addr[40013]= -1828428082;
assign addr[40014]= -1903957513;
assign addr[40015]= -1969828744;
assign addr[40016]= -2025707632;
assign addr[40017]= -2071310720;
assign addr[40018]= -2106406677;
assign addr[40019]= -2130817471;
assign addr[40020]= -2144419275;
assign addr[40021]= -2147143090;
assign addr[40022]= -2138975100;
assign addr[40023]= -2119956737;
assign addr[40024]= -2090184478;
assign addr[40025]= -2049809346;
assign addr[40026]= -1999036154;
assign addr[40027]= -1938122457;
assign addr[40028]= -1867377253;
assign addr[40029]= -1787159411;
assign addr[40030]= -1697875851;
assign addr[40031]= -1599979481;
assign addr[40032]= -1493966902;
assign addr[40033]= -1380375881;
assign addr[40034]= -1259782632;
assign addr[40035]= -1132798888;
assign addr[40036]= -1000068799;
assign addr[40037]= -862265664;
assign addr[40038]= -720088517;
assign addr[40039]= -574258580;
assign addr[40040]= -425515602;
assign addr[40041]= -274614114;
assign addr[40042]= -122319591;
assign addr[40043]= 30595422;
assign addr[40044]= 183355234;
assign addr[40045]= 335184940;
assign addr[40046]= 485314355;
assign addr[40047]= 632981917;
assign addr[40048]= 777438554;
assign addr[40049]= 917951481;
assign addr[40050]= 1053807919;
assign addr[40051]= 1184318708;
assign addr[40052]= 1308821808;
assign addr[40053]= 1426685652;
assign addr[40054]= 1537312353;
assign addr[40055]= 1640140734;
assign addr[40056]= 1734649179;
assign addr[40057]= 1820358275;
assign addr[40058]= 1896833245;
assign addr[40059]= 1963686155;
assign addr[40060]= 2020577882;
assign addr[40061]= 2067219829;
assign addr[40062]= 2103375398;
assign addr[40063]= 2128861181;
assign addr[40064]= 2143547897;
assign addr[40065]= 2147361045;
assign addr[40066]= 2140281282;
assign addr[40067]= 2122344521;
assign addr[40068]= 2093641749;
assign addr[40069]= 2054318569;
assign addr[40070]= 2004574453;
assign addr[40071]= 1944661739;
assign addr[40072]= 1874884346;
assign addr[40073]= 1795596234;
assign addr[40074]= 1707199606;
assign addr[40075]= 1610142873;
assign addr[40076]= 1504918373;
assign addr[40077]= 1392059879;
assign addr[40078]= 1272139887;
assign addr[40079]= 1145766716;
assign addr[40080]= 1013581418;
assign addr[40081]= 876254528;
assign addr[40082]= 734482665;
assign addr[40083]= 588984994;
assign addr[40084]= 440499581;
assign addr[40085]= 289779648;
assign addr[40086]= 137589750;
assign addr[40087]= -15298099;
assign addr[40088]= -168108346;
assign addr[40089]= -320065829;
assign addr[40090]= -470399716;
assign addr[40091]= -618347408;
assign addr[40092]= -763158411;
assign addr[40093]= -904098143;
assign addr[40094]= -1040451659;
assign addr[40095]= -1171527280;
assign addr[40096]= -1296660098;
assign addr[40097]= -1415215352;
assign addr[40098]= -1526591649;
assign addr[40099]= -1630224009;
assign addr[40100]= -1725586737;
assign addr[40101]= -1812196087;
assign addr[40102]= -1889612716;
assign addr[40103]= -1957443913;
assign addr[40104]= -2015345591;
assign addr[40105]= -2063024031;
assign addr[40106]= -2100237377;
assign addr[40107]= -2126796855;
assign addr[40108]= -2142567738;
assign addr[40109]= -2147470025;
assign addr[40110]= -2141478848;
assign addr[40111]= -2124624598;
assign addr[40112]= -2096992772;
assign addr[40113]= -2058723538;
assign addr[40114]= -2010011024;
assign addr[40115]= -1951102334;
assign addr[40116]= -1882296293;
assign addr[40117]= -1803941934;
assign addr[40118]= -1716436725;
assign addr[40119]= -1620224553;
assign addr[40120]= -1515793473;
assign addr[40121]= -1403673233;
assign addr[40122]= -1284432584;
assign addr[40123]= -1158676398;
assign addr[40124]= -1027042599;
assign addr[40125]= -890198924;
assign addr[40126]= -748839539;
assign addr[40127]= -603681519;
assign addr[40128]= -455461206;
assign addr[40129]= -304930476;
assign addr[40130]= -152852926;
assign addr[40131]= 0;
assign addr[40132]= 152852926;
assign addr[40133]= 304930476;
assign addr[40134]= 455461206;
assign addr[40135]= 603681519;
assign addr[40136]= 748839539;
assign addr[40137]= 890198924;
assign addr[40138]= 1027042599;
assign addr[40139]= 1158676398;
assign addr[40140]= 1284432584;
assign addr[40141]= 1403673233;
assign addr[40142]= 1515793473;
assign addr[40143]= 1620224553;
assign addr[40144]= 1716436725;
assign addr[40145]= 1803941934;
assign addr[40146]= 1882296293;
assign addr[40147]= 1951102334;
assign addr[40148]= 2010011024;
assign addr[40149]= 2058723538;
assign addr[40150]= 2096992772;
assign addr[40151]= 2124624598;
assign addr[40152]= 2141478848;
assign addr[40153]= 2147470025;
assign addr[40154]= 2142567738;
assign addr[40155]= 2126796855;
assign addr[40156]= 2100237377;
assign addr[40157]= 2063024031;
assign addr[40158]= 2015345591;
assign addr[40159]= 1957443913;
assign addr[40160]= 1889612716;
assign addr[40161]= 1812196087;
assign addr[40162]= 1725586737;
assign addr[40163]= 1630224009;
assign addr[40164]= 1526591649;
assign addr[40165]= 1415215352;
assign addr[40166]= 1296660098;
assign addr[40167]= 1171527280;
assign addr[40168]= 1040451659;
assign addr[40169]= 904098143;
assign addr[40170]= 763158411;
assign addr[40171]= 618347408;
assign addr[40172]= 470399716;
assign addr[40173]= 320065829;
assign addr[40174]= 168108346;
assign addr[40175]= 15298099;
assign addr[40176]= -137589750;
assign addr[40177]= -289779648;
assign addr[40178]= -440499581;
assign addr[40179]= -588984994;
assign addr[40180]= -734482665;
assign addr[40181]= -876254528;
assign addr[40182]= -1013581418;
assign addr[40183]= -1145766716;
assign addr[40184]= -1272139887;
assign addr[40185]= -1392059879;
assign addr[40186]= -1504918373;
assign addr[40187]= -1610142873;
assign addr[40188]= -1707199606;
assign addr[40189]= -1795596234;
assign addr[40190]= -1874884346;
assign addr[40191]= -1944661739;
assign addr[40192]= -2004574453;
assign addr[40193]= -2054318569;
assign addr[40194]= -2093641749;
assign addr[40195]= -2122344521;
assign addr[40196]= -2140281282;
assign addr[40197]= -2147361045;
assign addr[40198]= -2143547897;
assign addr[40199]= -2128861181;
assign addr[40200]= -2103375398;
assign addr[40201]= -2067219829;
assign addr[40202]= -2020577882;
assign addr[40203]= -1963686155;
assign addr[40204]= -1896833245;
assign addr[40205]= -1820358275;
assign addr[40206]= -1734649179;
assign addr[40207]= -1640140734;
assign addr[40208]= -1537312353;
assign addr[40209]= -1426685652;
assign addr[40210]= -1308821808;
assign addr[40211]= -1184318708;
assign addr[40212]= -1053807919;
assign addr[40213]= -917951481;
assign addr[40214]= -777438554;
assign addr[40215]= -632981917;
assign addr[40216]= -485314355;
assign addr[40217]= -335184940;
assign addr[40218]= -183355234;
assign addr[40219]= -30595422;
assign addr[40220]= 122319591;
assign addr[40221]= 274614114;
assign addr[40222]= 425515602;
assign addr[40223]= 574258580;
assign addr[40224]= 720088517;
assign addr[40225]= 862265664;
assign addr[40226]= 1000068799;
assign addr[40227]= 1132798888;
assign addr[40228]= 1259782632;
assign addr[40229]= 1380375881;
assign addr[40230]= 1493966902;
assign addr[40231]= 1599979481;
assign addr[40232]= 1697875851;
assign addr[40233]= 1787159411;
assign addr[40234]= 1867377253;
assign addr[40235]= 1938122457;
assign addr[40236]= 1999036154;
assign addr[40237]= 2049809346;
assign addr[40238]= 2090184478;
assign addr[40239]= 2119956737;
assign addr[40240]= 2138975100;
assign addr[40241]= 2147143090;
assign addr[40242]= 2144419275;
assign addr[40243]= 2130817471;
assign addr[40244]= 2106406677;
assign addr[40245]= 2071310720;
assign addr[40246]= 2025707632;
assign addr[40247]= 1969828744;
assign addr[40248]= 1903957513;
assign addr[40249]= 1828428082;
assign addr[40250]= 1743623590;
assign addr[40251]= 1649974225;
assign addr[40252]= 1547955041;
assign addr[40253]= 1438083551;
assign addr[40254]= 1320917099;
assign addr[40255]= 1197050035;
assign addr[40256]= 1067110699;
assign addr[40257]= 931758235;
assign addr[40258]= 791679244;
assign addr[40259]= 647584304;
assign addr[40260]= 500204365;
assign addr[40261]= 350287041;
assign addr[40262]= 198592817;
assign addr[40263]= 45891193;
assign addr[40264]= -107043224;
assign addr[40265]= -259434643;
assign addr[40266]= -410510029;
assign addr[40267]= -559503022;
assign addr[40268]= -705657826;
assign addr[40269]= -848233042;
assign addr[40270]= -986505429;
assign addr[40271]= -1119773573;
assign addr[40272]= -1247361445;
assign addr[40273]= -1368621831;
assign addr[40274]= -1482939614;
assign addr[40275]= -1589734894;
assign addr[40276]= -1688465931;
assign addr[40277]= -1778631892;
assign addr[40278]= -1859775393;
assign addr[40279]= -1931484818;
assign addr[40280]= -1993396407;
assign addr[40281]= -2045196100;
assign addr[40282]= -2086621133;
assign addr[40283]= -2117461370;
assign addr[40284]= -2137560369;
assign addr[40285]= -2146816171;
assign addr[40286]= -2145181827;
assign addr[40287]= -2132665626;
assign addr[40288]= -2109331059;
assign addr[40289]= -2075296495;
assign addr[40290]= -2030734582;
assign addr[40291]= -1975871368;
assign addr[40292]= -1910985158;
assign addr[40293]= -1836405100;
assign addr[40294]= -1752509516;
assign addr[40295]= -1659723983;
assign addr[40296]= -1558519173;
assign addr[40297]= -1449408469;
assign addr[40298]= -1332945355;
assign addr[40299]= -1209720613;
assign addr[40300]= -1080359326;
assign addr[40301]= -945517704;
assign addr[40302]= -805879757;
assign addr[40303]= -662153826;
assign addr[40304]= -515068990;
assign addr[40305]= -365371365;
assign addr[40306]= -213820322;
assign addr[40307]= -61184634;
assign addr[40308]= 91761426;
assign addr[40309]= 244242007;
assign addr[40310]= 395483624;
assign addr[40311]= 544719071;
assign addr[40312]= 691191324;
assign addr[40313]= 834157373;
assign addr[40314]= 972891995;
assign addr[40315]= 1106691431;
assign addr[40316]= 1234876957;
assign addr[40317]= 1356798326;
assign addr[40318]= 1471837070;
assign addr[40319]= 1579409630;
assign addr[40320]= 1678970324;
assign addr[40321]= 1770014111;
assign addr[40322]= 1852079154;
assign addr[40323]= 1924749160;
assign addr[40324]= 1987655498;
assign addr[40325]= 2040479063;
assign addr[40326]= 2082951896;
assign addr[40327]= 2114858546;
assign addr[40328]= 2136037160;
assign addr[40329]= 2146380306;
assign addr[40330]= 2145835515;
assign addr[40331]= 2134405552;
assign addr[40332]= 2112148396;
assign addr[40333]= 2079176953;
assign addr[40334]= 2035658475;
assign addr[40335]= 1981813720;
assign addr[40336]= 1917915825;
assign addr[40337]= 1844288924;
assign addr[40338]= 1761306505;
assign addr[40339]= 1669389513;
assign addr[40340]= 1569004214;
assign addr[40341]= 1460659832;
assign addr[40342]= 1344905966;
assign addr[40343]= 1222329801;
assign addr[40344]= 1093553126;
assign addr[40345]= 959229189;
assign addr[40346]= 820039373;
assign addr[40347]= 676689746;
assign addr[40348]= 529907477;
assign addr[40349]= 380437148;
assign addr[40350]= 229036977;
assign addr[40351]= 76474970;
assign addr[40352]= -76474970;
assign addr[40353]= -229036977;
assign addr[40354]= -380437148;
assign addr[40355]= -529907477;
assign addr[40356]= -676689746;
assign addr[40357]= -820039373;
assign addr[40358]= -959229189;
assign addr[40359]= -1093553126;
assign addr[40360]= -1222329801;
assign addr[40361]= -1344905966;
assign addr[40362]= -1460659832;
assign addr[40363]= -1569004214;
assign addr[40364]= -1669389513;
assign addr[40365]= -1761306505;
assign addr[40366]= -1844288924;
assign addr[40367]= -1917915825;
assign addr[40368]= -1981813720;
assign addr[40369]= -2035658475;
assign addr[40370]= -2079176953;
assign addr[40371]= -2112148396;
assign addr[40372]= -2134405552;
assign addr[40373]= -2145835515;
assign addr[40374]= -2146380306;
assign addr[40375]= -2136037160;
assign addr[40376]= -2114858546;
assign addr[40377]= -2082951896;
assign addr[40378]= -2040479063;
assign addr[40379]= -1987655498;
assign addr[40380]= -1924749160;
assign addr[40381]= -1852079154;
assign addr[40382]= -1770014111;
assign addr[40383]= -1678970324;
assign addr[40384]= -1579409630;
assign addr[40385]= -1471837070;
assign addr[40386]= -1356798326;
assign addr[40387]= -1234876957;
assign addr[40388]= -1106691431;
assign addr[40389]= -972891995;
assign addr[40390]= -834157373;
assign addr[40391]= -691191324;
assign addr[40392]= -544719071;
assign addr[40393]= -395483624;
assign addr[40394]= -244242007;
assign addr[40395]= -91761426;
assign addr[40396]= 61184634;
assign addr[40397]= 213820322;
assign addr[40398]= 365371365;
assign addr[40399]= 515068990;
assign addr[40400]= 662153826;
assign addr[40401]= 805879757;
assign addr[40402]= 945517704;
assign addr[40403]= 1080359326;
assign addr[40404]= 1209720613;
assign addr[40405]= 1332945355;
assign addr[40406]= 1449408469;
assign addr[40407]= 1558519173;
assign addr[40408]= 1659723983;
assign addr[40409]= 1752509516;
assign addr[40410]= 1836405100;
assign addr[40411]= 1910985158;
assign addr[40412]= 1975871368;
assign addr[40413]= 2030734582;
assign addr[40414]= 2075296495;
assign addr[40415]= 2109331059;
assign addr[40416]= 2132665626;
assign addr[40417]= 2145181827;
assign addr[40418]= 2146816171;
assign addr[40419]= 2137560369;
assign addr[40420]= 2117461370;
assign addr[40421]= 2086621133;
assign addr[40422]= 2045196100;
assign addr[40423]= 1993396407;
assign addr[40424]= 1931484818;
assign addr[40425]= 1859775393;
assign addr[40426]= 1778631892;
assign addr[40427]= 1688465931;
assign addr[40428]= 1589734894;
assign addr[40429]= 1482939614;
assign addr[40430]= 1368621831;
assign addr[40431]= 1247361445;
assign addr[40432]= 1119773573;
assign addr[40433]= 986505429;
assign addr[40434]= 848233042;
assign addr[40435]= 705657826;
assign addr[40436]= 559503022;
assign addr[40437]= 410510029;
assign addr[40438]= 259434643;
assign addr[40439]= 107043224;
assign addr[40440]= -45891193;
assign addr[40441]= -198592817;
assign addr[40442]= -350287041;
assign addr[40443]= -500204365;
assign addr[40444]= -647584304;
assign addr[40445]= -791679244;
assign addr[40446]= -931758235;
assign addr[40447]= -1067110699;
assign addr[40448]= -1197050035;
assign addr[40449]= -1320917099;
assign addr[40450]= -1438083551;
assign addr[40451]= -1547955041;
assign addr[40452]= -1649974225;
assign addr[40453]= -1743623590;
assign addr[40454]= -1828428082;
assign addr[40455]= -1903957513;
assign addr[40456]= -1969828744;
assign addr[40457]= -2025707632;
assign addr[40458]= -2071310720;
assign addr[40459]= -2106406677;
assign addr[40460]= -2130817471;
assign addr[40461]= -2144419275;
assign addr[40462]= -2147143090;
assign addr[40463]= -2138975100;
assign addr[40464]= -2119956737;
assign addr[40465]= -2090184478;
assign addr[40466]= -2049809346;
assign addr[40467]= -1999036154;
assign addr[40468]= -1938122457;
assign addr[40469]= -1867377253;
assign addr[40470]= -1787159411;
assign addr[40471]= -1697875851;
assign addr[40472]= -1599979481;
assign addr[40473]= -1493966902;
assign addr[40474]= -1380375881;
assign addr[40475]= -1259782632;
assign addr[40476]= -1132798888;
assign addr[40477]= -1000068799;
assign addr[40478]= -862265664;
assign addr[40479]= -720088517;
assign addr[40480]= -574258580;
assign addr[40481]= -425515602;
assign addr[40482]= -274614114;
assign addr[40483]= -122319591;
assign addr[40484]= 30595422;
assign addr[40485]= 183355234;
assign addr[40486]= 335184940;
assign addr[40487]= 485314355;
assign addr[40488]= 632981917;
assign addr[40489]= 777438554;
assign addr[40490]= 917951481;
assign addr[40491]= 1053807919;
assign addr[40492]= 1184318708;
assign addr[40493]= 1308821808;
assign addr[40494]= 1426685652;
assign addr[40495]= 1537312353;
assign addr[40496]= 1640140734;
assign addr[40497]= 1734649179;
assign addr[40498]= 1820358275;
assign addr[40499]= 1896833245;
assign addr[40500]= 1963686155;
assign addr[40501]= 2020577882;
assign addr[40502]= 2067219829;
assign addr[40503]= 2103375398;
assign addr[40504]= 2128861181;
assign addr[40505]= 2143547897;
assign addr[40506]= 2147361045;
assign addr[40507]= 2140281282;
assign addr[40508]= 2122344521;
assign addr[40509]= 2093641749;
assign addr[40510]= 2054318569;
assign addr[40511]= 2004574453;
assign addr[40512]= 1944661739;
assign addr[40513]= 1874884346;
assign addr[40514]= 1795596234;
assign addr[40515]= 1707199606;
assign addr[40516]= 1610142873;
assign addr[40517]= 1504918373;
assign addr[40518]= 1392059879;
assign addr[40519]= 1272139887;
assign addr[40520]= 1145766716;
assign addr[40521]= 1013581418;
assign addr[40522]= 876254528;
assign addr[40523]= 734482665;
assign addr[40524]= 588984994;
assign addr[40525]= 440499581;
assign addr[40526]= 289779648;
assign addr[40527]= 137589750;
assign addr[40528]= -15298099;
assign addr[40529]= -168108346;
assign addr[40530]= -320065829;
assign addr[40531]= -470399716;
assign addr[40532]= -618347408;
assign addr[40533]= -763158411;
assign addr[40534]= -904098143;
assign addr[40535]= -1040451659;
assign addr[40536]= -1171527280;
assign addr[40537]= -1296660098;
assign addr[40538]= -1415215352;
assign addr[40539]= -1526591649;
assign addr[40540]= -1630224009;
assign addr[40541]= -1725586737;
assign addr[40542]= -1812196087;
assign addr[40543]= -1889612716;
assign addr[40544]= -1957443913;
assign addr[40545]= -2015345591;
assign addr[40546]= -2063024031;
assign addr[40547]= -2100237377;
assign addr[40548]= -2126796855;
assign addr[40549]= -2142567738;
assign addr[40550]= -2147470025;
assign addr[40551]= -2141478848;
assign addr[40552]= -2124624598;
assign addr[40553]= -2096992772;
assign addr[40554]= -2058723538;
assign addr[40555]= -2010011024;
assign addr[40556]= -1951102334;
assign addr[40557]= -1882296293;
assign addr[40558]= -1803941934;
assign addr[40559]= -1716436725;
assign addr[40560]= -1620224553;
assign addr[40561]= -1515793473;
assign addr[40562]= -1403673233;
assign addr[40563]= -1284432584;
assign addr[40564]= -1158676398;
assign addr[40565]= -1027042599;
assign addr[40566]= -890198924;
assign addr[40567]= -748839539;
assign addr[40568]= -603681519;
assign addr[40569]= -455461206;
assign addr[40570]= -304930476;
assign addr[40571]= -152852926;
assign addr[40572]= 0;
assign addr[40573]= 152852926;
assign addr[40574]= 304930476;
assign addr[40575]= 455461206;
assign addr[40576]= 603681519;
assign addr[40577]= 748839539;
assign addr[40578]= 890198924;
assign addr[40579]= 1027042599;
assign addr[40580]= 1158676398;
assign addr[40581]= 1284432584;
assign addr[40582]= 1403673233;
assign addr[40583]= 1515793473;
assign addr[40584]= 1620224553;
assign addr[40585]= 1716436725;
assign addr[40586]= 1803941934;
assign addr[40587]= 1882296293;
assign addr[40588]= 1951102334;
assign addr[40589]= 2010011024;
assign addr[40590]= 2058723538;
assign addr[40591]= 2096992772;
assign addr[40592]= 2124624598;
assign addr[40593]= 2141478848;
assign addr[40594]= 2147470025;
assign addr[40595]= 2142567738;
assign addr[40596]= 2126796855;
assign addr[40597]= 2100237377;
assign addr[40598]= 2063024031;
assign addr[40599]= 2015345591;
assign addr[40600]= 1957443913;
assign addr[40601]= 1889612716;
assign addr[40602]= 1812196087;
assign addr[40603]= 1725586737;
assign addr[40604]= 1630224009;
assign addr[40605]= 1526591649;
assign addr[40606]= 1415215352;
assign addr[40607]= 1296660098;
assign addr[40608]= 1171527280;
assign addr[40609]= 1040451659;
assign addr[40610]= 904098143;
assign addr[40611]= 763158411;
assign addr[40612]= 618347408;
assign addr[40613]= 470399716;
assign addr[40614]= 320065829;
assign addr[40615]= 168108346;
assign addr[40616]= 15298099;
assign addr[40617]= -137589750;
assign addr[40618]= -289779648;
assign addr[40619]= -440499581;
assign addr[40620]= -588984994;
assign addr[40621]= -734482665;
assign addr[40622]= -876254528;
assign addr[40623]= -1013581418;
assign addr[40624]= -1145766716;
assign addr[40625]= -1272139887;
assign addr[40626]= -1392059879;
assign addr[40627]= -1504918373;
assign addr[40628]= -1610142873;
assign addr[40629]= -1707199606;
assign addr[40630]= -1795596234;
assign addr[40631]= -1874884346;
assign addr[40632]= -1944661739;
assign addr[40633]= -2004574453;
assign addr[40634]= -2054318569;
assign addr[40635]= -2093641749;
assign addr[40636]= -2122344521;
assign addr[40637]= -2140281282;
assign addr[40638]= -2147361045;
assign addr[40639]= -2143547897;
assign addr[40640]= -2128861181;
assign addr[40641]= -2103375398;
assign addr[40642]= -2067219829;
assign addr[40643]= -2020577882;
assign addr[40644]= -1963686155;
assign addr[40645]= -1896833245;
assign addr[40646]= -1820358275;
assign addr[40647]= -1734649179;
assign addr[40648]= -1640140734;
assign addr[40649]= -1537312353;
assign addr[40650]= -1426685652;
assign addr[40651]= -1308821808;
assign addr[40652]= -1184318708;
assign addr[40653]= -1053807919;
assign addr[40654]= -917951481;
assign addr[40655]= -777438554;
assign addr[40656]= -632981917;
assign addr[40657]= -485314355;
assign addr[40658]= -335184940;
assign addr[40659]= -183355234;
assign addr[40660]= -30595422;
assign addr[40661]= 122319591;
assign addr[40662]= 274614114;
assign addr[40663]= 425515602;
assign addr[40664]= 574258580;
assign addr[40665]= 720088517;
assign addr[40666]= 862265664;
assign addr[40667]= 1000068799;
assign addr[40668]= 1132798888;
assign addr[40669]= 1259782632;
assign addr[40670]= 1380375881;
assign addr[40671]= 1493966902;
assign addr[40672]= 1599979481;
assign addr[40673]= 1697875851;
assign addr[40674]= 1787159411;
assign addr[40675]= 1867377253;
assign addr[40676]= 1938122457;
assign addr[40677]= 1999036154;
assign addr[40678]= 2049809346;
assign addr[40679]= 2090184478;
assign addr[40680]= 2119956737;
assign addr[40681]= 2138975100;
assign addr[40682]= 2147143090;
assign addr[40683]= 2144419275;
assign addr[40684]= 2130817471;
assign addr[40685]= 2106406677;
assign addr[40686]= 2071310720;
assign addr[40687]= 2025707632;
assign addr[40688]= 1969828744;
assign addr[40689]= 1903957513;
assign addr[40690]= 1828428082;
assign addr[40691]= 1743623590;
assign addr[40692]= 1649974225;
assign addr[40693]= 1547955041;
assign addr[40694]= 1438083551;
assign addr[40695]= 1320917099;
assign addr[40696]= 1197050035;
assign addr[40697]= 1067110699;
assign addr[40698]= 931758235;
assign addr[40699]= 791679244;
assign addr[40700]= 647584304;
assign addr[40701]= 500204365;
assign addr[40702]= 350287041;
assign addr[40703]= 198592817;
assign addr[40704]= 45891193;
assign addr[40705]= -107043224;
assign addr[40706]= -259434643;
assign addr[40707]= -410510029;
assign addr[40708]= -559503022;
assign addr[40709]= -705657826;
assign addr[40710]= -848233042;
assign addr[40711]= -986505429;
assign addr[40712]= -1119773573;
assign addr[40713]= -1247361445;
assign addr[40714]= -1368621831;
assign addr[40715]= -1482939614;
assign addr[40716]= -1589734894;
assign addr[40717]= -1688465931;
assign addr[40718]= -1778631892;
assign addr[40719]= -1859775393;
assign addr[40720]= -1931484818;
assign addr[40721]= -1993396407;
assign addr[40722]= -2045196100;
assign addr[40723]= -2086621133;
assign addr[40724]= -2117461370;
assign addr[40725]= -2137560369;
assign addr[40726]= -2146816171;
assign addr[40727]= -2145181827;
assign addr[40728]= -2132665626;
assign addr[40729]= -2109331059;
assign addr[40730]= -2075296495;
assign addr[40731]= -2030734582;
assign addr[40732]= -1975871368;
assign addr[40733]= -1910985158;
assign addr[40734]= -1836405100;
assign addr[40735]= -1752509516;
assign addr[40736]= -1659723983;
assign addr[40737]= -1558519173;
assign addr[40738]= -1449408469;
assign addr[40739]= -1332945355;
assign addr[40740]= -1209720613;
assign addr[40741]= -1080359326;
assign addr[40742]= -945517704;
assign addr[40743]= -805879757;
assign addr[40744]= -662153826;
assign addr[40745]= -515068990;
assign addr[40746]= -365371365;
assign addr[40747]= -213820322;
assign addr[40748]= -61184634;
assign addr[40749]= 91761426;
assign addr[40750]= 244242007;
assign addr[40751]= 395483624;
assign addr[40752]= 544719071;
assign addr[40753]= 691191324;
assign addr[40754]= 834157373;
assign addr[40755]= 972891995;
assign addr[40756]= 1106691431;
assign addr[40757]= 1234876957;
assign addr[40758]= 1356798326;
assign addr[40759]= 1471837070;
assign addr[40760]= 1579409630;
assign addr[40761]= 1678970324;
assign addr[40762]= 1770014111;
assign addr[40763]= 1852079154;
assign addr[40764]= 1924749160;
assign addr[40765]= 1987655498;
assign addr[40766]= 2040479063;
assign addr[40767]= 2082951896;
assign addr[40768]= 2114858546;
assign addr[40769]= 2136037160;
assign addr[40770]= 2146380306;
assign addr[40771]= 2145835515;
assign addr[40772]= 2134405552;
assign addr[40773]= 2112148396;
assign addr[40774]= 2079176953;
assign addr[40775]= 2035658475;
assign addr[40776]= 1981813720;
assign addr[40777]= 1917915825;
assign addr[40778]= 1844288924;
assign addr[40779]= 1761306505;
assign addr[40780]= 1669389513;
assign addr[40781]= 1569004214;
assign addr[40782]= 1460659832;
assign addr[40783]= 1344905966;
assign addr[40784]= 1222329801;
assign addr[40785]= 1093553126;
assign addr[40786]= 959229189;
assign addr[40787]= 820039373;
assign addr[40788]= 676689746;
assign addr[40789]= 529907477;
assign addr[40790]= 380437148;
assign addr[40791]= 229036977;
assign addr[40792]= 76474970;
assign addr[40793]= -76474970;
assign addr[40794]= -229036977;
assign addr[40795]= -380437148;
assign addr[40796]= -529907477;
assign addr[40797]= -676689746;
assign addr[40798]= -820039373;
assign addr[40799]= -959229189;
assign addr[40800]= -1093553126;
assign addr[40801]= -1222329801;
assign addr[40802]= -1344905966;
assign addr[40803]= -1460659832;
assign addr[40804]= -1569004214;
assign addr[40805]= -1669389513;
assign addr[40806]= -1761306505;
assign addr[40807]= -1844288924;
assign addr[40808]= -1917915825;
assign addr[40809]= -1981813720;
assign addr[40810]= -2035658475;
assign addr[40811]= -2079176953;
assign addr[40812]= -2112148396;
assign addr[40813]= -2134405552;
assign addr[40814]= -2145835515;
assign addr[40815]= -2146380306;
assign addr[40816]= -2136037160;
assign addr[40817]= -2114858546;
assign addr[40818]= -2082951896;
assign addr[40819]= -2040479063;
assign addr[40820]= -1987655498;
assign addr[40821]= -1924749160;
assign addr[40822]= -1852079154;
assign addr[40823]= -1770014111;
assign addr[40824]= -1678970324;
assign addr[40825]= -1579409630;
assign addr[40826]= -1471837070;
assign addr[40827]= -1356798326;
assign addr[40828]= -1234876957;
assign addr[40829]= -1106691431;
assign addr[40830]= -972891995;
assign addr[40831]= -834157373;
assign addr[40832]= -691191324;
assign addr[40833]= -544719071;
assign addr[40834]= -395483624;
assign addr[40835]= -244242007;
assign addr[40836]= -91761426;
assign addr[40837]= 61184634;
assign addr[40838]= 213820322;
assign addr[40839]= 365371365;
assign addr[40840]= 515068990;
assign addr[40841]= 662153826;
assign addr[40842]= 805879757;
assign addr[40843]= 945517704;
assign addr[40844]= 1080359326;
assign addr[40845]= 1209720613;
assign addr[40846]= 1332945355;
assign addr[40847]= 1449408469;
assign addr[40848]= 1558519173;
assign addr[40849]= 1659723983;
assign addr[40850]= 1752509516;
assign addr[40851]= 1836405100;
assign addr[40852]= 1910985158;
assign addr[40853]= 1975871368;
assign addr[40854]= 2030734582;
assign addr[40855]= 2075296495;
assign addr[40856]= 2109331059;
assign addr[40857]= 2132665626;
assign addr[40858]= 2145181827;
assign addr[40859]= 2146816171;
assign addr[40860]= 2137560369;
assign addr[40861]= 2117461370;
assign addr[40862]= 2086621133;
assign addr[40863]= 2045196100;
assign addr[40864]= 1993396407;
assign addr[40865]= 1931484818;
assign addr[40866]= 1859775393;
assign addr[40867]= 1778631892;
assign addr[40868]= 1688465931;
assign addr[40869]= 1589734894;
assign addr[40870]= 1482939614;
assign addr[40871]= 1368621831;
assign addr[40872]= 1247361445;
assign addr[40873]= 1119773573;
assign addr[40874]= 986505429;
assign addr[40875]= 848233042;
assign addr[40876]= 705657826;
assign addr[40877]= 559503022;
assign addr[40878]= 410510029;
assign addr[40879]= 259434643;
assign addr[40880]= 107043224;
assign addr[40881]= -45891193;
assign addr[40882]= -198592817;
assign addr[40883]= -350287041;
assign addr[40884]= -500204365;
assign addr[40885]= -647584304;
assign addr[40886]= -791679244;
assign addr[40887]= -931758235;
assign addr[40888]= -1067110699;
assign addr[40889]= -1197050035;
assign addr[40890]= -1320917099;
assign addr[40891]= -1438083551;
assign addr[40892]= -1547955041;
assign addr[40893]= -1649974225;
assign addr[40894]= -1743623590;
assign addr[40895]= -1828428082;
assign addr[40896]= -1903957513;
assign addr[40897]= -1969828744;
assign addr[40898]= -2025707632;
assign addr[40899]= -2071310720;
assign addr[40900]= -2106406677;
assign addr[40901]= -2130817471;
assign addr[40902]= -2144419275;
assign addr[40903]= -2147143090;
assign addr[40904]= -2138975100;
assign addr[40905]= -2119956737;
assign addr[40906]= -2090184478;
assign addr[40907]= -2049809346;
assign addr[40908]= -1999036154;
assign addr[40909]= -1938122457;
assign addr[40910]= -1867377253;
assign addr[40911]= -1787159411;
assign addr[40912]= -1697875851;
assign addr[40913]= -1599979481;
assign addr[40914]= -1493966902;
assign addr[40915]= -1380375881;
assign addr[40916]= -1259782632;
assign addr[40917]= -1132798888;
assign addr[40918]= -1000068799;
assign addr[40919]= -862265664;
assign addr[40920]= -720088517;
assign addr[40921]= -574258580;
assign addr[40922]= -425515602;
assign addr[40923]= -274614114;
assign addr[40924]= -122319591;
assign addr[40925]= 30595422;
assign addr[40926]= 183355234;
assign addr[40927]= 335184940;
assign addr[40928]= 485314355;
assign addr[40929]= 632981917;
assign addr[40930]= 777438554;
assign addr[40931]= 917951481;
assign addr[40932]= 1053807919;
assign addr[40933]= 1184318708;
assign addr[40934]= 1308821808;
assign addr[40935]= 1426685652;
assign addr[40936]= 1537312353;
assign addr[40937]= 1640140734;
assign addr[40938]= 1734649179;
assign addr[40939]= 1820358275;
assign addr[40940]= 1896833245;
assign addr[40941]= 1963686155;
assign addr[40942]= 2020577882;
assign addr[40943]= 2067219829;
assign addr[40944]= 2103375398;
assign addr[40945]= 2128861181;
assign addr[40946]= 2143547897;
assign addr[40947]= 2147361045;
assign addr[40948]= 2140281282;
assign addr[40949]= 2122344521;
assign addr[40950]= 2093641749;
assign addr[40951]= 2054318569;
assign addr[40952]= 2004574453;
assign addr[40953]= 1944661739;
assign addr[40954]= 1874884346;
assign addr[40955]= 1795596234;
assign addr[40956]= 1707199606;
assign addr[40957]= 1610142873;
assign addr[40958]= 1504918373;
assign addr[40959]= 1392059879;
assign addr[40960]= 1272139887;
assign addr[40961]= 1145766716;
assign addr[40962]= 1013581418;
assign addr[40963]= 876254528;
assign addr[40964]= 734482665;
assign addr[40965]= 588984994;
assign addr[40966]= 440499581;
assign addr[40967]= 289779648;
assign addr[40968]= 137589750;
assign addr[40969]= -15298099;
assign addr[40970]= -168108346;
assign addr[40971]= -320065829;
assign addr[40972]= -470399716;
assign addr[40973]= -618347408;
assign addr[40974]= -763158411;
assign addr[40975]= -904098143;
assign addr[40976]= -1040451659;
assign addr[40977]= -1171527280;
assign addr[40978]= -1296660098;
assign addr[40979]= -1415215352;
assign addr[40980]= -1526591649;
assign addr[40981]= -1630224009;
assign addr[40982]= -1725586737;
assign addr[40983]= -1812196087;
assign addr[40984]= -1889612716;
assign addr[40985]= -1957443913;
assign addr[40986]= -2015345591;
assign addr[40987]= -2063024031;
assign addr[40988]= -2100237377;
assign addr[40989]= -2126796855;
assign addr[40990]= -2142567738;
assign addr[40991]= -2147470025;
assign addr[40992]= -2141478848;
assign addr[40993]= -2124624598;
assign addr[40994]= -2096992772;
assign addr[40995]= -2058723538;
assign addr[40996]= -2010011024;
assign addr[40997]= -1951102334;
assign addr[40998]= -1882296293;
assign addr[40999]= -1803941934;
assign addr[41000]= -1716436725;
assign addr[41001]= -1620224553;
assign addr[41002]= -1515793473;
assign addr[41003]= -1403673233;
assign addr[41004]= -1284432584;
assign addr[41005]= -1158676398;
assign addr[41006]= -1027042599;
assign addr[41007]= -890198924;
assign addr[41008]= -748839539;
assign addr[41009]= -603681519;
assign addr[41010]= -455461206;
assign addr[41011]= -304930476;
assign addr[41012]= -152852926;
assign addr[41013]= 0;
assign addr[41014]= 152852926;
assign addr[41015]= 304930476;
assign addr[41016]= 455461206;
assign addr[41017]= 603681519;
assign addr[41018]= 748839539;
assign addr[41019]= 890198924;
assign addr[41020]= 1027042599;
assign addr[41021]= 1158676398;
assign addr[41022]= 1284432584;
assign addr[41023]= 1403673233;
assign addr[41024]= 1515793473;
assign addr[41025]= 1620224553;
assign addr[41026]= 1716436725;
assign addr[41027]= 1803941934;
assign addr[41028]= 1882296293;
assign addr[41029]= 1951102334;
assign addr[41030]= 2010011024;
assign addr[41031]= 2058723538;
assign addr[41032]= 2096992772;
assign addr[41033]= 2124624598;
assign addr[41034]= 2141478848;
assign addr[41035]= 2147470025;
assign addr[41036]= 2142567738;
assign addr[41037]= 2126796855;
assign addr[41038]= 2100237377;
assign addr[41039]= 2063024031;
assign addr[41040]= 2015345591;
assign addr[41041]= 1957443913;
assign addr[41042]= 1889612716;
assign addr[41043]= 1812196087;
assign addr[41044]= 1725586737;
assign addr[41045]= 1630224009;
assign addr[41046]= 1526591649;
assign addr[41047]= 1415215352;
assign addr[41048]= 1296660098;
assign addr[41049]= 1171527280;
assign addr[41050]= 1040451659;
assign addr[41051]= 904098143;
assign addr[41052]= 763158411;
assign addr[41053]= 618347408;
assign addr[41054]= 470399716;
assign addr[41055]= 320065829;
assign addr[41056]= 168108346;
assign addr[41057]= 15298099;
assign addr[41058]= -137589750;
assign addr[41059]= -289779648;
assign addr[41060]= -440499581;
assign addr[41061]= -588984994;
assign addr[41062]= -734482665;
assign addr[41063]= -876254528;
assign addr[41064]= -1013581418;
assign addr[41065]= -1145766716;
assign addr[41066]= -1272139887;
assign addr[41067]= -1392059879;
assign addr[41068]= -1504918373;
assign addr[41069]= -1610142873;
assign addr[41070]= -1707199606;
assign addr[41071]= -1795596234;
assign addr[41072]= -1874884346;
assign addr[41073]= -1944661739;
assign addr[41074]= -2004574453;
assign addr[41075]= -2054318569;
assign addr[41076]= -2093641749;
assign addr[41077]= -2122344521;
assign addr[41078]= -2140281282;
assign addr[41079]= -2147361045;
assign addr[41080]= -2143547897;
assign addr[41081]= -2128861181;
assign addr[41082]= -2103375398;
assign addr[41083]= -2067219829;
assign addr[41084]= -2020577882;
assign addr[41085]= -1963686155;
assign addr[41086]= -1896833245;
assign addr[41087]= -1820358275;
assign addr[41088]= -1734649179;
assign addr[41089]= -1640140734;
assign addr[41090]= -1537312353;
assign addr[41091]= -1426685652;
assign addr[41092]= -1308821808;
assign addr[41093]= -1184318708;
assign addr[41094]= -1053807919;
assign addr[41095]= -917951481;
assign addr[41096]= -777438554;
assign addr[41097]= -632981917;
assign addr[41098]= -485314355;
assign addr[41099]= -335184940;
assign addr[41100]= -183355234;
assign addr[41101]= -30595422;
assign addr[41102]= 122319591;
assign addr[41103]= 274614114;
assign addr[41104]= 425515602;
assign addr[41105]= 574258580;
assign addr[41106]= 720088517;
assign addr[41107]= 862265664;
assign addr[41108]= 1000068799;
assign addr[41109]= 1132798888;
assign addr[41110]= 1259782632;
assign addr[41111]= 1380375881;
assign addr[41112]= 1493966902;
assign addr[41113]= 1599979481;
assign addr[41114]= 1697875851;
assign addr[41115]= 1787159411;
assign addr[41116]= 1867377253;
assign addr[41117]= 1938122457;
assign addr[41118]= 1999036154;
assign addr[41119]= 2049809346;
assign addr[41120]= 2090184478;
assign addr[41121]= 2119956737;
assign addr[41122]= 2138975100;
assign addr[41123]= 2147143090;
assign addr[41124]= 2144419275;
assign addr[41125]= 2130817471;
assign addr[41126]= 2106406677;
assign addr[41127]= 2071310720;
assign addr[41128]= 2025707632;
assign addr[41129]= 1969828744;
assign addr[41130]= 1903957513;
assign addr[41131]= 1828428082;
assign addr[41132]= 1743623590;
assign addr[41133]= 1649974225;
assign addr[41134]= 1547955041;
assign addr[41135]= 1438083551;
assign addr[41136]= 1320917099;
assign addr[41137]= 1197050035;
assign addr[41138]= 1067110699;
assign addr[41139]= 931758235;
assign addr[41140]= 791679244;
assign addr[41141]= 647584304;
assign addr[41142]= 500204365;
assign addr[41143]= 350287041;
assign addr[41144]= 198592817;
assign addr[41145]= 45891193;
assign addr[41146]= -107043224;
assign addr[41147]= -259434643;
assign addr[41148]= -410510029;
assign addr[41149]= -559503022;
assign addr[41150]= -705657826;
assign addr[41151]= -848233042;
assign addr[41152]= -986505429;
assign addr[41153]= -1119773573;
assign addr[41154]= -1247361445;
assign addr[41155]= -1368621831;
assign addr[41156]= -1482939614;
assign addr[41157]= -1589734894;
assign addr[41158]= -1688465931;
assign addr[41159]= -1778631892;
assign addr[41160]= -1859775393;
assign addr[41161]= -1931484818;
assign addr[41162]= -1993396407;
assign addr[41163]= -2045196100;
assign addr[41164]= -2086621133;
assign addr[41165]= -2117461370;
assign addr[41166]= -2137560369;
assign addr[41167]= -2146816171;
assign addr[41168]= -2145181827;
assign addr[41169]= -2132665626;
assign addr[41170]= -2109331059;
assign addr[41171]= -2075296495;
assign addr[41172]= -2030734582;
assign addr[41173]= -1975871368;
assign addr[41174]= -1910985158;
assign addr[41175]= -1836405100;
assign addr[41176]= -1752509516;
assign addr[41177]= -1659723983;
assign addr[41178]= -1558519173;
assign addr[41179]= -1449408469;
assign addr[41180]= -1332945355;
assign addr[41181]= -1209720613;
assign addr[41182]= -1080359326;
assign addr[41183]= -945517704;
assign addr[41184]= -805879757;
assign addr[41185]= -662153826;
assign addr[41186]= -515068990;
assign addr[41187]= -365371365;
assign addr[41188]= -213820322;
assign addr[41189]= -61184634;
assign addr[41190]= 91761426;
assign addr[41191]= 244242007;
assign addr[41192]= 395483624;
assign addr[41193]= 544719071;
assign addr[41194]= 691191324;
assign addr[41195]= 834157373;
assign addr[41196]= 972891995;
assign addr[41197]= 1106691431;
assign addr[41198]= 1234876957;
assign addr[41199]= 1356798326;
assign addr[41200]= 1471837070;
assign addr[41201]= 1579409630;
assign addr[41202]= 1678970324;
assign addr[41203]= 1770014111;
assign addr[41204]= 1852079154;
assign addr[41205]= 1924749160;
assign addr[41206]= 1987655498;
assign addr[41207]= 2040479063;
assign addr[41208]= 2082951896;
assign addr[41209]= 2114858546;
assign addr[41210]= 2136037160;
assign addr[41211]= 2146380306;
assign addr[41212]= 2145835515;
assign addr[41213]= 2134405552;
assign addr[41214]= 2112148396;
assign addr[41215]= 2079176953;
assign addr[41216]= 2035658475;
assign addr[41217]= 1981813720;
assign addr[41218]= 1917915825;
assign addr[41219]= 1844288924;
assign addr[41220]= 1761306505;
assign addr[41221]= 1669389513;
assign addr[41222]= 1569004214;
assign addr[41223]= 1460659832;
assign addr[41224]= 1344905966;
assign addr[41225]= 1222329801;
assign addr[41226]= 1093553126;
assign addr[41227]= 959229189;
assign addr[41228]= 820039373;
assign addr[41229]= 676689746;
assign addr[41230]= 529907477;
assign addr[41231]= 380437148;
assign addr[41232]= 229036977;
assign addr[41233]= 76474970;
assign addr[41234]= -76474970;
assign addr[41235]= -229036977;
assign addr[41236]= -380437148;
assign addr[41237]= -529907477;
assign addr[41238]= -676689746;
assign addr[41239]= -820039373;
assign addr[41240]= -959229189;
assign addr[41241]= -1093553126;
assign addr[41242]= -1222329801;
assign addr[41243]= -1344905966;
assign addr[41244]= -1460659832;
assign addr[41245]= -1569004214;
assign addr[41246]= -1669389513;
assign addr[41247]= -1761306505;
assign addr[41248]= -1844288924;
assign addr[41249]= -1917915825;
assign addr[41250]= -1981813720;
assign addr[41251]= -2035658475;
assign addr[41252]= -2079176953;
assign addr[41253]= -2112148396;
assign addr[41254]= -2134405552;
assign addr[41255]= -2145835515;
assign addr[41256]= -2146380306;
assign addr[41257]= -2136037160;
assign addr[41258]= -2114858546;
assign addr[41259]= -2082951896;
assign addr[41260]= -2040479063;
assign addr[41261]= -1987655498;
assign addr[41262]= -1924749160;
assign addr[41263]= -1852079154;
assign addr[41264]= -1770014111;
assign addr[41265]= -1678970324;
assign addr[41266]= -1579409630;
assign addr[41267]= -1471837070;
assign addr[41268]= -1356798326;
assign addr[41269]= -1234876957;
assign addr[41270]= -1106691431;
assign addr[41271]= -972891995;
assign addr[41272]= -834157373;
assign addr[41273]= -691191324;
assign addr[41274]= -544719071;
assign addr[41275]= -395483624;
assign addr[41276]= -244242007;
assign addr[41277]= -91761426;
assign addr[41278]= 61184634;
assign addr[41279]= 213820322;
assign addr[41280]= 365371365;
assign addr[41281]= 515068990;
assign addr[41282]= 662153826;
assign addr[41283]= 805879757;
assign addr[41284]= 945517704;
assign addr[41285]= 1080359326;
assign addr[41286]= 1209720613;
assign addr[41287]= 1332945355;
assign addr[41288]= 1449408469;
assign addr[41289]= 1558519173;
assign addr[41290]= 1659723983;
assign addr[41291]= 1752509516;
assign addr[41292]= 1836405100;
assign addr[41293]= 1910985158;
assign addr[41294]= 1975871368;
assign addr[41295]= 2030734582;
assign addr[41296]= 2075296495;
assign addr[41297]= 2109331059;
assign addr[41298]= 2132665626;
assign addr[41299]= 2145181827;
assign addr[41300]= 2146816171;
assign addr[41301]= 2137560369;
assign addr[41302]= 2117461370;
assign addr[41303]= 2086621133;
assign addr[41304]= 2045196100;
assign addr[41305]= 1993396407;
assign addr[41306]= 1931484818;
assign addr[41307]= 1859775393;
assign addr[41308]= 1778631892;
assign addr[41309]= 1688465931;
assign addr[41310]= 1589734894;
assign addr[41311]= 1482939614;
assign addr[41312]= 1368621831;
assign addr[41313]= 1247361445;
assign addr[41314]= 1119773573;
assign addr[41315]= 986505429;
assign addr[41316]= 848233042;
assign addr[41317]= 705657826;
assign addr[41318]= 559503022;
assign addr[41319]= 410510029;
assign addr[41320]= 259434643;
assign addr[41321]= 107043224;
assign addr[41322]= -45891193;
assign addr[41323]= -198592817;
assign addr[41324]= -350287041;
assign addr[41325]= -500204365;
assign addr[41326]= -647584304;
assign addr[41327]= -791679244;
assign addr[41328]= -931758235;
assign addr[41329]= -1067110699;
assign addr[41330]= -1197050035;
assign addr[41331]= -1320917099;
assign addr[41332]= -1438083551;
assign addr[41333]= -1547955041;
assign addr[41334]= -1649974225;
assign addr[41335]= -1743623590;
assign addr[41336]= -1828428082;
assign addr[41337]= -1903957513;
assign addr[41338]= -1969828744;
assign addr[41339]= -2025707632;
assign addr[41340]= -2071310720;
assign addr[41341]= -2106406677;
assign addr[41342]= -2130817471;
assign addr[41343]= -2144419275;
assign addr[41344]= -2147143090;
assign addr[41345]= -2138975100;
assign addr[41346]= -2119956737;
assign addr[41347]= -2090184478;
assign addr[41348]= -2049809346;
assign addr[41349]= -1999036154;
assign addr[41350]= -1938122457;
assign addr[41351]= -1867377253;
assign addr[41352]= -1787159411;
assign addr[41353]= -1697875851;
assign addr[41354]= -1599979481;
assign addr[41355]= -1493966902;
assign addr[41356]= -1380375881;
assign addr[41357]= -1259782632;
assign addr[41358]= -1132798888;
assign addr[41359]= -1000068799;
assign addr[41360]= -862265664;
assign addr[41361]= -720088517;
assign addr[41362]= -574258580;
assign addr[41363]= -425515602;
assign addr[41364]= -274614114;
assign addr[41365]= -122319591;
assign addr[41366]= 30595422;
assign addr[41367]= 183355234;
assign addr[41368]= 335184940;
assign addr[41369]= 485314355;
assign addr[41370]= 632981917;
assign addr[41371]= 777438554;
assign addr[41372]= 917951481;
assign addr[41373]= 1053807919;
assign addr[41374]= 1184318708;
assign addr[41375]= 1308821808;
assign addr[41376]= 1426685652;
assign addr[41377]= 1537312353;
assign addr[41378]= 1640140734;
assign addr[41379]= 1734649179;
assign addr[41380]= 1820358275;
assign addr[41381]= 1896833245;
assign addr[41382]= 1963686155;
assign addr[41383]= 2020577882;
assign addr[41384]= 2067219829;
assign addr[41385]= 2103375398;
assign addr[41386]= 2128861181;
assign addr[41387]= 2143547897;
assign addr[41388]= 2147361045;
assign addr[41389]= 2140281282;
assign addr[41390]= 2122344521;
assign addr[41391]= 2093641749;
assign addr[41392]= 2054318569;
assign addr[41393]= 2004574453;
assign addr[41394]= 1944661739;
assign addr[41395]= 1874884346;
assign addr[41396]= 1795596234;
assign addr[41397]= 1707199606;
assign addr[41398]= 1610142873;
assign addr[41399]= 1504918373;
assign addr[41400]= 1392059879;
assign addr[41401]= 1272139887;
assign addr[41402]= 1145766716;
assign addr[41403]= 1013581418;
assign addr[41404]= 876254528;
assign addr[41405]= 734482665;
assign addr[41406]= 588984994;
assign addr[41407]= 440499581;
assign addr[41408]= 289779648;
assign addr[41409]= 137589750;
assign addr[41410]= -15298099;
assign addr[41411]= -168108346;
assign addr[41412]= -320065829;
assign addr[41413]= -470399716;
assign addr[41414]= -618347408;
assign addr[41415]= -763158411;
assign addr[41416]= -904098143;
assign addr[41417]= -1040451659;
assign addr[41418]= -1171527280;
assign addr[41419]= -1296660098;
assign addr[41420]= -1415215352;
assign addr[41421]= -1526591649;
assign addr[41422]= -1630224009;
assign addr[41423]= -1725586737;
assign addr[41424]= -1812196087;
assign addr[41425]= -1889612716;
assign addr[41426]= -1957443913;
assign addr[41427]= -2015345591;
assign addr[41428]= -2063024031;
assign addr[41429]= -2100237377;
assign addr[41430]= -2126796855;
assign addr[41431]= -2142567738;
assign addr[41432]= -2147470025;
assign addr[41433]= -2141478848;
assign addr[41434]= -2124624598;
assign addr[41435]= -2096992772;
assign addr[41436]= -2058723538;
assign addr[41437]= -2010011024;
assign addr[41438]= -1951102334;
assign addr[41439]= -1882296293;
assign addr[41440]= -1803941934;
assign addr[41441]= -1716436725;
assign addr[41442]= -1620224553;
assign addr[41443]= -1515793473;
assign addr[41444]= -1403673233;
assign addr[41445]= -1284432584;
assign addr[41446]= -1158676398;
assign addr[41447]= -1027042599;
assign addr[41448]= -890198924;
assign addr[41449]= -748839539;
assign addr[41450]= -603681519;
assign addr[41451]= -455461206;
assign addr[41452]= -304930476;
assign addr[41453]= -152852926;
assign addr[41454]= 0;
assign addr[41455]= 152852926;
assign addr[41456]= 304930476;
assign addr[41457]= 455461206;
assign addr[41458]= 603681519;
assign addr[41459]= 748839539;
assign addr[41460]= 890198924;
assign addr[41461]= 1027042599;
assign addr[41462]= 1158676398;
assign addr[41463]= 1284432584;
assign addr[41464]= 1403673233;
assign addr[41465]= 1515793473;
assign addr[41466]= 1620224553;
assign addr[41467]= 1716436725;
assign addr[41468]= 1803941934;
assign addr[41469]= 1882296293;
assign addr[41470]= 1951102334;
assign addr[41471]= 2010011024;
assign addr[41472]= 2058723538;
assign addr[41473]= 2096992772;
assign addr[41474]= 2124624598;
assign addr[41475]= 2141478848;
assign addr[41476]= 2147470025;
assign addr[41477]= 2142567738;
assign addr[41478]= 2126796855;
assign addr[41479]= 2100237377;
assign addr[41480]= 2063024031;
assign addr[41481]= 2015345591;
assign addr[41482]= 1957443913;
assign addr[41483]= 1889612716;
assign addr[41484]= 1812196087;
assign addr[41485]= 1725586737;
assign addr[41486]= 1630224009;
assign addr[41487]= 1526591649;
assign addr[41488]= 1415215352;
assign addr[41489]= 1296660098;
assign addr[41490]= 1171527280;
assign addr[41491]= 1040451659;
assign addr[41492]= 904098143;
assign addr[41493]= 763158411;
assign addr[41494]= 618347408;
assign addr[41495]= 470399716;
assign addr[41496]= 320065829;
assign addr[41497]= 168108346;
assign addr[41498]= 15298099;
assign addr[41499]= -137589750;
assign addr[41500]= -289779648;
assign addr[41501]= -440499581;
assign addr[41502]= -588984994;
assign addr[41503]= -734482665;
assign addr[41504]= -876254528;
assign addr[41505]= -1013581418;
assign addr[41506]= -1145766716;
assign addr[41507]= -1272139887;
assign addr[41508]= -1392059879;
assign addr[41509]= -1504918373;
assign addr[41510]= -1610142873;
assign addr[41511]= -1707199606;
assign addr[41512]= -1795596234;
assign addr[41513]= -1874884346;
assign addr[41514]= -1944661739;
assign addr[41515]= -2004574453;
assign addr[41516]= -2054318569;
assign addr[41517]= -2093641749;
assign addr[41518]= -2122344521;
assign addr[41519]= -2140281282;
assign addr[41520]= -2147361045;
assign addr[41521]= -2143547897;
assign addr[41522]= -2128861181;
assign addr[41523]= -2103375398;
assign addr[41524]= -2067219829;
assign addr[41525]= -2020577882;
assign addr[41526]= -1963686155;
assign addr[41527]= -1896833245;
assign addr[41528]= -1820358275;
assign addr[41529]= -1734649179;
assign addr[41530]= -1640140734;
assign addr[41531]= -1537312353;
assign addr[41532]= -1426685652;
assign addr[41533]= -1308821808;
assign addr[41534]= -1184318708;
assign addr[41535]= -1053807919;
assign addr[41536]= -917951481;
assign addr[41537]= -777438554;
assign addr[41538]= -632981917;
assign addr[41539]= -485314355;
assign addr[41540]= -335184940;
assign addr[41541]= -183355234;
assign addr[41542]= -30595422;
assign addr[41543]= 122319591;
assign addr[41544]= 274614114;
assign addr[41545]= 425515602;
assign addr[41546]= 574258580;
assign addr[41547]= 720088517;
assign addr[41548]= 862265664;
assign addr[41549]= 1000068799;
assign addr[41550]= 1132798888;
assign addr[41551]= 1259782632;
assign addr[41552]= 1380375881;
assign addr[41553]= 1493966902;
assign addr[41554]= 1599979481;
assign addr[41555]= 1697875851;
assign addr[41556]= 1787159411;
assign addr[41557]= 1867377253;
assign addr[41558]= 1938122457;
assign addr[41559]= 1999036154;
assign addr[41560]= 2049809346;
assign addr[41561]= 2090184478;
assign addr[41562]= 2119956737;
assign addr[41563]= 2138975100;
assign addr[41564]= 2147143090;
assign addr[41565]= 2144419275;
assign addr[41566]= 2130817471;
assign addr[41567]= 2106406677;
assign addr[41568]= 2071310720;
assign addr[41569]= 2025707632;
assign addr[41570]= 1969828744;
assign addr[41571]= 1903957513;
assign addr[41572]= 1828428082;
assign addr[41573]= 1743623590;
assign addr[41574]= 1649974225;
assign addr[41575]= 1547955041;
assign addr[41576]= 1438083551;
assign addr[41577]= 1320917099;
assign addr[41578]= 1197050035;
assign addr[41579]= 1067110699;
assign addr[41580]= 931758235;
assign addr[41581]= 791679244;
assign addr[41582]= 647584304;
assign addr[41583]= 500204365;
assign addr[41584]= 350287041;
assign addr[41585]= 198592817;
assign addr[41586]= 45891193;
assign addr[41587]= -107043224;
assign addr[41588]= -259434643;
assign addr[41589]= -410510029;
assign addr[41590]= -559503022;
assign addr[41591]= -705657826;
assign addr[41592]= -848233042;
assign addr[41593]= -986505429;
assign addr[41594]= -1119773573;
assign addr[41595]= -1247361445;
assign addr[41596]= -1368621831;
assign addr[41597]= -1482939614;
assign addr[41598]= -1589734894;
assign addr[41599]= -1688465931;
assign addr[41600]= -1778631892;
assign addr[41601]= -1859775393;
assign addr[41602]= -1931484818;
assign addr[41603]= -1993396407;
assign addr[41604]= -2045196100;
assign addr[41605]= -2086621133;
assign addr[41606]= -2117461370;
assign addr[41607]= -2137560369;
assign addr[41608]= -2146816171;
assign addr[41609]= -2145181827;
assign addr[41610]= -2132665626;
assign addr[41611]= -2109331059;
assign addr[41612]= -2075296495;
assign addr[41613]= -2030734582;
assign addr[41614]= -1975871368;
assign addr[41615]= -1910985158;
assign addr[41616]= -1836405100;
assign addr[41617]= -1752509516;
assign addr[41618]= -1659723983;
assign addr[41619]= -1558519173;
assign addr[41620]= -1449408469;
assign addr[41621]= -1332945355;
assign addr[41622]= -1209720613;
assign addr[41623]= -1080359326;
assign addr[41624]= -945517704;
assign addr[41625]= -805879757;
assign addr[41626]= -662153826;
assign addr[41627]= -515068990;
assign addr[41628]= -365371365;
assign addr[41629]= -213820322;
assign addr[41630]= -61184634;
assign addr[41631]= 91761426;
assign addr[41632]= 244242007;
assign addr[41633]= 395483624;
assign addr[41634]= 544719071;
assign addr[41635]= 691191324;
assign addr[41636]= 834157373;
assign addr[41637]= 972891995;
assign addr[41638]= 1106691431;
assign addr[41639]= 1234876957;
assign addr[41640]= 1356798326;
assign addr[41641]= 1471837070;
assign addr[41642]= 1579409630;
assign addr[41643]= 1678970324;
assign addr[41644]= 1770014111;
assign addr[41645]= 1852079154;
assign addr[41646]= 1924749160;
assign addr[41647]= 1987655498;
assign addr[41648]= 2040479063;
assign addr[41649]= 2082951896;
assign addr[41650]= 2114858546;
assign addr[41651]= 2136037160;
assign addr[41652]= 2146380306;
assign addr[41653]= 2145835515;
assign addr[41654]= 2134405552;
assign addr[41655]= 2112148396;
assign addr[41656]= 2079176953;
assign addr[41657]= 2035658475;
assign addr[41658]= 1981813720;
assign addr[41659]= 1917915825;
assign addr[41660]= 1844288924;
assign addr[41661]= 1761306505;
assign addr[41662]= 1669389513;
assign addr[41663]= 1569004214;
assign addr[41664]= 1460659832;
assign addr[41665]= 1344905966;
assign addr[41666]= 1222329801;
assign addr[41667]= 1093553126;
assign addr[41668]= 959229189;
assign addr[41669]= 820039373;
assign addr[41670]= 676689746;
assign addr[41671]= 529907477;
assign addr[41672]= 380437148;
assign addr[41673]= 229036977;
assign addr[41674]= 76474970;
assign addr[41675]= -76474970;
assign addr[41676]= -229036977;
assign addr[41677]= -380437148;
assign addr[41678]= -529907477;
assign addr[41679]= -676689746;
assign addr[41680]= -820039373;
assign addr[41681]= -959229189;
assign addr[41682]= -1093553126;
assign addr[41683]= -1222329801;
assign addr[41684]= -1344905966;
assign addr[41685]= -1460659832;
assign addr[41686]= -1569004214;
assign addr[41687]= -1669389513;
assign addr[41688]= -1761306505;
assign addr[41689]= -1844288924;
assign addr[41690]= -1917915825;
assign addr[41691]= -1981813720;
assign addr[41692]= -2035658475;
assign addr[41693]= -2079176953;
assign addr[41694]= -2112148396;
assign addr[41695]= -2134405552;
assign addr[41696]= -2145835515;
assign addr[41697]= -2146380306;
assign addr[41698]= -2136037160;
assign addr[41699]= -2114858546;
assign addr[41700]= -2082951896;
assign addr[41701]= -2040479063;
assign addr[41702]= -1987655498;
assign addr[41703]= -1924749160;
assign addr[41704]= -1852079154;
assign addr[41705]= -1770014111;
assign addr[41706]= -1678970324;
assign addr[41707]= -1579409630;
assign addr[41708]= -1471837070;
assign addr[41709]= -1356798326;
assign addr[41710]= -1234876957;
assign addr[41711]= -1106691431;
assign addr[41712]= -972891995;
assign addr[41713]= -834157373;
assign addr[41714]= -691191324;
assign addr[41715]= -544719071;
assign addr[41716]= -395483624;
assign addr[41717]= -244242007;
assign addr[41718]= -91761426;
assign addr[41719]= 61184634;
assign addr[41720]= 213820322;
assign addr[41721]= 365371365;
assign addr[41722]= 515068990;
assign addr[41723]= 662153826;
assign addr[41724]= 805879757;
assign addr[41725]= 945517704;
assign addr[41726]= 1080359326;
assign addr[41727]= 1209720613;
assign addr[41728]= 1332945355;
assign addr[41729]= 1449408469;
assign addr[41730]= 1558519173;
assign addr[41731]= 1659723983;
assign addr[41732]= 1752509516;
assign addr[41733]= 1836405100;
assign addr[41734]= 1910985158;
assign addr[41735]= 1975871368;
assign addr[41736]= 2030734582;
assign addr[41737]= 2075296495;
assign addr[41738]= 2109331059;
assign addr[41739]= 2132665626;
assign addr[41740]= 2145181827;
assign addr[41741]= 2146816171;
assign addr[41742]= 2137560369;
assign addr[41743]= 2117461370;
assign addr[41744]= 2086621133;
assign addr[41745]= 2045196100;
assign addr[41746]= 1993396407;
assign addr[41747]= 1931484818;
assign addr[41748]= 1859775393;
assign addr[41749]= 1778631892;
assign addr[41750]= 1688465931;
assign addr[41751]= 1589734894;
assign addr[41752]= 1482939614;
assign addr[41753]= 1368621831;
assign addr[41754]= 1247361445;
assign addr[41755]= 1119773573;
assign addr[41756]= 986505429;
assign addr[41757]= 848233042;
assign addr[41758]= 705657826;
assign addr[41759]= 559503022;
assign addr[41760]= 410510029;
assign addr[41761]= 259434643;
assign addr[41762]= 107043224;
assign addr[41763]= -45891193;
assign addr[41764]= -198592817;
assign addr[41765]= -350287041;
assign addr[41766]= -500204365;
assign addr[41767]= -647584304;
assign addr[41768]= -791679244;
assign addr[41769]= -931758235;
assign addr[41770]= -1067110699;
assign addr[41771]= -1197050035;
assign addr[41772]= -1320917099;
assign addr[41773]= -1438083551;
assign addr[41774]= -1547955041;
assign addr[41775]= -1649974225;
assign addr[41776]= -1743623590;
assign addr[41777]= -1828428082;
assign addr[41778]= -1903957513;
assign addr[41779]= -1969828744;
assign addr[41780]= -2025707632;
assign addr[41781]= -2071310720;
assign addr[41782]= -2106406677;
assign addr[41783]= -2130817471;
assign addr[41784]= -2144419275;
assign addr[41785]= -2147143090;
assign addr[41786]= -2138975100;
assign addr[41787]= -2119956737;
assign addr[41788]= -2090184478;
assign addr[41789]= -2049809346;
assign addr[41790]= -1999036154;
assign addr[41791]= -1938122457;
assign addr[41792]= -1867377253;
assign addr[41793]= -1787159411;
assign addr[41794]= -1697875851;
assign addr[41795]= -1599979481;
assign addr[41796]= -1493966902;
assign addr[41797]= -1380375881;
assign addr[41798]= -1259782632;
assign addr[41799]= -1132798888;
assign addr[41800]= -1000068799;
assign addr[41801]= -862265664;
assign addr[41802]= -720088517;
assign addr[41803]= -574258580;
assign addr[41804]= -425515602;
assign addr[41805]= -274614114;
assign addr[41806]= -122319591;
assign addr[41807]= 30595422;
assign addr[41808]= 183355234;
assign addr[41809]= 335184940;
assign addr[41810]= 485314355;
assign addr[41811]= 632981917;
assign addr[41812]= 777438554;
assign addr[41813]= 917951481;
assign addr[41814]= 1053807919;
assign addr[41815]= 1184318708;
assign addr[41816]= 1308821808;
assign addr[41817]= 1426685652;
assign addr[41818]= 1537312353;
assign addr[41819]= 1640140734;
assign addr[41820]= 1734649179;
assign addr[41821]= 1820358275;
assign addr[41822]= 1896833245;
assign addr[41823]= 1963686155;
assign addr[41824]= 2020577882;
assign addr[41825]= 2067219829;
assign addr[41826]= 2103375398;
assign addr[41827]= 2128861181;
assign addr[41828]= 2143547897;
assign addr[41829]= 2147361045;
assign addr[41830]= 2140281282;
assign addr[41831]= 2122344521;
assign addr[41832]= 2093641749;
assign addr[41833]= 2054318569;
assign addr[41834]= 2004574453;
assign addr[41835]= 1944661739;
assign addr[41836]= 1874884346;
assign addr[41837]= 1795596234;
assign addr[41838]= 1707199606;
assign addr[41839]= 1610142873;
assign addr[41840]= 1504918373;
assign addr[41841]= 1392059879;
assign addr[41842]= 1272139887;
assign addr[41843]= 1145766716;
assign addr[41844]= 1013581418;
assign addr[41845]= 876254528;
assign addr[41846]= 734482665;
assign addr[41847]= 588984994;
assign addr[41848]= 440499581;
assign addr[41849]= 289779648;
assign addr[41850]= 137589750;
assign addr[41851]= -15298099;
assign addr[41852]= -168108346;
assign addr[41853]= -320065829;
assign addr[41854]= -470399716;
assign addr[41855]= -618347408;
assign addr[41856]= -763158411;
assign addr[41857]= -904098143;
assign addr[41858]= -1040451659;
assign addr[41859]= -1171527280;
assign addr[41860]= -1296660098;
assign addr[41861]= -1415215352;
assign addr[41862]= -1526591649;
assign addr[41863]= -1630224009;
assign addr[41864]= -1725586737;
assign addr[41865]= -1812196087;
assign addr[41866]= -1889612716;
assign addr[41867]= -1957443913;
assign addr[41868]= -2015345591;
assign addr[41869]= -2063024031;
assign addr[41870]= -2100237377;
assign addr[41871]= -2126796855;
assign addr[41872]= -2142567738;
assign addr[41873]= -2147470025;
assign addr[41874]= -2141478848;
assign addr[41875]= -2124624598;
assign addr[41876]= -2096992772;
assign addr[41877]= -2058723538;
assign addr[41878]= -2010011024;
assign addr[41879]= -1951102334;
assign addr[41880]= -1882296293;
assign addr[41881]= -1803941934;
assign addr[41882]= -1716436725;
assign addr[41883]= -1620224553;
assign addr[41884]= -1515793473;
assign addr[41885]= -1403673233;
assign addr[41886]= -1284432584;
assign addr[41887]= -1158676398;
assign addr[41888]= -1027042599;
assign addr[41889]= -890198924;
assign addr[41890]= -748839539;
assign addr[41891]= -603681519;
assign addr[41892]= -455461206;
assign addr[41893]= -304930476;
assign addr[41894]= -152852926;
assign addr[41895]= 0;
assign addr[41896]= 152852926;
assign addr[41897]= 304930476;
assign addr[41898]= 455461206;
assign addr[41899]= 603681519;
assign addr[41900]= 748839539;
assign addr[41901]= 890198924;
assign addr[41902]= 1027042599;
assign addr[41903]= 1158676398;
assign addr[41904]= 1284432584;
assign addr[41905]= 1403673233;
assign addr[41906]= 1515793473;
assign addr[41907]= 1620224553;
assign addr[41908]= 1716436725;
assign addr[41909]= 1803941934;
assign addr[41910]= 1882296293;
assign addr[41911]= 1951102334;
assign addr[41912]= 2010011024;
assign addr[41913]= 2058723538;
assign addr[41914]= 2096992772;
assign addr[41915]= 2124624598;
assign addr[41916]= 2141478848;
assign addr[41917]= 2147470025;
assign addr[41918]= 2142567738;
assign addr[41919]= 2126796855;
assign addr[41920]= 2100237377;
assign addr[41921]= 2063024031;
assign addr[41922]= 2015345591;
assign addr[41923]= 1957443913;
assign addr[41924]= 1889612716;
assign addr[41925]= 1812196087;
assign addr[41926]= 1725586737;
assign addr[41927]= 1630224009;
assign addr[41928]= 1526591649;
assign addr[41929]= 1415215352;
assign addr[41930]= 1296660098;
assign addr[41931]= 1171527280;
assign addr[41932]= 1040451659;
assign addr[41933]= 904098143;
assign addr[41934]= 763158411;
assign addr[41935]= 618347408;
assign addr[41936]= 470399716;
assign addr[41937]= 320065829;
assign addr[41938]= 168108346;
assign addr[41939]= 15298099;
assign addr[41940]= -137589750;
assign addr[41941]= -289779648;
assign addr[41942]= -440499581;
assign addr[41943]= -588984994;
assign addr[41944]= -734482665;
assign addr[41945]= -876254528;
assign addr[41946]= -1013581418;
assign addr[41947]= -1145766716;
assign addr[41948]= -1272139887;
assign addr[41949]= -1392059879;
assign addr[41950]= -1504918373;
assign addr[41951]= -1610142873;
assign addr[41952]= -1707199606;
assign addr[41953]= -1795596234;
assign addr[41954]= -1874884346;
assign addr[41955]= -1944661739;
assign addr[41956]= -2004574453;
assign addr[41957]= -2054318569;
assign addr[41958]= -2093641749;
assign addr[41959]= -2122344521;
assign addr[41960]= -2140281282;
assign addr[41961]= -2147361045;
assign addr[41962]= -2143547897;
assign addr[41963]= -2128861181;
assign addr[41964]= -2103375398;
assign addr[41965]= -2067219829;
assign addr[41966]= -2020577882;
assign addr[41967]= -1963686155;
assign addr[41968]= -1896833245;
assign addr[41969]= -1820358275;
assign addr[41970]= -1734649179;
assign addr[41971]= -1640140734;
assign addr[41972]= -1537312353;
assign addr[41973]= -1426685652;
assign addr[41974]= -1308821808;
assign addr[41975]= -1184318708;
assign addr[41976]= -1053807919;
assign addr[41977]= -917951481;
assign addr[41978]= -777438554;
assign addr[41979]= -632981917;
assign addr[41980]= -485314355;
assign addr[41981]= -335184940;
assign addr[41982]= -183355234;
assign addr[41983]= -30595422;
assign addr[41984]= 122319591;
assign addr[41985]= 274614114;
assign addr[41986]= 425515602;
assign addr[41987]= 574258580;
assign addr[41988]= 720088517;
assign addr[41989]= 862265664;
assign addr[41990]= 1000068799;
assign addr[41991]= 1132798888;
assign addr[41992]= 1259782632;
assign addr[41993]= 1380375881;
assign addr[41994]= 1493966902;
assign addr[41995]= 1599979481;
assign addr[41996]= 1697875851;
assign addr[41997]= 1787159411;
assign addr[41998]= 1867377253;
assign addr[41999]= 1938122457;
assign addr[42000]= 1999036154;
assign addr[42001]= 2049809346;
assign addr[42002]= 2090184478;
assign addr[42003]= 2119956737;
assign addr[42004]= 2138975100;
assign addr[42005]= 2147143090;
assign addr[42006]= 2144419275;
assign addr[42007]= 2130817471;
assign addr[42008]= 2106406677;
assign addr[42009]= 2071310720;
assign addr[42010]= 2025707632;
assign addr[42011]= 1969828744;
assign addr[42012]= 1903957513;
assign addr[42013]= 1828428082;
assign addr[42014]= 1743623590;
assign addr[42015]= 1649974225;
assign addr[42016]= 1547955041;
assign addr[42017]= 1438083551;
assign addr[42018]= 1320917099;
assign addr[42019]= 1197050035;
assign addr[42020]= 1067110699;
assign addr[42021]= 931758235;
assign addr[42022]= 791679244;
assign addr[42023]= 647584304;
assign addr[42024]= 500204365;
assign addr[42025]= 350287041;
assign addr[42026]= 198592817;
assign addr[42027]= 45891193;
assign addr[42028]= -107043224;
assign addr[42029]= -259434643;
assign addr[42030]= -410510029;
assign addr[42031]= -559503022;
assign addr[42032]= -705657826;
assign addr[42033]= -848233042;
assign addr[42034]= -986505429;
assign addr[42035]= -1119773573;
assign addr[42036]= -1247361445;
assign addr[42037]= -1368621831;
assign addr[42038]= -1482939614;
assign addr[42039]= -1589734894;
assign addr[42040]= -1688465931;
assign addr[42041]= -1778631892;
assign addr[42042]= -1859775393;
assign addr[42043]= -1931484818;
assign addr[42044]= -1993396407;
assign addr[42045]= -2045196100;
assign addr[42046]= -2086621133;
assign addr[42047]= -2117461370;
assign addr[42048]= -2137560369;
assign addr[42049]= -2146816171;
assign addr[42050]= -2145181827;
assign addr[42051]= -2132665626;
assign addr[42052]= -2109331059;
assign addr[42053]= -2075296495;
assign addr[42054]= -2030734582;
assign addr[42055]= -1975871368;
assign addr[42056]= -1910985158;
assign addr[42057]= -1836405100;
assign addr[42058]= -1752509516;
assign addr[42059]= -1659723983;
assign addr[42060]= -1558519173;
assign addr[42061]= -1449408469;
assign addr[42062]= -1332945355;
assign addr[42063]= -1209720613;
assign addr[42064]= -1080359326;
assign addr[42065]= -945517704;
assign addr[42066]= -805879757;
assign addr[42067]= -662153826;
assign addr[42068]= -515068990;
assign addr[42069]= -365371365;
assign addr[42070]= -213820322;
assign addr[42071]= -61184634;
assign addr[42072]= 91761426;
assign addr[42073]= 244242007;
assign addr[42074]= 395483624;
assign addr[42075]= 544719071;
assign addr[42076]= 691191324;
assign addr[42077]= 834157373;
assign addr[42078]= 972891995;
assign addr[42079]= 1106691431;
assign addr[42080]= 1234876957;
assign addr[42081]= 1356798326;
assign addr[42082]= 1471837070;
assign addr[42083]= 1579409630;
assign addr[42084]= 1678970324;
assign addr[42085]= 1770014111;
assign addr[42086]= 1852079154;
assign addr[42087]= 1924749160;
assign addr[42088]= 1987655498;
assign addr[42089]= 2040479063;
assign addr[42090]= 2082951896;
assign addr[42091]= 2114858546;
assign addr[42092]= 2136037160;
assign addr[42093]= 2146380306;
assign addr[42094]= 2145835515;
assign addr[42095]= 2134405552;
assign addr[42096]= 2112148396;
assign addr[42097]= 2079176953;
assign addr[42098]= 2035658475;
assign addr[42099]= 1981813720;
assign addr[42100]= 1917915825;
assign addr[42101]= 1844288924;
assign addr[42102]= 1761306505;
assign addr[42103]= 1669389513;
assign addr[42104]= 1569004214;
assign addr[42105]= 1460659832;
assign addr[42106]= 1344905966;
assign addr[42107]= 1222329801;
assign addr[42108]= 1093553126;
assign addr[42109]= 959229189;
assign addr[42110]= 820039373;
assign addr[42111]= 676689746;
assign addr[42112]= 529907477;
assign addr[42113]= 380437148;
assign addr[42114]= 229036977;
assign addr[42115]= 76474970;
assign addr[42116]= -76474970;
assign addr[42117]= -229036977;
assign addr[42118]= -380437148;
assign addr[42119]= -529907477;
assign addr[42120]= -676689746;
assign addr[42121]= -820039373;
assign addr[42122]= -959229189;
assign addr[42123]= -1093553126;
assign addr[42124]= -1222329801;
assign addr[42125]= -1344905966;
assign addr[42126]= -1460659832;
assign addr[42127]= -1569004214;
assign addr[42128]= -1669389513;
assign addr[42129]= -1761306505;
assign addr[42130]= -1844288924;
assign addr[42131]= -1917915825;
assign addr[42132]= -1981813720;
assign addr[42133]= -2035658475;
assign addr[42134]= -2079176953;
assign addr[42135]= -2112148396;
assign addr[42136]= -2134405552;
assign addr[42137]= -2145835515;
assign addr[42138]= -2146380306;
assign addr[42139]= -2136037160;
assign addr[42140]= -2114858546;
assign addr[42141]= -2082951896;
assign addr[42142]= -2040479063;
assign addr[42143]= -1987655498;
assign addr[42144]= -1924749160;
assign addr[42145]= -1852079154;
assign addr[42146]= -1770014111;
assign addr[42147]= -1678970324;
assign addr[42148]= -1579409630;
assign addr[42149]= -1471837070;
assign addr[42150]= -1356798326;
assign addr[42151]= -1234876957;
assign addr[42152]= -1106691431;
assign addr[42153]= -972891995;
assign addr[42154]= -834157373;
assign addr[42155]= -691191324;
assign addr[42156]= -544719071;
assign addr[42157]= -395483624;
assign addr[42158]= -244242007;
assign addr[42159]= -91761426;
assign addr[42160]= 61184634;
assign addr[42161]= 213820322;
assign addr[42162]= 365371365;
assign addr[42163]= 515068990;
assign addr[42164]= 662153826;
assign addr[42165]= 805879757;
assign addr[42166]= 945517704;
assign addr[42167]= 1080359326;
assign addr[42168]= 1209720613;
assign addr[42169]= 1332945355;
assign addr[42170]= 1449408469;
assign addr[42171]= 1558519173;
assign addr[42172]= 1659723983;
assign addr[42173]= 1752509516;
assign addr[42174]= 1836405100;
assign addr[42175]= 1910985158;
assign addr[42176]= 1975871368;
assign addr[42177]= 2030734582;
assign addr[42178]= 2075296495;
assign addr[42179]= 2109331059;
assign addr[42180]= 2132665626;
assign addr[42181]= 2145181827;
assign addr[42182]= 2146816171;
assign addr[42183]= 2137560369;
assign addr[42184]= 2117461370;
assign addr[42185]= 2086621133;
assign addr[42186]= 2045196100;
assign addr[42187]= 1993396407;
assign addr[42188]= 1931484818;
assign addr[42189]= 1859775393;
assign addr[42190]= 1778631892;
assign addr[42191]= 1688465931;
assign addr[42192]= 1589734894;
assign addr[42193]= 1482939614;
assign addr[42194]= 1368621831;
assign addr[42195]= 1247361445;
assign addr[42196]= 1119773573;
assign addr[42197]= 986505429;
assign addr[42198]= 848233042;
assign addr[42199]= 705657826;
assign addr[42200]= 559503022;
assign addr[42201]= 410510029;
assign addr[42202]= 259434643;
assign addr[42203]= 107043224;
assign addr[42204]= -45891193;
assign addr[42205]= -198592817;
assign addr[42206]= -350287041;
assign addr[42207]= -500204365;
assign addr[42208]= -647584304;
assign addr[42209]= -791679244;
assign addr[42210]= -931758235;
assign addr[42211]= -1067110699;
assign addr[42212]= -1197050035;
assign addr[42213]= -1320917099;
assign addr[42214]= -1438083551;
assign addr[42215]= -1547955041;
assign addr[42216]= -1649974225;
assign addr[42217]= -1743623590;
assign addr[42218]= -1828428082;
assign addr[42219]= -1903957513;
assign addr[42220]= -1969828744;
assign addr[42221]= -2025707632;
assign addr[42222]= -2071310720;
assign addr[42223]= -2106406677;
assign addr[42224]= -2130817471;
assign addr[42225]= -2144419275;
assign addr[42226]= -2147143090;
assign addr[42227]= -2138975100;
assign addr[42228]= -2119956737;
assign addr[42229]= -2090184478;
assign addr[42230]= -2049809346;
assign addr[42231]= -1999036154;
assign addr[42232]= -1938122457;
assign addr[42233]= -1867377253;
assign addr[42234]= -1787159411;
assign addr[42235]= -1697875851;
assign addr[42236]= -1599979481;
assign addr[42237]= -1493966902;
assign addr[42238]= -1380375881;
assign addr[42239]= -1259782632;
assign addr[42240]= -1132798888;
assign addr[42241]= -1000068799;
assign addr[42242]= -862265664;
assign addr[42243]= -720088517;
assign addr[42244]= -574258580;
assign addr[42245]= -425515602;
assign addr[42246]= -274614114;
assign addr[42247]= -122319591;
assign addr[42248]= 30595422;
assign addr[42249]= 183355234;
assign addr[42250]= 335184940;
assign addr[42251]= 485314355;
assign addr[42252]= 632981917;
assign addr[42253]= 777438554;
assign addr[42254]= 917951481;
assign addr[42255]= 1053807919;
assign addr[42256]= 1184318708;
assign addr[42257]= 1308821808;
assign addr[42258]= 1426685652;
assign addr[42259]= 1537312353;
assign addr[42260]= 1640140734;
assign addr[42261]= 1734649179;
assign addr[42262]= 1820358275;
assign addr[42263]= 1896833245;
assign addr[42264]= 1963686155;
assign addr[42265]= 2020577882;
assign addr[42266]= 2067219829;
assign addr[42267]= 2103375398;
assign addr[42268]= 2128861181;
assign addr[42269]= 2143547897;
assign addr[42270]= 2147361045;
assign addr[42271]= 2140281282;
assign addr[42272]= 2122344521;
assign addr[42273]= 2093641749;
assign addr[42274]= 2054318569;
assign addr[42275]= 2004574453;
assign addr[42276]= 1944661739;
assign addr[42277]= 1874884346;
assign addr[42278]= 1795596234;
assign addr[42279]= 1707199606;
assign addr[42280]= 1610142873;
assign addr[42281]= 1504918373;
assign addr[42282]= 1392059879;
assign addr[42283]= 1272139887;
assign addr[42284]= 1145766716;
assign addr[42285]= 1013581418;
assign addr[42286]= 876254528;
assign addr[42287]= 734482665;
assign addr[42288]= 588984994;
assign addr[42289]= 440499581;
assign addr[42290]= 289779648;
assign addr[42291]= 137589750;
assign addr[42292]= -15298099;
assign addr[42293]= -168108346;
assign addr[42294]= -320065829;
assign addr[42295]= -470399716;
assign addr[42296]= -618347408;
assign addr[42297]= -763158411;
assign addr[42298]= -904098143;
assign addr[42299]= -1040451659;
assign addr[42300]= -1171527280;
assign addr[42301]= -1296660098;
assign addr[42302]= -1415215352;
assign addr[42303]= -1526591649;
assign addr[42304]= -1630224009;
assign addr[42305]= -1725586737;
assign addr[42306]= -1812196087;
assign addr[42307]= -1889612716;
assign addr[42308]= -1957443913;
assign addr[42309]= -2015345591;
assign addr[42310]= -2063024031;
assign addr[42311]= -2100237377;
assign addr[42312]= -2126796855;
assign addr[42313]= -2142567738;
assign addr[42314]= -2147470025;
assign addr[42315]= -2141478848;
assign addr[42316]= -2124624598;
assign addr[42317]= -2096992772;
assign addr[42318]= -2058723538;
assign addr[42319]= -2010011024;
assign addr[42320]= -1951102334;
assign addr[42321]= -1882296293;
assign addr[42322]= -1803941934;
assign addr[42323]= -1716436725;
assign addr[42324]= -1620224553;
assign addr[42325]= -1515793473;
assign addr[42326]= -1403673233;
assign addr[42327]= -1284432584;
assign addr[42328]= -1158676398;
assign addr[42329]= -1027042599;
assign addr[42330]= -890198924;
assign addr[42331]= -748839539;
assign addr[42332]= -603681519;
assign addr[42333]= -455461206;
assign addr[42334]= -304930476;
assign addr[42335]= -152852926;
assign addr[42336]= 0;
assign addr[42337]= 152852926;
assign addr[42338]= 304930476;
assign addr[42339]= 455461206;
assign addr[42340]= 603681519;
assign addr[42341]= 748839539;
assign addr[42342]= 890198924;
assign addr[42343]= 1027042599;
assign addr[42344]= 1158676398;
assign addr[42345]= 1284432584;
assign addr[42346]= 1403673233;
assign addr[42347]= 1515793473;
assign addr[42348]= 1620224553;
assign addr[42349]= 1716436725;
assign addr[42350]= 1803941934;
assign addr[42351]= 1882296293;
assign addr[42352]= 1951102334;
assign addr[42353]= 2010011024;
assign addr[42354]= 2058723538;
assign addr[42355]= 2096992772;
assign addr[42356]= 2124624598;
assign addr[42357]= 2141478848;
assign addr[42358]= 2147470025;
assign addr[42359]= 2142567738;
assign addr[42360]= 2126796855;
assign addr[42361]= 2100237377;
assign addr[42362]= 2063024031;
assign addr[42363]= 2015345591;
assign addr[42364]= 1957443913;
assign addr[42365]= 1889612716;
assign addr[42366]= 1812196087;
assign addr[42367]= 1725586737;
assign addr[42368]= 1630224009;
assign addr[42369]= 1526591649;
assign addr[42370]= 1415215352;
assign addr[42371]= 1296660098;
assign addr[42372]= 1171527280;
assign addr[42373]= 1040451659;
assign addr[42374]= 904098143;
assign addr[42375]= 763158411;
assign addr[42376]= 618347408;
assign addr[42377]= 470399716;
assign addr[42378]= 320065829;
assign addr[42379]= 168108346;
assign addr[42380]= 15298099;
assign addr[42381]= -137589750;
assign addr[42382]= -289779648;
assign addr[42383]= -440499581;
assign addr[42384]= -588984994;
assign addr[42385]= -734482665;
assign addr[42386]= -876254528;
assign addr[42387]= -1013581418;
assign addr[42388]= -1145766716;
assign addr[42389]= -1272139887;
assign addr[42390]= -1392059879;
assign addr[42391]= -1504918373;
assign addr[42392]= -1610142873;
assign addr[42393]= -1707199606;
assign addr[42394]= -1795596234;
assign addr[42395]= -1874884346;
assign addr[42396]= -1944661739;
assign addr[42397]= -2004574453;
assign addr[42398]= -2054318569;
assign addr[42399]= -2093641749;
assign addr[42400]= -2122344521;
assign addr[42401]= -2140281282;
assign addr[42402]= -2147361045;
assign addr[42403]= -2143547897;
assign addr[42404]= -2128861181;
assign addr[42405]= -2103375398;
assign addr[42406]= -2067219829;
assign addr[42407]= -2020577882;
assign addr[42408]= -1963686155;
assign addr[42409]= -1896833245;
assign addr[42410]= -1820358275;
assign addr[42411]= -1734649179;
assign addr[42412]= -1640140734;
assign addr[42413]= -1537312353;
assign addr[42414]= -1426685652;
assign addr[42415]= -1308821808;
assign addr[42416]= -1184318708;
assign addr[42417]= -1053807919;
assign addr[42418]= -917951481;
assign addr[42419]= -777438554;
assign addr[42420]= -632981917;
assign addr[42421]= -485314355;
assign addr[42422]= -335184940;
assign addr[42423]= -183355234;
assign addr[42424]= -30595422;
assign addr[42425]= 122319591;
assign addr[42426]= 274614114;
assign addr[42427]= 425515602;
assign addr[42428]= 574258580;
assign addr[42429]= 720088517;
assign addr[42430]= 862265664;
assign addr[42431]= 1000068799;
assign addr[42432]= 1132798888;
assign addr[42433]= 1259782632;
assign addr[42434]= 1380375881;
assign addr[42435]= 1493966902;
assign addr[42436]= 1599979481;
assign addr[42437]= 1697875851;
assign addr[42438]= 1787159411;
assign addr[42439]= 1867377253;
assign addr[42440]= 1938122457;
assign addr[42441]= 1999036154;
assign addr[42442]= 2049809346;
assign addr[42443]= 2090184478;
assign addr[42444]= 2119956737;
assign addr[42445]= 2138975100;
assign addr[42446]= 2147143090;
assign addr[42447]= 2144419275;
assign addr[42448]= 2130817471;
assign addr[42449]= 2106406677;
assign addr[42450]= 2071310720;
assign addr[42451]= 2025707632;
assign addr[42452]= 1969828744;
assign addr[42453]= 1903957513;
assign addr[42454]= 1828428082;
assign addr[42455]= 1743623590;
assign addr[42456]= 1649974225;
assign addr[42457]= 1547955041;
assign addr[42458]= 1438083551;
assign addr[42459]= 1320917099;
assign addr[42460]= 1197050035;
assign addr[42461]= 1067110699;
assign addr[42462]= 931758235;
assign addr[42463]= 791679244;
assign addr[42464]= 647584304;
assign addr[42465]= 500204365;
assign addr[42466]= 350287041;
assign addr[42467]= 198592817;
assign addr[42468]= 45891193;
assign addr[42469]= -107043224;
assign addr[42470]= -259434643;
assign addr[42471]= -410510029;
assign addr[42472]= -559503022;
assign addr[42473]= -705657826;
assign addr[42474]= -848233042;
assign addr[42475]= -986505429;
assign addr[42476]= -1119773573;
assign addr[42477]= -1247361445;
assign addr[42478]= -1368621831;
assign addr[42479]= -1482939614;
assign addr[42480]= -1589734894;
assign addr[42481]= -1688465931;
assign addr[42482]= -1778631892;
assign addr[42483]= -1859775393;
assign addr[42484]= -1931484818;
assign addr[42485]= -1993396407;
assign addr[42486]= -2045196100;
assign addr[42487]= -2086621133;
assign addr[42488]= -2117461370;
assign addr[42489]= -2137560369;
assign addr[42490]= -2146816171;
assign addr[42491]= -2145181827;
assign addr[42492]= -2132665626;
assign addr[42493]= -2109331059;
assign addr[42494]= -2075296495;
assign addr[42495]= -2030734582;
assign addr[42496]= -1975871368;
assign addr[42497]= -1910985158;
assign addr[42498]= -1836405100;
assign addr[42499]= -1752509516;
assign addr[42500]= -1659723983;
assign addr[42501]= -1558519173;
assign addr[42502]= -1449408469;
assign addr[42503]= -1332945355;
assign addr[42504]= -1209720613;
assign addr[42505]= -1080359326;
assign addr[42506]= -945517704;
assign addr[42507]= -805879757;
assign addr[42508]= -662153826;
assign addr[42509]= -515068990;
assign addr[42510]= -365371365;
assign addr[42511]= -213820322;
assign addr[42512]= -61184634;
assign addr[42513]= 91761426;
assign addr[42514]= 244242007;
assign addr[42515]= 395483624;
assign addr[42516]= 544719071;
assign addr[42517]= 691191324;
assign addr[42518]= 834157373;
assign addr[42519]= 972891995;
assign addr[42520]= 1106691431;
assign addr[42521]= 1234876957;
assign addr[42522]= 1356798326;
assign addr[42523]= 1471837070;
assign addr[42524]= 1579409630;
assign addr[42525]= 1678970324;
assign addr[42526]= 1770014111;
assign addr[42527]= 1852079154;
assign addr[42528]= 1924749160;
assign addr[42529]= 1987655498;
assign addr[42530]= 2040479063;
assign addr[42531]= 2082951896;
assign addr[42532]= 2114858546;
assign addr[42533]= 2136037160;
assign addr[42534]= 2146380306;
assign addr[42535]= 2145835515;
assign addr[42536]= 2134405552;
assign addr[42537]= 2112148396;
assign addr[42538]= 2079176953;
assign addr[42539]= 2035658475;
assign addr[42540]= 1981813720;
assign addr[42541]= 1917915825;
assign addr[42542]= 1844288924;
assign addr[42543]= 1761306505;
assign addr[42544]= 1669389513;
assign addr[42545]= 1569004214;
assign addr[42546]= 1460659832;
assign addr[42547]= 1344905966;
assign addr[42548]= 1222329801;
assign addr[42549]= 1093553126;
assign addr[42550]= 959229189;
assign addr[42551]= 820039373;
assign addr[42552]= 676689746;
assign addr[42553]= 529907477;
assign addr[42554]= 380437148;
assign addr[42555]= 229036977;
assign addr[42556]= 76474970;
assign addr[42557]= -76474970;
assign addr[42558]= -229036977;
assign addr[42559]= -380437148;
assign addr[42560]= -529907477;
assign addr[42561]= -676689746;
assign addr[42562]= -820039373;
assign addr[42563]= -959229189;
assign addr[42564]= -1093553126;
assign addr[42565]= -1222329801;
assign addr[42566]= -1344905966;
assign addr[42567]= -1460659832;
assign addr[42568]= -1569004214;
assign addr[42569]= -1669389513;
assign addr[42570]= -1761306505;
assign addr[42571]= -1844288924;
assign addr[42572]= -1917915825;
assign addr[42573]= -1981813720;
assign addr[42574]= -2035658475;
assign addr[42575]= -2079176953;
assign addr[42576]= -2112148396;
assign addr[42577]= -2134405552;
assign addr[42578]= -2145835515;
assign addr[42579]= -2146380306;
assign addr[42580]= -2136037160;
assign addr[42581]= -2114858546;
assign addr[42582]= -2082951896;
assign addr[42583]= -2040479063;
assign addr[42584]= -1987655498;
assign addr[42585]= -1924749160;
assign addr[42586]= -1852079154;
assign addr[42587]= -1770014111;
assign addr[42588]= -1678970324;
assign addr[42589]= -1579409630;
assign addr[42590]= -1471837070;
assign addr[42591]= -1356798326;
assign addr[42592]= -1234876957;
assign addr[42593]= -1106691431;
assign addr[42594]= -972891995;
assign addr[42595]= -834157373;
assign addr[42596]= -691191324;
assign addr[42597]= -544719071;
assign addr[42598]= -395483624;
assign addr[42599]= -244242007;
assign addr[42600]= -91761426;
assign addr[42601]= 61184634;
assign addr[42602]= 213820322;
assign addr[42603]= 365371365;
assign addr[42604]= 515068990;
assign addr[42605]= 662153826;
assign addr[42606]= 805879757;
assign addr[42607]= 945517704;
assign addr[42608]= 1080359326;
assign addr[42609]= 1209720613;
assign addr[42610]= 1332945355;
assign addr[42611]= 1449408469;
assign addr[42612]= 1558519173;
assign addr[42613]= 1659723983;
assign addr[42614]= 1752509516;
assign addr[42615]= 1836405100;
assign addr[42616]= 1910985158;
assign addr[42617]= 1975871368;
assign addr[42618]= 2030734582;
assign addr[42619]= 2075296495;
assign addr[42620]= 2109331059;
assign addr[42621]= 2132665626;
assign addr[42622]= 2145181827;
assign addr[42623]= 2146816171;
assign addr[42624]= 2137560369;
assign addr[42625]= 2117461370;
assign addr[42626]= 2086621133;
assign addr[42627]= 2045196100;
assign addr[42628]= 1993396407;
assign addr[42629]= 1931484818;
assign addr[42630]= 1859775393;
assign addr[42631]= 1778631892;
assign addr[42632]= 1688465931;
assign addr[42633]= 1589734894;
assign addr[42634]= 1482939614;
assign addr[42635]= 1368621831;
assign addr[42636]= 1247361445;
assign addr[42637]= 1119773573;
assign addr[42638]= 986505429;
assign addr[42639]= 848233042;
assign addr[42640]= 705657826;
assign addr[42641]= 559503022;
assign addr[42642]= 410510029;
assign addr[42643]= 259434643;
assign addr[42644]= 107043224;
assign addr[42645]= -45891193;
assign addr[42646]= -198592817;
assign addr[42647]= -350287041;
assign addr[42648]= -500204365;
assign addr[42649]= -647584304;
assign addr[42650]= -791679244;
assign addr[42651]= -931758235;
assign addr[42652]= -1067110699;
assign addr[42653]= -1197050035;
assign addr[42654]= -1320917099;
assign addr[42655]= -1438083551;
assign addr[42656]= -1547955041;
assign addr[42657]= -1649974225;
assign addr[42658]= -1743623590;
assign addr[42659]= -1828428082;
assign addr[42660]= -1903957513;
assign addr[42661]= -1969828744;
assign addr[42662]= -2025707632;
assign addr[42663]= -2071310720;
assign addr[42664]= -2106406677;
assign addr[42665]= -2130817471;
assign addr[42666]= -2144419275;
assign addr[42667]= -2147143090;
assign addr[42668]= -2138975100;
assign addr[42669]= -2119956737;
assign addr[42670]= -2090184478;
assign addr[42671]= -2049809346;
assign addr[42672]= -1999036154;
assign addr[42673]= -1938122457;
assign addr[42674]= -1867377253;
assign addr[42675]= -1787159411;
assign addr[42676]= -1697875851;
assign addr[42677]= -1599979481;
assign addr[42678]= -1493966902;
assign addr[42679]= -1380375881;
assign addr[42680]= -1259782632;
assign addr[42681]= -1132798888;
assign addr[42682]= -1000068799;
assign addr[42683]= -862265664;
assign addr[42684]= -720088517;
assign addr[42685]= -574258580;
assign addr[42686]= -425515602;
assign addr[42687]= -274614114;
assign addr[42688]= -122319591;
assign addr[42689]= 30595422;
assign addr[42690]= 183355234;
assign addr[42691]= 335184940;
assign addr[42692]= 485314355;
assign addr[42693]= 632981917;
assign addr[42694]= 777438554;
assign addr[42695]= 917951481;
assign addr[42696]= 1053807919;
assign addr[42697]= 1184318708;
assign addr[42698]= 1308821808;
assign addr[42699]= 1426685652;
assign addr[42700]= 1537312353;
assign addr[42701]= 1640140734;
assign addr[42702]= 1734649179;
assign addr[42703]= 1820358275;
assign addr[42704]= 1896833245;
assign addr[42705]= 1963686155;
assign addr[42706]= 2020577882;
assign addr[42707]= 2067219829;
assign addr[42708]= 2103375398;
assign addr[42709]= 2128861181;
assign addr[42710]= 2143547897;
assign addr[42711]= 2147361045;
assign addr[42712]= 2140281282;
assign addr[42713]= 2122344521;
assign addr[42714]= 2093641749;
assign addr[42715]= 2054318569;
assign addr[42716]= 2004574453;
assign addr[42717]= 1944661739;
assign addr[42718]= 1874884346;
assign addr[42719]= 1795596234;
assign addr[42720]= 1707199606;
assign addr[42721]= 1610142873;
assign addr[42722]= 1504918373;
assign addr[42723]= 1392059879;
assign addr[42724]= 1272139887;
assign addr[42725]= 1145766716;
assign addr[42726]= 1013581418;
assign addr[42727]= 876254528;
assign addr[42728]= 734482665;
assign addr[42729]= 588984994;
assign addr[42730]= 440499581;
assign addr[42731]= 289779648;
assign addr[42732]= 137589750;
assign addr[42733]= -15298099;
assign addr[42734]= -168108346;
assign addr[42735]= -320065829;
assign addr[42736]= -470399716;
assign addr[42737]= -618347408;
assign addr[42738]= -763158411;
assign addr[42739]= -904098143;
assign addr[42740]= -1040451659;
assign addr[42741]= -1171527280;
assign addr[42742]= -1296660098;
assign addr[42743]= -1415215352;
assign addr[42744]= -1526591649;
assign addr[42745]= -1630224009;
assign addr[42746]= -1725586737;
assign addr[42747]= -1812196087;
assign addr[42748]= -1889612716;
assign addr[42749]= -1957443913;
assign addr[42750]= -2015345591;
assign addr[42751]= -2063024031;
assign addr[42752]= -2100237377;
assign addr[42753]= -2126796855;
assign addr[42754]= -2142567738;
assign addr[42755]= -2147470025;
assign addr[42756]= -2141478848;
assign addr[42757]= -2124624598;
assign addr[42758]= -2096992772;
assign addr[42759]= -2058723538;
assign addr[42760]= -2010011024;
assign addr[42761]= -1951102334;
assign addr[42762]= -1882296293;
assign addr[42763]= -1803941934;
assign addr[42764]= -1716436725;
assign addr[42765]= -1620224553;
assign addr[42766]= -1515793473;
assign addr[42767]= -1403673233;
assign addr[42768]= -1284432584;
assign addr[42769]= -1158676398;
assign addr[42770]= -1027042599;
assign addr[42771]= -890198924;
assign addr[42772]= -748839539;
assign addr[42773]= -603681519;
assign addr[42774]= -455461206;
assign addr[42775]= -304930476;
assign addr[42776]= -152852926;
assign addr[42777]= 0;
assign addr[42778]= 152852926;
assign addr[42779]= 304930476;
assign addr[42780]= 455461206;
assign addr[42781]= 603681519;
assign addr[42782]= 748839539;
assign addr[42783]= 890198924;
assign addr[42784]= 1027042599;
assign addr[42785]= 1158676398;
assign addr[42786]= 1284432584;
assign addr[42787]= 1403673233;
assign addr[42788]= 1515793473;
assign addr[42789]= 1620224553;
assign addr[42790]= 1716436725;
assign addr[42791]= 1803941934;
assign addr[42792]= 1882296293;
assign addr[42793]= 1951102334;
assign addr[42794]= 2010011024;
assign addr[42795]= 2058723538;
assign addr[42796]= 2096992772;
assign addr[42797]= 2124624598;
assign addr[42798]= 2141478848;
assign addr[42799]= 2147470025;
assign addr[42800]= 2142567738;
assign addr[42801]= 2126796855;
assign addr[42802]= 2100237377;
assign addr[42803]= 2063024031;
assign addr[42804]= 2015345591;
assign addr[42805]= 1957443913;
assign addr[42806]= 1889612716;
assign addr[42807]= 1812196087;
assign addr[42808]= 1725586737;
assign addr[42809]= 1630224009;
assign addr[42810]= 1526591649;
assign addr[42811]= 1415215352;
assign addr[42812]= 1296660098;
assign addr[42813]= 1171527280;
assign addr[42814]= 1040451659;
assign addr[42815]= 904098143;
assign addr[42816]= 763158411;
assign addr[42817]= 618347408;
assign addr[42818]= 470399716;
assign addr[42819]= 320065829;
assign addr[42820]= 168108346;
assign addr[42821]= 15298099;
assign addr[42822]= -137589750;
assign addr[42823]= -289779648;
assign addr[42824]= -440499581;
assign addr[42825]= -588984994;
assign addr[42826]= -734482665;
assign addr[42827]= -876254528;
assign addr[42828]= -1013581418;
assign addr[42829]= -1145766716;
assign addr[42830]= -1272139887;
assign addr[42831]= -1392059879;
assign addr[42832]= -1504918373;
assign addr[42833]= -1610142873;
assign addr[42834]= -1707199606;
assign addr[42835]= -1795596234;
assign addr[42836]= -1874884346;
assign addr[42837]= -1944661739;
assign addr[42838]= -2004574453;
assign addr[42839]= -2054318569;
assign addr[42840]= -2093641749;
assign addr[42841]= -2122344521;
assign addr[42842]= -2140281282;
assign addr[42843]= -2147361045;
assign addr[42844]= -2143547897;
assign addr[42845]= -2128861181;
assign addr[42846]= -2103375398;
assign addr[42847]= -2067219829;
assign addr[42848]= -2020577882;
assign addr[42849]= -1963686155;
assign addr[42850]= -1896833245;
assign addr[42851]= -1820358275;
assign addr[42852]= -1734649179;
assign addr[42853]= -1640140734;
assign addr[42854]= -1537312353;
assign addr[42855]= -1426685652;
assign addr[42856]= -1308821808;
assign addr[42857]= -1184318708;
assign addr[42858]= -1053807919;
assign addr[42859]= -917951481;
assign addr[42860]= -777438554;
assign addr[42861]= -632981917;
assign addr[42862]= -485314355;
assign addr[42863]= -335184940;
assign addr[42864]= -183355234;
assign addr[42865]= -30595422;
assign addr[42866]= 122319591;
assign addr[42867]= 274614114;
assign addr[42868]= 425515602;
assign addr[42869]= 574258580;
assign addr[42870]= 720088517;
assign addr[42871]= 862265664;
assign addr[42872]= 1000068799;
assign addr[42873]= 1132798888;
assign addr[42874]= 1259782632;
assign addr[42875]= 1380375881;
assign addr[42876]= 1493966902;
assign addr[42877]= 1599979481;
assign addr[42878]= 1697875851;
assign addr[42879]= 1787159411;
assign addr[42880]= 1867377253;
assign addr[42881]= 1938122457;
assign addr[42882]= 1999036154;
assign addr[42883]= 2049809346;
assign addr[42884]= 2090184478;
assign addr[42885]= 2119956737;
assign addr[42886]= 2138975100;
assign addr[42887]= 2147143090;
assign addr[42888]= 2144419275;
assign addr[42889]= 2130817471;
assign addr[42890]= 2106406677;
assign addr[42891]= 2071310720;
assign addr[42892]= 2025707632;
assign addr[42893]= 1969828744;
assign addr[42894]= 1903957513;
assign addr[42895]= 1828428082;
assign addr[42896]= 1743623590;
assign addr[42897]= 1649974225;
assign addr[42898]= 1547955041;
assign addr[42899]= 1438083551;
assign addr[42900]= 1320917099;
assign addr[42901]= 1197050035;
assign addr[42902]= 1067110699;
assign addr[42903]= 931758235;
assign addr[42904]= 791679244;
assign addr[42905]= 647584304;
assign addr[42906]= 500204365;
assign addr[42907]= 350287041;
assign addr[42908]= 198592817;
assign addr[42909]= 45891193;
assign addr[42910]= -107043224;
assign addr[42911]= -259434643;
assign addr[42912]= -410510029;
assign addr[42913]= -559503022;
assign addr[42914]= -705657826;
assign addr[42915]= -848233042;
assign addr[42916]= -986505429;
assign addr[42917]= -1119773573;
assign addr[42918]= -1247361445;
assign addr[42919]= -1368621831;
assign addr[42920]= -1482939614;
assign addr[42921]= -1589734894;
assign addr[42922]= -1688465931;
assign addr[42923]= -1778631892;
assign addr[42924]= -1859775393;
assign addr[42925]= -1931484818;
assign addr[42926]= -1993396407;
assign addr[42927]= -2045196100;
assign addr[42928]= -2086621133;
assign addr[42929]= -2117461370;
assign addr[42930]= -2137560369;
assign addr[42931]= -2146816171;
assign addr[42932]= -2145181827;
assign addr[42933]= -2132665626;
assign addr[42934]= -2109331059;
assign addr[42935]= -2075296495;
assign addr[42936]= -2030734582;
assign addr[42937]= -1975871368;
assign addr[42938]= -1910985158;
assign addr[42939]= -1836405100;
assign addr[42940]= -1752509516;
assign addr[42941]= -1659723983;
assign addr[42942]= -1558519173;
assign addr[42943]= -1449408469;
assign addr[42944]= -1332945355;
assign addr[42945]= -1209720613;
assign addr[42946]= -1080359326;
assign addr[42947]= -945517704;
assign addr[42948]= -805879757;
assign addr[42949]= -662153826;
assign addr[42950]= -515068990;
assign addr[42951]= -365371365;
assign addr[42952]= -213820322;
assign addr[42953]= -61184634;
assign addr[42954]= 91761426;
assign addr[42955]= 244242007;
assign addr[42956]= 395483624;
assign addr[42957]= 544719071;
assign addr[42958]= 691191324;
assign addr[42959]= 834157373;
assign addr[42960]= 972891995;
assign addr[42961]= 1106691431;
assign addr[42962]= 1234876957;
assign addr[42963]= 1356798326;
assign addr[42964]= 1471837070;
assign addr[42965]= 1579409630;
assign addr[42966]= 1678970324;
assign addr[42967]= 1770014111;
assign addr[42968]= 1852079154;
assign addr[42969]= 1924749160;
assign addr[42970]= 1987655498;
assign addr[42971]= 2040479063;
assign addr[42972]= 2082951896;
assign addr[42973]= 2114858546;
assign addr[42974]= 2136037160;
assign addr[42975]= 2146380306;
assign addr[42976]= 2145835515;
assign addr[42977]= 2134405552;
assign addr[42978]= 2112148396;
assign addr[42979]= 2079176953;
assign addr[42980]= 2035658475;
assign addr[42981]= 1981813720;
assign addr[42982]= 1917915825;
assign addr[42983]= 1844288924;
assign addr[42984]= 1761306505;
assign addr[42985]= 1669389513;
assign addr[42986]= 1569004214;
assign addr[42987]= 1460659832;
assign addr[42988]= 1344905966;
assign addr[42989]= 1222329801;
assign addr[42990]= 1093553126;
assign addr[42991]= 959229189;
assign addr[42992]= 820039373;
assign addr[42993]= 676689746;
assign addr[42994]= 529907477;
assign addr[42995]= 380437148;
assign addr[42996]= 229036977;
assign addr[42997]= 76474970;
assign addr[42998]= -76474970;
assign addr[42999]= -229036977;
assign addr[43000]= -380437148;
assign addr[43001]= -529907477;
assign addr[43002]= -676689746;
assign addr[43003]= -820039373;
assign addr[43004]= -959229189;
assign addr[43005]= -1093553126;
assign addr[43006]= -1222329801;
assign addr[43007]= -1344905966;
assign addr[43008]= -1460659832;
assign addr[43009]= -1569004214;
assign addr[43010]= -1669389513;
assign addr[43011]= -1761306505;
assign addr[43012]= -1844288924;
assign addr[43013]= -1917915825;
assign addr[43014]= -1981813720;
assign addr[43015]= -2035658475;
assign addr[43016]= -2079176953;
assign addr[43017]= -2112148396;
assign addr[43018]= -2134405552;
assign addr[43019]= -2145835515;
assign addr[43020]= -2146380306;
assign addr[43021]= -2136037160;
assign addr[43022]= -2114858546;
assign addr[43023]= -2082951896;
assign addr[43024]= -2040479063;
assign addr[43025]= -1987655498;
assign addr[43026]= -1924749160;
assign addr[43027]= -1852079154;
assign addr[43028]= -1770014111;
assign addr[43029]= -1678970324;
assign addr[43030]= -1579409630;
assign addr[43031]= -1471837070;
assign addr[43032]= -1356798326;
assign addr[43033]= -1234876957;
assign addr[43034]= -1106691431;
assign addr[43035]= -972891995;
assign addr[43036]= -834157373;
assign addr[43037]= -691191324;
assign addr[43038]= -544719071;
assign addr[43039]= -395483624;
assign addr[43040]= -244242007;
assign addr[43041]= -91761426;
assign addr[43042]= 61184634;
assign addr[43043]= 213820322;
assign addr[43044]= 365371365;
assign addr[43045]= 515068990;
assign addr[43046]= 662153826;
assign addr[43047]= 805879757;
assign addr[43048]= 945517704;
assign addr[43049]= 1080359326;
assign addr[43050]= 1209720613;
assign addr[43051]= 1332945355;
assign addr[43052]= 1449408469;
assign addr[43053]= 1558519173;
assign addr[43054]= 1659723983;
assign addr[43055]= 1752509516;
assign addr[43056]= 1836405100;
assign addr[43057]= 1910985158;
assign addr[43058]= 1975871368;
assign addr[43059]= 2030734582;
assign addr[43060]= 2075296495;
assign addr[43061]= 2109331059;
assign addr[43062]= 2132665626;
assign addr[43063]= 2145181827;
assign addr[43064]= 2146816171;
assign addr[43065]= 2137560369;
assign addr[43066]= 2117461370;
assign addr[43067]= 2086621133;
assign addr[43068]= 2045196100;
assign addr[43069]= 1993396407;
assign addr[43070]= 1931484818;
assign addr[43071]= 1859775393;
assign addr[43072]= 1778631892;
assign addr[43073]= 1688465931;
assign addr[43074]= 1589734894;
assign addr[43075]= 1482939614;
assign addr[43076]= 1368621831;
assign addr[43077]= 1247361445;
assign addr[43078]= 1119773573;
assign addr[43079]= 986505429;
assign addr[43080]= 848233042;
assign addr[43081]= 705657826;
assign addr[43082]= 559503022;
assign addr[43083]= 410510029;
assign addr[43084]= 259434643;
assign addr[43085]= 107043224;
assign addr[43086]= -45891193;
assign addr[43087]= -198592817;
assign addr[43088]= -350287041;
assign addr[43089]= -500204365;
assign addr[43090]= -647584304;
assign addr[43091]= -791679244;
assign addr[43092]= -931758235;
assign addr[43093]= -1067110699;
assign addr[43094]= -1197050035;
assign addr[43095]= -1320917099;
assign addr[43096]= -1438083551;
assign addr[43097]= -1547955041;
assign addr[43098]= -1649974225;
assign addr[43099]= -1743623590;
assign addr[43100]= -1828428082;
assign addr[43101]= -1903957513;
assign addr[43102]= -1969828744;
assign addr[43103]= -2025707632;
assign addr[43104]= -2071310720;
assign addr[43105]= -2106406677;
assign addr[43106]= -2130817471;
assign addr[43107]= -2144419275;
assign addr[43108]= -2147143090;
assign addr[43109]= -2138975100;
assign addr[43110]= -2119956737;
assign addr[43111]= -2090184478;
assign addr[43112]= -2049809346;
assign addr[43113]= -1999036154;
assign addr[43114]= -1938122457;
assign addr[43115]= -1867377253;
assign addr[43116]= -1787159411;
assign addr[43117]= -1697875851;
assign addr[43118]= -1599979481;
assign addr[43119]= -1493966902;
assign addr[43120]= -1380375881;
assign addr[43121]= -1259782632;
assign addr[43122]= -1132798888;
assign addr[43123]= -1000068799;
assign addr[43124]= -862265664;
assign addr[43125]= -720088517;
assign addr[43126]= -574258580;
assign addr[43127]= -425515602;
assign addr[43128]= -274614114;
assign addr[43129]= -122319591;
assign addr[43130]= 30595422;
assign addr[43131]= 183355234;
assign addr[43132]= 335184940;
assign addr[43133]= 485314355;
assign addr[43134]= 632981917;
assign addr[43135]= 777438554;
assign addr[43136]= 917951481;
assign addr[43137]= 1053807919;
assign addr[43138]= 1184318708;
assign addr[43139]= 1308821808;
assign addr[43140]= 1426685652;
assign addr[43141]= 1537312353;
assign addr[43142]= 1640140734;
assign addr[43143]= 1734649179;
assign addr[43144]= 1820358275;
assign addr[43145]= 1896833245;
assign addr[43146]= 1963686155;
assign addr[43147]= 2020577882;
assign addr[43148]= 2067219829;
assign addr[43149]= 2103375398;
assign addr[43150]= 2128861181;
assign addr[43151]= 2143547897;
assign addr[43152]= 2147361045;
assign addr[43153]= 2140281282;
assign addr[43154]= 2122344521;
assign addr[43155]= 2093641749;
assign addr[43156]= 2054318569;
assign addr[43157]= 2004574453;
assign addr[43158]= 1944661739;
assign addr[43159]= 1874884346;
assign addr[43160]= 1795596234;
assign addr[43161]= 1707199606;
assign addr[43162]= 1610142873;
assign addr[43163]= 1504918373;
assign addr[43164]= 1392059879;
assign addr[43165]= 1272139887;
assign addr[43166]= 1145766716;
assign addr[43167]= 1013581418;
assign addr[43168]= 876254528;
assign addr[43169]= 734482665;
assign addr[43170]= 588984994;
assign addr[43171]= 440499581;
assign addr[43172]= 289779648;
assign addr[43173]= 137589750;
assign addr[43174]= -15298099;
assign addr[43175]= -168108346;
assign addr[43176]= -320065829;
assign addr[43177]= -470399716;
assign addr[43178]= -618347408;
assign addr[43179]= -763158411;
assign addr[43180]= -904098143;
assign addr[43181]= -1040451659;
assign addr[43182]= -1171527280;
assign addr[43183]= -1296660098;
assign addr[43184]= -1415215352;
assign addr[43185]= -1526591649;
assign addr[43186]= -1630224009;
assign addr[43187]= -1725586737;
assign addr[43188]= -1812196087;
assign addr[43189]= -1889612716;
assign addr[43190]= -1957443913;
assign addr[43191]= -2015345591;
assign addr[43192]= -2063024031;
assign addr[43193]= -2100237377;
assign addr[43194]= -2126796855;
assign addr[43195]= -2142567738;
assign addr[43196]= -2147470025;
assign addr[43197]= -2141478848;
assign addr[43198]= -2124624598;
assign addr[43199]= -2096992772;
assign addr[43200]= -2058723538;
assign addr[43201]= -2010011024;
assign addr[43202]= -1951102334;
assign addr[43203]= -1882296293;
assign addr[43204]= -1803941934;
assign addr[43205]= -1716436725;
assign addr[43206]= -1620224553;
assign addr[43207]= -1515793473;
assign addr[43208]= -1403673233;
assign addr[43209]= -1284432584;
assign addr[43210]= -1158676398;
assign addr[43211]= -1027042599;
assign addr[43212]= -890198924;
assign addr[43213]= -748839539;
assign addr[43214]= -603681519;
assign addr[43215]= -455461206;
assign addr[43216]= -304930476;
assign addr[43217]= -152852926;
assign addr[43218]= 0;
assign addr[43219]= 152852926;
assign addr[43220]= 304930476;
assign addr[43221]= 455461206;
assign addr[43222]= 603681519;
assign addr[43223]= 748839539;
assign addr[43224]= 890198924;
assign addr[43225]= 1027042599;
assign addr[43226]= 1158676398;
assign addr[43227]= 1284432584;
assign addr[43228]= 1403673233;
assign addr[43229]= 1515793473;
assign addr[43230]= 1620224553;
assign addr[43231]= 1716436725;
assign addr[43232]= 1803941934;
assign addr[43233]= 1882296293;
assign addr[43234]= 1951102334;
assign addr[43235]= 2010011024;
assign addr[43236]= 2058723538;
assign addr[43237]= 2096992772;
assign addr[43238]= 2124624598;
assign addr[43239]= 2141478848;
assign addr[43240]= 2147470025;
assign addr[43241]= 2142567738;
assign addr[43242]= 2126796855;
assign addr[43243]= 2100237377;
assign addr[43244]= 2063024031;
assign addr[43245]= 2015345591;
assign addr[43246]= 1957443913;
assign addr[43247]= 1889612716;
assign addr[43248]= 1812196087;
assign addr[43249]= 1725586737;
assign addr[43250]= 1630224009;
assign addr[43251]= 1526591649;
assign addr[43252]= 1415215352;
assign addr[43253]= 1296660098;
assign addr[43254]= 1171527280;
assign addr[43255]= 1040451659;
assign addr[43256]= 904098143;
assign addr[43257]= 763158411;
assign addr[43258]= 618347408;
assign addr[43259]= 470399716;
assign addr[43260]= 320065829;
assign addr[43261]= 168108346;
assign addr[43262]= 15298099;
assign addr[43263]= -137589750;
assign addr[43264]= -289779648;
assign addr[43265]= -440499581;
assign addr[43266]= -588984994;
assign addr[43267]= -734482665;
assign addr[43268]= -876254528;
assign addr[43269]= -1013581418;
assign addr[43270]= -1145766716;
assign addr[43271]= -1272139887;
assign addr[43272]= -1392059879;
assign addr[43273]= -1504918373;
assign addr[43274]= -1610142873;
assign addr[43275]= -1707199606;
assign addr[43276]= -1795596234;
assign addr[43277]= -1874884346;
assign addr[43278]= -1944661739;
assign addr[43279]= -2004574453;
assign addr[43280]= -2054318569;
assign addr[43281]= -2093641749;
assign addr[43282]= -2122344521;
assign addr[43283]= -2140281282;
assign addr[43284]= -2147361045;
assign addr[43285]= -2143547897;
assign addr[43286]= -2128861181;
assign addr[43287]= -2103375398;
assign addr[43288]= -2067219829;
assign addr[43289]= -2020577882;
assign addr[43290]= -1963686155;
assign addr[43291]= -1896833245;
assign addr[43292]= -1820358275;
assign addr[43293]= -1734649179;
assign addr[43294]= -1640140734;
assign addr[43295]= -1537312353;
assign addr[43296]= -1426685652;
assign addr[43297]= -1308821808;
assign addr[43298]= -1184318708;
assign addr[43299]= -1053807919;
assign addr[43300]= -917951481;
assign addr[43301]= -777438554;
assign addr[43302]= -632981917;
assign addr[43303]= -485314355;
assign addr[43304]= -335184940;
assign addr[43305]= -183355234;
assign addr[43306]= -30595422;
assign addr[43307]= 122319591;
assign addr[43308]= 274614114;
assign addr[43309]= 425515602;
assign addr[43310]= 574258580;
assign addr[43311]= 720088517;
assign addr[43312]= 862265664;
assign addr[43313]= 1000068799;
assign addr[43314]= 1132798888;
assign addr[43315]= 1259782632;
assign addr[43316]= 1380375881;
assign addr[43317]= 1493966902;
assign addr[43318]= 1599979481;
assign addr[43319]= 1697875851;
assign addr[43320]= 1787159411;
assign addr[43321]= 1867377253;
assign addr[43322]= 1938122457;
assign addr[43323]= 1999036154;
assign addr[43324]= 2049809346;
assign addr[43325]= 2090184478;
assign addr[43326]= 2119956737;
assign addr[43327]= 2138975100;
assign addr[43328]= 2147143090;
assign addr[43329]= 2144419275;
assign addr[43330]= 2130817471;
assign addr[43331]= 2106406677;
assign addr[43332]= 2071310720;
assign addr[43333]= 2025707632;
assign addr[43334]= 1969828744;
assign addr[43335]= 1903957513;
assign addr[43336]= 1828428082;
assign addr[43337]= 1743623590;
assign addr[43338]= 1649974225;
assign addr[43339]= 1547955041;
assign addr[43340]= 1438083551;
assign addr[43341]= 1320917099;
assign addr[43342]= 1197050035;
assign addr[43343]= 1067110699;
assign addr[43344]= 931758235;
assign addr[43345]= 791679244;
assign addr[43346]= 647584304;
assign addr[43347]= 500204365;
assign addr[43348]= 350287041;
assign addr[43349]= 198592817;
assign addr[43350]= 45891193;
assign addr[43351]= -107043224;
assign addr[43352]= -259434643;
assign addr[43353]= -410510029;
assign addr[43354]= -559503022;
assign addr[43355]= -705657826;
assign addr[43356]= -848233042;
assign addr[43357]= -986505429;
assign addr[43358]= -1119773573;
assign addr[43359]= -1247361445;
assign addr[43360]= -1368621831;
assign addr[43361]= -1482939614;
assign addr[43362]= -1589734894;
assign addr[43363]= -1688465931;
assign addr[43364]= -1778631892;
assign addr[43365]= -1859775393;
assign addr[43366]= -1931484818;
assign addr[43367]= -1993396407;
assign addr[43368]= -2045196100;
assign addr[43369]= -2086621133;
assign addr[43370]= -2117461370;
assign addr[43371]= -2137560369;
assign addr[43372]= -2146816171;
assign addr[43373]= -2145181827;
assign addr[43374]= -2132665626;
assign addr[43375]= -2109331059;
assign addr[43376]= -2075296495;
assign addr[43377]= -2030734582;
assign addr[43378]= -1975871368;
assign addr[43379]= -1910985158;
assign addr[43380]= -1836405100;
assign addr[43381]= -1752509516;
assign addr[43382]= -1659723983;
assign addr[43383]= -1558519173;
assign addr[43384]= -1449408469;
assign addr[43385]= -1332945355;
assign addr[43386]= -1209720613;
assign addr[43387]= -1080359326;
assign addr[43388]= -945517704;
assign addr[43389]= -805879757;
assign addr[43390]= -662153826;
assign addr[43391]= -515068990;
assign addr[43392]= -365371365;
assign addr[43393]= -213820322;
assign addr[43394]= -61184634;
assign addr[43395]= 91761426;
assign addr[43396]= 244242007;
assign addr[43397]= 395483624;
assign addr[43398]= 544719071;
assign addr[43399]= 691191324;
assign addr[43400]= 834157373;
assign addr[43401]= 972891995;
assign addr[43402]= 1106691431;
assign addr[43403]= 1234876957;
assign addr[43404]= 1356798326;
assign addr[43405]= 1471837070;
assign addr[43406]= 1579409630;
assign addr[43407]= 1678970324;
assign addr[43408]= 1770014111;
assign addr[43409]= 1852079154;
assign addr[43410]= 1924749160;
assign addr[43411]= 1987655498;
assign addr[43412]= 2040479063;
assign addr[43413]= 2082951896;
assign addr[43414]= 2114858546;
assign addr[43415]= 2136037160;
assign addr[43416]= 2146380306;
assign addr[43417]= 2145835515;
assign addr[43418]= 2134405552;
assign addr[43419]= 2112148396;
assign addr[43420]= 2079176953;
assign addr[43421]= 2035658475;
assign addr[43422]= 1981813720;
assign addr[43423]= 1917915825;
assign addr[43424]= 1844288924;
assign addr[43425]= 1761306505;
assign addr[43426]= 1669389513;
assign addr[43427]= 1569004214;
assign addr[43428]= 1460659832;
assign addr[43429]= 1344905966;
assign addr[43430]= 1222329801;
assign addr[43431]= 1093553126;
assign addr[43432]= 959229189;
assign addr[43433]= 820039373;
assign addr[43434]= 676689746;
assign addr[43435]= 529907477;
assign addr[43436]= 380437148;
assign addr[43437]= 229036977;
assign addr[43438]= 76474970;
assign addr[43439]= -76474970;
assign addr[43440]= -229036977;
assign addr[43441]= -380437148;
assign addr[43442]= -529907477;
assign addr[43443]= -676689746;
assign addr[43444]= -820039373;
assign addr[43445]= -959229189;
assign addr[43446]= -1093553126;
assign addr[43447]= -1222329801;
assign addr[43448]= -1344905966;
assign addr[43449]= -1460659832;
assign addr[43450]= -1569004214;
assign addr[43451]= -1669389513;
assign addr[43452]= -1761306505;
assign addr[43453]= -1844288924;
assign addr[43454]= -1917915825;
assign addr[43455]= -1981813720;
assign addr[43456]= -2035658475;
assign addr[43457]= -2079176953;
assign addr[43458]= -2112148396;
assign addr[43459]= -2134405552;
assign addr[43460]= -2145835515;
assign addr[43461]= -2146380306;
assign addr[43462]= -2136037160;
assign addr[43463]= -2114858546;
assign addr[43464]= -2082951896;
assign addr[43465]= -2040479063;
assign addr[43466]= -1987655498;
assign addr[43467]= -1924749160;
assign addr[43468]= -1852079154;
assign addr[43469]= -1770014111;
assign addr[43470]= -1678970324;
assign addr[43471]= -1579409630;
assign addr[43472]= -1471837070;
assign addr[43473]= -1356798326;
assign addr[43474]= -1234876957;
assign addr[43475]= -1106691431;
assign addr[43476]= -972891995;
assign addr[43477]= -834157373;
assign addr[43478]= -691191324;
assign addr[43479]= -544719071;
assign addr[43480]= -395483624;
assign addr[43481]= -244242007;
assign addr[43482]= -91761426;
assign addr[43483]= 61184634;
assign addr[43484]= 213820322;
assign addr[43485]= 365371365;
assign addr[43486]= 515068990;
assign addr[43487]= 662153826;
assign addr[43488]= 805879757;
assign addr[43489]= 945517704;
assign addr[43490]= 1080359326;
assign addr[43491]= 1209720613;
assign addr[43492]= 1332945355;
assign addr[43493]= 1449408469;
assign addr[43494]= 1558519173;
assign addr[43495]= 1659723983;
assign addr[43496]= 1752509516;
assign addr[43497]= 1836405100;
assign addr[43498]= 1910985158;
assign addr[43499]= 1975871368;
assign addr[43500]= 2030734582;
assign addr[43501]= 2075296495;
assign addr[43502]= 2109331059;
assign addr[43503]= 2132665626;
assign addr[43504]= 2145181827;
assign addr[43505]= 2146816171;
assign addr[43506]= 2137560369;
assign addr[43507]= 2117461370;
assign addr[43508]= 2086621133;
assign addr[43509]= 2045196100;
assign addr[43510]= 1993396407;
assign addr[43511]= 1931484818;
assign addr[43512]= 1859775393;
assign addr[43513]= 1778631892;
assign addr[43514]= 1688465931;
assign addr[43515]= 1589734894;
assign addr[43516]= 1482939614;
assign addr[43517]= 1368621831;
assign addr[43518]= 1247361445;
assign addr[43519]= 1119773573;
assign addr[43520]= 986505429;
assign addr[43521]= 848233042;
assign addr[43522]= 705657826;
assign addr[43523]= 559503022;
assign addr[43524]= 410510029;
assign addr[43525]= 259434643;
assign addr[43526]= 107043224;
assign addr[43527]= -45891193;
assign addr[43528]= -198592817;
assign addr[43529]= -350287041;
assign addr[43530]= -500204365;
assign addr[43531]= -647584304;
assign addr[43532]= -791679244;
assign addr[43533]= -931758235;
assign addr[43534]= -1067110699;
assign addr[43535]= -1197050035;
assign addr[43536]= -1320917099;
assign addr[43537]= -1438083551;
assign addr[43538]= -1547955041;
assign addr[43539]= -1649974225;
assign addr[43540]= -1743623590;
assign addr[43541]= -1828428082;
assign addr[43542]= -1903957513;
assign addr[43543]= -1969828744;
assign addr[43544]= -2025707632;
assign addr[43545]= -2071310720;
assign addr[43546]= -2106406677;
assign addr[43547]= -2130817471;
assign addr[43548]= -2144419275;
assign addr[43549]= -2147143090;
assign addr[43550]= -2138975100;
assign addr[43551]= -2119956737;
assign addr[43552]= -2090184478;
assign addr[43553]= -2049809346;
assign addr[43554]= -1999036154;
assign addr[43555]= -1938122457;
assign addr[43556]= -1867377253;
assign addr[43557]= -1787159411;
assign addr[43558]= -1697875851;
assign addr[43559]= -1599979481;
assign addr[43560]= -1493966902;
assign addr[43561]= -1380375881;
assign addr[43562]= -1259782632;
assign addr[43563]= -1132798888;
assign addr[43564]= -1000068799;
assign addr[43565]= -862265664;
assign addr[43566]= -720088517;
assign addr[43567]= -574258580;
assign addr[43568]= -425515602;
assign addr[43569]= -274614114;
assign addr[43570]= -122319591;
assign addr[43571]= 30595422;
assign addr[43572]= 183355234;
assign addr[43573]= 335184940;
assign addr[43574]= 485314355;
assign addr[43575]= 632981917;
assign addr[43576]= 777438554;
assign addr[43577]= 917951481;
assign addr[43578]= 1053807919;
assign addr[43579]= 1184318708;
assign addr[43580]= 1308821808;
assign addr[43581]= 1426685652;
assign addr[43582]= 1537312353;
assign addr[43583]= 1640140734;
assign addr[43584]= 1734649179;
assign addr[43585]= 1820358275;
assign addr[43586]= 1896833245;
assign addr[43587]= 1963686155;
assign addr[43588]= 2020577882;
assign addr[43589]= 2067219829;
assign addr[43590]= 2103375398;
assign addr[43591]= 2128861181;
assign addr[43592]= 2143547897;
assign addr[43593]= 2147361045;
assign addr[43594]= 2140281282;
assign addr[43595]= 2122344521;
assign addr[43596]= 2093641749;
assign addr[43597]= 2054318569;
assign addr[43598]= 2004574453;
assign addr[43599]= 1944661739;
assign addr[43600]= 1874884346;
assign addr[43601]= 1795596234;
assign addr[43602]= 1707199606;
assign addr[43603]= 1610142873;
assign addr[43604]= 1504918373;
assign addr[43605]= 1392059879;
assign addr[43606]= 1272139887;
assign addr[43607]= 1145766716;
assign addr[43608]= 1013581418;
assign addr[43609]= 876254528;
assign addr[43610]= 734482665;
assign addr[43611]= 588984994;
assign addr[43612]= 440499581;
assign addr[43613]= 289779648;
assign addr[43614]= 137589750;
assign addr[43615]= -15298099;
assign addr[43616]= -168108346;
assign addr[43617]= -320065829;
assign addr[43618]= -470399716;
assign addr[43619]= -618347408;
assign addr[43620]= -763158411;
assign addr[43621]= -904098143;
assign addr[43622]= -1040451659;
assign addr[43623]= -1171527280;
assign addr[43624]= -1296660098;
assign addr[43625]= -1415215352;
assign addr[43626]= -1526591649;
assign addr[43627]= -1630224009;
assign addr[43628]= -1725586737;
assign addr[43629]= -1812196087;
assign addr[43630]= -1889612716;
assign addr[43631]= -1957443913;
assign addr[43632]= -2015345591;
assign addr[43633]= -2063024031;
assign addr[43634]= -2100237377;
assign addr[43635]= -2126796855;
assign addr[43636]= -2142567738;
assign addr[43637]= -2147470025;
assign addr[43638]= -2141478848;
assign addr[43639]= -2124624598;
assign addr[43640]= -2096992772;
assign addr[43641]= -2058723538;
assign addr[43642]= -2010011024;
assign addr[43643]= -1951102334;
assign addr[43644]= -1882296293;
assign addr[43645]= -1803941934;
assign addr[43646]= -1716436725;
assign addr[43647]= -1620224553;
assign addr[43648]= -1515793473;
assign addr[43649]= -1403673233;
assign addr[43650]= -1284432584;
assign addr[43651]= -1158676398;
assign addr[43652]= -1027042599;
assign addr[43653]= -890198924;
assign addr[43654]= -748839539;
assign addr[43655]= -603681519;
assign addr[43656]= -455461206;
assign addr[43657]= -304930476;
assign addr[43658]= -152852926;
assign addr[43659]= 0;
assign addr[43660]= 152852926;
assign addr[43661]= 304930476;
assign addr[43662]= 455461206;
assign addr[43663]= 603681519;
assign addr[43664]= 748839539;
assign addr[43665]= 890198924;
assign addr[43666]= 1027042599;
assign addr[43667]= 1158676398;
assign addr[43668]= 1284432584;
assign addr[43669]= 1403673233;
assign addr[43670]= 1515793473;
assign addr[43671]= 1620224553;
assign addr[43672]= 1716436725;
assign addr[43673]= 1803941934;
assign addr[43674]= 1882296293;
assign addr[43675]= 1951102334;
assign addr[43676]= 2010011024;
assign addr[43677]= 2058723538;
assign addr[43678]= 2096992772;
assign addr[43679]= 2124624598;
assign addr[43680]= 2141478848;
assign addr[43681]= 2147470025;
assign addr[43682]= 2142567738;
assign addr[43683]= 2126796855;
assign addr[43684]= 2100237377;
assign addr[43685]= 2063024031;
assign addr[43686]= 2015345591;
assign addr[43687]= 1957443913;
assign addr[43688]= 1889612716;
assign addr[43689]= 1812196087;
assign addr[43690]= 1725586737;
assign addr[43691]= 1630224009;
assign addr[43692]= 1526591649;
assign addr[43693]= 1415215352;
assign addr[43694]= 1296660098;
assign addr[43695]= 1171527280;
assign addr[43696]= 1040451659;
assign addr[43697]= 904098143;
assign addr[43698]= 763158411;
assign addr[43699]= 618347408;
assign addr[43700]= 470399716;
assign addr[43701]= 320065829;
assign addr[43702]= 168108346;
assign addr[43703]= 15298099;
assign addr[43704]= -137589750;
assign addr[43705]= -289779648;
assign addr[43706]= -440499581;
assign addr[43707]= -588984994;
assign addr[43708]= -734482665;
assign addr[43709]= -876254528;
assign addr[43710]= -1013581418;
assign addr[43711]= -1145766716;
assign addr[43712]= -1272139887;
assign addr[43713]= -1392059879;
assign addr[43714]= -1504918373;
assign addr[43715]= -1610142873;
assign addr[43716]= -1707199606;
assign addr[43717]= -1795596234;
assign addr[43718]= -1874884346;
assign addr[43719]= -1944661739;
assign addr[43720]= -2004574453;
assign addr[43721]= -2054318569;
assign addr[43722]= -2093641749;
assign addr[43723]= -2122344521;
assign addr[43724]= -2140281282;
assign addr[43725]= -2147361045;
assign addr[43726]= -2143547897;
assign addr[43727]= -2128861181;
assign addr[43728]= -2103375398;
assign addr[43729]= -2067219829;
assign addr[43730]= -2020577882;
assign addr[43731]= -1963686155;
assign addr[43732]= -1896833245;
assign addr[43733]= -1820358275;
assign addr[43734]= -1734649179;
assign addr[43735]= -1640140734;
assign addr[43736]= -1537312353;
assign addr[43737]= -1426685652;
assign addr[43738]= -1308821808;
assign addr[43739]= -1184318708;
assign addr[43740]= -1053807919;
assign addr[43741]= -917951481;
assign addr[43742]= -777438554;
assign addr[43743]= -632981917;
assign addr[43744]= -485314355;
assign addr[43745]= -335184940;
assign addr[43746]= -183355234;
assign addr[43747]= -30595422;
assign addr[43748]= 122319591;
assign addr[43749]= 274614114;
assign addr[43750]= 425515602;
assign addr[43751]= 574258580;
assign addr[43752]= 720088517;
assign addr[43753]= 862265664;
assign addr[43754]= 1000068799;
assign addr[43755]= 1132798888;
assign addr[43756]= 1259782632;
assign addr[43757]= 1380375881;
assign addr[43758]= 1493966902;
assign addr[43759]= 1599979481;
assign addr[43760]= 1697875851;
assign addr[43761]= 1787159411;
assign addr[43762]= 1867377253;
assign addr[43763]= 1938122457;
assign addr[43764]= 1999036154;
assign addr[43765]= 2049809346;
assign addr[43766]= 2090184478;
assign addr[43767]= 2119956737;
assign addr[43768]= 2138975100;
assign addr[43769]= 2147143090;
assign addr[43770]= 2144419275;
assign addr[43771]= 2130817471;
assign addr[43772]= 2106406677;
assign addr[43773]= 2071310720;
assign addr[43774]= 2025707632;
assign addr[43775]= 1969828744;
assign addr[43776]= 1903957513;
assign addr[43777]= 1828428082;
assign addr[43778]= 1743623590;
assign addr[43779]= 1649974225;
assign addr[43780]= 1547955041;
assign addr[43781]= 1438083551;
assign addr[43782]= 1320917099;
assign addr[43783]= 1197050035;
assign addr[43784]= 1067110699;
assign addr[43785]= 931758235;
assign addr[43786]= 791679244;
assign addr[43787]= 647584304;
assign addr[43788]= 500204365;
assign addr[43789]= 350287041;
assign addr[43790]= 198592817;
assign addr[43791]= 45891193;
assign addr[43792]= -107043224;
assign addr[43793]= -259434643;
assign addr[43794]= -410510029;
assign addr[43795]= -559503022;
assign addr[43796]= -705657826;
assign addr[43797]= -848233042;
assign addr[43798]= -986505429;
assign addr[43799]= -1119773573;
assign addr[43800]= -1247361445;
assign addr[43801]= -1368621831;
assign addr[43802]= -1482939614;
assign addr[43803]= -1589734894;
assign addr[43804]= -1688465931;
assign addr[43805]= -1778631892;
assign addr[43806]= -1859775393;
assign addr[43807]= -1931484818;
assign addr[43808]= -1993396407;
assign addr[43809]= -2045196100;
assign addr[43810]= -2086621133;
assign addr[43811]= -2117461370;
assign addr[43812]= -2137560369;
assign addr[43813]= -2146816171;
assign addr[43814]= -2145181827;
assign addr[43815]= -2132665626;
assign addr[43816]= -2109331059;
assign addr[43817]= -2075296495;
assign addr[43818]= -2030734582;
assign addr[43819]= -1975871368;
assign addr[43820]= -1910985158;
assign addr[43821]= -1836405100;
assign addr[43822]= -1752509516;
assign addr[43823]= -1659723983;
assign addr[43824]= -1558519173;
assign addr[43825]= -1449408469;
assign addr[43826]= -1332945355;
assign addr[43827]= -1209720613;
assign addr[43828]= -1080359326;
assign addr[43829]= -945517704;
assign addr[43830]= -805879757;
assign addr[43831]= -662153826;
assign addr[43832]= -515068990;
assign addr[43833]= -365371365;
assign addr[43834]= -213820322;
assign addr[43835]= -61184634;
assign addr[43836]= 91761426;
assign addr[43837]= 244242007;
assign addr[43838]= 395483624;
assign addr[43839]= 544719071;
assign addr[43840]= 691191324;
assign addr[43841]= 834157373;
assign addr[43842]= 972891995;
assign addr[43843]= 1106691431;
assign addr[43844]= 1234876957;
assign addr[43845]= 1356798326;
assign addr[43846]= 1471837070;
assign addr[43847]= 1579409630;
assign addr[43848]= 1678970324;
assign addr[43849]= 1770014111;
assign addr[43850]= 1852079154;
assign addr[43851]= 1924749160;
assign addr[43852]= 1987655498;
assign addr[43853]= 2040479063;
assign addr[43854]= 2082951896;
assign addr[43855]= 2114858546;
assign addr[43856]= 2136037160;
assign addr[43857]= 2146380306;
assign addr[43858]= 2145835515;
assign addr[43859]= 2134405552;
assign addr[43860]= 2112148396;
assign addr[43861]= 2079176953;
assign addr[43862]= 2035658475;
assign addr[43863]= 1981813720;
assign addr[43864]= 1917915825;
assign addr[43865]= 1844288924;
assign addr[43866]= 1761306505;
assign addr[43867]= 1669389513;
assign addr[43868]= 1569004214;
assign addr[43869]= 1460659832;
assign addr[43870]= 1344905966;
assign addr[43871]= 1222329801;
assign addr[43872]= 1093553126;
assign addr[43873]= 959229189;
assign addr[43874]= 820039373;
assign addr[43875]= 676689746;
assign addr[43876]= 529907477;
assign addr[43877]= 380437148;
assign addr[43878]= 229036977;
assign addr[43879]= 76474970;
assign addr[43880]= -76474970;
assign addr[43881]= -229036977;
assign addr[43882]= -380437148;
assign addr[43883]= -529907477;
assign addr[43884]= -676689746;
assign addr[43885]= -820039373;
assign addr[43886]= -959229189;
assign addr[43887]= -1093553126;
assign addr[43888]= -1222329801;
assign addr[43889]= -1344905966;
assign addr[43890]= -1460659832;
assign addr[43891]= -1569004214;
assign addr[43892]= -1669389513;
assign addr[43893]= -1761306505;
assign addr[43894]= -1844288924;
assign addr[43895]= -1917915825;
assign addr[43896]= -1981813720;
assign addr[43897]= -2035658475;
assign addr[43898]= -2079176953;
assign addr[43899]= -2112148396;
assign addr[43900]= -2134405552;
assign addr[43901]= -2145835515;
assign addr[43902]= -2146380306;
assign addr[43903]= -2136037160;
assign addr[43904]= -2114858546;
assign addr[43905]= -2082951896;
assign addr[43906]= -2040479063;
assign addr[43907]= -1987655498;
assign addr[43908]= -1924749160;
assign addr[43909]= -1852079154;
assign addr[43910]= -1770014111;
assign addr[43911]= -1678970324;
assign addr[43912]= -1579409630;
assign addr[43913]= -1471837070;
assign addr[43914]= -1356798326;
assign addr[43915]= -1234876957;
assign addr[43916]= -1106691431;
assign addr[43917]= -972891995;
assign addr[43918]= -834157373;
assign addr[43919]= -691191324;
assign addr[43920]= -544719071;
assign addr[43921]= -395483624;
assign addr[43922]= -244242007;
assign addr[43923]= -91761426;
assign addr[43924]= 61184634;
assign addr[43925]= 213820322;
assign addr[43926]= 365371365;
assign addr[43927]= 515068990;
assign addr[43928]= 662153826;
assign addr[43929]= 805879757;
assign addr[43930]= 945517704;
assign addr[43931]= 1080359326;
assign addr[43932]= 1209720613;
assign addr[43933]= 1332945355;
assign addr[43934]= 1449408469;
assign addr[43935]= 1558519173;
assign addr[43936]= 1659723983;
assign addr[43937]= 1752509516;
assign addr[43938]= 1836405100;
assign addr[43939]= 1910985158;
assign addr[43940]= 1975871368;
assign addr[43941]= 2030734582;
assign addr[43942]= 2075296495;
assign addr[43943]= 2109331059;
assign addr[43944]= 2132665626;
assign addr[43945]= 2145181827;
assign addr[43946]= 2146816171;
assign addr[43947]= 2137560369;
assign addr[43948]= 2117461370;
assign addr[43949]= 2086621133;
assign addr[43950]= 2045196100;
assign addr[43951]= 1993396407;
assign addr[43952]= 1931484818;
assign addr[43953]= 1859775393;
assign addr[43954]= 1778631892;
assign addr[43955]= 1688465931;
assign addr[43956]= 1589734894;
assign addr[43957]= 1482939614;
assign addr[43958]= 1368621831;
assign addr[43959]= 1247361445;
assign addr[43960]= 1119773573;
assign addr[43961]= 986505429;
assign addr[43962]= 848233042;
assign addr[43963]= 705657826;
assign addr[43964]= 559503022;
assign addr[43965]= 410510029;
assign addr[43966]= 259434643;
assign addr[43967]= 107043224;
assign addr[43968]= -45891193;
assign addr[43969]= -198592817;
assign addr[43970]= -350287041;
assign addr[43971]= -500204365;
assign addr[43972]= -647584304;
assign addr[43973]= -791679244;
assign addr[43974]= -931758235;
assign addr[43975]= -1067110699;
assign addr[43976]= -1197050035;
assign addr[43977]= -1320917099;
assign addr[43978]= -1438083551;
assign addr[43979]= -1547955041;
assign addr[43980]= -1649974225;
assign addr[43981]= -1743623590;
assign addr[43982]= -1828428082;
assign addr[43983]= -1903957513;
assign addr[43984]= -1969828744;
assign addr[43985]= -2025707632;
assign addr[43986]= -2071310720;
assign addr[43987]= -2106406677;
assign addr[43988]= -2130817471;
assign addr[43989]= -2144419275;
assign addr[43990]= -2147143090;
assign addr[43991]= -2138975100;
assign addr[43992]= -2119956737;
assign addr[43993]= -2090184478;
assign addr[43994]= -2049809346;
assign addr[43995]= -1999036154;
assign addr[43996]= -1938122457;
assign addr[43997]= -1867377253;
assign addr[43998]= -1787159411;
assign addr[43999]= -1697875851;
assign addr[44000]= -1599979481;
assign addr[44001]= -1493966902;
assign addr[44002]= -1380375881;
assign addr[44003]= -1259782632;
assign addr[44004]= -1132798888;
assign addr[44005]= -1000068799;
assign addr[44006]= -862265664;
assign addr[44007]= -720088517;
assign addr[44008]= -574258580;
assign addr[44009]= -425515602;
assign addr[44010]= -274614114;
assign addr[44011]= -122319591;
assign addr[44012]= 30595422;
assign addr[44013]= 183355234;
assign addr[44014]= 335184940;
assign addr[44015]= 485314355;
assign addr[44016]= 632981917;
assign addr[44017]= 777438554;
assign addr[44018]= 917951481;
assign addr[44019]= 1053807919;
assign addr[44020]= 1184318708;
assign addr[44021]= 1308821808;
assign addr[44022]= 1426685652;
assign addr[44023]= 1537312353;
assign addr[44024]= 1640140734;
assign addr[44025]= 1734649179;
assign addr[44026]= 1820358275;
assign addr[44027]= 1896833245;
assign addr[44028]= 1963686155;
assign addr[44029]= 2020577882;
assign addr[44030]= 2067219829;
assign addr[44031]= 2103375398;
assign addr[44032]= 2128861181;
assign addr[44033]= 2143547897;
assign addr[44034]= 2147361045;
assign addr[44035]= 2140281282;
assign addr[44036]= 2122344521;
assign addr[44037]= 2093641749;
assign addr[44038]= 2054318569;
assign addr[44039]= 2004574453;
assign addr[44040]= 1944661739;
assign addr[44041]= 1874884346;
assign addr[44042]= 1795596234;
assign addr[44043]= 1707199606;
assign addr[44044]= 1610142873;
assign addr[44045]= 1504918373;
assign addr[44046]= 1392059879;
assign addr[44047]= 1272139887;
assign addr[44048]= 1145766716;
assign addr[44049]= 1013581418;
assign addr[44050]= 876254528;
assign addr[44051]= 734482665;
assign addr[44052]= 588984994;
assign addr[44053]= 440499581;
assign addr[44054]= 289779648;
assign addr[44055]= 137589750;
assign addr[44056]= -15298099;
assign addr[44057]= -168108346;
assign addr[44058]= -320065829;
assign addr[44059]= -470399716;
assign addr[44060]= -618347408;
assign addr[44061]= -763158411;
assign addr[44062]= -904098143;
assign addr[44063]= -1040451659;
assign addr[44064]= -1171527280;
assign addr[44065]= -1296660098;
assign addr[44066]= -1415215352;
assign addr[44067]= -1526591649;
assign addr[44068]= -1630224009;
assign addr[44069]= -1725586737;
assign addr[44070]= -1812196087;
assign addr[44071]= -1889612716;
assign addr[44072]= -1957443913;
assign addr[44073]= -2015345591;
assign addr[44074]= -2063024031;
assign addr[44075]= -2100237377;
assign addr[44076]= -2126796855;
assign addr[44077]= -2142567738;
assign addr[44078]= -2147470025;
assign addr[44079]= -2141478848;
assign addr[44080]= -2124624598;
assign addr[44081]= -2096992772;
assign addr[44082]= -2058723538;
assign addr[44083]= -2010011024;
assign addr[44084]= -1951102334;
assign addr[44085]= -1882296293;
assign addr[44086]= -1803941934;
assign addr[44087]= -1716436725;
assign addr[44088]= -1620224553;
assign addr[44089]= -1515793473;
assign addr[44090]= -1403673233;
assign addr[44091]= -1284432584;
assign addr[44092]= -1158676398;
assign addr[44093]= -1027042599;
assign addr[44094]= -890198924;
assign addr[44095]= -748839539;
assign addr[44096]= -603681519;
assign addr[44097]= -455461206;
assign addr[44098]= -304930476;
assign addr[44099]= -152852926;
assign addr[44100]= 0;
assign addr[44101]= 152852926;
assign addr[44102]= 304930476;
assign addr[44103]= 455461206;
assign addr[44104]= 603681519;
assign addr[44105]= 748839539;
assign addr[44106]= 890198924;
assign addr[44107]= 1027042599;
assign addr[44108]= 1158676398;
assign addr[44109]= 1284432584;
assign addr[44110]= 1403673233;
assign addr[44111]= 1515793473;
assign addr[44112]= 1620224553;
assign addr[44113]= 1716436725;
assign addr[44114]= 1803941934;
assign addr[44115]= 1882296293;
assign addr[44116]= 1951102334;
assign addr[44117]= 2010011024;
assign addr[44118]= 2058723538;
assign addr[44119]= 2096992772;
assign addr[44120]= 2124624598;
assign addr[44121]= 2141478848;
assign addr[44122]= 2147470025;
assign addr[44123]= 2142567738;
assign addr[44124]= 2126796855;
assign addr[44125]= 2100237377;
assign addr[44126]= 2063024031;
assign addr[44127]= 2015345591;
assign addr[44128]= 1957443913;
assign addr[44129]= 1889612716;
assign addr[44130]= 1812196087;
assign addr[44131]= 1725586737;
assign addr[44132]= 1630224009;
assign addr[44133]= 1526591649;
assign addr[44134]= 1415215352;
assign addr[44135]= 1296660098;
assign addr[44136]= 1171527280;
assign addr[44137]= 1040451659;
assign addr[44138]= 904098143;
assign addr[44139]= 763158411;
assign addr[44140]= 618347408;
assign addr[44141]= 470399716;
assign addr[44142]= 320065829;
assign addr[44143]= 168108346;
assign addr[44144]= 15298099;
assign addr[44145]= -137589750;
assign addr[44146]= -289779648;
assign addr[44147]= -440499581;
assign addr[44148]= -588984994;
assign addr[44149]= -734482665;
assign addr[44150]= -876254528;
assign addr[44151]= -1013581418;
assign addr[44152]= -1145766716;
assign addr[44153]= -1272139887;
assign addr[44154]= -1392059879;
assign addr[44155]= -1504918373;
assign addr[44156]= -1610142873;
assign addr[44157]= -1707199606;
assign addr[44158]= -1795596234;
assign addr[44159]= -1874884346;
assign addr[44160]= -1944661739;
assign addr[44161]= -2004574453;
assign addr[44162]= -2054318569;
assign addr[44163]= -2093641749;
assign addr[44164]= -2122344521;
assign addr[44165]= -2140281282;
assign addr[44166]= -2147361045;
assign addr[44167]= -2143547897;
assign addr[44168]= -2128861181;
assign addr[44169]= -2103375398;
assign addr[44170]= -2067219829;
assign addr[44171]= -2020577882;
assign addr[44172]= -1963686155;
assign addr[44173]= -1896833245;
assign addr[44174]= -1820358275;
assign addr[44175]= -1734649179;
assign addr[44176]= -1640140734;
assign addr[44177]= -1537312353;
assign addr[44178]= -1426685652;
assign addr[44179]= -1308821808;
assign addr[44180]= -1184318708;
assign addr[44181]= -1053807919;
assign addr[44182]= -917951481;
assign addr[44183]= -777438554;
assign addr[44184]= -632981917;
assign addr[44185]= -485314355;
assign addr[44186]= -335184940;
assign addr[44187]= -183355234;
assign addr[44188]= -30595422;
assign addr[44189]= 122319591;
assign addr[44190]= 274614114;
assign addr[44191]= 425515602;
assign addr[44192]= 574258580;
assign addr[44193]= 720088517;
assign addr[44194]= 862265664;
assign addr[44195]= 1000068799;
assign addr[44196]= 1132798888;
assign addr[44197]= 1259782632;
assign addr[44198]= 1380375881;
assign addr[44199]= 1493966902;
assign addr[44200]= 1599979481;
assign addr[44201]= 1697875851;
assign addr[44202]= 1787159411;
assign addr[44203]= 1867377253;
assign addr[44204]= 1938122457;
assign addr[44205]= 1999036154;
assign addr[44206]= 2049809346;
assign addr[44207]= 2090184478;
assign addr[44208]= 2119956737;
assign addr[44209]= 2138975100;
assign addr[44210]= 2147143090;
assign addr[44211]= 2144419275;
assign addr[44212]= 2130817471;
assign addr[44213]= 2106406677;
assign addr[44214]= 2071310720;
assign addr[44215]= 2025707632;
assign addr[44216]= 1969828744;
assign addr[44217]= 1903957513;
assign addr[44218]= 1828428082;
assign addr[44219]= 1743623590;
assign addr[44220]= 1649974225;
assign addr[44221]= 1547955041;
assign addr[44222]= 1438083551;
assign addr[44223]= 1320917099;
assign addr[44224]= 1197050035;
assign addr[44225]= 1067110699;
assign addr[44226]= 931758235;
assign addr[44227]= 791679244;
assign addr[44228]= 647584304;
assign addr[44229]= 500204365;
assign addr[44230]= 350287041;
assign addr[44231]= 198592817;
assign addr[44232]= 45891193;
assign addr[44233]= -107043224;
assign addr[44234]= -259434643;
assign addr[44235]= -410510029;
assign addr[44236]= -559503022;
assign addr[44237]= -705657826;
assign addr[44238]= -848233042;
assign addr[44239]= -986505429;
assign addr[44240]= -1119773573;
assign addr[44241]= -1247361445;
assign addr[44242]= -1368621831;
assign addr[44243]= -1482939614;
assign addr[44244]= -1589734894;
assign addr[44245]= -1688465931;
assign addr[44246]= -1778631892;
assign addr[44247]= -1859775393;
assign addr[44248]= -1931484818;
assign addr[44249]= -1993396407;
assign addr[44250]= -2045196100;
assign addr[44251]= -2086621133;
assign addr[44252]= -2117461370;
assign addr[44253]= -2137560369;
assign addr[44254]= -2146816171;
assign addr[44255]= -2145181827;
assign addr[44256]= -2132665626;
assign addr[44257]= -2109331059;
assign addr[44258]= -2075296495;
assign addr[44259]= -2030734582;
assign addr[44260]= -1975871368;
assign addr[44261]= -1910985158;
assign addr[44262]= -1836405100;
assign addr[44263]= -1752509516;
assign addr[44264]= -1659723983;
assign addr[44265]= -1558519173;
assign addr[44266]= -1449408469;
assign addr[44267]= -1332945355;
assign addr[44268]= -1209720613;
assign addr[44269]= -1080359326;
assign addr[44270]= -945517704;
assign addr[44271]= -805879757;
assign addr[44272]= -662153826;
assign addr[44273]= -515068990;
assign addr[44274]= -365371365;
assign addr[44275]= -213820322;
assign addr[44276]= -61184634;
assign addr[44277]= 91761426;
assign addr[44278]= 244242007;
assign addr[44279]= 395483624;
assign addr[44280]= 544719071;
assign addr[44281]= 691191324;
assign addr[44282]= 834157373;
assign addr[44283]= 972891995;
assign addr[44284]= 1106691431;
assign addr[44285]= 1234876957;
assign addr[44286]= 1356798326;
assign addr[44287]= 1471837070;
assign addr[44288]= 1579409630;
assign addr[44289]= 1678970324;
assign addr[44290]= 1770014111;
assign addr[44291]= 1852079154;
assign addr[44292]= 1924749160;
assign addr[44293]= 1987655498;
assign addr[44294]= 2040479063;
assign addr[44295]= 2082951896;
assign addr[44296]= 2114858546;
assign addr[44297]= 2136037160;
assign addr[44298]= 2146380306;
assign addr[44299]= 2145835515;
assign addr[44300]= 2134405552;
assign addr[44301]= 2112148396;
assign addr[44302]= 2079176953;
assign addr[44303]= 2035658475;
assign addr[44304]= 1981813720;
assign addr[44305]= 1917915825;
assign addr[44306]= 1844288924;
assign addr[44307]= 1761306505;
assign addr[44308]= 1669389513;
assign addr[44309]= 1569004214;
assign addr[44310]= 1460659832;
assign addr[44311]= 1344905966;
assign addr[44312]= 1222329801;
assign addr[44313]= 1093553126;
assign addr[44314]= 959229189;
assign addr[44315]= 820039373;
assign addr[44316]= 676689746;
assign addr[44317]= 529907477;
assign addr[44318]= 380437148;
assign addr[44319]= 229036977;
assign addr[44320]= 76474970;
assign addr[44321]= -76474970;
assign addr[44322]= -229036977;
assign addr[44323]= -380437148;
assign addr[44324]= -529907477;
assign addr[44325]= -676689746;
assign addr[44326]= -820039373;
assign addr[44327]= -959229189;
assign addr[44328]= -1093553126;
assign addr[44329]= -1222329801;
assign addr[44330]= -1344905966;
assign addr[44331]= -1460659832;
assign addr[44332]= -1569004214;
assign addr[44333]= -1669389513;
assign addr[44334]= -1761306505;
assign addr[44335]= -1844288924;
assign addr[44336]= -1917915825;
assign addr[44337]= -1981813720;
assign addr[44338]= -2035658475;
assign addr[44339]= -2079176953;
assign addr[44340]= -2112148396;
assign addr[44341]= -2134405552;
assign addr[44342]= -2145835515;
assign addr[44343]= -2146380306;
assign addr[44344]= -2136037160;
assign addr[44345]= -2114858546;
assign addr[44346]= -2082951896;
assign addr[44347]= -2040479063;
assign addr[44348]= -1987655498;
assign addr[44349]= -1924749160;
assign addr[44350]= -1852079154;
assign addr[44351]= -1770014111;
assign addr[44352]= -1678970324;
assign addr[44353]= -1579409630;
assign addr[44354]= -1471837070;
assign addr[44355]= -1356798326;
assign addr[44356]= -1234876957;
assign addr[44357]= -1106691431;
assign addr[44358]= -972891995;
assign addr[44359]= -834157373;
assign addr[44360]= -691191324;
assign addr[44361]= -544719071;
assign addr[44362]= -395483624;
assign addr[44363]= -244242007;
assign addr[44364]= -91761426;
assign addr[44365]= 61184634;
assign addr[44366]= 213820322;
assign addr[44367]= 365371365;
assign addr[44368]= 515068990;
assign addr[44369]= 662153826;
assign addr[44370]= 805879757;
assign addr[44371]= 945517704;
assign addr[44372]= 1080359326;
assign addr[44373]= 1209720613;
assign addr[44374]= 1332945355;
assign addr[44375]= 1449408469;
assign addr[44376]= 1558519173;
assign addr[44377]= 1659723983;
assign addr[44378]= 1752509516;
assign addr[44379]= 1836405100;
assign addr[44380]= 1910985158;
assign addr[44381]= 1975871368;
assign addr[44382]= 2030734582;
assign addr[44383]= 2075296495;
assign addr[44384]= 2109331059;
assign addr[44385]= 2132665626;
assign addr[44386]= 2145181827;
assign addr[44387]= 2146816171;
assign addr[44388]= 2137560369;
assign addr[44389]= 2117461370;
assign addr[44390]= 2086621133;
assign addr[44391]= 2045196100;
assign addr[44392]= 1993396407;
assign addr[44393]= 1931484818;
assign addr[44394]= 1859775393;
assign addr[44395]= 1778631892;
assign addr[44396]= 1688465931;
assign addr[44397]= 1589734894;
assign addr[44398]= 1482939614;
assign addr[44399]= 1368621831;
assign addr[44400]= 1247361445;
assign addr[44401]= 1119773573;
assign addr[44402]= 986505429;
assign addr[44403]= 848233042;
assign addr[44404]= 705657826;
assign addr[44405]= 559503022;
assign addr[44406]= 410510029;
assign addr[44407]= 259434643;
assign addr[44408]= 107043224;
assign addr[44409]= -45891193;
assign addr[44410]= -198592817;
assign addr[44411]= -350287041;
assign addr[44412]= -500204365;
assign addr[44413]= -647584304;
assign addr[44414]= -791679244;
assign addr[44415]= -931758235;
assign addr[44416]= -1067110699;
assign addr[44417]= -1197050035;
assign addr[44418]= -1320917099;
assign addr[44419]= -1438083551;
assign addr[44420]= -1547955041;
assign addr[44421]= -1649974225;
assign addr[44422]= -1743623590;
assign addr[44423]= -1828428082;
assign addr[44424]= -1903957513;
assign addr[44425]= -1969828744;
assign addr[44426]= -2025707632;
assign addr[44427]= -2071310720;
assign addr[44428]= -2106406677;
assign addr[44429]= -2130817471;
assign addr[44430]= -2144419275;
assign addr[44431]= -2147143090;
assign addr[44432]= -2138975100;
assign addr[44433]= -2119956737;
assign addr[44434]= -2090184478;
assign addr[44435]= -2049809346;
assign addr[44436]= -1999036154;
assign addr[44437]= -1938122457;
assign addr[44438]= -1867377253;
assign addr[44439]= -1787159411;
assign addr[44440]= -1697875851;
assign addr[44441]= -1599979481;
assign addr[44442]= -1493966902;
assign addr[44443]= -1380375881;
assign addr[44444]= -1259782632;
assign addr[44445]= -1132798888;
assign addr[44446]= -1000068799;
assign addr[44447]= -862265664;
assign addr[44448]= -720088517;
assign addr[44449]= -574258580;
assign addr[44450]= -425515602;
assign addr[44451]= -274614114;
assign addr[44452]= -122319591;
assign addr[44453]= 30595422;
assign addr[44454]= 183355234;
assign addr[44455]= 335184940;
assign addr[44456]= 485314355;
assign addr[44457]= 632981917;
assign addr[44458]= 777438554;
assign addr[44459]= 917951481;
assign addr[44460]= 1053807919;
assign addr[44461]= 1184318708;
assign addr[44462]= 1308821808;
assign addr[44463]= 1426685652;
assign addr[44464]= 1537312353;
assign addr[44465]= 1640140734;
assign addr[44466]= 1734649179;
assign addr[44467]= 1820358275;
assign addr[44468]= 1896833245;
assign addr[44469]= 1963686155;
assign addr[44470]= 2020577882;
assign addr[44471]= 2067219829;
assign addr[44472]= 2103375398;
assign addr[44473]= 2128861181;
assign addr[44474]= 2143547897;
assign addr[44475]= 2147361045;
assign addr[44476]= 2140281282;
assign addr[44477]= 2122344521;
assign addr[44478]= 2093641749;
assign addr[44479]= 2054318569;
assign addr[44480]= 2004574453;
assign addr[44481]= 1944661739;
assign addr[44482]= 1874884346;
assign addr[44483]= 1795596234;
assign addr[44484]= 1707199606;
assign addr[44485]= 1610142873;
assign addr[44486]= 1504918373;
assign addr[44487]= 1392059879;
assign addr[44488]= 1272139887;
assign addr[44489]= 1145766716;
assign addr[44490]= 1013581418;
assign addr[44491]= 876254528;
assign addr[44492]= 734482665;
assign addr[44493]= 588984994;
assign addr[44494]= 440499581;
assign addr[44495]= 289779648;
assign addr[44496]= 137589750;
assign addr[44497]= -15298099;
assign addr[44498]= -168108346;
assign addr[44499]= -320065829;
assign addr[44500]= -470399716;
assign addr[44501]= -618347408;
assign addr[44502]= -763158411;
assign addr[44503]= -904098143;
assign addr[44504]= -1040451659;
assign addr[44505]= -1171527280;
assign addr[44506]= -1296660098;
assign addr[44507]= -1415215352;
assign addr[44508]= -1526591649;
assign addr[44509]= -1630224009;
assign addr[44510]= -1725586737;
assign addr[44511]= -1812196087;
assign addr[44512]= -1889612716;
assign addr[44513]= -1957443913;
assign addr[44514]= -2015345591;
assign addr[44515]= -2063024031;
assign addr[44516]= -2100237377;
assign addr[44517]= -2126796855;
assign addr[44518]= -2142567738;
assign addr[44519]= -2147470025;
assign addr[44520]= -2141478848;
assign addr[44521]= -2124624598;
assign addr[44522]= -2096992772;
assign addr[44523]= -2058723538;
assign addr[44524]= -2010011024;
assign addr[44525]= -1951102334;
assign addr[44526]= -1882296293;
assign addr[44527]= -1803941934;
assign addr[44528]= -1716436725;
assign addr[44529]= -1620224553;
assign addr[44530]= -1515793473;
assign addr[44531]= -1403673233;
assign addr[44532]= -1284432584;
assign addr[44533]= -1158676398;
assign addr[44534]= -1027042599;
assign addr[44535]= -890198924;
assign addr[44536]= -748839539;
assign addr[44537]= -603681519;
assign addr[44538]= -455461206;
assign addr[44539]= -304930476;
assign addr[44540]= -152852926;
assign addr[44541]= 0;
assign addr[44542]= 152852926;
assign addr[44543]= 304930476;
assign addr[44544]= 455461206;
assign addr[44545]= 603681519;
assign addr[44546]= 748839539;
assign addr[44547]= 890198924;
assign addr[44548]= 1027042599;
assign addr[44549]= 1158676398;
assign addr[44550]= 1284432584;
assign addr[44551]= 1403673233;
assign addr[44552]= 1515793473;
assign addr[44553]= 1620224553;
assign addr[44554]= 1716436725;
assign addr[44555]= 1803941934;
assign addr[44556]= 1882296293;
assign addr[44557]= 1951102334;
assign addr[44558]= 2010011024;
assign addr[44559]= 2058723538;
assign addr[44560]= 2096992772;
assign addr[44561]= 2124624598;
assign addr[44562]= 2141478848;
assign addr[44563]= 2147470025;
assign addr[44564]= 2142567738;
assign addr[44565]= 2126796855;
assign addr[44566]= 2100237377;
assign addr[44567]= 2063024031;
assign addr[44568]= 2015345591;
assign addr[44569]= 1957443913;
assign addr[44570]= 1889612716;
assign addr[44571]= 1812196087;
assign addr[44572]= 1725586737;
assign addr[44573]= 1630224009;
assign addr[44574]= 1526591649;
assign addr[44575]= 1415215352;
assign addr[44576]= 1296660098;
assign addr[44577]= 1171527280;
assign addr[44578]= 1040451659;
assign addr[44579]= 904098143;
assign addr[44580]= 763158411;
assign addr[44581]= 618347408;
assign addr[44582]= 470399716;
assign addr[44583]= 320065829;
assign addr[44584]= 168108346;
assign addr[44585]= 15298099;
assign addr[44586]= -137589750;
assign addr[44587]= -289779648;
assign addr[44588]= -440499581;
assign addr[44589]= -588984994;
assign addr[44590]= -734482665;
assign addr[44591]= -876254528;
assign addr[44592]= -1013581418;
assign addr[44593]= -1145766716;
assign addr[44594]= -1272139887;
assign addr[44595]= -1392059879;
assign addr[44596]= -1504918373;
assign addr[44597]= -1610142873;
assign addr[44598]= -1707199606;
assign addr[44599]= -1795596234;
assign addr[44600]= -1874884346;
assign addr[44601]= -1944661739;
assign addr[44602]= -2004574453;
assign addr[44603]= -2054318569;
assign addr[44604]= -2093641749;
assign addr[44605]= -2122344521;
assign addr[44606]= -2140281282;
assign addr[44607]= -2147361045;
assign addr[44608]= -2143547897;
assign addr[44609]= -2128861181;
assign addr[44610]= -2103375398;
assign addr[44611]= -2067219829;
assign addr[44612]= -2020577882;
assign addr[44613]= -1963686155;
assign addr[44614]= -1896833245;
assign addr[44615]= -1820358275;
assign addr[44616]= -1734649179;
assign addr[44617]= -1640140734;
assign addr[44618]= -1537312353;
assign addr[44619]= -1426685652;
assign addr[44620]= -1308821808;
assign addr[44621]= -1184318708;
assign addr[44622]= -1053807919;
assign addr[44623]= -917951481;
assign addr[44624]= -777438554;
assign addr[44625]= -632981917;
assign addr[44626]= -485314355;
assign addr[44627]= -335184940;
assign addr[44628]= -183355234;
assign addr[44629]= -30595422;
assign addr[44630]= 122319591;
assign addr[44631]= 274614114;
assign addr[44632]= 425515602;
assign addr[44633]= 574258580;
assign addr[44634]= 720088517;
assign addr[44635]= 862265664;
assign addr[44636]= 1000068799;
assign addr[44637]= 1132798888;
assign addr[44638]= 1259782632;
assign addr[44639]= 1380375881;
assign addr[44640]= 1493966902;
assign addr[44641]= 1599979481;
assign addr[44642]= 1697875851;
assign addr[44643]= 1787159411;
assign addr[44644]= 1867377253;
assign addr[44645]= 1938122457;
assign addr[44646]= 1999036154;
assign addr[44647]= 2049809346;
assign addr[44648]= 2090184478;
assign addr[44649]= 2119956737;
assign addr[44650]= 2138975100;
assign addr[44651]= 2147143090;
assign addr[44652]= 2144419275;
assign addr[44653]= 2130817471;
assign addr[44654]= 2106406677;
assign addr[44655]= 2071310720;
assign addr[44656]= 2025707632;
assign addr[44657]= 1969828744;
assign addr[44658]= 1903957513;
assign addr[44659]= 1828428082;
assign addr[44660]= 1743623590;
assign addr[44661]= 1649974225;
assign addr[44662]= 1547955041;
assign addr[44663]= 1438083551;
assign addr[44664]= 1320917099;
assign addr[44665]= 1197050035;
assign addr[44666]= 1067110699;
assign addr[44667]= 931758235;
assign addr[44668]= 791679244;
assign addr[44669]= 647584304;
assign addr[44670]= 500204365;
assign addr[44671]= 350287041;
assign addr[44672]= 198592817;
assign addr[44673]= 45891193;
assign addr[44674]= -107043224;
assign addr[44675]= -259434643;
assign addr[44676]= -410510029;
assign addr[44677]= -559503022;
assign addr[44678]= -705657826;
assign addr[44679]= -848233042;
assign addr[44680]= -986505429;
assign addr[44681]= -1119773573;
assign addr[44682]= -1247361445;
assign addr[44683]= -1368621831;
assign addr[44684]= -1482939614;
assign addr[44685]= -1589734894;
assign addr[44686]= -1688465931;
assign addr[44687]= -1778631892;
assign addr[44688]= -1859775393;
assign addr[44689]= -1931484818;
assign addr[44690]= -1993396407;
assign addr[44691]= -2045196100;
assign addr[44692]= -2086621133;
assign addr[44693]= -2117461370;
assign addr[44694]= -2137560369;
assign addr[44695]= -2146816171;
assign addr[44696]= -2145181827;
assign addr[44697]= -2132665626;
assign addr[44698]= -2109331059;
assign addr[44699]= -2075296495;
assign addr[44700]= -2030734582;
assign addr[44701]= -1975871368;
assign addr[44702]= -1910985158;
assign addr[44703]= -1836405100;
assign addr[44704]= -1752509516;
assign addr[44705]= -1659723983;
assign addr[44706]= -1558519173;
assign addr[44707]= -1449408469;
assign addr[44708]= -1332945355;
assign addr[44709]= -1209720613;
assign addr[44710]= -1080359326;
assign addr[44711]= -945517704;
assign addr[44712]= -805879757;
assign addr[44713]= -662153826;
assign addr[44714]= -515068990;
assign addr[44715]= -365371365;
assign addr[44716]= -213820322;
assign addr[44717]= -61184634;
assign addr[44718]= 91761426;
assign addr[44719]= 244242007;
assign addr[44720]= 395483624;
assign addr[44721]= 544719071;
assign addr[44722]= 691191324;
assign addr[44723]= 834157373;
assign addr[44724]= 972891995;
assign addr[44725]= 1106691431;
assign addr[44726]= 1234876957;
assign addr[44727]= 1356798326;
assign addr[44728]= 1471837070;
assign addr[44729]= 1579409630;
assign addr[44730]= 1678970324;
assign addr[44731]= 1770014111;
assign addr[44732]= 1852079154;
assign addr[44733]= 1924749160;
assign addr[44734]= 1987655498;
assign addr[44735]= 2040479063;
assign addr[44736]= 2082951896;
assign addr[44737]= 2114858546;
assign addr[44738]= 2136037160;
assign addr[44739]= 2146380306;
assign addr[44740]= 2145835515;
assign addr[44741]= 2134405552;
assign addr[44742]= 2112148396;
assign addr[44743]= 2079176953;
assign addr[44744]= 2035658475;
assign addr[44745]= 1981813720;
assign addr[44746]= 1917915825;
assign addr[44747]= 1844288924;
assign addr[44748]= 1761306505;
assign addr[44749]= 1669389513;
assign addr[44750]= 1569004214;
assign addr[44751]= 1460659832;
assign addr[44752]= 1344905966;
assign addr[44753]= 1222329801;
assign addr[44754]= 1093553126;
assign addr[44755]= 959229189;
assign addr[44756]= 820039373;
assign addr[44757]= 676689746;
assign addr[44758]= 529907477;
assign addr[44759]= 380437148;
assign addr[44760]= 229036977;
assign addr[44761]= 76474970;
assign addr[44762]= -76474970;
assign addr[44763]= -229036977;
assign addr[44764]= -380437148;
assign addr[44765]= -529907477;
assign addr[44766]= -676689746;
assign addr[44767]= -820039373;
assign addr[44768]= -959229189;
assign addr[44769]= -1093553126;
assign addr[44770]= -1222329801;
assign addr[44771]= -1344905966;
assign addr[44772]= -1460659832;
assign addr[44773]= -1569004214;
assign addr[44774]= -1669389513;
assign addr[44775]= -1761306505;
assign addr[44776]= -1844288924;
assign addr[44777]= -1917915825;
assign addr[44778]= -1981813720;
assign addr[44779]= -2035658475;
assign addr[44780]= -2079176953;
assign addr[44781]= -2112148396;
assign addr[44782]= -2134405552;
assign addr[44783]= -2145835515;
assign addr[44784]= -2146380306;
assign addr[44785]= -2136037160;
assign addr[44786]= -2114858546;
assign addr[44787]= -2082951896;
assign addr[44788]= -2040479063;
assign addr[44789]= -1987655498;
assign addr[44790]= -1924749160;
assign addr[44791]= -1852079154;
assign addr[44792]= -1770014111;
assign addr[44793]= -1678970324;
assign addr[44794]= -1579409630;
assign addr[44795]= -1471837070;
assign addr[44796]= -1356798326;
assign addr[44797]= -1234876957;
assign addr[44798]= -1106691431;
assign addr[44799]= -972891995;
assign addr[44800]= -834157373;
assign addr[44801]= -691191324;
assign addr[44802]= -544719071;
assign addr[44803]= -395483624;
assign addr[44804]= -244242007;
assign addr[44805]= -91761426;
assign addr[44806]= 61184634;
assign addr[44807]= 213820322;
assign addr[44808]= 365371365;
assign addr[44809]= 515068990;
assign addr[44810]= 662153826;
assign addr[44811]= 805879757;
assign addr[44812]= 945517704;
assign addr[44813]= 1080359326;
assign addr[44814]= 1209720613;
assign addr[44815]= 1332945355;
assign addr[44816]= 1449408469;
assign addr[44817]= 1558519173;
assign addr[44818]= 1659723983;
assign addr[44819]= 1752509516;
assign addr[44820]= 1836405100;
assign addr[44821]= 1910985158;
assign addr[44822]= 1975871368;
assign addr[44823]= 2030734582;
assign addr[44824]= 2075296495;
assign addr[44825]= 2109331059;
assign addr[44826]= 2132665626;
assign addr[44827]= 2145181827;
assign addr[44828]= 2146816171;
assign addr[44829]= 2137560369;
assign addr[44830]= 2117461370;
assign addr[44831]= 2086621133;
assign addr[44832]= 2045196100;
assign addr[44833]= 1993396407;
assign addr[44834]= 1931484818;
assign addr[44835]= 1859775393;
assign addr[44836]= 1778631892;
assign addr[44837]= 1688465931;
assign addr[44838]= 1589734894;
assign addr[44839]= 1482939614;
assign addr[44840]= 1368621831;
assign addr[44841]= 1247361445;
assign addr[44842]= 1119773573;
assign addr[44843]= 986505429;
assign addr[44844]= 848233042;
assign addr[44845]= 705657826;
assign addr[44846]= 559503022;
assign addr[44847]= 410510029;
assign addr[44848]= 259434643;
assign addr[44849]= 107043224;
assign addr[44850]= -45891193;
assign addr[44851]= -198592817;
assign addr[44852]= -350287041;
assign addr[44853]= -500204365;
assign addr[44854]= -647584304;
assign addr[44855]= -791679244;
assign addr[44856]= -931758235;
assign addr[44857]= -1067110699;
assign addr[44858]= -1197050035;
assign addr[44859]= -1320917099;
assign addr[44860]= -1438083551;
assign addr[44861]= -1547955041;
assign addr[44862]= -1649974225;
assign addr[44863]= -1743623590;
assign addr[44864]= -1828428082;
assign addr[44865]= -1903957513;
assign addr[44866]= -1969828744;
assign addr[44867]= -2025707632;
assign addr[44868]= -2071310720;
assign addr[44869]= -2106406677;
assign addr[44870]= -2130817471;
assign addr[44871]= -2144419275;
assign addr[44872]= -2147143090;
assign addr[44873]= -2138975100;
assign addr[44874]= -2119956737;
assign addr[44875]= -2090184478;
assign addr[44876]= -2049809346;
assign addr[44877]= -1999036154;
assign addr[44878]= -1938122457;
assign addr[44879]= -1867377253;
assign addr[44880]= -1787159411;
assign addr[44881]= -1697875851;
assign addr[44882]= -1599979481;
assign addr[44883]= -1493966902;
assign addr[44884]= -1380375881;
assign addr[44885]= -1259782632;
assign addr[44886]= -1132798888;
assign addr[44887]= -1000068799;
assign addr[44888]= -862265664;
assign addr[44889]= -720088517;
assign addr[44890]= -574258580;
assign addr[44891]= -425515602;
assign addr[44892]= -274614114;
assign addr[44893]= -122319591;
assign addr[44894]= 30595422;
assign addr[44895]= 183355234;
assign addr[44896]= 335184940;
assign addr[44897]= 485314355;
assign addr[44898]= 632981917;
assign addr[44899]= 777438554;
assign addr[44900]= 917951481;
assign addr[44901]= 1053807919;
assign addr[44902]= 1184318708;
assign addr[44903]= 1308821808;
assign addr[44904]= 1426685652;
assign addr[44905]= 1537312353;
assign addr[44906]= 1640140734;
assign addr[44907]= 1734649179;
assign addr[44908]= 1820358275;
assign addr[44909]= 1896833245;
assign addr[44910]= 1963686155;
assign addr[44911]= 2020577882;
assign addr[44912]= 2067219829;
assign addr[44913]= 2103375398;
assign addr[44914]= 2128861181;
assign addr[44915]= 2143547897;
assign addr[44916]= 2147361045;
assign addr[44917]= 2140281282;
assign addr[44918]= 2122344521;
assign addr[44919]= 2093641749;
assign addr[44920]= 2054318569;
assign addr[44921]= 2004574453;
assign addr[44922]= 1944661739;
assign addr[44923]= 1874884346;
assign addr[44924]= 1795596234;
assign addr[44925]= 1707199606;
assign addr[44926]= 1610142873;
assign addr[44927]= 1504918373;
assign addr[44928]= 1392059879;
assign addr[44929]= 1272139887;
assign addr[44930]= 1145766716;
assign addr[44931]= 1013581418;
assign addr[44932]= 876254528;
assign addr[44933]= 734482665;
assign addr[44934]= 588984994;
assign addr[44935]= 440499581;
assign addr[44936]= 289779648;
assign addr[44937]= 137589750;
assign addr[44938]= -15298099;
assign addr[44939]= -168108346;
assign addr[44940]= -320065829;
assign addr[44941]= -470399716;
assign addr[44942]= -618347408;
assign addr[44943]= -763158411;
assign addr[44944]= -904098143;
assign addr[44945]= -1040451659;
assign addr[44946]= -1171527280;
assign addr[44947]= -1296660098;
assign addr[44948]= -1415215352;
assign addr[44949]= -1526591649;
assign addr[44950]= -1630224009;
assign addr[44951]= -1725586737;
assign addr[44952]= -1812196087;
assign addr[44953]= -1889612716;
assign addr[44954]= -1957443913;
assign addr[44955]= -2015345591;
assign addr[44956]= -2063024031;
assign addr[44957]= -2100237377;
assign addr[44958]= -2126796855;
assign addr[44959]= -2142567738;
assign addr[44960]= -2147470025;
assign addr[44961]= -2141478848;
assign addr[44962]= -2124624598;
assign addr[44963]= -2096992772;
assign addr[44964]= -2058723538;
assign addr[44965]= -2010011024;
assign addr[44966]= -1951102334;
assign addr[44967]= -1882296293;
assign addr[44968]= -1803941934;
assign addr[44969]= -1716436725;
assign addr[44970]= -1620224553;
assign addr[44971]= -1515793473;
assign addr[44972]= -1403673233;
assign addr[44973]= -1284432584;
assign addr[44974]= -1158676398;
assign addr[44975]= -1027042599;
assign addr[44976]= -890198924;
assign addr[44977]= -748839539;
assign addr[44978]= -603681519;
assign addr[44979]= -455461206;
assign addr[44980]= -304930476;
assign addr[44981]= -152852926;
assign addr[44982]= 0;
assign addr[44983]= 152852926;
assign addr[44984]= 304930476;
assign addr[44985]= 455461206;
assign addr[44986]= 603681519;
assign addr[44987]= 748839539;
assign addr[44988]= 890198924;
assign addr[44989]= 1027042599;
assign addr[44990]= 1158676398;
assign addr[44991]= 1284432584;
assign addr[44992]= 1403673233;
assign addr[44993]= 1515793473;
assign addr[44994]= 1620224553;
assign addr[44995]= 1716436725;
assign addr[44996]= 1803941934;
assign addr[44997]= 1882296293;
assign addr[44998]= 1951102334;
assign addr[44999]= 2010011024;
assign addr[45000]= 2058723538;
assign addr[45001]= 2096992772;
assign addr[45002]= 2124624598;
assign addr[45003]= 2141478848;
assign addr[45004]= 2147470025;
assign addr[45005]= 2142567738;
assign addr[45006]= 2126796855;
assign addr[45007]= 2100237377;
assign addr[45008]= 2063024031;
assign addr[45009]= 2015345591;
assign addr[45010]= 1957443913;
assign addr[45011]= 1889612716;
assign addr[45012]= 1812196087;
assign addr[45013]= 1725586737;
assign addr[45014]= 1630224009;
assign addr[45015]= 1526591649;
assign addr[45016]= 1415215352;
assign addr[45017]= 1296660098;
assign addr[45018]= 1171527280;
assign addr[45019]= 1040451659;
assign addr[45020]= 904098143;
assign addr[45021]= 763158411;
assign addr[45022]= 618347408;
assign addr[45023]= 470399716;
assign addr[45024]= 320065829;
assign addr[45025]= 168108346;
assign addr[45026]= 15298099;
assign addr[45027]= -137589750;
assign addr[45028]= -289779648;
assign addr[45029]= -440499581;
assign addr[45030]= -588984994;
assign addr[45031]= -734482665;
assign addr[45032]= -876254528;
assign addr[45033]= -1013581418;
assign addr[45034]= -1145766716;
assign addr[45035]= -1272139887;
assign addr[45036]= -1392059879;
assign addr[45037]= -1504918373;
assign addr[45038]= -1610142873;
assign addr[45039]= -1707199606;
assign addr[45040]= -1795596234;
assign addr[45041]= -1874884346;
assign addr[45042]= -1944661739;
assign addr[45043]= -2004574453;
assign addr[45044]= -2054318569;
assign addr[45045]= -2093641749;
assign addr[45046]= -2122344521;
assign addr[45047]= -2140281282;
assign addr[45048]= -2147361045;
assign addr[45049]= -2143547897;
assign addr[45050]= -2128861181;
assign addr[45051]= -2103375398;
assign addr[45052]= -2067219829;
assign addr[45053]= -2020577882;
assign addr[45054]= -1963686155;
assign addr[45055]= -1896833245;
assign addr[45056]= -1820358275;
assign addr[45057]= -1734649179;
assign addr[45058]= -1640140734;
assign addr[45059]= -1537312353;
assign addr[45060]= -1426685652;
assign addr[45061]= -1308821808;
assign addr[45062]= -1184318708;
assign addr[45063]= -1053807919;
assign addr[45064]= -917951481;
assign addr[45065]= -777438554;
assign addr[45066]= -632981917;
assign addr[45067]= -485314355;
assign addr[45068]= -335184940;
assign addr[45069]= -183355234;
assign addr[45070]= -30595422;
assign addr[45071]= 122319591;
assign addr[45072]= 274614114;
assign addr[45073]= 425515602;
assign addr[45074]= 574258580;
assign addr[45075]= 720088517;
assign addr[45076]= 862265664;
assign addr[45077]= 1000068799;
assign addr[45078]= 1132798888;
assign addr[45079]= 1259782632;
assign addr[45080]= 1380375881;
assign addr[45081]= 1493966902;
assign addr[45082]= 1599979481;
assign addr[45083]= 1697875851;
assign addr[45084]= 1787159411;
assign addr[45085]= 1867377253;
assign addr[45086]= 1938122457;
assign addr[45087]= 1999036154;
assign addr[45088]= 2049809346;
assign addr[45089]= 2090184478;
assign addr[45090]= 2119956737;
assign addr[45091]= 2138975100;
assign addr[45092]= 2147143090;
assign addr[45093]= 2144419275;
assign addr[45094]= 2130817471;
assign addr[45095]= 2106406677;
assign addr[45096]= 2071310720;
assign addr[45097]= 2025707632;
assign addr[45098]= 1969828744;
assign addr[45099]= 1903957513;
assign addr[45100]= 1828428082;
assign addr[45101]= 1743623590;
assign addr[45102]= 1649974225;
assign addr[45103]= 1547955041;
assign addr[45104]= 1438083551;
assign addr[45105]= 1320917099;
assign addr[45106]= 1197050035;
assign addr[45107]= 1067110699;
assign addr[45108]= 931758235;
assign addr[45109]= 791679244;
assign addr[45110]= 647584304;
assign addr[45111]= 500204365;
assign addr[45112]= 350287041;
assign addr[45113]= 198592817;
assign addr[45114]= 45891193;
assign addr[45115]= -107043224;
assign addr[45116]= -259434643;
assign addr[45117]= -410510029;
assign addr[45118]= -559503022;
assign addr[45119]= -705657826;
assign addr[45120]= -848233042;
assign addr[45121]= -986505429;
assign addr[45122]= -1119773573;
assign addr[45123]= -1247361445;
assign addr[45124]= -1368621831;
assign addr[45125]= -1482939614;
assign addr[45126]= -1589734894;
assign addr[45127]= -1688465931;
assign addr[45128]= -1778631892;
assign addr[45129]= -1859775393;
assign addr[45130]= -1931484818;
assign addr[45131]= -1993396407;
assign addr[45132]= -2045196100;
assign addr[45133]= -2086621133;
assign addr[45134]= -2117461370;
assign addr[45135]= -2137560369;
assign addr[45136]= -2146816171;
assign addr[45137]= -2145181827;
assign addr[45138]= -2132665626;
assign addr[45139]= -2109331059;
assign addr[45140]= -2075296495;
assign addr[45141]= -2030734582;
assign addr[45142]= -1975871368;
assign addr[45143]= -1910985158;
assign addr[45144]= -1836405100;
assign addr[45145]= -1752509516;
assign addr[45146]= -1659723983;
assign addr[45147]= -1558519173;
assign addr[45148]= -1449408469;
assign addr[45149]= -1332945355;
assign addr[45150]= -1209720613;
assign addr[45151]= -1080359326;
assign addr[45152]= -945517704;
assign addr[45153]= -805879757;
assign addr[45154]= -662153826;
assign addr[45155]= -515068990;
assign addr[45156]= -365371365;
assign addr[45157]= -213820322;
assign addr[45158]= -61184634;
assign addr[45159]= 91761426;
assign addr[45160]= 244242007;
assign addr[45161]= 395483624;
assign addr[45162]= 544719071;
assign addr[45163]= 691191324;
assign addr[45164]= 834157373;
assign addr[45165]= 972891995;
assign addr[45166]= 1106691431;
assign addr[45167]= 1234876957;
assign addr[45168]= 1356798326;
assign addr[45169]= 1471837070;
assign addr[45170]= 1579409630;
assign addr[45171]= 1678970324;
assign addr[45172]= 1770014111;
assign addr[45173]= 1852079154;
assign addr[45174]= 1924749160;
assign addr[45175]= 1987655498;
assign addr[45176]= 2040479063;
assign addr[45177]= 2082951896;
assign addr[45178]= 2114858546;
assign addr[45179]= 2136037160;
assign addr[45180]= 2146380306;
assign addr[45181]= 2145835515;
assign addr[45182]= 2134405552;
assign addr[45183]= 2112148396;
assign addr[45184]= 2079176953;
assign addr[45185]= 2035658475;
assign addr[45186]= 1981813720;
assign addr[45187]= 1917915825;
assign addr[45188]= 1844288924;
assign addr[45189]= 1761306505;
assign addr[45190]= 1669389513;
assign addr[45191]= 1569004214;
assign addr[45192]= 1460659832;
assign addr[45193]= 1344905966;
assign addr[45194]= 1222329801;
assign addr[45195]= 1093553126;
assign addr[45196]= 959229189;
assign addr[45197]= 820039373;
assign addr[45198]= 676689746;
assign addr[45199]= 529907477;
assign addr[45200]= 380437148;
assign addr[45201]= 229036977;
assign addr[45202]= 76474970;
assign addr[45203]= -76474970;
assign addr[45204]= -229036977;
assign addr[45205]= -380437148;
assign addr[45206]= -529907477;
assign addr[45207]= -676689746;
assign addr[45208]= -820039373;
assign addr[45209]= -959229189;
assign addr[45210]= -1093553126;
assign addr[45211]= -1222329801;
assign addr[45212]= -1344905966;
assign addr[45213]= -1460659832;
assign addr[45214]= -1569004214;
assign addr[45215]= -1669389513;
assign addr[45216]= -1761306505;
assign addr[45217]= -1844288924;
assign addr[45218]= -1917915825;
assign addr[45219]= -1981813720;
assign addr[45220]= -2035658475;
assign addr[45221]= -2079176953;
assign addr[45222]= -2112148396;
assign addr[45223]= -2134405552;
assign addr[45224]= -2145835515;
assign addr[45225]= -2146380306;
assign addr[45226]= -2136037160;
assign addr[45227]= -2114858546;
assign addr[45228]= -2082951896;
assign addr[45229]= -2040479063;
assign addr[45230]= -1987655498;
assign addr[45231]= -1924749160;
assign addr[45232]= -1852079154;
assign addr[45233]= -1770014111;
assign addr[45234]= -1678970324;
assign addr[45235]= -1579409630;
assign addr[45236]= -1471837070;
assign addr[45237]= -1356798326;
assign addr[45238]= -1234876957;
assign addr[45239]= -1106691431;
assign addr[45240]= -972891995;
assign addr[45241]= -834157373;
assign addr[45242]= -691191324;
assign addr[45243]= -544719071;
assign addr[45244]= -395483624;
assign addr[45245]= -244242007;
assign addr[45246]= -91761426;
assign addr[45247]= 61184634;
assign addr[45248]= 213820322;
assign addr[45249]= 365371365;
assign addr[45250]= 515068990;
assign addr[45251]= 662153826;
assign addr[45252]= 805879757;
assign addr[45253]= 945517704;
assign addr[45254]= 1080359326;
assign addr[45255]= 1209720613;
assign addr[45256]= 1332945355;
assign addr[45257]= 1449408469;
assign addr[45258]= 1558519173;
assign addr[45259]= 1659723983;
assign addr[45260]= 1752509516;
assign addr[45261]= 1836405100;
assign addr[45262]= 1910985158;
assign addr[45263]= 1975871368;
assign addr[45264]= 2030734582;
assign addr[45265]= 2075296495;
assign addr[45266]= 2109331059;
assign addr[45267]= 2132665626;
assign addr[45268]= 2145181827;
assign addr[45269]= 2146816171;
assign addr[45270]= 2137560369;
assign addr[45271]= 2117461370;
assign addr[45272]= 2086621133;
assign addr[45273]= 2045196100;
assign addr[45274]= 1993396407;
assign addr[45275]= 1931484818;
assign addr[45276]= 1859775393;
assign addr[45277]= 1778631892;
assign addr[45278]= 1688465931;
assign addr[45279]= 1589734894;
assign addr[45280]= 1482939614;
assign addr[45281]= 1368621831;
assign addr[45282]= 1247361445;
assign addr[45283]= 1119773573;
assign addr[45284]= 986505429;
assign addr[45285]= 848233042;
assign addr[45286]= 705657826;
assign addr[45287]= 559503022;
assign addr[45288]= 410510029;
assign addr[45289]= 259434643;
assign addr[45290]= 107043224;
assign addr[45291]= -45891193;
assign addr[45292]= -198592817;
assign addr[45293]= -350287041;
assign addr[45294]= -500204365;
assign addr[45295]= -647584304;
assign addr[45296]= -791679244;
assign addr[45297]= -931758235;
assign addr[45298]= -1067110699;
assign addr[45299]= -1197050035;
assign addr[45300]= -1320917099;
assign addr[45301]= -1438083551;
assign addr[45302]= -1547955041;
assign addr[45303]= -1649974225;
assign addr[45304]= -1743623590;
assign addr[45305]= -1828428082;
assign addr[45306]= -1903957513;
assign addr[45307]= -1969828744;
assign addr[45308]= -2025707632;
assign addr[45309]= -2071310720;
assign addr[45310]= -2106406677;
assign addr[45311]= -2130817471;
assign addr[45312]= -2144419275;
assign addr[45313]= -2147143090;
assign addr[45314]= -2138975100;
assign addr[45315]= -2119956737;
assign addr[45316]= -2090184478;
assign addr[45317]= -2049809346;
assign addr[45318]= -1999036154;
assign addr[45319]= -1938122457;
assign addr[45320]= -1867377253;
assign addr[45321]= -1787159411;
assign addr[45322]= -1697875851;
assign addr[45323]= -1599979481;
assign addr[45324]= -1493966902;
assign addr[45325]= -1380375881;
assign addr[45326]= -1259782632;
assign addr[45327]= -1132798888;
assign addr[45328]= -1000068799;
assign addr[45329]= -862265664;
assign addr[45330]= -720088517;
assign addr[45331]= -574258580;
assign addr[45332]= -425515602;
assign addr[45333]= -274614114;
assign addr[45334]= -122319591;
assign addr[45335]= 30595422;
assign addr[45336]= 183355234;
assign addr[45337]= 335184940;
assign addr[45338]= 485314355;
assign addr[45339]= 632981917;
assign addr[45340]= 777438554;
assign addr[45341]= 917951481;
assign addr[45342]= 1053807919;
assign addr[45343]= 1184318708;
assign addr[45344]= 1308821808;
assign addr[45345]= 1426685652;
assign addr[45346]= 1537312353;
assign addr[45347]= 1640140734;
assign addr[45348]= 1734649179;
assign addr[45349]= 1820358275;
assign addr[45350]= 1896833245;
assign addr[45351]= 1963686155;
assign addr[45352]= 2020577882;
assign addr[45353]= 2067219829;
assign addr[45354]= 2103375398;
assign addr[45355]= 2128861181;
assign addr[45356]= 2143547897;
assign addr[45357]= 2147361045;
assign addr[45358]= 2140281282;
assign addr[45359]= 2122344521;
assign addr[45360]= 2093641749;
assign addr[45361]= 2054318569;
assign addr[45362]= 2004574453;
assign addr[45363]= 1944661739;
assign addr[45364]= 1874884346;
assign addr[45365]= 1795596234;
assign addr[45366]= 1707199606;
assign addr[45367]= 1610142873;
assign addr[45368]= 1504918373;
assign addr[45369]= 1392059879;
assign addr[45370]= 1272139887;
assign addr[45371]= 1145766716;
assign addr[45372]= 1013581418;
assign addr[45373]= 876254528;
assign addr[45374]= 734482665;
assign addr[45375]= 588984994;
assign addr[45376]= 440499581;
assign addr[45377]= 289779648;
assign addr[45378]= 137589750;
assign addr[45379]= -15298099;
assign addr[45380]= -168108346;
assign addr[45381]= -320065829;
assign addr[45382]= -470399716;
assign addr[45383]= -618347408;
assign addr[45384]= -763158411;
assign addr[45385]= -904098143;
assign addr[45386]= -1040451659;
assign addr[45387]= -1171527280;
assign addr[45388]= -1296660098;
assign addr[45389]= -1415215352;
assign addr[45390]= -1526591649;
assign addr[45391]= -1630224009;
assign addr[45392]= -1725586737;
assign addr[45393]= -1812196087;
assign addr[45394]= -1889612716;
assign addr[45395]= -1957443913;
assign addr[45396]= -2015345591;
assign addr[45397]= -2063024031;
assign addr[45398]= -2100237377;
assign addr[45399]= -2126796855;
assign addr[45400]= -2142567738;
assign addr[45401]= -2147470025;
assign addr[45402]= -2141478848;
assign addr[45403]= -2124624598;
assign addr[45404]= -2096992772;
assign addr[45405]= -2058723538;
assign addr[45406]= -2010011024;
assign addr[45407]= -1951102334;
assign addr[45408]= -1882296293;
assign addr[45409]= -1803941934;
assign addr[45410]= -1716436725;
assign addr[45411]= -1620224553;
assign addr[45412]= -1515793473;
assign addr[45413]= -1403673233;
assign addr[45414]= -1284432584;
assign addr[45415]= -1158676398;
assign addr[45416]= -1027042599;
assign addr[45417]= -890198924;
assign addr[45418]= -748839539;
assign addr[45419]= -603681519;
assign addr[45420]= -455461206;
assign addr[45421]= -304930476;
assign addr[45422]= -152852926;
assign addr[45423]= 0;
assign addr[45424]= 152852926;
assign addr[45425]= 304930476;
assign addr[45426]= 455461206;
assign addr[45427]= 603681519;
assign addr[45428]= 748839539;
assign addr[45429]= 890198924;
assign addr[45430]= 1027042599;
assign addr[45431]= 1158676398;
assign addr[45432]= 1284432584;
assign addr[45433]= 1403673233;
assign addr[45434]= 1515793473;
assign addr[45435]= 1620224553;
assign addr[45436]= 1716436725;
assign addr[45437]= 1803941934;
assign addr[45438]= 1882296293;
assign addr[45439]= 1951102334;
assign addr[45440]= 2010011024;
assign addr[45441]= 2058723538;
assign addr[45442]= 2096992772;
assign addr[45443]= 2124624598;
assign addr[45444]= 2141478848;
assign addr[45445]= 2147470025;
assign addr[45446]= 2142567738;
assign addr[45447]= 2126796855;
assign addr[45448]= 2100237377;
assign addr[45449]= 2063024031;
assign addr[45450]= 2015345591;
assign addr[45451]= 1957443913;
assign addr[45452]= 1889612716;
assign addr[45453]= 1812196087;
assign addr[45454]= 1725586737;
assign addr[45455]= 1630224009;
assign addr[45456]= 1526591649;
assign addr[45457]= 1415215352;
assign addr[45458]= 1296660098;
assign addr[45459]= 1171527280;
assign addr[45460]= 1040451659;
assign addr[45461]= 904098143;
assign addr[45462]= 763158411;
assign addr[45463]= 618347408;
assign addr[45464]= 470399716;
assign addr[45465]= 320065829;
assign addr[45466]= 168108346;
assign addr[45467]= 15298099;
assign addr[45468]= -137589750;
assign addr[45469]= -289779648;
assign addr[45470]= -440499581;
assign addr[45471]= -588984994;
assign addr[45472]= -734482665;
assign addr[45473]= -876254528;
assign addr[45474]= -1013581418;
assign addr[45475]= -1145766716;
assign addr[45476]= -1272139887;
assign addr[45477]= -1392059879;
assign addr[45478]= -1504918373;
assign addr[45479]= -1610142873;
assign addr[45480]= -1707199606;
assign addr[45481]= -1795596234;
assign addr[45482]= -1874884346;
assign addr[45483]= -1944661739;
assign addr[45484]= -2004574453;
assign addr[45485]= -2054318569;
assign addr[45486]= -2093641749;
assign addr[45487]= -2122344521;
assign addr[45488]= -2140281282;
assign addr[45489]= -2147361045;
assign addr[45490]= -2143547897;
assign addr[45491]= -2128861181;
assign addr[45492]= -2103375398;
assign addr[45493]= -2067219829;
assign addr[45494]= -2020577882;
assign addr[45495]= -1963686155;
assign addr[45496]= -1896833245;
assign addr[45497]= -1820358275;
assign addr[45498]= -1734649179;
assign addr[45499]= -1640140734;
assign addr[45500]= -1537312353;
assign addr[45501]= -1426685652;
assign addr[45502]= -1308821808;
assign addr[45503]= -1184318708;
assign addr[45504]= -1053807919;
assign addr[45505]= -917951481;
assign addr[45506]= -777438554;
assign addr[45507]= -632981917;
assign addr[45508]= -485314355;
assign addr[45509]= -335184940;
assign addr[45510]= -183355234;
assign addr[45511]= -30595422;
assign addr[45512]= 122319591;
assign addr[45513]= 274614114;
assign addr[45514]= 425515602;
assign addr[45515]= 574258580;
assign addr[45516]= 720088517;
assign addr[45517]= 862265664;
assign addr[45518]= 1000068799;
assign addr[45519]= 1132798888;
assign addr[45520]= 1259782632;
assign addr[45521]= 1380375881;
assign addr[45522]= 1493966902;
assign addr[45523]= 1599979481;
assign addr[45524]= 1697875851;
assign addr[45525]= 1787159411;
assign addr[45526]= 1867377253;
assign addr[45527]= 1938122457;
assign addr[45528]= 1999036154;
assign addr[45529]= 2049809346;
assign addr[45530]= 2090184478;
assign addr[45531]= 2119956737;
assign addr[45532]= 2138975100;
assign addr[45533]= 2147143090;
assign addr[45534]= 2144419275;
assign addr[45535]= 2130817471;
assign addr[45536]= 2106406677;
assign addr[45537]= 2071310720;
assign addr[45538]= 2025707632;
assign addr[45539]= 1969828744;
assign addr[45540]= 1903957513;
assign addr[45541]= 1828428082;
assign addr[45542]= 1743623590;
assign addr[45543]= 1649974225;
assign addr[45544]= 1547955041;
assign addr[45545]= 1438083551;
assign addr[45546]= 1320917099;
assign addr[45547]= 1197050035;
assign addr[45548]= 1067110699;
assign addr[45549]= 931758235;
assign addr[45550]= 791679244;
assign addr[45551]= 647584304;
assign addr[45552]= 500204365;
assign addr[45553]= 350287041;
assign addr[45554]= 198592817;
assign addr[45555]= 45891193;
assign addr[45556]= -107043224;
assign addr[45557]= -259434643;
assign addr[45558]= -410510029;
assign addr[45559]= -559503022;
assign addr[45560]= -705657826;
assign addr[45561]= -848233042;
assign addr[45562]= -986505429;
assign addr[45563]= -1119773573;
assign addr[45564]= -1247361445;
assign addr[45565]= -1368621831;
assign addr[45566]= -1482939614;
assign addr[45567]= -1589734894;
assign addr[45568]= -1688465931;
assign addr[45569]= -1778631892;
assign addr[45570]= -1859775393;
assign addr[45571]= -1931484818;
assign addr[45572]= -1993396407;
assign addr[45573]= -2045196100;
assign addr[45574]= -2086621133;
assign addr[45575]= -2117461370;
assign addr[45576]= -2137560369;
assign addr[45577]= -2146816171;
assign addr[45578]= -2145181827;
assign addr[45579]= -2132665626;
assign addr[45580]= -2109331059;
assign addr[45581]= -2075296495;
assign addr[45582]= -2030734582;
assign addr[45583]= -1975871368;
assign addr[45584]= -1910985158;
assign addr[45585]= -1836405100;
assign addr[45586]= -1752509516;
assign addr[45587]= -1659723983;
assign addr[45588]= -1558519173;
assign addr[45589]= -1449408469;
assign addr[45590]= -1332945355;
assign addr[45591]= -1209720613;
assign addr[45592]= -1080359326;
assign addr[45593]= -945517704;
assign addr[45594]= -805879757;
assign addr[45595]= -662153826;
assign addr[45596]= -515068990;
assign addr[45597]= -365371365;
assign addr[45598]= -213820322;
assign addr[45599]= -61184634;
assign addr[45600]= 91761426;
assign addr[45601]= 244242007;
assign addr[45602]= 395483624;
assign addr[45603]= 544719071;
assign addr[45604]= 691191324;
assign addr[45605]= 834157373;
assign addr[45606]= 972891995;
assign addr[45607]= 1106691431;
assign addr[45608]= 1234876957;
assign addr[45609]= 1356798326;
assign addr[45610]= 1471837070;
assign addr[45611]= 1579409630;
assign addr[45612]= 1678970324;
assign addr[45613]= 1770014111;
assign addr[45614]= 1852079154;
assign addr[45615]= 1924749160;
assign addr[45616]= 1987655498;
assign addr[45617]= 2040479063;
assign addr[45618]= 2082951896;
assign addr[45619]= 2114858546;
assign addr[45620]= 2136037160;
assign addr[45621]= 2146380306;
assign addr[45622]= 2145835515;
assign addr[45623]= 2134405552;
assign addr[45624]= 2112148396;
assign addr[45625]= 2079176953;
assign addr[45626]= 2035658475;
assign addr[45627]= 1981813720;
assign addr[45628]= 1917915825;
assign addr[45629]= 1844288924;
assign addr[45630]= 1761306505;
assign addr[45631]= 1669389513;
assign addr[45632]= 1569004214;
assign addr[45633]= 1460659832;
assign addr[45634]= 1344905966;
assign addr[45635]= 1222329801;
assign addr[45636]= 1093553126;
assign addr[45637]= 959229189;
assign addr[45638]= 820039373;
assign addr[45639]= 676689746;
assign addr[45640]= 529907477;
assign addr[45641]= 380437148;
assign addr[45642]= 229036977;
assign addr[45643]= 76474970;
assign addr[45644]= -76474970;
assign addr[45645]= -229036977;
assign addr[45646]= -380437148;
assign addr[45647]= -529907477;
assign addr[45648]= -676689746;
assign addr[45649]= -820039373;
assign addr[45650]= -959229189;
assign addr[45651]= -1093553126;
assign addr[45652]= -1222329801;
assign addr[45653]= -1344905966;
assign addr[45654]= -1460659832;
assign addr[45655]= -1569004214;
assign addr[45656]= -1669389513;
assign addr[45657]= -1761306505;
assign addr[45658]= -1844288924;
assign addr[45659]= -1917915825;
assign addr[45660]= -1981813720;
assign addr[45661]= -2035658475;
assign addr[45662]= -2079176953;
assign addr[45663]= -2112148396;
assign addr[45664]= -2134405552;
assign addr[45665]= -2145835515;
assign addr[45666]= -2146380306;
assign addr[45667]= -2136037160;
assign addr[45668]= -2114858546;
assign addr[45669]= -2082951896;
assign addr[45670]= -2040479063;
assign addr[45671]= -1987655498;
assign addr[45672]= -1924749160;
assign addr[45673]= -1852079154;
assign addr[45674]= -1770014111;
assign addr[45675]= -1678970324;
assign addr[45676]= -1579409630;
assign addr[45677]= -1471837070;
assign addr[45678]= -1356798326;
assign addr[45679]= -1234876957;
assign addr[45680]= -1106691431;
assign addr[45681]= -972891995;
assign addr[45682]= -834157373;
assign addr[45683]= -691191324;
assign addr[45684]= -544719071;
assign addr[45685]= -395483624;
assign addr[45686]= -244242007;
assign addr[45687]= -91761426;
assign addr[45688]= 61184634;
assign addr[45689]= 213820322;
assign addr[45690]= 365371365;
assign addr[45691]= 515068990;
assign addr[45692]= 662153826;
assign addr[45693]= 805879757;
assign addr[45694]= 945517704;
assign addr[45695]= 1080359326;
assign addr[45696]= 1209720613;
assign addr[45697]= 1332945355;
assign addr[45698]= 1449408469;
assign addr[45699]= 1558519173;
assign addr[45700]= 1659723983;
assign addr[45701]= 1752509516;
assign addr[45702]= 1836405100;
assign addr[45703]= 1910985158;
assign addr[45704]= 1975871368;
assign addr[45705]= 2030734582;
assign addr[45706]= 2075296495;
assign addr[45707]= 2109331059;
assign addr[45708]= 2132665626;
assign addr[45709]= 2145181827;
assign addr[45710]= 2146816171;
assign addr[45711]= 2137560369;
assign addr[45712]= 2117461370;
assign addr[45713]= 2086621133;
assign addr[45714]= 2045196100;
assign addr[45715]= 1993396407;
assign addr[45716]= 1931484818;
assign addr[45717]= 1859775393;
assign addr[45718]= 1778631892;
assign addr[45719]= 1688465931;
assign addr[45720]= 1589734894;
assign addr[45721]= 1482939614;
assign addr[45722]= 1368621831;
assign addr[45723]= 1247361445;
assign addr[45724]= 1119773573;
assign addr[45725]= 986505429;
assign addr[45726]= 848233042;
assign addr[45727]= 705657826;
assign addr[45728]= 559503022;
assign addr[45729]= 410510029;
assign addr[45730]= 259434643;
assign addr[45731]= 107043224;
assign addr[45732]= -45891193;
assign addr[45733]= -198592817;
assign addr[45734]= -350287041;
assign addr[45735]= -500204365;
assign addr[45736]= -647584304;
assign addr[45737]= -791679244;
assign addr[45738]= -931758235;
assign addr[45739]= -1067110699;
assign addr[45740]= -1197050035;
assign addr[45741]= -1320917099;
assign addr[45742]= -1438083551;
assign addr[45743]= -1547955041;
assign addr[45744]= -1649974225;
assign addr[45745]= -1743623590;
assign addr[45746]= -1828428082;
assign addr[45747]= -1903957513;
assign addr[45748]= -1969828744;
assign addr[45749]= -2025707632;
assign addr[45750]= -2071310720;
assign addr[45751]= -2106406677;
assign addr[45752]= -2130817471;
assign addr[45753]= -2144419275;
assign addr[45754]= -2147143090;
assign addr[45755]= -2138975100;
assign addr[45756]= -2119956737;
assign addr[45757]= -2090184478;
assign addr[45758]= -2049809346;
assign addr[45759]= -1999036154;
assign addr[45760]= -1938122457;
assign addr[45761]= -1867377253;
assign addr[45762]= -1787159411;
assign addr[45763]= -1697875851;
assign addr[45764]= -1599979481;
assign addr[45765]= -1493966902;
assign addr[45766]= -1380375881;
assign addr[45767]= -1259782632;
assign addr[45768]= -1132798888;
assign addr[45769]= -1000068799;
assign addr[45770]= -862265664;
assign addr[45771]= -720088517;
assign addr[45772]= -574258580;
assign addr[45773]= -425515602;
assign addr[45774]= -274614114;
assign addr[45775]= -122319591;
assign addr[45776]= 30595422;
assign addr[45777]= 183355234;
assign addr[45778]= 335184940;
assign addr[45779]= 485314355;
assign addr[45780]= 632981917;
assign addr[45781]= 777438554;
assign addr[45782]= 917951481;
assign addr[45783]= 1053807919;
assign addr[45784]= 1184318708;
assign addr[45785]= 1308821808;
assign addr[45786]= 1426685652;
assign addr[45787]= 1537312353;
assign addr[45788]= 1640140734;
assign addr[45789]= 1734649179;
assign addr[45790]= 1820358275;
assign addr[45791]= 1896833245;
assign addr[45792]= 1963686155;
assign addr[45793]= 2020577882;
assign addr[45794]= 2067219829;
assign addr[45795]= 2103375398;
assign addr[45796]= 2128861181;
assign addr[45797]= 2143547897;
assign addr[45798]= 2147361045;
assign addr[45799]= 2140281282;
assign addr[45800]= 2122344521;
assign addr[45801]= 2093641749;
assign addr[45802]= 2054318569;
assign addr[45803]= 2004574453;
assign addr[45804]= 1944661739;
assign addr[45805]= 1874884346;
assign addr[45806]= 1795596234;
assign addr[45807]= 1707199606;
assign addr[45808]= 1610142873;
assign addr[45809]= 1504918373;
assign addr[45810]= 1392059879;
assign addr[45811]= 1272139887;
assign addr[45812]= 1145766716;
assign addr[45813]= 1013581418;
assign addr[45814]= 876254528;
assign addr[45815]= 734482665;
assign addr[45816]= 588984994;
assign addr[45817]= 440499581;
assign addr[45818]= 289779648;
assign addr[45819]= 137589750;
assign addr[45820]= -15298099;
assign addr[45821]= -168108346;
assign addr[45822]= -320065829;
assign addr[45823]= -470399716;
assign addr[45824]= -618347408;
assign addr[45825]= -763158411;
assign addr[45826]= -904098143;
assign addr[45827]= -1040451659;
assign addr[45828]= -1171527280;
assign addr[45829]= -1296660098;
assign addr[45830]= -1415215352;
assign addr[45831]= -1526591649;
assign addr[45832]= -1630224009;
assign addr[45833]= -1725586737;
assign addr[45834]= -1812196087;
assign addr[45835]= -1889612716;
assign addr[45836]= -1957443913;
assign addr[45837]= -2015345591;
assign addr[45838]= -2063024031;
assign addr[45839]= -2100237377;
assign addr[45840]= -2126796855;
assign addr[45841]= -2142567738;
assign addr[45842]= -2147470025;
assign addr[45843]= -2141478848;
assign addr[45844]= -2124624598;
assign addr[45845]= -2096992772;
assign addr[45846]= -2058723538;
assign addr[45847]= -2010011024;
assign addr[45848]= -1951102334;
assign addr[45849]= -1882296293;
assign addr[45850]= -1803941934;
assign addr[45851]= -1716436725;
assign addr[45852]= -1620224553;
assign addr[45853]= -1515793473;
assign addr[45854]= -1403673233;
assign addr[45855]= -1284432584;
assign addr[45856]= -1158676398;
assign addr[45857]= -1027042599;
assign addr[45858]= -890198924;
assign addr[45859]= -748839539;
assign addr[45860]= -603681519;
assign addr[45861]= -455461206;
assign addr[45862]= -304930476;
assign addr[45863]= -152852926;
assign addr[45864]= 0;
assign addr[45865]= 152852926;
assign addr[45866]= 304930476;
assign addr[45867]= 455461206;
assign addr[45868]= 603681519;
assign addr[45869]= 748839539;
assign addr[45870]= 890198924;
assign addr[45871]= 1027042599;
assign addr[45872]= 1158676398;
assign addr[45873]= 1284432584;
assign addr[45874]= 1403673233;
assign addr[45875]= 1515793473;
assign addr[45876]= 1620224553;
assign addr[45877]= 1716436725;
assign addr[45878]= 1803941934;
assign addr[45879]= 1882296293;
assign addr[45880]= 1951102334;
assign addr[45881]= 2010011024;
assign addr[45882]= 2058723538;
assign addr[45883]= 2096992772;
assign addr[45884]= 2124624598;
assign addr[45885]= 2141478848;
assign addr[45886]= 2147470025;
assign addr[45887]= 2142567738;
assign addr[45888]= 2126796855;
assign addr[45889]= 2100237377;
assign addr[45890]= 2063024031;
assign addr[45891]= 2015345591;
assign addr[45892]= 1957443913;
assign addr[45893]= 1889612716;
assign addr[45894]= 1812196087;
assign addr[45895]= 1725586737;
assign addr[45896]= 1630224009;
assign addr[45897]= 1526591649;
assign addr[45898]= 1415215352;
assign addr[45899]= 1296660098;
assign addr[45900]= 1171527280;
assign addr[45901]= 1040451659;
assign addr[45902]= 904098143;
assign addr[45903]= 763158411;
assign addr[45904]= 618347408;
assign addr[45905]= 470399716;
assign addr[45906]= 320065829;
assign addr[45907]= 168108346;
assign addr[45908]= 15298099;
assign addr[45909]= -137589750;
assign addr[45910]= -289779648;
assign addr[45911]= -440499581;
assign addr[45912]= -588984994;
assign addr[45913]= -734482665;
assign addr[45914]= -876254528;
assign addr[45915]= -1013581418;
assign addr[45916]= -1145766716;
assign addr[45917]= -1272139887;
assign addr[45918]= -1392059879;
assign addr[45919]= -1504918373;
assign addr[45920]= -1610142873;
assign addr[45921]= -1707199606;
assign addr[45922]= -1795596234;
assign addr[45923]= -1874884346;
assign addr[45924]= -1944661739;
assign addr[45925]= -2004574453;
assign addr[45926]= -2054318569;
assign addr[45927]= -2093641749;
assign addr[45928]= -2122344521;
assign addr[45929]= -2140281282;
assign addr[45930]= -2147361045;
assign addr[45931]= -2143547897;
assign addr[45932]= -2128861181;
assign addr[45933]= -2103375398;
assign addr[45934]= -2067219829;
assign addr[45935]= -2020577882;
assign addr[45936]= -1963686155;
assign addr[45937]= -1896833245;
assign addr[45938]= -1820358275;
assign addr[45939]= -1734649179;
assign addr[45940]= -1640140734;
assign addr[45941]= -1537312353;
assign addr[45942]= -1426685652;
assign addr[45943]= -1308821808;
assign addr[45944]= -1184318708;
assign addr[45945]= -1053807919;
assign addr[45946]= -917951481;
assign addr[45947]= -777438554;
assign addr[45948]= -632981917;
assign addr[45949]= -485314355;
assign addr[45950]= -335184940;
assign addr[45951]= -183355234;
assign addr[45952]= -30595422;
assign addr[45953]= 122319591;
assign addr[45954]= 274614114;
assign addr[45955]= 425515602;
assign addr[45956]= 574258580;
assign addr[45957]= 720088517;
assign addr[45958]= 862265664;
assign addr[45959]= 1000068799;
assign addr[45960]= 1132798888;
assign addr[45961]= 1259782632;
assign addr[45962]= 1380375881;
assign addr[45963]= 1493966902;
assign addr[45964]= 1599979481;
assign addr[45965]= 1697875851;
assign addr[45966]= 1787159411;
assign addr[45967]= 1867377253;
assign addr[45968]= 1938122457;
assign addr[45969]= 1999036154;
assign addr[45970]= 2049809346;
assign addr[45971]= 2090184478;
assign addr[45972]= 2119956737;
assign addr[45973]= 2138975100;
assign addr[45974]= 2147143090;
assign addr[45975]= 2144419275;
assign addr[45976]= 2130817471;
assign addr[45977]= 2106406677;
assign addr[45978]= 2071310720;
assign addr[45979]= 2025707632;
assign addr[45980]= 1969828744;
assign addr[45981]= 1903957513;
assign addr[45982]= 1828428082;
assign addr[45983]= 1743623590;
assign addr[45984]= 1649974225;
assign addr[45985]= 1547955041;
assign addr[45986]= 1438083551;
assign addr[45987]= 1320917099;
assign addr[45988]= 1197050035;
assign addr[45989]= 1067110699;
assign addr[45990]= 931758235;
assign addr[45991]= 791679244;
assign addr[45992]= 647584304;
assign addr[45993]= 500204365;
assign addr[45994]= 350287041;
assign addr[45995]= 198592817;
assign addr[45996]= 45891193;
assign addr[45997]= -107043224;
assign addr[45998]= -259434643;
assign addr[45999]= -410510029;
assign addr[46000]= -559503022;
assign addr[46001]= -705657826;
assign addr[46002]= -848233042;
assign addr[46003]= -986505429;
assign addr[46004]= -1119773573;
assign addr[46005]= -1247361445;
assign addr[46006]= -1368621831;
assign addr[46007]= -1482939614;
assign addr[46008]= -1589734894;
assign addr[46009]= -1688465931;
assign addr[46010]= -1778631892;
assign addr[46011]= -1859775393;
assign addr[46012]= -1931484818;
assign addr[46013]= -1993396407;
assign addr[46014]= -2045196100;
assign addr[46015]= -2086621133;
assign addr[46016]= -2117461370;
assign addr[46017]= -2137560369;
assign addr[46018]= -2146816171;
assign addr[46019]= -2145181827;
assign addr[46020]= -2132665626;
assign addr[46021]= -2109331059;
assign addr[46022]= -2075296495;
assign addr[46023]= -2030734582;
assign addr[46024]= -1975871368;
assign addr[46025]= -1910985158;
assign addr[46026]= -1836405100;
assign addr[46027]= -1752509516;
assign addr[46028]= -1659723983;
assign addr[46029]= -1558519173;
assign addr[46030]= -1449408469;
assign addr[46031]= -1332945355;
assign addr[46032]= -1209720613;
assign addr[46033]= -1080359326;
assign addr[46034]= -945517704;
assign addr[46035]= -805879757;
assign addr[46036]= -662153826;
assign addr[46037]= -515068990;
assign addr[46038]= -365371365;
assign addr[46039]= -213820322;
assign addr[46040]= -61184634;
assign addr[46041]= 91761426;
assign addr[46042]= 244242007;
assign addr[46043]= 395483624;
assign addr[46044]= 544719071;
assign addr[46045]= 691191324;
assign addr[46046]= 834157373;
assign addr[46047]= 972891995;
assign addr[46048]= 1106691431;
assign addr[46049]= 1234876957;
assign addr[46050]= 1356798326;
assign addr[46051]= 1471837070;
assign addr[46052]= 1579409630;
assign addr[46053]= 1678970324;
assign addr[46054]= 1770014111;
assign addr[46055]= 1852079154;
assign addr[46056]= 1924749160;
assign addr[46057]= 1987655498;
assign addr[46058]= 2040479063;
assign addr[46059]= 2082951896;
assign addr[46060]= 2114858546;
assign addr[46061]= 2136037160;
assign addr[46062]= 2146380306;
assign addr[46063]= 2145835515;
assign addr[46064]= 2134405552;
assign addr[46065]= 2112148396;
assign addr[46066]= 2079176953;
assign addr[46067]= 2035658475;
assign addr[46068]= 1981813720;
assign addr[46069]= 1917915825;
assign addr[46070]= 1844288924;
assign addr[46071]= 1761306505;
assign addr[46072]= 1669389513;
assign addr[46073]= 1569004214;
assign addr[46074]= 1460659832;
assign addr[46075]= 1344905966;
assign addr[46076]= 1222329801;
assign addr[46077]= 1093553126;
assign addr[46078]= 959229189;
assign addr[46079]= 820039373;
assign addr[46080]= 676689746;
assign addr[46081]= 529907477;
assign addr[46082]= 380437148;
assign addr[46083]= 229036977;
assign addr[46084]= 76474970;
assign addr[46085]= -76474970;
assign addr[46086]= -229036977;
assign addr[46087]= -380437148;
assign addr[46088]= -529907477;
assign addr[46089]= -676689746;
assign addr[46090]= -820039373;
assign addr[46091]= -959229189;
assign addr[46092]= -1093553126;
assign addr[46093]= -1222329801;
assign addr[46094]= -1344905966;
assign addr[46095]= -1460659832;
assign addr[46096]= -1569004214;
assign addr[46097]= -1669389513;
assign addr[46098]= -1761306505;
assign addr[46099]= -1844288924;
assign addr[46100]= -1917915825;
assign addr[46101]= -1981813720;
assign addr[46102]= -2035658475;
assign addr[46103]= -2079176953;
assign addr[46104]= -2112148396;
assign addr[46105]= -2134405552;
assign addr[46106]= -2145835515;
assign addr[46107]= -2146380306;
assign addr[46108]= -2136037160;
assign addr[46109]= -2114858546;
assign addr[46110]= -2082951896;
assign addr[46111]= -2040479063;
assign addr[46112]= -1987655498;
assign addr[46113]= -1924749160;
assign addr[46114]= -1852079154;
assign addr[46115]= -1770014111;
assign addr[46116]= -1678970324;
assign addr[46117]= -1579409630;
assign addr[46118]= -1471837070;
assign addr[46119]= -1356798326;
assign addr[46120]= -1234876957;
assign addr[46121]= -1106691431;
assign addr[46122]= -972891995;
assign addr[46123]= -834157373;
assign addr[46124]= -691191324;
assign addr[46125]= -544719071;
assign addr[46126]= -395483624;
assign addr[46127]= -244242007;
assign addr[46128]= -91761426;
assign addr[46129]= 61184634;
assign addr[46130]= 213820322;
assign addr[46131]= 365371365;
assign addr[46132]= 515068990;
assign addr[46133]= 662153826;
assign addr[46134]= 805879757;
assign addr[46135]= 945517704;
assign addr[46136]= 1080359326;
assign addr[46137]= 1209720613;
assign addr[46138]= 1332945355;
assign addr[46139]= 1449408469;
assign addr[46140]= 1558519173;
assign addr[46141]= 1659723983;
assign addr[46142]= 1752509516;
assign addr[46143]= 1836405100;
assign addr[46144]= 1910985158;
assign addr[46145]= 1975871368;
assign addr[46146]= 2030734582;
assign addr[46147]= 2075296495;
assign addr[46148]= 2109331059;
assign addr[46149]= 2132665626;
assign addr[46150]= 2145181827;
assign addr[46151]= 2146816171;
assign addr[46152]= 2137560369;
assign addr[46153]= 2117461370;
assign addr[46154]= 2086621133;
assign addr[46155]= 2045196100;
assign addr[46156]= 1993396407;
assign addr[46157]= 1931484818;
assign addr[46158]= 1859775393;
assign addr[46159]= 1778631892;
assign addr[46160]= 1688465931;
assign addr[46161]= 1589734894;
assign addr[46162]= 1482939614;
assign addr[46163]= 1368621831;
assign addr[46164]= 1247361445;
assign addr[46165]= 1119773573;
assign addr[46166]= 986505429;
assign addr[46167]= 848233042;
assign addr[46168]= 705657826;
assign addr[46169]= 559503022;
assign addr[46170]= 410510029;
assign addr[46171]= 259434643;
assign addr[46172]= 107043224;
assign addr[46173]= -45891193;
assign addr[46174]= -198592817;
assign addr[46175]= -350287041;
assign addr[46176]= -500204365;
assign addr[46177]= -647584304;
assign addr[46178]= -791679244;
assign addr[46179]= -931758235;
assign addr[46180]= -1067110699;
assign addr[46181]= -1197050035;
assign addr[46182]= -1320917099;
assign addr[46183]= -1438083551;
assign addr[46184]= -1547955041;
assign addr[46185]= -1649974225;
assign addr[46186]= -1743623590;
assign addr[46187]= -1828428082;
assign addr[46188]= -1903957513;
assign addr[46189]= -1969828744;
assign addr[46190]= -2025707632;
assign addr[46191]= -2071310720;
assign addr[46192]= -2106406677;
assign addr[46193]= -2130817471;
assign addr[46194]= -2144419275;
assign addr[46195]= -2147143090;
assign addr[46196]= -2138975100;
assign addr[46197]= -2119956737;
assign addr[46198]= -2090184478;
assign addr[46199]= -2049809346;
assign addr[46200]= -1999036154;
assign addr[46201]= -1938122457;
assign addr[46202]= -1867377253;
assign addr[46203]= -1787159411;
assign addr[46204]= -1697875851;
assign addr[46205]= -1599979481;
assign addr[46206]= -1493966902;
assign addr[46207]= -1380375881;
assign addr[46208]= -1259782632;
assign addr[46209]= -1132798888;
assign addr[46210]= -1000068799;
assign addr[46211]= -862265664;
assign addr[46212]= -720088517;
assign addr[46213]= -574258580;
assign addr[46214]= -425515602;
assign addr[46215]= -274614114;
assign addr[46216]= -122319591;
assign addr[46217]= 30595422;
assign addr[46218]= 183355234;
assign addr[46219]= 335184940;
assign addr[46220]= 485314355;
assign addr[46221]= 632981917;
assign addr[46222]= 777438554;
assign addr[46223]= 917951481;
assign addr[46224]= 1053807919;
assign addr[46225]= 1184318708;
assign addr[46226]= 1308821808;
assign addr[46227]= 1426685652;
assign addr[46228]= 1537312353;
assign addr[46229]= 1640140734;
assign addr[46230]= 1734649179;
assign addr[46231]= 1820358275;
assign addr[46232]= 1896833245;
assign addr[46233]= 1963686155;
assign addr[46234]= 2020577882;
assign addr[46235]= 2067219829;
assign addr[46236]= 2103375398;
assign addr[46237]= 2128861181;
assign addr[46238]= 2143547897;
assign addr[46239]= 2147361045;
assign addr[46240]= 2140281282;
assign addr[46241]= 2122344521;
assign addr[46242]= 2093641749;
assign addr[46243]= 2054318569;
assign addr[46244]= 2004574453;
assign addr[46245]= 1944661739;
assign addr[46246]= 1874884346;
assign addr[46247]= 1795596234;
assign addr[46248]= 1707199606;
assign addr[46249]= 1610142873;
assign addr[46250]= 1504918373;
assign addr[46251]= 1392059879;
assign addr[46252]= 1272139887;
assign addr[46253]= 1145766716;
assign addr[46254]= 1013581418;
assign addr[46255]= 876254528;
assign addr[46256]= 734482665;
assign addr[46257]= 588984994;
assign addr[46258]= 440499581;
assign addr[46259]= 289779648;
assign addr[46260]= 137589750;
assign addr[46261]= -15298099;
assign addr[46262]= -168108346;
assign addr[46263]= -320065829;
assign addr[46264]= -470399716;
assign addr[46265]= -618347408;
assign addr[46266]= -763158411;
assign addr[46267]= -904098143;
assign addr[46268]= -1040451659;
assign addr[46269]= -1171527280;
assign addr[46270]= -1296660098;
assign addr[46271]= -1415215352;
assign addr[46272]= -1526591649;
assign addr[46273]= -1630224009;
assign addr[46274]= -1725586737;
assign addr[46275]= -1812196087;
assign addr[46276]= -1889612716;
assign addr[46277]= -1957443913;
assign addr[46278]= -2015345591;
assign addr[46279]= -2063024031;
assign addr[46280]= -2100237377;
assign addr[46281]= -2126796855;
assign addr[46282]= -2142567738;
assign addr[46283]= -2147470025;
assign addr[46284]= -2141478848;
assign addr[46285]= -2124624598;
assign addr[46286]= -2096992772;
assign addr[46287]= -2058723538;
assign addr[46288]= -2010011024;
assign addr[46289]= -1951102334;
assign addr[46290]= -1882296293;
assign addr[46291]= -1803941934;
assign addr[46292]= -1716436725;
assign addr[46293]= -1620224553;
assign addr[46294]= -1515793473;
assign addr[46295]= -1403673233;
assign addr[46296]= -1284432584;
assign addr[46297]= -1158676398;
assign addr[46298]= -1027042599;
assign addr[46299]= -890198924;
assign addr[46300]= -748839539;
assign addr[46301]= -603681519;
assign addr[46302]= -455461206;
assign addr[46303]= -304930476;
assign addr[46304]= -152852926;
assign addr[46305]= 0;
assign addr[46306]= 152852926;
assign addr[46307]= 304930476;
assign addr[46308]= 455461206;
assign addr[46309]= 603681519;
assign addr[46310]= 748839539;
assign addr[46311]= 890198924;
assign addr[46312]= 1027042599;
assign addr[46313]= 1158676398;
assign addr[46314]= 1284432584;
assign addr[46315]= 1403673233;
assign addr[46316]= 1515793473;
assign addr[46317]= 1620224553;
assign addr[46318]= 1716436725;
assign addr[46319]= 1803941934;
assign addr[46320]= 1882296293;
assign addr[46321]= 1951102334;
assign addr[46322]= 2010011024;
assign addr[46323]= 2058723538;
assign addr[46324]= 2096992772;
assign addr[46325]= 2124624598;
assign addr[46326]= 2141478848;
assign addr[46327]= 2147470025;
assign addr[46328]= 2142567738;
assign addr[46329]= 2126796855;
assign addr[46330]= 2100237377;
assign addr[46331]= 2063024031;
assign addr[46332]= 2015345591;
assign addr[46333]= 1957443913;
assign addr[46334]= 1889612716;
assign addr[46335]= 1812196087;
assign addr[46336]= 1725586737;
assign addr[46337]= 1630224009;
assign addr[46338]= 1526591649;
assign addr[46339]= 1415215352;
assign addr[46340]= 1296660098;
assign addr[46341]= 1171527280;
assign addr[46342]= 1040451659;
assign addr[46343]= 904098143;
assign addr[46344]= 763158411;
assign addr[46345]= 618347408;
assign addr[46346]= 470399716;
assign addr[46347]= 320065829;
assign addr[46348]= 168108346;
assign addr[46349]= 15298099;
assign addr[46350]= -137589750;
assign addr[46351]= -289779648;
assign addr[46352]= -440499581;
assign addr[46353]= -588984994;
assign addr[46354]= -734482665;
assign addr[46355]= -876254528;
assign addr[46356]= -1013581418;
assign addr[46357]= -1145766716;
assign addr[46358]= -1272139887;
assign addr[46359]= -1392059879;
assign addr[46360]= -1504918373;
assign addr[46361]= -1610142873;
assign addr[46362]= -1707199606;
assign addr[46363]= -1795596234;
assign addr[46364]= -1874884346;
assign addr[46365]= -1944661739;
assign addr[46366]= -2004574453;
assign addr[46367]= -2054318569;
assign addr[46368]= -2093641749;
assign addr[46369]= -2122344521;
assign addr[46370]= -2140281282;
assign addr[46371]= -2147361045;
assign addr[46372]= -2143547897;
assign addr[46373]= -2128861181;
assign addr[46374]= -2103375398;
assign addr[46375]= -2067219829;
assign addr[46376]= -2020577882;
assign addr[46377]= -1963686155;
assign addr[46378]= -1896833245;
assign addr[46379]= -1820358275;
assign addr[46380]= -1734649179;
assign addr[46381]= -1640140734;
assign addr[46382]= -1537312353;
assign addr[46383]= -1426685652;
assign addr[46384]= -1308821808;
assign addr[46385]= -1184318708;
assign addr[46386]= -1053807919;
assign addr[46387]= -917951481;
assign addr[46388]= -777438554;
assign addr[46389]= -632981917;
assign addr[46390]= -485314355;
assign addr[46391]= -335184940;
assign addr[46392]= -183355234;
assign addr[46393]= -30595422;
assign addr[46394]= 122319591;
assign addr[46395]= 274614114;
assign addr[46396]= 425515602;
assign addr[46397]= 574258580;
assign addr[46398]= 720088517;
assign addr[46399]= 862265664;
assign addr[46400]= 1000068799;
assign addr[46401]= 1132798888;
assign addr[46402]= 1259782632;
assign addr[46403]= 1380375881;
assign addr[46404]= 1493966902;
assign addr[46405]= 1599979481;
assign addr[46406]= 1697875851;
assign addr[46407]= 1787159411;
assign addr[46408]= 1867377253;
assign addr[46409]= 1938122457;
assign addr[46410]= 1999036154;
assign addr[46411]= 2049809346;
assign addr[46412]= 2090184478;
assign addr[46413]= 2119956737;
assign addr[46414]= 2138975100;
assign addr[46415]= 2147143090;
assign addr[46416]= 2144419275;
assign addr[46417]= 2130817471;
assign addr[46418]= 2106406677;
assign addr[46419]= 2071310720;
assign addr[46420]= 2025707632;
assign addr[46421]= 1969828744;
assign addr[46422]= 1903957513;
assign addr[46423]= 1828428082;
assign addr[46424]= 1743623590;
assign addr[46425]= 1649974225;
assign addr[46426]= 1547955041;
assign addr[46427]= 1438083551;
assign addr[46428]= 1320917099;
assign addr[46429]= 1197050035;
assign addr[46430]= 1067110699;
assign addr[46431]= 931758235;
assign addr[46432]= 791679244;
assign addr[46433]= 647584304;
assign addr[46434]= 500204365;
assign addr[46435]= 350287041;
assign addr[46436]= 198592817;
assign addr[46437]= 45891193;
assign addr[46438]= -107043224;
assign addr[46439]= -259434643;
assign addr[46440]= -410510029;
assign addr[46441]= -559503022;
assign addr[46442]= -705657826;
assign addr[46443]= -848233042;
assign addr[46444]= -986505429;
assign addr[46445]= -1119773573;
assign addr[46446]= -1247361445;
assign addr[46447]= -1368621831;
assign addr[46448]= -1482939614;
assign addr[46449]= -1589734894;
assign addr[46450]= -1688465931;
assign addr[46451]= -1778631892;
assign addr[46452]= -1859775393;
assign addr[46453]= -1931484818;
assign addr[46454]= -1993396407;
assign addr[46455]= -2045196100;
assign addr[46456]= -2086621133;
assign addr[46457]= -2117461370;
assign addr[46458]= -2137560369;
assign addr[46459]= -2146816171;
assign addr[46460]= -2145181827;
assign addr[46461]= -2132665626;
assign addr[46462]= -2109331059;
assign addr[46463]= -2075296495;
assign addr[46464]= -2030734582;
assign addr[46465]= -1975871368;
assign addr[46466]= -1910985158;
assign addr[46467]= -1836405100;
assign addr[46468]= -1752509516;
assign addr[46469]= -1659723983;
assign addr[46470]= -1558519173;
assign addr[46471]= -1449408469;
assign addr[46472]= -1332945355;
assign addr[46473]= -1209720613;
assign addr[46474]= -1080359326;
assign addr[46475]= -945517704;
assign addr[46476]= -805879757;
assign addr[46477]= -662153826;
assign addr[46478]= -515068990;
assign addr[46479]= -365371365;
assign addr[46480]= -213820322;
assign addr[46481]= -61184634;
assign addr[46482]= 91761426;
assign addr[46483]= 244242007;
assign addr[46484]= 395483624;
assign addr[46485]= 544719071;
assign addr[46486]= 691191324;
assign addr[46487]= 834157373;
assign addr[46488]= 972891995;
assign addr[46489]= 1106691431;
assign addr[46490]= 1234876957;
assign addr[46491]= 1356798326;
assign addr[46492]= 1471837070;
assign addr[46493]= 1579409630;
assign addr[46494]= 1678970324;
assign addr[46495]= 1770014111;
assign addr[46496]= 1852079154;
assign addr[46497]= 1924749160;
assign addr[46498]= 1987655498;
assign addr[46499]= 2040479063;
assign addr[46500]= 2082951896;
assign addr[46501]= 2114858546;
assign addr[46502]= 2136037160;
assign addr[46503]= 2146380306;
assign addr[46504]= 2145835515;
assign addr[46505]= 2134405552;
assign addr[46506]= 2112148396;
assign addr[46507]= 2079176953;
assign addr[46508]= 2035658475;
assign addr[46509]= 1981813720;
assign addr[46510]= 1917915825;
assign addr[46511]= 1844288924;
assign addr[46512]= 1761306505;
assign addr[46513]= 1669389513;
assign addr[46514]= 1569004214;
assign addr[46515]= 1460659832;
assign addr[46516]= 1344905966;
assign addr[46517]= 1222329801;
assign addr[46518]= 1093553126;
assign addr[46519]= 959229189;
assign addr[46520]= 820039373;
assign addr[46521]= 676689746;
assign addr[46522]= 529907477;
assign addr[46523]= 380437148;
assign addr[46524]= 229036977;
assign addr[46525]= 76474970;
assign addr[46526]= -76474970;
assign addr[46527]= -229036977;
assign addr[46528]= -380437148;
assign addr[46529]= -529907477;
assign addr[46530]= -676689746;
assign addr[46531]= -820039373;
assign addr[46532]= -959229189;
assign addr[46533]= -1093553126;
assign addr[46534]= -1222329801;
assign addr[46535]= -1344905966;
assign addr[46536]= -1460659832;
assign addr[46537]= -1569004214;
assign addr[46538]= -1669389513;
assign addr[46539]= -1761306505;
assign addr[46540]= -1844288924;
assign addr[46541]= -1917915825;
assign addr[46542]= -1981813720;
assign addr[46543]= -2035658475;
assign addr[46544]= -2079176953;
assign addr[46545]= -2112148396;
assign addr[46546]= -2134405552;
assign addr[46547]= -2145835515;
assign addr[46548]= -2146380306;
assign addr[46549]= -2136037160;
assign addr[46550]= -2114858546;
assign addr[46551]= -2082951896;
assign addr[46552]= -2040479063;
assign addr[46553]= -1987655498;
assign addr[46554]= -1924749160;
assign addr[46555]= -1852079154;
assign addr[46556]= -1770014111;
assign addr[46557]= -1678970324;
assign addr[46558]= -1579409630;
assign addr[46559]= -1471837070;
assign addr[46560]= -1356798326;
assign addr[46561]= -1234876957;
assign addr[46562]= -1106691431;
assign addr[46563]= -972891995;
assign addr[46564]= -834157373;
assign addr[46565]= -691191324;
assign addr[46566]= -544719071;
assign addr[46567]= -395483624;
assign addr[46568]= -244242007;
assign addr[46569]= -91761426;
assign addr[46570]= 61184634;
assign addr[46571]= 213820322;
assign addr[46572]= 365371365;
assign addr[46573]= 515068990;
assign addr[46574]= 662153826;
assign addr[46575]= 805879757;
assign addr[46576]= 945517704;
assign addr[46577]= 1080359326;
assign addr[46578]= 1209720613;
assign addr[46579]= 1332945355;
assign addr[46580]= 1449408469;
assign addr[46581]= 1558519173;
assign addr[46582]= 1659723983;
assign addr[46583]= 1752509516;
assign addr[46584]= 1836405100;
assign addr[46585]= 1910985158;
assign addr[46586]= 1975871368;
assign addr[46587]= 2030734582;
assign addr[46588]= 2075296495;
assign addr[46589]= 2109331059;
assign addr[46590]= 2132665626;
assign addr[46591]= 2145181827;
assign addr[46592]= 2146816171;
assign addr[46593]= 2137560369;
assign addr[46594]= 2117461370;
assign addr[46595]= 2086621133;
assign addr[46596]= 2045196100;
assign addr[46597]= 1993396407;
assign addr[46598]= 1931484818;
assign addr[46599]= 1859775393;
assign addr[46600]= 1778631892;
assign addr[46601]= 1688465931;
assign addr[46602]= 1589734894;
assign addr[46603]= 1482939614;
assign addr[46604]= 1368621831;
assign addr[46605]= 1247361445;
assign addr[46606]= 1119773573;
assign addr[46607]= 986505429;
assign addr[46608]= 848233042;
assign addr[46609]= 705657826;
assign addr[46610]= 559503022;
assign addr[46611]= 410510029;
assign addr[46612]= 259434643;
assign addr[46613]= 107043224;
assign addr[46614]= -45891193;
assign addr[46615]= -198592817;
assign addr[46616]= -350287041;
assign addr[46617]= -500204365;
assign addr[46618]= -647584304;
assign addr[46619]= -791679244;
assign addr[46620]= -931758235;
assign addr[46621]= -1067110699;
assign addr[46622]= -1197050035;
assign addr[46623]= -1320917099;
assign addr[46624]= -1438083551;
assign addr[46625]= -1547955041;
assign addr[46626]= -1649974225;
assign addr[46627]= -1743623590;
assign addr[46628]= -1828428082;
assign addr[46629]= -1903957513;
assign addr[46630]= -1969828744;
assign addr[46631]= -2025707632;
assign addr[46632]= -2071310720;
assign addr[46633]= -2106406677;
assign addr[46634]= -2130817471;
assign addr[46635]= -2144419275;
assign addr[46636]= -2147143090;
assign addr[46637]= -2138975100;
assign addr[46638]= -2119956737;
assign addr[46639]= -2090184478;
assign addr[46640]= -2049809346;
assign addr[46641]= -1999036154;
assign addr[46642]= -1938122457;
assign addr[46643]= -1867377253;
assign addr[46644]= -1787159411;
assign addr[46645]= -1697875851;
assign addr[46646]= -1599979481;
assign addr[46647]= -1493966902;
assign addr[46648]= -1380375881;
assign addr[46649]= -1259782632;
assign addr[46650]= -1132798888;
assign addr[46651]= -1000068799;
assign addr[46652]= -862265664;
assign addr[46653]= -720088517;
assign addr[46654]= -574258580;
assign addr[46655]= -425515602;
assign addr[46656]= -274614114;
assign addr[46657]= -122319591;
assign addr[46658]= 30595422;
assign addr[46659]= 183355234;
assign addr[46660]= 335184940;
assign addr[46661]= 485314355;
assign addr[46662]= 632981917;
assign addr[46663]= 777438554;
assign addr[46664]= 917951481;
assign addr[46665]= 1053807919;
assign addr[46666]= 1184318708;
assign addr[46667]= 1308821808;
assign addr[46668]= 1426685652;
assign addr[46669]= 1537312353;
assign addr[46670]= 1640140734;
assign addr[46671]= 1734649179;
assign addr[46672]= 1820358275;
assign addr[46673]= 1896833245;
assign addr[46674]= 1963686155;
assign addr[46675]= 2020577882;
assign addr[46676]= 2067219829;
assign addr[46677]= 2103375398;
assign addr[46678]= 2128861181;
assign addr[46679]= 2143547897;
assign addr[46680]= 2147361045;
assign addr[46681]= 2140281282;
assign addr[46682]= 2122344521;
assign addr[46683]= 2093641749;
assign addr[46684]= 2054318569;
assign addr[46685]= 2004574453;
assign addr[46686]= 1944661739;
assign addr[46687]= 1874884346;
assign addr[46688]= 1795596234;
assign addr[46689]= 1707199606;
assign addr[46690]= 1610142873;
assign addr[46691]= 1504918373;
assign addr[46692]= 1392059879;
assign addr[46693]= 1272139887;
assign addr[46694]= 1145766716;
assign addr[46695]= 1013581418;
assign addr[46696]= 876254528;
assign addr[46697]= 734482665;
assign addr[46698]= 588984994;
assign addr[46699]= 440499581;
assign addr[46700]= 289779648;
assign addr[46701]= 137589750;
assign addr[46702]= -15298099;
assign addr[46703]= -168108346;
assign addr[46704]= -320065829;
assign addr[46705]= -470399716;
assign addr[46706]= -618347408;
assign addr[46707]= -763158411;
assign addr[46708]= -904098143;
assign addr[46709]= -1040451659;
assign addr[46710]= -1171527280;
assign addr[46711]= -1296660098;
assign addr[46712]= -1415215352;
assign addr[46713]= -1526591649;
assign addr[46714]= -1630224009;
assign addr[46715]= -1725586737;
assign addr[46716]= -1812196087;
assign addr[46717]= -1889612716;
assign addr[46718]= -1957443913;
assign addr[46719]= -2015345591;
assign addr[46720]= -2063024031;
assign addr[46721]= -2100237377;
assign addr[46722]= -2126796855;
assign addr[46723]= -2142567738;
assign addr[46724]= -2147470025;
assign addr[46725]= -2141478848;
assign addr[46726]= -2124624598;
assign addr[46727]= -2096992772;
assign addr[46728]= -2058723538;
assign addr[46729]= -2010011024;
assign addr[46730]= -1951102334;
assign addr[46731]= -1882296293;
assign addr[46732]= -1803941934;
assign addr[46733]= -1716436725;
assign addr[46734]= -1620224553;
assign addr[46735]= -1515793473;
assign addr[46736]= -1403673233;
assign addr[46737]= -1284432584;
assign addr[46738]= -1158676398;
assign addr[46739]= -1027042599;
assign addr[46740]= -890198924;
assign addr[46741]= -748839539;
assign addr[46742]= -603681519;
assign addr[46743]= -455461206;
assign addr[46744]= -304930476;
assign addr[46745]= -152852926;
assign addr[46746]= 0;
assign addr[46747]= 152852926;
assign addr[46748]= 304930476;
assign addr[46749]= 455461206;
assign addr[46750]= 603681519;
assign addr[46751]= 748839539;
assign addr[46752]= 890198924;
assign addr[46753]= 1027042599;
assign addr[46754]= 1158676398;
assign addr[46755]= 1284432584;
assign addr[46756]= 1403673233;
assign addr[46757]= 1515793473;
assign addr[46758]= 1620224553;
assign addr[46759]= 1716436725;
assign addr[46760]= 1803941934;
assign addr[46761]= 1882296293;
assign addr[46762]= 1951102334;
assign addr[46763]= 2010011024;
assign addr[46764]= 2058723538;
assign addr[46765]= 2096992772;
assign addr[46766]= 2124624598;
assign addr[46767]= 2141478848;
assign addr[46768]= 2147470025;
assign addr[46769]= 2142567738;
assign addr[46770]= 2126796855;
assign addr[46771]= 2100237377;
assign addr[46772]= 2063024031;
assign addr[46773]= 2015345591;
assign addr[46774]= 1957443913;
assign addr[46775]= 1889612716;
assign addr[46776]= 1812196087;
assign addr[46777]= 1725586737;
assign addr[46778]= 1630224009;
assign addr[46779]= 1526591649;
assign addr[46780]= 1415215352;
assign addr[46781]= 1296660098;
assign addr[46782]= 1171527280;
assign addr[46783]= 1040451659;
assign addr[46784]= 904098143;
assign addr[46785]= 763158411;
assign addr[46786]= 618347408;
assign addr[46787]= 470399716;
assign addr[46788]= 320065829;
assign addr[46789]= 168108346;
assign addr[46790]= 15298099;
assign addr[46791]= -137589750;
assign addr[46792]= -289779648;
assign addr[46793]= -440499581;
assign addr[46794]= -588984994;
assign addr[46795]= -734482665;
assign addr[46796]= -876254528;
assign addr[46797]= -1013581418;
assign addr[46798]= -1145766716;
assign addr[46799]= -1272139887;
assign addr[46800]= -1392059879;
assign addr[46801]= -1504918373;
assign addr[46802]= -1610142873;
assign addr[46803]= -1707199606;
assign addr[46804]= -1795596234;
assign addr[46805]= -1874884346;
assign addr[46806]= -1944661739;
assign addr[46807]= -2004574453;
assign addr[46808]= -2054318569;
assign addr[46809]= -2093641749;
assign addr[46810]= -2122344521;
assign addr[46811]= -2140281282;
assign addr[46812]= -2147361045;
assign addr[46813]= -2143547897;
assign addr[46814]= -2128861181;
assign addr[46815]= -2103375398;
assign addr[46816]= -2067219829;
assign addr[46817]= -2020577882;
assign addr[46818]= -1963686155;
assign addr[46819]= -1896833245;
assign addr[46820]= -1820358275;
assign addr[46821]= -1734649179;
assign addr[46822]= -1640140734;
assign addr[46823]= -1537312353;
assign addr[46824]= -1426685652;
assign addr[46825]= -1308821808;
assign addr[46826]= -1184318708;
assign addr[46827]= -1053807919;
assign addr[46828]= -917951481;
assign addr[46829]= -777438554;
assign addr[46830]= -632981917;
assign addr[46831]= -485314355;
assign addr[46832]= -335184940;
assign addr[46833]= -183355234;
assign addr[46834]= -30595422;
assign addr[46835]= 122319591;
assign addr[46836]= 274614114;
assign addr[46837]= 425515602;
assign addr[46838]= 574258580;
assign addr[46839]= 720088517;
assign addr[46840]= 862265664;
assign addr[46841]= 1000068799;
assign addr[46842]= 1132798888;
assign addr[46843]= 1259782632;
assign addr[46844]= 1380375881;
assign addr[46845]= 1493966902;
assign addr[46846]= 1599979481;
assign addr[46847]= 1697875851;
assign addr[46848]= 1787159411;
assign addr[46849]= 1867377253;
assign addr[46850]= 1938122457;
assign addr[46851]= 1999036154;
assign addr[46852]= 2049809346;
assign addr[46853]= 2090184478;
assign addr[46854]= 2119956737;
assign addr[46855]= 2138975100;
assign addr[46856]= 2147143090;
assign addr[46857]= 2144419275;
assign addr[46858]= 2130817471;
assign addr[46859]= 2106406677;
assign addr[46860]= 2071310720;
assign addr[46861]= 2025707632;
assign addr[46862]= 1969828744;
assign addr[46863]= 1903957513;
assign addr[46864]= 1828428082;
assign addr[46865]= 1743623590;
assign addr[46866]= 1649974225;
assign addr[46867]= 1547955041;
assign addr[46868]= 1438083551;
assign addr[46869]= 1320917099;
assign addr[46870]= 1197050035;
assign addr[46871]= 1067110699;
assign addr[46872]= 931758235;
assign addr[46873]= 791679244;
assign addr[46874]= 647584304;
assign addr[46875]= 500204365;
assign addr[46876]= 350287041;
assign addr[46877]= 198592817;
assign addr[46878]= 45891193;
assign addr[46879]= -107043224;
assign addr[46880]= -259434643;
assign addr[46881]= -410510029;
assign addr[46882]= -559503022;
assign addr[46883]= -705657826;
assign addr[46884]= -848233042;
assign addr[46885]= -986505429;
assign addr[46886]= -1119773573;
assign addr[46887]= -1247361445;
assign addr[46888]= -1368621831;
assign addr[46889]= -1482939614;
assign addr[46890]= -1589734894;
assign addr[46891]= -1688465931;
assign addr[46892]= -1778631892;
assign addr[46893]= -1859775393;
assign addr[46894]= -1931484818;
assign addr[46895]= -1993396407;
assign addr[46896]= -2045196100;
assign addr[46897]= -2086621133;
assign addr[46898]= -2117461370;
assign addr[46899]= -2137560369;
assign addr[46900]= -2146816171;
assign addr[46901]= -2145181827;
assign addr[46902]= -2132665626;
assign addr[46903]= -2109331059;
assign addr[46904]= -2075296495;
assign addr[46905]= -2030734582;
assign addr[46906]= -1975871368;
assign addr[46907]= -1910985158;
assign addr[46908]= -1836405100;
assign addr[46909]= -1752509516;
assign addr[46910]= -1659723983;
assign addr[46911]= -1558519173;
assign addr[46912]= -1449408469;
assign addr[46913]= -1332945355;
assign addr[46914]= -1209720613;
assign addr[46915]= -1080359326;
assign addr[46916]= -945517704;
assign addr[46917]= -805879757;
assign addr[46918]= -662153826;
assign addr[46919]= -515068990;
assign addr[46920]= -365371365;
assign addr[46921]= -213820322;
assign addr[46922]= -61184634;
assign addr[46923]= 91761426;
assign addr[46924]= 244242007;
assign addr[46925]= 395483624;
assign addr[46926]= 544719071;
assign addr[46927]= 691191324;
assign addr[46928]= 834157373;
assign addr[46929]= 972891995;
assign addr[46930]= 1106691431;
assign addr[46931]= 1234876957;
assign addr[46932]= 1356798326;
assign addr[46933]= 1471837070;
assign addr[46934]= 1579409630;
assign addr[46935]= 1678970324;
assign addr[46936]= 1770014111;
assign addr[46937]= 1852079154;
assign addr[46938]= 1924749160;
assign addr[46939]= 1987655498;
assign addr[46940]= 2040479063;
assign addr[46941]= 2082951896;
assign addr[46942]= 2114858546;
assign addr[46943]= 2136037160;
assign addr[46944]= 2146380306;
assign addr[46945]= 2145835515;
assign addr[46946]= 2134405552;
assign addr[46947]= 2112148396;
assign addr[46948]= 2079176953;
assign addr[46949]= 2035658475;
assign addr[46950]= 1981813720;
assign addr[46951]= 1917915825;
assign addr[46952]= 1844288924;
assign addr[46953]= 1761306505;
assign addr[46954]= 1669389513;
assign addr[46955]= 1569004214;
assign addr[46956]= 1460659832;
assign addr[46957]= 1344905966;
assign addr[46958]= 1222329801;
assign addr[46959]= 1093553126;
assign addr[46960]= 959229189;
assign addr[46961]= 820039373;
assign addr[46962]= 676689746;
assign addr[46963]= 529907477;
assign addr[46964]= 380437148;
assign addr[46965]= 229036977;
assign addr[46966]= 76474970;
assign addr[46967]= -76474970;
assign addr[46968]= -229036977;
assign addr[46969]= -380437148;
assign addr[46970]= -529907477;
assign addr[46971]= -676689746;
assign addr[46972]= -820039373;
assign addr[46973]= -959229189;
assign addr[46974]= -1093553126;
assign addr[46975]= -1222329801;
assign addr[46976]= -1344905966;
assign addr[46977]= -1460659832;
assign addr[46978]= -1569004214;
assign addr[46979]= -1669389513;
assign addr[46980]= -1761306505;
assign addr[46981]= -1844288924;
assign addr[46982]= -1917915825;
assign addr[46983]= -1981813720;
assign addr[46984]= -2035658475;
assign addr[46985]= -2079176953;
assign addr[46986]= -2112148396;
assign addr[46987]= -2134405552;
assign addr[46988]= -2145835515;
assign addr[46989]= -2146380306;
assign addr[46990]= -2136037160;
assign addr[46991]= -2114858546;
assign addr[46992]= -2082951896;
assign addr[46993]= -2040479063;
assign addr[46994]= -1987655498;
assign addr[46995]= -1924749160;
assign addr[46996]= -1852079154;
assign addr[46997]= -1770014111;
assign addr[46998]= -1678970324;
assign addr[46999]= -1579409630;
assign addr[47000]= -1471837070;
assign addr[47001]= -1356798326;
assign addr[47002]= -1234876957;
assign addr[47003]= -1106691431;
assign addr[47004]= -972891995;
assign addr[47005]= -834157373;
assign addr[47006]= -691191324;
assign addr[47007]= -544719071;
assign addr[47008]= -395483624;
assign addr[47009]= -244242007;
assign addr[47010]= -91761426;
assign addr[47011]= 61184634;
assign addr[47012]= 213820322;
assign addr[47013]= 365371365;
assign addr[47014]= 515068990;
assign addr[47015]= 662153826;
assign addr[47016]= 805879757;
assign addr[47017]= 945517704;
assign addr[47018]= 1080359326;
assign addr[47019]= 1209720613;
assign addr[47020]= 1332945355;
assign addr[47021]= 1449408469;
assign addr[47022]= 1558519173;
assign addr[47023]= 1659723983;
assign addr[47024]= 1752509516;
assign addr[47025]= 1836405100;
assign addr[47026]= 1910985158;
assign addr[47027]= 1975871368;
assign addr[47028]= 2030734582;
assign addr[47029]= 2075296495;
assign addr[47030]= 2109331059;
assign addr[47031]= 2132665626;
assign addr[47032]= 2145181827;
assign addr[47033]= 2146816171;
assign addr[47034]= 2137560369;
assign addr[47035]= 2117461370;
assign addr[47036]= 2086621133;
assign addr[47037]= 2045196100;
assign addr[47038]= 1993396407;
assign addr[47039]= 1931484818;
assign addr[47040]= 1859775393;
assign addr[47041]= 1778631892;
assign addr[47042]= 1688465931;
assign addr[47043]= 1589734894;
assign addr[47044]= 1482939614;
assign addr[47045]= 1368621831;
assign addr[47046]= 1247361445;
assign addr[47047]= 1119773573;
assign addr[47048]= 986505429;
assign addr[47049]= 848233042;
assign addr[47050]= 705657826;
assign addr[47051]= 559503022;
assign addr[47052]= 410510029;
assign addr[47053]= 259434643;
assign addr[47054]= 107043224;
assign addr[47055]= -45891193;
assign addr[47056]= -198592817;
assign addr[47057]= -350287041;
assign addr[47058]= -500204365;
assign addr[47059]= -647584304;
assign addr[47060]= -791679244;
assign addr[47061]= -931758235;
assign addr[47062]= -1067110699;
assign addr[47063]= -1197050035;
assign addr[47064]= -1320917099;
assign addr[47065]= -1438083551;
assign addr[47066]= -1547955041;
assign addr[47067]= -1649974225;
assign addr[47068]= -1743623590;
assign addr[47069]= -1828428082;
assign addr[47070]= -1903957513;
assign addr[47071]= -1969828744;
assign addr[47072]= -2025707632;
assign addr[47073]= -2071310720;
assign addr[47074]= -2106406677;
assign addr[47075]= -2130817471;
assign addr[47076]= -2144419275;
assign addr[47077]= -2147143090;
assign addr[47078]= -2138975100;
assign addr[47079]= -2119956737;
assign addr[47080]= -2090184478;
assign addr[47081]= -2049809346;
assign addr[47082]= -1999036154;
assign addr[47083]= -1938122457;
assign addr[47084]= -1867377253;
assign addr[47085]= -1787159411;
assign addr[47086]= -1697875851;
assign addr[47087]= -1599979481;
assign addr[47088]= -1493966902;
assign addr[47089]= -1380375881;
assign addr[47090]= -1259782632;
assign addr[47091]= -1132798888;
assign addr[47092]= -1000068799;
assign addr[47093]= -862265664;
assign addr[47094]= -720088517;
assign addr[47095]= -574258580;
assign addr[47096]= -425515602;
assign addr[47097]= -274614114;
assign addr[47098]= -122319591;
assign addr[47099]= 30595422;
assign addr[47100]= 183355234;
assign addr[47101]= 335184940;
assign addr[47102]= 485314355;
assign addr[47103]= 632981917;
assign addr[47104]= 777438554;
assign addr[47105]= 917951481;
assign addr[47106]= 1053807919;
assign addr[47107]= 1184318708;
assign addr[47108]= 1308821808;
assign addr[47109]= 1426685652;
assign addr[47110]= 1537312353;
assign addr[47111]= 1640140734;
assign addr[47112]= 1734649179;
assign addr[47113]= 1820358275;
assign addr[47114]= 1896833245;
assign addr[47115]= 1963686155;
assign addr[47116]= 2020577882;
assign addr[47117]= 2067219829;
assign addr[47118]= 2103375398;
assign addr[47119]= 2128861181;
assign addr[47120]= 2143547897;
assign addr[47121]= 2147361045;
assign addr[47122]= 2140281282;
assign addr[47123]= 2122344521;
assign addr[47124]= 2093641749;
assign addr[47125]= 2054318569;
assign addr[47126]= 2004574453;
assign addr[47127]= 1944661739;
assign addr[47128]= 1874884346;
assign addr[47129]= 1795596234;
assign addr[47130]= 1707199606;
assign addr[47131]= 1610142873;
assign addr[47132]= 1504918373;
assign addr[47133]= 1392059879;
assign addr[47134]= 1272139887;
assign addr[47135]= 1145766716;
assign addr[47136]= 1013581418;
assign addr[47137]= 876254528;
assign addr[47138]= 734482665;
assign addr[47139]= 588984994;
assign addr[47140]= 440499581;
assign addr[47141]= 289779648;
assign addr[47142]= 137589750;
assign addr[47143]= -15298099;
assign addr[47144]= -168108346;
assign addr[47145]= -320065829;
assign addr[47146]= -470399716;
assign addr[47147]= -618347408;
assign addr[47148]= -763158411;
assign addr[47149]= -904098143;
assign addr[47150]= -1040451659;
assign addr[47151]= -1171527280;
assign addr[47152]= -1296660098;
assign addr[47153]= -1415215352;
assign addr[47154]= -1526591649;
assign addr[47155]= -1630224009;
assign addr[47156]= -1725586737;
assign addr[47157]= -1812196087;
assign addr[47158]= -1889612716;
assign addr[47159]= -1957443913;
assign addr[47160]= -2015345591;
assign addr[47161]= -2063024031;
assign addr[47162]= -2100237377;
assign addr[47163]= -2126796855;
assign addr[47164]= -2142567738;
assign addr[47165]= -2147470025;
assign addr[47166]= -2141478848;
assign addr[47167]= -2124624598;
assign addr[47168]= -2096992772;
assign addr[47169]= -2058723538;
assign addr[47170]= -2010011024;
assign addr[47171]= -1951102334;
assign addr[47172]= -1882296293;
assign addr[47173]= -1803941934;
assign addr[47174]= -1716436725;
assign addr[47175]= -1620224553;
assign addr[47176]= -1515793473;
assign addr[47177]= -1403673233;
assign addr[47178]= -1284432584;
assign addr[47179]= -1158676398;
assign addr[47180]= -1027042599;
assign addr[47181]= -890198924;
assign addr[47182]= -748839539;
assign addr[47183]= -603681519;
assign addr[47184]= -455461206;
assign addr[47185]= -304930476;
assign addr[47186]= -152852926;
assign addr[47187]= 0;
assign addr[47188]= 152852926;
assign addr[47189]= 304930476;
assign addr[47190]= 455461206;
assign addr[47191]= 603681519;
assign addr[47192]= 748839539;
assign addr[47193]= 890198924;
assign addr[47194]= 1027042599;
assign addr[47195]= 1158676398;
assign addr[47196]= 1284432584;
assign addr[47197]= 1403673233;
assign addr[47198]= 1515793473;
assign addr[47199]= 1620224553;
assign addr[47200]= 1716436725;
assign addr[47201]= 1803941934;
assign addr[47202]= 1882296293;
assign addr[47203]= 1951102334;
assign addr[47204]= 2010011024;
assign addr[47205]= 2058723538;
assign addr[47206]= 2096992772;
assign addr[47207]= 2124624598;
assign addr[47208]= 2141478848;
assign addr[47209]= 2147470025;
assign addr[47210]= 2142567738;
assign addr[47211]= 2126796855;
assign addr[47212]= 2100237377;
assign addr[47213]= 2063024031;
assign addr[47214]= 2015345591;
assign addr[47215]= 1957443913;
assign addr[47216]= 1889612716;
assign addr[47217]= 1812196087;
assign addr[47218]= 1725586737;
assign addr[47219]= 1630224009;
assign addr[47220]= 1526591649;
assign addr[47221]= 1415215352;
assign addr[47222]= 1296660098;
assign addr[47223]= 1171527280;
assign addr[47224]= 1040451659;
assign addr[47225]= 904098143;
assign addr[47226]= 763158411;
assign addr[47227]= 618347408;
assign addr[47228]= 470399716;
assign addr[47229]= 320065829;
assign addr[47230]= 168108346;
assign addr[47231]= 15298099;
assign addr[47232]= -137589750;
assign addr[47233]= -289779648;
assign addr[47234]= -440499581;
assign addr[47235]= -588984994;
assign addr[47236]= -734482665;
assign addr[47237]= -876254528;
assign addr[47238]= -1013581418;
assign addr[47239]= -1145766716;
assign addr[47240]= -1272139887;
assign addr[47241]= -1392059879;
assign addr[47242]= -1504918373;
assign addr[47243]= -1610142873;
assign addr[47244]= -1707199606;
assign addr[47245]= -1795596234;
assign addr[47246]= -1874884346;
assign addr[47247]= -1944661739;
assign addr[47248]= -2004574453;
assign addr[47249]= -2054318569;
assign addr[47250]= -2093641749;
assign addr[47251]= -2122344521;
assign addr[47252]= -2140281282;
assign addr[47253]= -2147361045;
assign addr[47254]= -2143547897;
assign addr[47255]= -2128861181;
assign addr[47256]= -2103375398;
assign addr[47257]= -2067219829;
assign addr[47258]= -2020577882;
assign addr[47259]= -1963686155;
assign addr[47260]= -1896833245;
assign addr[47261]= -1820358275;
assign addr[47262]= -1734649179;
assign addr[47263]= -1640140734;
assign addr[47264]= -1537312353;
assign addr[47265]= -1426685652;
assign addr[47266]= -1308821808;
assign addr[47267]= -1184318708;
assign addr[47268]= -1053807919;
assign addr[47269]= -917951481;
assign addr[47270]= -777438554;
assign addr[47271]= -632981917;
assign addr[47272]= -485314355;
assign addr[47273]= -335184940;
assign addr[47274]= -183355234;
assign addr[47275]= -30595422;
assign addr[47276]= 122319591;
assign addr[47277]= 274614114;
assign addr[47278]= 425515602;
assign addr[47279]= 574258580;
assign addr[47280]= 720088517;
assign addr[47281]= 862265664;
assign addr[47282]= 1000068799;
assign addr[47283]= 1132798888;
assign addr[47284]= 1259782632;
assign addr[47285]= 1380375881;
assign addr[47286]= 1493966902;
assign addr[47287]= 1599979481;
assign addr[47288]= 1697875851;
assign addr[47289]= 1787159411;
assign addr[47290]= 1867377253;
assign addr[47291]= 1938122457;
assign addr[47292]= 1999036154;
assign addr[47293]= 2049809346;
assign addr[47294]= 2090184478;
assign addr[47295]= 2119956737;
assign addr[47296]= 2138975100;
assign addr[47297]= 2147143090;
assign addr[47298]= 2144419275;
assign addr[47299]= 2130817471;
assign addr[47300]= 2106406677;
assign addr[47301]= 2071310720;
assign addr[47302]= 2025707632;
assign addr[47303]= 1969828744;
assign addr[47304]= 1903957513;
assign addr[47305]= 1828428082;
assign addr[47306]= 1743623590;
assign addr[47307]= 1649974225;
assign addr[47308]= 1547955041;
assign addr[47309]= 1438083551;
assign addr[47310]= 1320917099;
assign addr[47311]= 1197050035;
assign addr[47312]= 1067110699;
assign addr[47313]= 931758235;
assign addr[47314]= 791679244;
assign addr[47315]= 647584304;
assign addr[47316]= 500204365;
assign addr[47317]= 350287041;
assign addr[47318]= 198592817;
assign addr[47319]= 45891193;
assign addr[47320]= -107043224;
assign addr[47321]= -259434643;
assign addr[47322]= -410510029;
assign addr[47323]= -559503022;
assign addr[47324]= -705657826;
assign addr[47325]= -848233042;
assign addr[47326]= -986505429;
assign addr[47327]= -1119773573;
assign addr[47328]= -1247361445;
assign addr[47329]= -1368621831;
assign addr[47330]= -1482939614;
assign addr[47331]= -1589734894;
assign addr[47332]= -1688465931;
assign addr[47333]= -1778631892;
assign addr[47334]= -1859775393;
assign addr[47335]= -1931484818;
assign addr[47336]= -1993396407;
assign addr[47337]= -2045196100;
assign addr[47338]= -2086621133;
assign addr[47339]= -2117461370;
assign addr[47340]= -2137560369;
assign addr[47341]= -2146816171;
assign addr[47342]= -2145181827;
assign addr[47343]= -2132665626;
assign addr[47344]= -2109331059;
assign addr[47345]= -2075296495;
assign addr[47346]= -2030734582;
assign addr[47347]= -1975871368;
assign addr[47348]= -1910985158;
assign addr[47349]= -1836405100;
assign addr[47350]= -1752509516;
assign addr[47351]= -1659723983;
assign addr[47352]= -1558519173;
assign addr[47353]= -1449408469;
assign addr[47354]= -1332945355;
assign addr[47355]= -1209720613;
assign addr[47356]= -1080359326;
assign addr[47357]= -945517704;
assign addr[47358]= -805879757;
assign addr[47359]= -662153826;
assign addr[47360]= -515068990;
assign addr[47361]= -365371365;
assign addr[47362]= -213820322;
assign addr[47363]= -61184634;
assign addr[47364]= 91761426;
assign addr[47365]= 244242007;
assign addr[47366]= 395483624;
assign addr[47367]= 544719071;
assign addr[47368]= 691191324;
assign addr[47369]= 834157373;
assign addr[47370]= 972891995;
assign addr[47371]= 1106691431;
assign addr[47372]= 1234876957;
assign addr[47373]= 1356798326;
assign addr[47374]= 1471837070;
assign addr[47375]= 1579409630;
assign addr[47376]= 1678970324;
assign addr[47377]= 1770014111;
assign addr[47378]= 1852079154;
assign addr[47379]= 1924749160;
assign addr[47380]= 1987655498;
assign addr[47381]= 2040479063;
assign addr[47382]= 2082951896;
assign addr[47383]= 2114858546;
assign addr[47384]= 2136037160;
assign addr[47385]= 2146380306;
assign addr[47386]= 2145835515;
assign addr[47387]= 2134405552;
assign addr[47388]= 2112148396;
assign addr[47389]= 2079176953;
assign addr[47390]= 2035658475;
assign addr[47391]= 1981813720;
assign addr[47392]= 1917915825;
assign addr[47393]= 1844288924;
assign addr[47394]= 1761306505;
assign addr[47395]= 1669389513;
assign addr[47396]= 1569004214;
assign addr[47397]= 1460659832;
assign addr[47398]= 1344905966;
assign addr[47399]= 1222329801;
assign addr[47400]= 1093553126;
assign addr[47401]= 959229189;
assign addr[47402]= 820039373;
assign addr[47403]= 676689746;
assign addr[47404]= 529907477;
assign addr[47405]= 380437148;
assign addr[47406]= 229036977;
assign addr[47407]= 76474970;
assign addr[47408]= -76474970;
assign addr[47409]= -229036977;
assign addr[47410]= -380437148;
assign addr[47411]= -529907477;
assign addr[47412]= -676689746;
assign addr[47413]= -820039373;
assign addr[47414]= -959229189;
assign addr[47415]= -1093553126;
assign addr[47416]= -1222329801;
assign addr[47417]= -1344905966;
assign addr[47418]= -1460659832;
assign addr[47419]= -1569004214;
assign addr[47420]= -1669389513;
assign addr[47421]= -1761306505;
assign addr[47422]= -1844288924;
assign addr[47423]= -1917915825;
assign addr[47424]= -1981813720;
assign addr[47425]= -2035658475;
assign addr[47426]= -2079176953;
assign addr[47427]= -2112148396;
assign addr[47428]= -2134405552;
assign addr[47429]= -2145835515;
assign addr[47430]= -2146380306;
assign addr[47431]= -2136037160;
assign addr[47432]= -2114858546;
assign addr[47433]= -2082951896;
assign addr[47434]= -2040479063;
assign addr[47435]= -1987655498;
assign addr[47436]= -1924749160;
assign addr[47437]= -1852079154;
assign addr[47438]= -1770014111;
assign addr[47439]= -1678970324;
assign addr[47440]= -1579409630;
assign addr[47441]= -1471837070;
assign addr[47442]= -1356798326;
assign addr[47443]= -1234876957;
assign addr[47444]= -1106691431;
assign addr[47445]= -972891995;
assign addr[47446]= -834157373;
assign addr[47447]= -691191324;
assign addr[47448]= -544719071;
assign addr[47449]= -395483624;
assign addr[47450]= -244242007;
assign addr[47451]= -91761426;
assign addr[47452]= 61184634;
assign addr[47453]= 213820322;
assign addr[47454]= 365371365;
assign addr[47455]= 515068990;
assign addr[47456]= 662153826;
assign addr[47457]= 805879757;
assign addr[47458]= 945517704;
assign addr[47459]= 1080359326;
assign addr[47460]= 1209720613;
assign addr[47461]= 1332945355;
assign addr[47462]= 1449408469;
assign addr[47463]= 1558519173;
assign addr[47464]= 1659723983;
assign addr[47465]= 1752509516;
assign addr[47466]= 1836405100;
assign addr[47467]= 1910985158;
assign addr[47468]= 1975871368;
assign addr[47469]= 2030734582;
assign addr[47470]= 2075296495;
assign addr[47471]= 2109331059;
assign addr[47472]= 2132665626;
assign addr[47473]= 2145181827;
assign addr[47474]= 2146816171;
assign addr[47475]= 2137560369;
assign addr[47476]= 2117461370;
assign addr[47477]= 2086621133;
assign addr[47478]= 2045196100;
assign addr[47479]= 1993396407;
assign addr[47480]= 1931484818;
assign addr[47481]= 1859775393;
assign addr[47482]= 1778631892;
assign addr[47483]= 1688465931;
assign addr[47484]= 1589734894;
assign addr[47485]= 1482939614;
assign addr[47486]= 1368621831;
assign addr[47487]= 1247361445;
assign addr[47488]= 1119773573;
assign addr[47489]= 986505429;
assign addr[47490]= 848233042;
assign addr[47491]= 705657826;
assign addr[47492]= 559503022;
assign addr[47493]= 410510029;
assign addr[47494]= 259434643;
assign addr[47495]= 107043224;
assign addr[47496]= -45891193;
assign addr[47497]= -198592817;
assign addr[47498]= -350287041;
assign addr[47499]= -500204365;
assign addr[47500]= -647584304;
assign addr[47501]= -791679244;
assign addr[47502]= -931758235;
assign addr[47503]= -1067110699;
assign addr[47504]= -1197050035;
assign addr[47505]= -1320917099;
assign addr[47506]= -1438083551;
assign addr[47507]= -1547955041;
assign addr[47508]= -1649974225;
assign addr[47509]= -1743623590;
assign addr[47510]= -1828428082;
assign addr[47511]= -1903957513;
assign addr[47512]= -1969828744;
assign addr[47513]= -2025707632;
assign addr[47514]= -2071310720;
assign addr[47515]= -2106406677;
assign addr[47516]= -2130817471;
assign addr[47517]= -2144419275;
assign addr[47518]= -2147143090;
assign addr[47519]= -2138975100;
assign addr[47520]= -2119956737;
assign addr[47521]= -2090184478;
assign addr[47522]= -2049809346;
assign addr[47523]= -1999036154;
assign addr[47524]= -1938122457;
assign addr[47525]= -1867377253;
assign addr[47526]= -1787159411;
assign addr[47527]= -1697875851;
assign addr[47528]= -1599979481;
assign addr[47529]= -1493966902;
assign addr[47530]= -1380375881;
assign addr[47531]= -1259782632;
assign addr[47532]= -1132798888;
assign addr[47533]= -1000068799;
assign addr[47534]= -862265664;
assign addr[47535]= -720088517;
assign addr[47536]= -574258580;
assign addr[47537]= -425515602;
assign addr[47538]= -274614114;
assign addr[47539]= -122319591;
assign addr[47540]= 30595422;
assign addr[47541]= 183355234;
assign addr[47542]= 335184940;
assign addr[47543]= 485314355;
assign addr[47544]= 632981917;
assign addr[47545]= 777438554;
assign addr[47546]= 917951481;
assign addr[47547]= 1053807919;
assign addr[47548]= 1184318708;
assign addr[47549]= 1308821808;
assign addr[47550]= 1426685652;
assign addr[47551]= 1537312353;
assign addr[47552]= 1640140734;
assign addr[47553]= 1734649179;
assign addr[47554]= 1820358275;
assign addr[47555]= 1896833245;
assign addr[47556]= 1963686155;
assign addr[47557]= 2020577882;
assign addr[47558]= 2067219829;
assign addr[47559]= 2103375398;
assign addr[47560]= 2128861181;
assign addr[47561]= 2143547897;
assign addr[47562]= 2147361045;
assign addr[47563]= 2140281282;
assign addr[47564]= 2122344521;
assign addr[47565]= 2093641749;
assign addr[47566]= 2054318569;
assign addr[47567]= 2004574453;
assign addr[47568]= 1944661739;
assign addr[47569]= 1874884346;
assign addr[47570]= 1795596234;
assign addr[47571]= 1707199606;
assign addr[47572]= 1610142873;
assign addr[47573]= 1504918373;
assign addr[47574]= 1392059879;
assign addr[47575]= 1272139887;
assign addr[47576]= 1145766716;
assign addr[47577]= 1013581418;
assign addr[47578]= 876254528;
assign addr[47579]= 734482665;
assign addr[47580]= 588984994;
assign addr[47581]= 440499581;
assign addr[47582]= 289779648;
assign addr[47583]= 137589750;
assign addr[47584]= -15298099;
assign addr[47585]= -168108346;
assign addr[47586]= -320065829;
assign addr[47587]= -470399716;
assign addr[47588]= -618347408;
assign addr[47589]= -763158411;
assign addr[47590]= -904098143;
assign addr[47591]= -1040451659;
assign addr[47592]= -1171527280;
assign addr[47593]= -1296660098;
assign addr[47594]= -1415215352;
assign addr[47595]= -1526591649;
assign addr[47596]= -1630224009;
assign addr[47597]= -1725586737;
assign addr[47598]= -1812196087;
assign addr[47599]= -1889612716;
assign addr[47600]= -1957443913;
assign addr[47601]= -2015345591;
assign addr[47602]= -2063024031;
assign addr[47603]= -2100237377;
assign addr[47604]= -2126796855;
assign addr[47605]= -2142567738;
assign addr[47606]= -2147470025;
assign addr[47607]= -2141478848;
assign addr[47608]= -2124624598;
assign addr[47609]= -2096992772;
assign addr[47610]= -2058723538;
assign addr[47611]= -2010011024;
assign addr[47612]= -1951102334;
assign addr[47613]= -1882296293;
assign addr[47614]= -1803941934;
assign addr[47615]= -1716436725;
assign addr[47616]= -1620224553;
assign addr[47617]= -1515793473;
assign addr[47618]= -1403673233;
assign addr[47619]= -1284432584;
assign addr[47620]= -1158676398;
assign addr[47621]= -1027042599;
assign addr[47622]= -890198924;
assign addr[47623]= -748839539;
assign addr[47624]= -603681519;
assign addr[47625]= -455461206;
assign addr[47626]= -304930476;
assign addr[47627]= -152852926;
assign addr[47628]= 0;
assign addr[47629]= 152852926;
assign addr[47630]= 304930476;
assign addr[47631]= 455461206;
assign addr[47632]= 603681519;
assign addr[47633]= 748839539;
assign addr[47634]= 890198924;
assign addr[47635]= 1027042599;
assign addr[47636]= 1158676398;
assign addr[47637]= 1284432584;
assign addr[47638]= 1403673233;
assign addr[47639]= 1515793473;
assign addr[47640]= 1620224553;
assign addr[47641]= 1716436725;
assign addr[47642]= 1803941934;
assign addr[47643]= 1882296293;
assign addr[47644]= 1951102334;
assign addr[47645]= 2010011024;
assign addr[47646]= 2058723538;
assign addr[47647]= 2096992772;
assign addr[47648]= 2124624598;
assign addr[47649]= 2141478848;
assign addr[47650]= 2147470025;
assign addr[47651]= 2142567738;
assign addr[47652]= 2126796855;
assign addr[47653]= 2100237377;
assign addr[47654]= 2063024031;
assign addr[47655]= 2015345591;
assign addr[47656]= 1957443913;
assign addr[47657]= 1889612716;
assign addr[47658]= 1812196087;
assign addr[47659]= 1725586737;
assign addr[47660]= 1630224009;
assign addr[47661]= 1526591649;
assign addr[47662]= 1415215352;
assign addr[47663]= 1296660098;
assign addr[47664]= 1171527280;
assign addr[47665]= 1040451659;
assign addr[47666]= 904098143;
assign addr[47667]= 763158411;
assign addr[47668]= 618347408;
assign addr[47669]= 470399716;
assign addr[47670]= 320065829;
assign addr[47671]= 168108346;
assign addr[47672]= 15298099;
assign addr[47673]= -137589750;
assign addr[47674]= -289779648;
assign addr[47675]= -440499581;
assign addr[47676]= -588984994;
assign addr[47677]= -734482665;
assign addr[47678]= -876254528;
assign addr[47679]= -1013581418;
assign addr[47680]= -1145766716;
assign addr[47681]= -1272139887;
assign addr[47682]= -1392059879;
assign addr[47683]= -1504918373;
assign addr[47684]= -1610142873;
assign addr[47685]= -1707199606;
assign addr[47686]= -1795596234;
assign addr[47687]= -1874884346;
assign addr[47688]= -1944661739;
assign addr[47689]= -2004574453;
assign addr[47690]= -2054318569;
assign addr[47691]= -2093641749;
assign addr[47692]= -2122344521;
assign addr[47693]= -2140281282;
assign addr[47694]= -2147361045;
assign addr[47695]= -2143547897;
assign addr[47696]= -2128861181;
assign addr[47697]= -2103375398;
assign addr[47698]= -2067219829;
assign addr[47699]= -2020577882;
assign addr[47700]= -1963686155;
assign addr[47701]= -1896833245;
assign addr[47702]= -1820358275;
assign addr[47703]= -1734649179;
assign addr[47704]= -1640140734;
assign addr[47705]= -1537312353;
assign addr[47706]= -1426685652;
assign addr[47707]= -1308821808;
assign addr[47708]= -1184318708;
assign addr[47709]= -1053807919;
assign addr[47710]= -917951481;
assign addr[47711]= -777438554;
assign addr[47712]= -632981917;
assign addr[47713]= -485314355;
assign addr[47714]= -335184940;
assign addr[47715]= -183355234;
assign addr[47716]= -30595422;
assign addr[47717]= 122319591;
assign addr[47718]= 274614114;
assign addr[47719]= 425515602;
assign addr[47720]= 574258580;
assign addr[47721]= 720088517;
assign addr[47722]= 862265664;
assign addr[47723]= 1000068799;
assign addr[47724]= 1132798888;
assign addr[47725]= 1259782632;
assign addr[47726]= 1380375881;
assign addr[47727]= 1493966902;
assign addr[47728]= 1599979481;
assign addr[47729]= 1697875851;
assign addr[47730]= 1787159411;
assign addr[47731]= 1867377253;
assign addr[47732]= 1938122457;
assign addr[47733]= 1999036154;
assign addr[47734]= 2049809346;
assign addr[47735]= 2090184478;
assign addr[47736]= 2119956737;
assign addr[47737]= 2138975100;
assign addr[47738]= 2147143090;
assign addr[47739]= 2144419275;
assign addr[47740]= 2130817471;
assign addr[47741]= 2106406677;
assign addr[47742]= 2071310720;
assign addr[47743]= 2025707632;
assign addr[47744]= 1969828744;
assign addr[47745]= 1903957513;
assign addr[47746]= 1828428082;
assign addr[47747]= 1743623590;
assign addr[47748]= 1649974225;
assign addr[47749]= 1547955041;
assign addr[47750]= 1438083551;
assign addr[47751]= 1320917099;
assign addr[47752]= 1197050035;
assign addr[47753]= 1067110699;
assign addr[47754]= 931758235;
assign addr[47755]= 791679244;
assign addr[47756]= 647584304;
assign addr[47757]= 500204365;
assign addr[47758]= 350287041;
assign addr[47759]= 198592817;
assign addr[47760]= 45891193;
assign addr[47761]= -107043224;
assign addr[47762]= -259434643;
assign addr[47763]= -410510029;
assign addr[47764]= -559503022;
assign addr[47765]= -705657826;
assign addr[47766]= -848233042;
assign addr[47767]= -986505429;
assign addr[47768]= -1119773573;
assign addr[47769]= -1247361445;
assign addr[47770]= -1368621831;
assign addr[47771]= -1482939614;
assign addr[47772]= -1589734894;
assign addr[47773]= -1688465931;
assign addr[47774]= -1778631892;
assign addr[47775]= -1859775393;
assign addr[47776]= -1931484818;
assign addr[47777]= -1993396407;
assign addr[47778]= -2045196100;
assign addr[47779]= -2086621133;
assign addr[47780]= -2117461370;
assign addr[47781]= -2137560369;
assign addr[47782]= -2146816171;
assign addr[47783]= -2145181827;
assign addr[47784]= -2132665626;
assign addr[47785]= -2109331059;
assign addr[47786]= -2075296495;
assign addr[47787]= -2030734582;
assign addr[47788]= -1975871368;
assign addr[47789]= -1910985158;
assign addr[47790]= -1836405100;
assign addr[47791]= -1752509516;
assign addr[47792]= -1659723983;
assign addr[47793]= -1558519173;
assign addr[47794]= -1449408469;
assign addr[47795]= -1332945355;
assign addr[47796]= -1209720613;
assign addr[47797]= -1080359326;
assign addr[47798]= -945517704;
assign addr[47799]= -805879757;
assign addr[47800]= -662153826;
assign addr[47801]= -515068990;
assign addr[47802]= -365371365;
assign addr[47803]= -213820322;
assign addr[47804]= -61184634;
assign addr[47805]= 91761426;
assign addr[47806]= 244242007;
assign addr[47807]= 395483624;
assign addr[47808]= 544719071;
assign addr[47809]= 691191324;
assign addr[47810]= 834157373;
assign addr[47811]= 972891995;
assign addr[47812]= 1106691431;
assign addr[47813]= 1234876957;
assign addr[47814]= 1356798326;
assign addr[47815]= 1471837070;
assign addr[47816]= 1579409630;
assign addr[47817]= 1678970324;
assign addr[47818]= 1770014111;
assign addr[47819]= 1852079154;
assign addr[47820]= 1924749160;
assign addr[47821]= 1987655498;
assign addr[47822]= 2040479063;
assign addr[47823]= 2082951896;
assign addr[47824]= 2114858546;
assign addr[47825]= 2136037160;
assign addr[47826]= 2146380306;
assign addr[47827]= 2145835515;
assign addr[47828]= 2134405552;
assign addr[47829]= 2112148396;
assign addr[47830]= 2079176953;
assign addr[47831]= 2035658475;
assign addr[47832]= 1981813720;
assign addr[47833]= 1917915825;
assign addr[47834]= 1844288924;
assign addr[47835]= 1761306505;
assign addr[47836]= 1669389513;
assign addr[47837]= 1569004214;
assign addr[47838]= 1460659832;
assign addr[47839]= 1344905966;
assign addr[47840]= 1222329801;
assign addr[47841]= 1093553126;
assign addr[47842]= 959229189;
assign addr[47843]= 820039373;
assign addr[47844]= 676689746;
assign addr[47845]= 529907477;
assign addr[47846]= 380437148;
assign addr[47847]= 229036977;
assign addr[47848]= 76474970;
assign addr[47849]= -76474970;
assign addr[47850]= -229036977;
assign addr[47851]= -380437148;
assign addr[47852]= -529907477;
assign addr[47853]= -676689746;
assign addr[47854]= -820039373;
assign addr[47855]= -959229189;
assign addr[47856]= -1093553126;
assign addr[47857]= -1222329801;
assign addr[47858]= -1344905966;
assign addr[47859]= -1460659832;
assign addr[47860]= -1569004214;
assign addr[47861]= -1669389513;
assign addr[47862]= -1761306505;
assign addr[47863]= -1844288924;
assign addr[47864]= -1917915825;
assign addr[47865]= -1981813720;
assign addr[47866]= -2035658475;
assign addr[47867]= -2079176953;
assign addr[47868]= -2112148396;
assign addr[47869]= -2134405552;
assign addr[47870]= -2145835515;
assign addr[47871]= -2146380306;
assign addr[47872]= -2136037160;
assign addr[47873]= -2114858546;
assign addr[47874]= -2082951896;
assign addr[47875]= -2040479063;
assign addr[47876]= -1987655498;
assign addr[47877]= -1924749160;
assign addr[47878]= -1852079154;
assign addr[47879]= -1770014111;
assign addr[47880]= -1678970324;
assign addr[47881]= -1579409630;
assign addr[47882]= -1471837070;
assign addr[47883]= -1356798326;
assign addr[47884]= -1234876957;
assign addr[47885]= -1106691431;
assign addr[47886]= -972891995;
assign addr[47887]= -834157373;
assign addr[47888]= -691191324;
assign addr[47889]= -544719071;
assign addr[47890]= -395483624;
assign addr[47891]= -244242007;
assign addr[47892]= -91761426;
assign addr[47893]= 61184634;
assign addr[47894]= 213820322;
assign addr[47895]= 365371365;
assign addr[47896]= 515068990;
assign addr[47897]= 662153826;
assign addr[47898]= 805879757;
assign addr[47899]= 945517704;
assign addr[47900]= 1080359326;
assign addr[47901]= 1209720613;
assign addr[47902]= 1332945355;
assign addr[47903]= 1449408469;
assign addr[47904]= 1558519173;
assign addr[47905]= 1659723983;
assign addr[47906]= 1752509516;
assign addr[47907]= 1836405100;
assign addr[47908]= 1910985158;
assign addr[47909]= 1975871368;
assign addr[47910]= 2030734582;
assign addr[47911]= 2075296495;
assign addr[47912]= 2109331059;
assign addr[47913]= 2132665626;
assign addr[47914]= 2145181827;
assign addr[47915]= 2146816171;
assign addr[47916]= 2137560369;
assign addr[47917]= 2117461370;
assign addr[47918]= 2086621133;
assign addr[47919]= 2045196100;
assign addr[47920]= 1993396407;
assign addr[47921]= 1931484818;
assign addr[47922]= 1859775393;
assign addr[47923]= 1778631892;
assign addr[47924]= 1688465931;
assign addr[47925]= 1589734894;
assign addr[47926]= 1482939614;
assign addr[47927]= 1368621831;
assign addr[47928]= 1247361445;
assign addr[47929]= 1119773573;
assign addr[47930]= 986505429;
assign addr[47931]= 848233042;
assign addr[47932]= 705657826;
assign addr[47933]= 559503022;
assign addr[47934]= 410510029;
assign addr[47935]= 259434643;
assign addr[47936]= 107043224;
assign addr[47937]= -45891193;
assign addr[47938]= -198592817;
assign addr[47939]= -350287041;
assign addr[47940]= -500204365;
assign addr[47941]= -647584304;
assign addr[47942]= -791679244;
assign addr[47943]= -931758235;
assign addr[47944]= -1067110699;
assign addr[47945]= -1197050035;
assign addr[47946]= -1320917099;
assign addr[47947]= -1438083551;
assign addr[47948]= -1547955041;
assign addr[47949]= -1649974225;
assign addr[47950]= -1743623590;
assign addr[47951]= -1828428082;
assign addr[47952]= -1903957513;
assign addr[47953]= -1969828744;
assign addr[47954]= -2025707632;
assign addr[47955]= -2071310720;
assign addr[47956]= -2106406677;
assign addr[47957]= -2130817471;
assign addr[47958]= -2144419275;
assign addr[47959]= -2147143090;
assign addr[47960]= -2138975100;
assign addr[47961]= -2119956737;
assign addr[47962]= -2090184478;
assign addr[47963]= -2049809346;
assign addr[47964]= -1999036154;
assign addr[47965]= -1938122457;
assign addr[47966]= -1867377253;
assign addr[47967]= -1787159411;
assign addr[47968]= -1697875851;
assign addr[47969]= -1599979481;
assign addr[47970]= -1493966902;
assign addr[47971]= -1380375881;
assign addr[47972]= -1259782632;
assign addr[47973]= -1132798888;
assign addr[47974]= -1000068799;
assign addr[47975]= -862265664;
assign addr[47976]= -720088517;
assign addr[47977]= -574258580;
assign addr[47978]= -425515602;
assign addr[47979]= -274614114;
assign addr[47980]= -122319591;
assign addr[47981]= 30595422;
assign addr[47982]= 183355234;
assign addr[47983]= 335184940;
assign addr[47984]= 485314355;
assign addr[47985]= 632981917;
assign addr[47986]= 777438554;
assign addr[47987]= 917951481;
assign addr[47988]= 1053807919;
assign addr[47989]= 1184318708;
assign addr[47990]= 1308821808;
assign addr[47991]= 1426685652;
assign addr[47992]= 1537312353;
assign addr[47993]= 1640140734;
assign addr[47994]= 1734649179;
assign addr[47995]= 1820358275;
assign addr[47996]= 1896833245;
assign addr[47997]= 1963686155;
assign addr[47998]= 2020577882;
assign addr[47999]= 2067219829;
assign addr[48000]= 2103375398;
assign addr[48001]= 2128861181;
assign addr[48002]= 2143547897;
assign addr[48003]= 2147361045;
assign addr[48004]= 2140281282;
assign addr[48005]= 2122344521;
assign addr[48006]= 2093641749;
assign addr[48007]= 2054318569;
assign addr[48008]= 2004574453;
assign addr[48009]= 1944661739;
assign addr[48010]= 1874884346;
assign addr[48011]= 1795596234;
assign addr[48012]= 1707199606;
assign addr[48013]= 1610142873;
assign addr[48014]= 1504918373;
assign addr[48015]= 1392059879;
assign addr[48016]= 1272139887;
assign addr[48017]= 1145766716;
assign addr[48018]= 1013581418;
assign addr[48019]= 876254528;
assign addr[48020]= 734482665;
assign addr[48021]= 588984994;
assign addr[48022]= 440499581;
assign addr[48023]= 289779648;
assign addr[48024]= 137589750;
assign addr[48025]= -15298099;
assign addr[48026]= -168108346;
assign addr[48027]= -320065829;
assign addr[48028]= -470399716;
assign addr[48029]= -618347408;
assign addr[48030]= -763158411;
assign addr[48031]= -904098143;
assign addr[48032]= -1040451659;
assign addr[48033]= -1171527280;
assign addr[48034]= -1296660098;
assign addr[48035]= -1415215352;
assign addr[48036]= -1526591649;
assign addr[48037]= -1630224009;
assign addr[48038]= -1725586737;
assign addr[48039]= -1812196087;
assign addr[48040]= -1889612716;
assign addr[48041]= -1957443913;
assign addr[48042]= -2015345591;
assign addr[48043]= -2063024031;
assign addr[48044]= -2100237377;
assign addr[48045]= -2126796855;
assign addr[48046]= -2142567738;
assign addr[48047]= -2147470025;
assign addr[48048]= -2141478848;
assign addr[48049]= -2124624598;
assign addr[48050]= -2096992772;
assign addr[48051]= -2058723538;
assign addr[48052]= -2010011024;
assign addr[48053]= -1951102334;
assign addr[48054]= -1882296293;
assign addr[48055]= -1803941934;
assign addr[48056]= -1716436725;
assign addr[48057]= -1620224553;
assign addr[48058]= -1515793473;
assign addr[48059]= -1403673233;
assign addr[48060]= -1284432584;
assign addr[48061]= -1158676398;
assign addr[48062]= -1027042599;
assign addr[48063]= -890198924;
assign addr[48064]= -748839539;
assign addr[48065]= -603681519;
assign addr[48066]= -455461206;
assign addr[48067]= -304930476;
assign addr[48068]= -152852926;
assign addr[48069]= 0;
assign addr[48070]= 152852926;
assign addr[48071]= 304930476;
assign addr[48072]= 455461206;
assign addr[48073]= 603681519;
assign addr[48074]= 748839539;
assign addr[48075]= 890198924;
assign addr[48076]= 1027042599;
assign addr[48077]= 1158676398;
assign addr[48078]= 1284432584;
assign addr[48079]= 1403673233;
assign addr[48080]= 1515793473;
assign addr[48081]= 1620224553;
assign addr[48082]= 1716436725;
assign addr[48083]= 1803941934;
assign addr[48084]= 1882296293;
assign addr[48085]= 1951102334;
assign addr[48086]= 2010011024;
assign addr[48087]= 2058723538;
assign addr[48088]= 2096992772;
assign addr[48089]= 2124624598;
assign addr[48090]= 2141478848;
assign addr[48091]= 2147470025;
assign addr[48092]= 2142567738;
assign addr[48093]= 2126796855;
assign addr[48094]= 2100237377;
assign addr[48095]= 2063024031;
assign addr[48096]= 2015345591;
assign addr[48097]= 1957443913;
assign addr[48098]= 1889612716;
assign addr[48099]= 1812196087;
assign addr[48100]= 1725586737;
assign addr[48101]= 1630224009;
assign addr[48102]= 1526591649;
assign addr[48103]= 1415215352;
assign addr[48104]= 1296660098;
assign addr[48105]= 1171527280;
assign addr[48106]= 1040451659;
assign addr[48107]= 904098143;
assign addr[48108]= 763158411;
assign addr[48109]= 618347408;
assign addr[48110]= 470399716;
assign addr[48111]= 320065829;
assign addr[48112]= 168108346;
assign addr[48113]= 15298099;
assign addr[48114]= -137589750;
assign addr[48115]= -289779648;
assign addr[48116]= -440499581;
assign addr[48117]= -588984994;
assign addr[48118]= -734482665;
assign addr[48119]= -876254528;
assign addr[48120]= -1013581418;
assign addr[48121]= -1145766716;
assign addr[48122]= -1272139887;
assign addr[48123]= -1392059879;
assign addr[48124]= -1504918373;
assign addr[48125]= -1610142873;
assign addr[48126]= -1707199606;
assign addr[48127]= -1795596234;
assign addr[48128]= -1874884346;
assign addr[48129]= -1944661739;
assign addr[48130]= -2004574453;
assign addr[48131]= -2054318569;
assign addr[48132]= -2093641749;
assign addr[48133]= -2122344521;
assign addr[48134]= -2140281282;
assign addr[48135]= -2147361045;
assign addr[48136]= -2143547897;
assign addr[48137]= -2128861181;
assign addr[48138]= -2103375398;
assign addr[48139]= -2067219829;
assign addr[48140]= -2020577882;
assign addr[48141]= -1963686155;
assign addr[48142]= -1896833245;
assign addr[48143]= -1820358275;
assign addr[48144]= -1734649179;
assign addr[48145]= -1640140734;
assign addr[48146]= -1537312353;
assign addr[48147]= -1426685652;
assign addr[48148]= -1308821808;
assign addr[48149]= -1184318708;
assign addr[48150]= -1053807919;
assign addr[48151]= -917951481;
assign addr[48152]= -777438554;
assign addr[48153]= -632981917;
assign addr[48154]= -485314355;
assign addr[48155]= -335184940;
assign addr[48156]= -183355234;
assign addr[48157]= -30595422;
assign addr[48158]= 122319591;
assign addr[48159]= 274614114;
assign addr[48160]= 425515602;
assign addr[48161]= 574258580;
assign addr[48162]= 720088517;
assign addr[48163]= 862265664;
assign addr[48164]= 1000068799;
assign addr[48165]= 1132798888;
assign addr[48166]= 1259782632;
assign addr[48167]= 1380375881;
assign addr[48168]= 1493966902;
assign addr[48169]= 1599979481;
assign addr[48170]= 1697875851;
assign addr[48171]= 1787159411;
assign addr[48172]= 1867377253;
assign addr[48173]= 1938122457;
assign addr[48174]= 1999036154;
assign addr[48175]= 2049809346;
assign addr[48176]= 2090184478;
assign addr[48177]= 2119956737;
assign addr[48178]= 2138975100;
assign addr[48179]= 2147143090;
assign addr[48180]= 2144419275;
assign addr[48181]= 2130817471;
assign addr[48182]= 2106406677;
assign addr[48183]= 2071310720;
assign addr[48184]= 2025707632;
assign addr[48185]= 1969828744;
assign addr[48186]= 1903957513;
assign addr[48187]= 1828428082;
assign addr[48188]= 1743623590;
assign addr[48189]= 1649974225;
assign addr[48190]= 1547955041;
assign addr[48191]= 1438083551;
assign addr[48192]= 1320917099;
assign addr[48193]= 1197050035;
assign addr[48194]= 1067110699;
assign addr[48195]= 931758235;
assign addr[48196]= 791679244;
assign addr[48197]= 647584304;
assign addr[48198]= 500204365;
assign addr[48199]= 350287041;
assign addr[48200]= 198592817;
assign addr[48201]= 45891193;
assign addr[48202]= -107043224;
assign addr[48203]= -259434643;
assign addr[48204]= -410510029;
assign addr[48205]= -559503022;
assign addr[48206]= -705657826;
assign addr[48207]= -848233042;
assign addr[48208]= -986505429;
assign addr[48209]= -1119773573;
assign addr[48210]= -1247361445;
assign addr[48211]= -1368621831;
assign addr[48212]= -1482939614;
assign addr[48213]= -1589734894;
assign addr[48214]= -1688465931;
assign addr[48215]= -1778631892;
assign addr[48216]= -1859775393;
assign addr[48217]= -1931484818;
assign addr[48218]= -1993396407;
assign addr[48219]= -2045196100;
assign addr[48220]= -2086621133;
assign addr[48221]= -2117461370;
assign addr[48222]= -2137560369;
assign addr[48223]= -2146816171;
assign addr[48224]= -2145181827;
assign addr[48225]= -2132665626;
assign addr[48226]= -2109331059;
assign addr[48227]= -2075296495;
assign addr[48228]= -2030734582;
assign addr[48229]= -1975871368;
assign addr[48230]= -1910985158;
assign addr[48231]= -1836405100;
assign addr[48232]= -1752509516;
assign addr[48233]= -1659723983;
assign addr[48234]= -1558519173;
assign addr[48235]= -1449408469;
assign addr[48236]= -1332945355;
assign addr[48237]= -1209720613;
assign addr[48238]= -1080359326;
assign addr[48239]= -945517704;
assign addr[48240]= -805879757;
assign addr[48241]= -662153826;
assign addr[48242]= -515068990;
assign addr[48243]= -365371365;
assign addr[48244]= -213820322;
assign addr[48245]= -61184634;
assign addr[48246]= 91761426;
assign addr[48247]= 244242007;
assign addr[48248]= 395483624;
assign addr[48249]= 544719071;
assign addr[48250]= 691191324;
assign addr[48251]= 834157373;
assign addr[48252]= 972891995;
assign addr[48253]= 1106691431;
assign addr[48254]= 1234876957;
assign addr[48255]= 1356798326;
assign addr[48256]= 1471837070;
assign addr[48257]= 1579409630;
assign addr[48258]= 1678970324;
assign addr[48259]= 1770014111;
assign addr[48260]= 1852079154;
assign addr[48261]= 1924749160;
assign addr[48262]= 1987655498;
assign addr[48263]= 2040479063;
assign addr[48264]= 2082951896;
assign addr[48265]= 2114858546;
assign addr[48266]= 2136037160;
assign addr[48267]= 2146380306;
assign addr[48268]= 2145835515;
assign addr[48269]= 2134405552;
assign addr[48270]= 2112148396;
assign addr[48271]= 2079176953;
assign addr[48272]= 2035658475;
assign addr[48273]= 1981813720;
assign addr[48274]= 1917915825;
assign addr[48275]= 1844288924;
assign addr[48276]= 1761306505;
assign addr[48277]= 1669389513;
assign addr[48278]= 1569004214;
assign addr[48279]= 1460659832;
assign addr[48280]= 1344905966;
assign addr[48281]= 1222329801;
assign addr[48282]= 1093553126;
assign addr[48283]= 959229189;
assign addr[48284]= 820039373;
assign addr[48285]= 676689746;
assign addr[48286]= 529907477;
assign addr[48287]= 380437148;
assign addr[48288]= 229036977;
assign addr[48289]= 76474970;
assign addr[48290]= -76474970;
assign addr[48291]= -229036977;
assign addr[48292]= -380437148;
assign addr[48293]= -529907477;
assign addr[48294]= -676689746;
assign addr[48295]= -820039373;
assign addr[48296]= -959229189;
assign addr[48297]= -1093553126;
assign addr[48298]= -1222329801;
assign addr[48299]= -1344905966;
assign addr[48300]= -1460659832;
assign addr[48301]= -1569004214;
assign addr[48302]= -1669389513;
assign addr[48303]= -1761306505;
assign addr[48304]= -1844288924;
assign addr[48305]= -1917915825;
assign addr[48306]= -1981813720;
assign addr[48307]= -2035658475;
assign addr[48308]= -2079176953;
assign addr[48309]= -2112148396;
assign addr[48310]= -2134405552;
assign addr[48311]= -2145835515;
assign addr[48312]= -2146380306;
assign addr[48313]= -2136037160;
assign addr[48314]= -2114858546;
assign addr[48315]= -2082951896;
assign addr[48316]= -2040479063;
assign addr[48317]= -1987655498;
assign addr[48318]= -1924749160;
assign addr[48319]= -1852079154;
assign addr[48320]= -1770014111;
assign addr[48321]= -1678970324;
assign addr[48322]= -1579409630;
assign addr[48323]= -1471837070;
assign addr[48324]= -1356798326;
assign addr[48325]= -1234876957;
assign addr[48326]= -1106691431;
assign addr[48327]= -972891995;
assign addr[48328]= -834157373;
assign addr[48329]= -691191324;
assign addr[48330]= -544719071;
assign addr[48331]= -395483624;
assign addr[48332]= -244242007;
assign addr[48333]= -91761426;
assign addr[48334]= 61184634;
assign addr[48335]= 213820322;
assign addr[48336]= 365371365;
assign addr[48337]= 515068990;
assign addr[48338]= 662153826;
assign addr[48339]= 805879757;
assign addr[48340]= 945517704;
assign addr[48341]= 1080359326;
assign addr[48342]= 1209720613;
assign addr[48343]= 1332945355;
assign addr[48344]= 1449408469;
assign addr[48345]= 1558519173;
assign addr[48346]= 1659723983;
assign addr[48347]= 1752509516;
assign addr[48348]= 1836405100;
assign addr[48349]= 1910985158;
assign addr[48350]= 1975871368;
assign addr[48351]= 2030734582;
assign addr[48352]= 2075296495;
assign addr[48353]= 2109331059;
assign addr[48354]= 2132665626;
assign addr[48355]= 2145181827;
assign addr[48356]= 2146816171;
assign addr[48357]= 2137560369;
assign addr[48358]= 2117461370;
assign addr[48359]= 2086621133;
assign addr[48360]= 2045196100;
assign addr[48361]= 1993396407;
assign addr[48362]= 1931484818;
assign addr[48363]= 1859775393;
assign addr[48364]= 1778631892;
assign addr[48365]= 1688465931;
assign addr[48366]= 1589734894;
assign addr[48367]= 1482939614;
assign addr[48368]= 1368621831;
assign addr[48369]= 1247361445;
assign addr[48370]= 1119773573;
assign addr[48371]= 986505429;
assign addr[48372]= 848233042;
assign addr[48373]= 705657826;
assign addr[48374]= 559503022;
assign addr[48375]= 410510029;
assign addr[48376]= 259434643;
assign addr[48377]= 107043224;
assign addr[48378]= -45891193;
assign addr[48379]= -198592817;
assign addr[48380]= -350287041;
assign addr[48381]= -500204365;
assign addr[48382]= -647584304;
assign addr[48383]= -791679244;
assign addr[48384]= -931758235;
assign addr[48385]= -1067110699;
assign addr[48386]= -1197050035;
assign addr[48387]= -1320917099;
assign addr[48388]= -1438083551;
assign addr[48389]= -1547955041;
assign addr[48390]= -1649974225;
assign addr[48391]= -1743623590;
assign addr[48392]= -1828428082;
assign addr[48393]= -1903957513;
assign addr[48394]= -1969828744;
assign addr[48395]= -2025707632;
assign addr[48396]= -2071310720;
assign addr[48397]= -2106406677;
assign addr[48398]= -2130817471;
assign addr[48399]= -2144419275;
assign addr[48400]= -2147143090;
assign addr[48401]= -2138975100;
assign addr[48402]= -2119956737;
assign addr[48403]= -2090184478;
assign addr[48404]= -2049809346;
assign addr[48405]= -1999036154;
assign addr[48406]= -1938122457;
assign addr[48407]= -1867377253;
assign addr[48408]= -1787159411;
assign addr[48409]= -1697875851;
assign addr[48410]= -1599979481;
assign addr[48411]= -1493966902;
assign addr[48412]= -1380375881;
assign addr[48413]= -1259782632;
assign addr[48414]= -1132798888;
assign addr[48415]= -1000068799;
assign addr[48416]= -862265664;
assign addr[48417]= -720088517;
assign addr[48418]= -574258580;
assign addr[48419]= -425515602;
assign addr[48420]= -274614114;
assign addr[48421]= -122319591;
assign addr[48422]= 30595422;
assign addr[48423]= 183355234;
assign addr[48424]= 335184940;
assign addr[48425]= 485314355;
assign addr[48426]= 632981917;
assign addr[48427]= 777438554;
assign addr[48428]= 917951481;
assign addr[48429]= 1053807919;
assign addr[48430]= 1184318708;
assign addr[48431]= 1308821808;
assign addr[48432]= 1426685652;
assign addr[48433]= 1537312353;
assign addr[48434]= 1640140734;
assign addr[48435]= 1734649179;
assign addr[48436]= 1820358275;
assign addr[48437]= 1896833245;
assign addr[48438]= 1963686155;
assign addr[48439]= 2020577882;
assign addr[48440]= 2067219829;
assign addr[48441]= 2103375398;
assign addr[48442]= 2128861181;
assign addr[48443]= 2143547897;
assign addr[48444]= 2147361045;
assign addr[48445]= 2140281282;
assign addr[48446]= 2122344521;
assign addr[48447]= 2093641749;
assign addr[48448]= 2054318569;
assign addr[48449]= 2004574453;
assign addr[48450]= 1944661739;
assign addr[48451]= 1874884346;
assign addr[48452]= 1795596234;
assign addr[48453]= 1707199606;
assign addr[48454]= 1610142873;
assign addr[48455]= 1504918373;
assign addr[48456]= 1392059879;
assign addr[48457]= 1272139887;
assign addr[48458]= 1145766716;
assign addr[48459]= 1013581418;
assign addr[48460]= 876254528;
assign addr[48461]= 734482665;
assign addr[48462]= 588984994;
assign addr[48463]= 440499581;
assign addr[48464]= 289779648;
assign addr[48465]= 137589750;
assign addr[48466]= -15298099;
assign addr[48467]= -168108346;
assign addr[48468]= -320065829;
assign addr[48469]= -470399716;
assign addr[48470]= -618347408;
assign addr[48471]= -763158411;
assign addr[48472]= -904098143;
assign addr[48473]= -1040451659;
assign addr[48474]= -1171527280;
assign addr[48475]= -1296660098;
assign addr[48476]= -1415215352;
assign addr[48477]= -1526591649;
assign addr[48478]= -1630224009;
assign addr[48479]= -1725586737;
assign addr[48480]= -1812196087;
assign addr[48481]= -1889612716;
assign addr[48482]= -1957443913;
assign addr[48483]= -2015345591;
assign addr[48484]= -2063024031;
assign addr[48485]= -2100237377;
assign addr[48486]= -2126796855;
assign addr[48487]= -2142567738;
assign addr[48488]= -2147470025;
assign addr[48489]= -2141478848;
assign addr[48490]= -2124624598;
assign addr[48491]= -2096992772;
assign addr[48492]= -2058723538;
assign addr[48493]= -2010011024;
assign addr[48494]= -1951102334;
assign addr[48495]= -1882296293;
assign addr[48496]= -1803941934;
assign addr[48497]= -1716436725;
assign addr[48498]= -1620224553;
assign addr[48499]= -1515793473;
assign addr[48500]= -1403673233;
assign addr[48501]= -1284432584;
assign addr[48502]= -1158676398;
assign addr[48503]= -1027042599;
assign addr[48504]= -890198924;
assign addr[48505]= -748839539;
assign addr[48506]= -603681519;
assign addr[48507]= -455461206;
assign addr[48508]= -304930476;
assign addr[48509]= -152852926;
assign addr[48510]= 0;
assign addr[48511]= 152852926;
assign addr[48512]= 304930476;
assign addr[48513]= 455461206;
assign addr[48514]= 603681519;
assign addr[48515]= 748839539;
assign addr[48516]= 890198924;
assign addr[48517]= 1027042599;
assign addr[48518]= 1158676398;
assign addr[48519]= 1284432584;
assign addr[48520]= 1403673233;
assign addr[48521]= 1515793473;
assign addr[48522]= 1620224553;
assign addr[48523]= 1716436725;
assign addr[48524]= 1803941934;
assign addr[48525]= 1882296293;
assign addr[48526]= 1951102334;
assign addr[48527]= 2010011024;
assign addr[48528]= 2058723538;
assign addr[48529]= 2096992772;
assign addr[48530]= 2124624598;
assign addr[48531]= 2141478848;
assign addr[48532]= 2147470025;
assign addr[48533]= 2142567738;
assign addr[48534]= 2126796855;
assign addr[48535]= 2100237377;
assign addr[48536]= 2063024031;
assign addr[48537]= 2015345591;
assign addr[48538]= 1957443913;
assign addr[48539]= 1889612716;
assign addr[48540]= 1812196087;
assign addr[48541]= 1725586737;
assign addr[48542]= 1630224009;
assign addr[48543]= 1526591649;
assign addr[48544]= 1415215352;
assign addr[48545]= 1296660098;
assign addr[48546]= 1171527280;
assign addr[48547]= 1040451659;
assign addr[48548]= 904098143;
assign addr[48549]= 763158411;
assign addr[48550]= 618347408;
assign addr[48551]= 470399716;
assign addr[48552]= 320065829;
assign addr[48553]= 168108346;
assign addr[48554]= 15298099;
assign addr[48555]= -137589750;
assign addr[48556]= -289779648;
assign addr[48557]= -440499581;
assign addr[48558]= -588984994;
assign addr[48559]= -734482665;
assign addr[48560]= -876254528;
assign addr[48561]= -1013581418;
assign addr[48562]= -1145766716;
assign addr[48563]= -1272139887;
assign addr[48564]= -1392059879;
assign addr[48565]= -1504918373;
assign addr[48566]= -1610142873;
assign addr[48567]= -1707199606;
assign addr[48568]= -1795596234;
assign addr[48569]= -1874884346;
assign addr[48570]= -1944661739;
assign addr[48571]= -2004574453;
assign addr[48572]= -2054318569;
assign addr[48573]= -2093641749;
assign addr[48574]= -2122344521;
assign addr[48575]= -2140281282;
assign addr[48576]= -2147361045;
assign addr[48577]= -2143547897;
assign addr[48578]= -2128861181;
assign addr[48579]= -2103375398;
assign addr[48580]= -2067219829;
assign addr[48581]= -2020577882;
assign addr[48582]= -1963686155;
assign addr[48583]= -1896833245;
assign addr[48584]= -1820358275;
assign addr[48585]= -1734649179;
assign addr[48586]= -1640140734;
assign addr[48587]= -1537312353;
assign addr[48588]= -1426685652;
assign addr[48589]= -1308821808;
assign addr[48590]= -1184318708;
assign addr[48591]= -1053807919;
assign addr[48592]= -917951481;
assign addr[48593]= -777438554;
assign addr[48594]= -632981917;
assign addr[48595]= -485314355;
assign addr[48596]= -335184940;
assign addr[48597]= -183355234;
assign addr[48598]= -30595422;
assign addr[48599]= 122319591;
assign addr[48600]= 274614114;
assign addr[48601]= 425515602;
assign addr[48602]= 574258580;
assign addr[48603]= 720088517;
assign addr[48604]= 862265664;
assign addr[48605]= 1000068799;
assign addr[48606]= 1132798888;
assign addr[48607]= 1259782632;
assign addr[48608]= 1380375881;
assign addr[48609]= 1493966902;
assign addr[48610]= 1599979481;
assign addr[48611]= 1697875851;
assign addr[48612]= 1787159411;
assign addr[48613]= 1867377253;
assign addr[48614]= 1938122457;
assign addr[48615]= 1999036154;
assign addr[48616]= 2049809346;
assign addr[48617]= 2090184478;
assign addr[48618]= 2119956737;
assign addr[48619]= 2138975100;
assign addr[48620]= 2147143090;
assign addr[48621]= 2144419275;
assign addr[48622]= 2130817471;
assign addr[48623]= 2106406677;
assign addr[48624]= 2071310720;
assign addr[48625]= 2025707632;
assign addr[48626]= 1969828744;
assign addr[48627]= 1903957513;
assign addr[48628]= 1828428082;
assign addr[48629]= 1743623590;
assign addr[48630]= 1649974225;
assign addr[48631]= 1547955041;
assign addr[48632]= 1438083551;
assign addr[48633]= 1320917099;
assign addr[48634]= 1197050035;
assign addr[48635]= 1067110699;
assign addr[48636]= 931758235;
assign addr[48637]= 791679244;
assign addr[48638]= 647584304;
assign addr[48639]= 500204365;
assign addr[48640]= 350287041;
assign addr[48641]= 198592817;
assign addr[48642]= 45891193;
assign addr[48643]= -107043224;
assign addr[48644]= -259434643;
assign addr[48645]= -410510029;
assign addr[48646]= -559503022;
assign addr[48647]= -705657826;
assign addr[48648]= -848233042;
assign addr[48649]= -986505429;
assign addr[48650]= -1119773573;
assign addr[48651]= -1247361445;
assign addr[48652]= -1368621831;
assign addr[48653]= -1482939614;
assign addr[48654]= -1589734894;
assign addr[48655]= -1688465931;
assign addr[48656]= -1778631892;
assign addr[48657]= -1859775393;
assign addr[48658]= -1931484818;
assign addr[48659]= -1993396407;
assign addr[48660]= -2045196100;
assign addr[48661]= -2086621133;
assign addr[48662]= -2117461370;
assign addr[48663]= -2137560369;
assign addr[48664]= -2146816171;
assign addr[48665]= -2145181827;
assign addr[48666]= -2132665626;
assign addr[48667]= -2109331059;
assign addr[48668]= -2075296495;
assign addr[48669]= -2030734582;
assign addr[48670]= -1975871368;
assign addr[48671]= -1910985158;
assign addr[48672]= -1836405100;
assign addr[48673]= -1752509516;
assign addr[48674]= -1659723983;
assign addr[48675]= -1558519173;
assign addr[48676]= -1449408469;
assign addr[48677]= -1332945355;
assign addr[48678]= -1209720613;
assign addr[48679]= -1080359326;
assign addr[48680]= -945517704;
assign addr[48681]= -805879757;
assign addr[48682]= -662153826;
assign addr[48683]= -515068990;
assign addr[48684]= -365371365;
assign addr[48685]= -213820322;
assign addr[48686]= -61184634;
assign addr[48687]= 91761426;
assign addr[48688]= 244242007;
assign addr[48689]= 395483624;
assign addr[48690]= 544719071;
assign addr[48691]= 691191324;
assign addr[48692]= 834157373;
assign addr[48693]= 972891995;
assign addr[48694]= 1106691431;
assign addr[48695]= 1234876957;
assign addr[48696]= 1356798326;
assign addr[48697]= 1471837070;
assign addr[48698]= 1579409630;
assign addr[48699]= 1678970324;
assign addr[48700]= 1770014111;
assign addr[48701]= 1852079154;
assign addr[48702]= 1924749160;
assign addr[48703]= 1987655498;
assign addr[48704]= 2040479063;
assign addr[48705]= 2082951896;
assign addr[48706]= 2114858546;
assign addr[48707]= 2136037160;
assign addr[48708]= 2146380306;
assign addr[48709]= 2145835515;
assign addr[48710]= 2134405552;
assign addr[48711]= 2112148396;
assign addr[48712]= 2079176953;
assign addr[48713]= 2035658475;
assign addr[48714]= 1981813720;
assign addr[48715]= 1917915825;
assign addr[48716]= 1844288924;
assign addr[48717]= 1761306505;
assign addr[48718]= 1669389513;
assign addr[48719]= 1569004214;
assign addr[48720]= 1460659832;
assign addr[48721]= 1344905966;
assign addr[48722]= 1222329801;
assign addr[48723]= 1093553126;
assign addr[48724]= 959229189;
assign addr[48725]= 820039373;
assign addr[48726]= 676689746;
assign addr[48727]= 529907477;
assign addr[48728]= 380437148;
assign addr[48729]= 229036977;
assign addr[48730]= 76474970;
assign addr[48731]= -76474970;
assign addr[48732]= -229036977;
assign addr[48733]= -380437148;
assign addr[48734]= -529907477;
assign addr[48735]= -676689746;
assign addr[48736]= -820039373;
assign addr[48737]= -959229189;
assign addr[48738]= -1093553126;
assign addr[48739]= -1222329801;
assign addr[48740]= -1344905966;
assign addr[48741]= -1460659832;
assign addr[48742]= -1569004214;
assign addr[48743]= -1669389513;
assign addr[48744]= -1761306505;
assign addr[48745]= -1844288924;
assign addr[48746]= -1917915825;
assign addr[48747]= -1981813720;
assign addr[48748]= -2035658475;
assign addr[48749]= -2079176953;
assign addr[48750]= -2112148396;
assign addr[48751]= -2134405552;
assign addr[48752]= -2145835515;
assign addr[48753]= -2146380306;
assign addr[48754]= -2136037160;
assign addr[48755]= -2114858546;
assign addr[48756]= -2082951896;
assign addr[48757]= -2040479063;
assign addr[48758]= -1987655498;
assign addr[48759]= -1924749160;
assign addr[48760]= -1852079154;
assign addr[48761]= -1770014111;
assign addr[48762]= -1678970324;
assign addr[48763]= -1579409630;
assign addr[48764]= -1471837070;
assign addr[48765]= -1356798326;
assign addr[48766]= -1234876957;
assign addr[48767]= -1106691431;
assign addr[48768]= -972891995;
assign addr[48769]= -834157373;
assign addr[48770]= -691191324;
assign addr[48771]= -544719071;
assign addr[48772]= -395483624;
assign addr[48773]= -244242007;
assign addr[48774]= -91761426;
assign addr[48775]= 61184634;
assign addr[48776]= 213820322;
assign addr[48777]= 365371365;
assign addr[48778]= 515068990;
assign addr[48779]= 662153826;
assign addr[48780]= 805879757;
assign addr[48781]= 945517704;
assign addr[48782]= 1080359326;
assign addr[48783]= 1209720613;
assign addr[48784]= 1332945355;
assign addr[48785]= 1449408469;
assign addr[48786]= 1558519173;
assign addr[48787]= 1659723983;
assign addr[48788]= 1752509516;
assign addr[48789]= 1836405100;
assign addr[48790]= 1910985158;
assign addr[48791]= 1975871368;
assign addr[48792]= 2030734582;
assign addr[48793]= 2075296495;
assign addr[48794]= 2109331059;
assign addr[48795]= 2132665626;
assign addr[48796]= 2145181827;
assign addr[48797]= 2146816171;
assign addr[48798]= 2137560369;
assign addr[48799]= 2117461370;
assign addr[48800]= 2086621133;
assign addr[48801]= 2045196100;
assign addr[48802]= 1993396407;
assign addr[48803]= 1931484818;
assign addr[48804]= 1859775393;
assign addr[48805]= 1778631892;
assign addr[48806]= 1688465931;
assign addr[48807]= 1589734894;
assign addr[48808]= 1482939614;
assign addr[48809]= 1368621831;
assign addr[48810]= 1247361445;
assign addr[48811]= 1119773573;
assign addr[48812]= 986505429;
assign addr[48813]= 848233042;
assign addr[48814]= 705657826;
assign addr[48815]= 559503022;
assign addr[48816]= 410510029;
assign addr[48817]= 259434643;
assign addr[48818]= 107043224;
assign addr[48819]= -45891193;
assign addr[48820]= -198592817;
assign addr[48821]= -350287041;
assign addr[48822]= -500204365;
assign addr[48823]= -647584304;
assign addr[48824]= -791679244;
assign addr[48825]= -931758235;
assign addr[48826]= -1067110699;
assign addr[48827]= -1197050035;
assign addr[48828]= -1320917099;
assign addr[48829]= -1438083551;
assign addr[48830]= -1547955041;
assign addr[48831]= -1649974225;
assign addr[48832]= -1743623590;
assign addr[48833]= -1828428082;
assign addr[48834]= -1903957513;
assign addr[48835]= -1969828744;
assign addr[48836]= -2025707632;
assign addr[48837]= -2071310720;
assign addr[48838]= -2106406677;
assign addr[48839]= -2130817471;
assign addr[48840]= -2144419275;
assign addr[48841]= -2147143090;
assign addr[48842]= -2138975100;
assign addr[48843]= -2119956737;
assign addr[48844]= -2090184478;
assign addr[48845]= -2049809346;
assign addr[48846]= -1999036154;
assign addr[48847]= -1938122457;
assign addr[48848]= -1867377253;
assign addr[48849]= -1787159411;
assign addr[48850]= -1697875851;
assign addr[48851]= -1599979481;
assign addr[48852]= -1493966902;
assign addr[48853]= -1380375881;
assign addr[48854]= -1259782632;
assign addr[48855]= -1132798888;
assign addr[48856]= -1000068799;
assign addr[48857]= -862265664;
assign addr[48858]= -720088517;
assign addr[48859]= -574258580;
assign addr[48860]= -425515602;
assign addr[48861]= -274614114;
assign addr[48862]= -122319591;
assign addr[48863]= 30595422;
assign addr[48864]= 183355234;
assign addr[48865]= 335184940;
assign addr[48866]= 485314355;
assign addr[48867]= 632981917;
assign addr[48868]= 777438554;
assign addr[48869]= 917951481;
assign addr[48870]= 1053807919;
assign addr[48871]= 1184318708;
assign addr[48872]= 1308821808;
assign addr[48873]= 1426685652;
assign addr[48874]= 1537312353;
assign addr[48875]= 1640140734;
assign addr[48876]= 1734649179;
assign addr[48877]= 1820358275;
assign addr[48878]= 1896833245;
assign addr[48879]= 1963686155;
assign addr[48880]= 2020577882;
assign addr[48881]= 2067219829;
assign addr[48882]= 2103375398;
assign addr[48883]= 2128861181;
assign addr[48884]= 2143547897;
assign addr[48885]= 2147361045;
assign addr[48886]= 2140281282;
assign addr[48887]= 2122344521;
assign addr[48888]= 2093641749;
assign addr[48889]= 2054318569;
assign addr[48890]= 2004574453;
assign addr[48891]= 1944661739;
assign addr[48892]= 1874884346;
assign addr[48893]= 1795596234;
assign addr[48894]= 1707199606;
assign addr[48895]= 1610142873;
assign addr[48896]= 1504918373;
assign addr[48897]= 1392059879;
assign addr[48898]= 1272139887;
assign addr[48899]= 1145766716;
assign addr[48900]= 1013581418;
assign addr[48901]= 876254528;
assign addr[48902]= 734482665;
assign addr[48903]= 588984994;
assign addr[48904]= 440499581;
assign addr[48905]= 289779648;
assign addr[48906]= 137589750;
assign addr[48907]= -15298099;
assign addr[48908]= -168108346;
assign addr[48909]= -320065829;
assign addr[48910]= -470399716;
assign addr[48911]= -618347408;
assign addr[48912]= -763158411;
assign addr[48913]= -904098143;
assign addr[48914]= -1040451659;
assign addr[48915]= -1171527280;
assign addr[48916]= -1296660098;
assign addr[48917]= -1415215352;
assign addr[48918]= -1526591649;
assign addr[48919]= -1630224009;
assign addr[48920]= -1725586737;
assign addr[48921]= -1812196087;
assign addr[48922]= -1889612716;
assign addr[48923]= -1957443913;
assign addr[48924]= -2015345591;
assign addr[48925]= -2063024031;
assign addr[48926]= -2100237377;
assign addr[48927]= -2126796855;
assign addr[48928]= -2142567738;
assign addr[48929]= -2147470025;
assign addr[48930]= -2141478848;
assign addr[48931]= -2124624598;
assign addr[48932]= -2096992772;
assign addr[48933]= -2058723538;
assign addr[48934]= -2010011024;
assign addr[48935]= -1951102334;
assign addr[48936]= -1882296293;
assign addr[48937]= -1803941934;
assign addr[48938]= -1716436725;
assign addr[48939]= -1620224553;
assign addr[48940]= -1515793473;
assign addr[48941]= -1403673233;
assign addr[48942]= -1284432584;
assign addr[48943]= -1158676398;
assign addr[48944]= -1027042599;
assign addr[48945]= -890198924;
assign addr[48946]= -748839539;
assign addr[48947]= -603681519;
assign addr[48948]= -455461206;
assign addr[48949]= -304930476;
assign addr[48950]= -152852926;
assign addr[48951]= 0;
assign addr[48952]= 152852926;
assign addr[48953]= 304930476;
assign addr[48954]= 455461206;
assign addr[48955]= 603681519;
assign addr[48956]= 748839539;
assign addr[48957]= 890198924;
assign addr[48958]= 1027042599;
assign addr[48959]= 1158676398;
assign addr[48960]= 1284432584;
assign addr[48961]= 1403673233;
assign addr[48962]= 1515793473;
assign addr[48963]= 1620224553;
assign addr[48964]= 1716436725;
assign addr[48965]= 1803941934;
assign addr[48966]= 1882296293;
assign addr[48967]= 1951102334;
assign addr[48968]= 2010011024;
assign addr[48969]= 2058723538;
assign addr[48970]= 2096992772;
assign addr[48971]= 2124624598;
assign addr[48972]= 2141478848;
assign addr[48973]= 2147470025;
assign addr[48974]= 2142567738;
assign addr[48975]= 2126796855;
assign addr[48976]= 2100237377;
assign addr[48977]= 2063024031;
assign addr[48978]= 2015345591;
assign addr[48979]= 1957443913;
assign addr[48980]= 1889612716;
assign addr[48981]= 1812196087;
assign addr[48982]= 1725586737;
assign addr[48983]= 1630224009;
assign addr[48984]= 1526591649;
assign addr[48985]= 1415215352;
assign addr[48986]= 1296660098;
assign addr[48987]= 1171527280;
assign addr[48988]= 1040451659;
assign addr[48989]= 904098143;
assign addr[48990]= 763158411;
assign addr[48991]= 618347408;
assign addr[48992]= 470399716;
assign addr[48993]= 320065829;
assign addr[48994]= 168108346;
assign addr[48995]= 15298099;
assign addr[48996]= -137589750;
assign addr[48997]= -289779648;
assign addr[48998]= -440499581;
assign addr[48999]= -588984994;
assign addr[49000]= -734482665;
assign addr[49001]= -876254528;
assign addr[49002]= -1013581418;
assign addr[49003]= -1145766716;
assign addr[49004]= -1272139887;
assign addr[49005]= -1392059879;
assign addr[49006]= -1504918373;
assign addr[49007]= -1610142873;
assign addr[49008]= -1707199606;
assign addr[49009]= -1795596234;
assign addr[49010]= -1874884346;
assign addr[49011]= -1944661739;
assign addr[49012]= -2004574453;
assign addr[49013]= -2054318569;
assign addr[49014]= -2093641749;
assign addr[49015]= -2122344521;
assign addr[49016]= -2140281282;
assign addr[49017]= -2147361045;
assign addr[49018]= -2143547897;
assign addr[49019]= -2128861181;
assign addr[49020]= -2103375398;
assign addr[49021]= -2067219829;
assign addr[49022]= -2020577882;
assign addr[49023]= -1963686155;
assign addr[49024]= -1896833245;
assign addr[49025]= -1820358275;
assign addr[49026]= -1734649179;
assign addr[49027]= -1640140734;
assign addr[49028]= -1537312353;
assign addr[49029]= -1426685652;
assign addr[49030]= -1308821808;
assign addr[49031]= -1184318708;
assign addr[49032]= -1053807919;
assign addr[49033]= -917951481;
assign addr[49034]= -777438554;
assign addr[49035]= -632981917;
assign addr[49036]= -485314355;
assign addr[49037]= -335184940;
assign addr[49038]= -183355234;
assign addr[49039]= -30595422;
assign addr[49040]= 122319591;
assign addr[49041]= 274614114;
assign addr[49042]= 425515602;
assign addr[49043]= 574258580;
assign addr[49044]= 720088517;
assign addr[49045]= 862265664;
assign addr[49046]= 1000068799;
assign addr[49047]= 1132798888;
assign addr[49048]= 1259782632;
assign addr[49049]= 1380375881;
assign addr[49050]= 1493966902;
assign addr[49051]= 1599979481;
assign addr[49052]= 1697875851;
assign addr[49053]= 1787159411;
assign addr[49054]= 1867377253;
assign addr[49055]= 1938122457;
assign addr[49056]= 1999036154;
assign addr[49057]= 2049809346;
assign addr[49058]= 2090184478;
assign addr[49059]= 2119956737;
assign addr[49060]= 2138975100;
assign addr[49061]= 2147143090;
assign addr[49062]= 2144419275;
assign addr[49063]= 2130817471;
assign addr[49064]= 2106406677;
assign addr[49065]= 2071310720;
assign addr[49066]= 2025707632;
assign addr[49067]= 1969828744;
assign addr[49068]= 1903957513;
assign addr[49069]= 1828428082;
assign addr[49070]= 1743623590;
assign addr[49071]= 1649974225;
assign addr[49072]= 1547955041;
assign addr[49073]= 1438083551;
assign addr[49074]= 1320917099;
assign addr[49075]= 1197050035;
assign addr[49076]= 1067110699;
assign addr[49077]= 931758235;
assign addr[49078]= 791679244;
assign addr[49079]= 647584304;
assign addr[49080]= 500204365;
assign addr[49081]= 350287041;
assign addr[49082]= 198592817;
assign addr[49083]= 45891193;
assign addr[49084]= -107043224;
assign addr[49085]= -259434643;
assign addr[49086]= -410510029;
assign addr[49087]= -559503022;
assign addr[49088]= -705657826;
assign addr[49089]= -848233042;
assign addr[49090]= -986505429;
assign addr[49091]= -1119773573;
assign addr[49092]= -1247361445;
assign addr[49093]= -1368621831;
assign addr[49094]= -1482939614;
assign addr[49095]= -1589734894;
assign addr[49096]= -1688465931;
assign addr[49097]= -1778631892;
assign addr[49098]= -1859775393;
assign addr[49099]= -1931484818;
assign addr[49100]= -1993396407;
assign addr[49101]= -2045196100;
assign addr[49102]= -2086621133;
assign addr[49103]= -2117461370;
assign addr[49104]= -2137560369;
assign addr[49105]= -2146816171;
assign addr[49106]= -2145181827;
assign addr[49107]= -2132665626;
assign addr[49108]= -2109331059;
assign addr[49109]= -2075296495;
assign addr[49110]= -2030734582;
assign addr[49111]= -1975871368;
assign addr[49112]= -1910985158;
assign addr[49113]= -1836405100;
assign addr[49114]= -1752509516;
assign addr[49115]= -1659723983;
assign addr[49116]= -1558519173;
assign addr[49117]= -1449408469;
assign addr[49118]= -1332945355;
assign addr[49119]= -1209720613;
assign addr[49120]= -1080359326;
assign addr[49121]= -945517704;
assign addr[49122]= -805879757;
assign addr[49123]= -662153826;
assign addr[49124]= -515068990;
assign addr[49125]= -365371365;
assign addr[49126]= -213820322;
assign addr[49127]= -61184634;
assign addr[49128]= 91761426;
assign addr[49129]= 244242007;
assign addr[49130]= 395483624;
assign addr[49131]= 544719071;
assign addr[49132]= 691191324;
assign addr[49133]= 834157373;
assign addr[49134]= 972891995;
assign addr[49135]= 1106691431;
assign addr[49136]= 1234876957;
assign addr[49137]= 1356798326;
assign addr[49138]= 1471837070;
assign addr[49139]= 1579409630;
assign addr[49140]= 1678970324;
assign addr[49141]= 1770014111;
assign addr[49142]= 1852079154;
assign addr[49143]= 1924749160;
assign addr[49144]= 1987655498;
assign addr[49145]= 2040479063;
assign addr[49146]= 2082951896;
assign addr[49147]= 2114858546;
assign addr[49148]= 2136037160;
assign addr[49149]= 2146380306;
assign addr[49150]= 2145835515;
assign addr[49151]= 2134405552;
assign addr[49152]= 2112148396;
assign addr[49153]= 2079176953;
assign addr[49154]= 2035658475;
assign addr[49155]= 1981813720;
assign addr[49156]= 1917915825;
assign addr[49157]= 1844288924;
assign addr[49158]= 1761306505;
assign addr[49159]= 1669389513;
assign addr[49160]= 1569004214;
assign addr[49161]= 1460659832;
assign addr[49162]= 1344905966;
assign addr[49163]= 1222329801;
assign addr[49164]= 1093553126;
assign addr[49165]= 959229189;
assign addr[49166]= 820039373;
assign addr[49167]= 676689746;
assign addr[49168]= 529907477;
assign addr[49169]= 380437148;
assign addr[49170]= 229036977;
assign addr[49171]= 76474970;
assign addr[49172]= -76474970;
assign addr[49173]= -229036977;
assign addr[49174]= -380437148;
assign addr[49175]= -529907477;
assign addr[49176]= -676689746;
assign addr[49177]= -820039373;
assign addr[49178]= -959229189;
assign addr[49179]= -1093553126;
assign addr[49180]= -1222329801;
assign addr[49181]= -1344905966;
assign addr[49182]= -1460659832;
assign addr[49183]= -1569004214;
assign addr[49184]= -1669389513;
assign addr[49185]= -1761306505;
assign addr[49186]= -1844288924;
assign addr[49187]= -1917915825;
assign addr[49188]= -1981813720;
assign addr[49189]= -2035658475;
assign addr[49190]= -2079176953;
assign addr[49191]= -2112148396;
assign addr[49192]= -2134405552;
assign addr[49193]= -2145835515;
assign addr[49194]= -2146380306;
assign addr[49195]= -2136037160;
assign addr[49196]= -2114858546;
assign addr[49197]= -2082951896;
assign addr[49198]= -2040479063;
assign addr[49199]= -1987655498;
assign addr[49200]= -1924749160;
assign addr[49201]= -1852079154;
assign addr[49202]= -1770014111;
assign addr[49203]= -1678970324;
assign addr[49204]= -1579409630;
assign addr[49205]= -1471837070;
assign addr[49206]= -1356798326;
assign addr[49207]= -1234876957;
assign addr[49208]= -1106691431;
assign addr[49209]= -972891995;
assign addr[49210]= -834157373;
assign addr[49211]= -691191324;
assign addr[49212]= -544719071;
assign addr[49213]= -395483624;
assign addr[49214]= -244242007;
assign addr[49215]= -91761426;
assign addr[49216]= 61184634;
assign addr[49217]= 213820322;
assign addr[49218]= 365371365;
assign addr[49219]= 515068990;
assign addr[49220]= 662153826;
assign addr[49221]= 805879757;
assign addr[49222]= 945517704;
assign addr[49223]= 1080359326;
assign addr[49224]= 1209720613;
assign addr[49225]= 1332945355;
assign addr[49226]= 1449408469;
assign addr[49227]= 1558519173;
assign addr[49228]= 1659723983;
assign addr[49229]= 1752509516;
assign addr[49230]= 1836405100;
assign addr[49231]= 1910985158;
assign addr[49232]= 1975871368;
assign addr[49233]= 2030734582;
assign addr[49234]= 2075296495;
assign addr[49235]= 2109331059;
assign addr[49236]= 2132665626;
assign addr[49237]= 2145181827;
assign addr[49238]= 2146816171;
assign addr[49239]= 2137560369;
assign addr[49240]= 2117461370;
assign addr[49241]= 2086621133;
assign addr[49242]= 2045196100;
assign addr[49243]= 1993396407;
assign addr[49244]= 1931484818;
assign addr[49245]= 1859775393;
assign addr[49246]= 1778631892;
assign addr[49247]= 1688465931;
assign addr[49248]= 1589734894;
assign addr[49249]= 1482939614;
assign addr[49250]= 1368621831;
assign addr[49251]= 1247361445;
assign addr[49252]= 1119773573;
assign addr[49253]= 986505429;
assign addr[49254]= 848233042;
assign addr[49255]= 705657826;
assign addr[49256]= 559503022;
assign addr[49257]= 410510029;
assign addr[49258]= 259434643;
assign addr[49259]= 107043224;
assign addr[49260]= -45891193;
assign addr[49261]= -198592817;
assign addr[49262]= -350287041;
assign addr[49263]= -500204365;
assign addr[49264]= -647584304;
assign addr[49265]= -791679244;
assign addr[49266]= -931758235;
assign addr[49267]= -1067110699;
assign addr[49268]= -1197050035;
assign addr[49269]= -1320917099;
assign addr[49270]= -1438083551;
assign addr[49271]= -1547955041;
assign addr[49272]= -1649974225;
assign addr[49273]= -1743623590;
assign addr[49274]= -1828428082;
assign addr[49275]= -1903957513;
assign addr[49276]= -1969828744;
assign addr[49277]= -2025707632;
assign addr[49278]= -2071310720;
assign addr[49279]= -2106406677;
assign addr[49280]= -2130817471;
assign addr[49281]= -2144419275;
assign addr[49282]= -2147143090;
assign addr[49283]= -2138975100;
assign addr[49284]= -2119956737;
assign addr[49285]= -2090184478;
assign addr[49286]= -2049809346;
assign addr[49287]= -1999036154;
assign addr[49288]= -1938122457;
assign addr[49289]= -1867377253;
assign addr[49290]= -1787159411;
assign addr[49291]= -1697875851;
assign addr[49292]= -1599979481;
assign addr[49293]= -1493966902;
assign addr[49294]= -1380375881;
assign addr[49295]= -1259782632;
assign addr[49296]= -1132798888;
assign addr[49297]= -1000068799;
assign addr[49298]= -862265664;
assign addr[49299]= -720088517;
assign addr[49300]= -574258580;
assign addr[49301]= -425515602;
assign addr[49302]= -274614114;
assign addr[49303]= -122319591;
assign addr[49304]= 30595422;
assign addr[49305]= 183355234;
assign addr[49306]= 335184940;
assign addr[49307]= 485314355;
assign addr[49308]= 632981917;
assign addr[49309]= 777438554;
assign addr[49310]= 917951481;
assign addr[49311]= 1053807919;
assign addr[49312]= 1184318708;
assign addr[49313]= 1308821808;
assign addr[49314]= 1426685652;
assign addr[49315]= 1537312353;
assign addr[49316]= 1640140734;
assign addr[49317]= 1734649179;
assign addr[49318]= 1820358275;
assign addr[49319]= 1896833245;
assign addr[49320]= 1963686155;
assign addr[49321]= 2020577882;
assign addr[49322]= 2067219829;
assign addr[49323]= 2103375398;
assign addr[49324]= 2128861181;
assign addr[49325]= 2143547897;
assign addr[49326]= 2147361045;
assign addr[49327]= 2140281282;
assign addr[49328]= 2122344521;
assign addr[49329]= 2093641749;
assign addr[49330]= 2054318569;
assign addr[49331]= 2004574453;
assign addr[49332]= 1944661739;
assign addr[49333]= 1874884346;
assign addr[49334]= 1795596234;
assign addr[49335]= 1707199606;
assign addr[49336]= 1610142873;
assign addr[49337]= 1504918373;
assign addr[49338]= 1392059879;
assign addr[49339]= 1272139887;
assign addr[49340]= 1145766716;
assign addr[49341]= 1013581418;
assign addr[49342]= 876254528;
assign addr[49343]= 734482665;
assign addr[49344]= 588984994;
assign addr[49345]= 440499581;
assign addr[49346]= 289779648;
assign addr[49347]= 137589750;
assign addr[49348]= -15298099;
assign addr[49349]= -168108346;
assign addr[49350]= -320065829;
assign addr[49351]= -470399716;
assign addr[49352]= -618347408;
assign addr[49353]= -763158411;
assign addr[49354]= -904098143;
assign addr[49355]= -1040451659;
assign addr[49356]= -1171527280;
assign addr[49357]= -1296660098;
assign addr[49358]= -1415215352;
assign addr[49359]= -1526591649;
assign addr[49360]= -1630224009;
assign addr[49361]= -1725586737;
assign addr[49362]= -1812196087;
assign addr[49363]= -1889612716;
assign addr[49364]= -1957443913;
assign addr[49365]= -2015345591;
assign addr[49366]= -2063024031;
assign addr[49367]= -2100237377;
assign addr[49368]= -2126796855;
assign addr[49369]= -2142567738;
assign addr[49370]= -2147470025;
assign addr[49371]= -2141478848;
assign addr[49372]= -2124624598;
assign addr[49373]= -2096992772;
assign addr[49374]= -2058723538;
assign addr[49375]= -2010011024;
assign addr[49376]= -1951102334;
assign addr[49377]= -1882296293;
assign addr[49378]= -1803941934;
assign addr[49379]= -1716436725;
assign addr[49380]= -1620224553;
assign addr[49381]= -1515793473;
assign addr[49382]= -1403673233;
assign addr[49383]= -1284432584;
assign addr[49384]= -1158676398;
assign addr[49385]= -1027042599;
assign addr[49386]= -890198924;
assign addr[49387]= -748839539;
assign addr[49388]= -603681519;
assign addr[49389]= -455461206;
assign addr[49390]= -304930476;
assign addr[49391]= -152852926;
assign addr[49392]= 0;
assign addr[49393]= 152852926;
assign addr[49394]= 304930476;
assign addr[49395]= 455461206;
assign addr[49396]= 603681519;
assign addr[49397]= 748839539;
assign addr[49398]= 890198924;
assign addr[49399]= 1027042599;
assign addr[49400]= 1158676398;
assign addr[49401]= 1284432584;
assign addr[49402]= 1403673233;
assign addr[49403]= 1515793473;
assign addr[49404]= 1620224553;
assign addr[49405]= 1716436725;
assign addr[49406]= 1803941934;
assign addr[49407]= 1882296293;
assign addr[49408]= 1951102334;
assign addr[49409]= 2010011024;
assign addr[49410]= 2058723538;
assign addr[49411]= 2096992772;
assign addr[49412]= 2124624598;
assign addr[49413]= 2141478848;
assign addr[49414]= 2147470025;
assign addr[49415]= 2142567738;
assign addr[49416]= 2126796855;
assign addr[49417]= 2100237377;
assign addr[49418]= 2063024031;
assign addr[49419]= 2015345591;
assign addr[49420]= 1957443913;
assign addr[49421]= 1889612716;
assign addr[49422]= 1812196087;
assign addr[49423]= 1725586737;
assign addr[49424]= 1630224009;
assign addr[49425]= 1526591649;
assign addr[49426]= 1415215352;
assign addr[49427]= 1296660098;
assign addr[49428]= 1171527280;
assign addr[49429]= 1040451659;
assign addr[49430]= 904098143;
assign addr[49431]= 763158411;
assign addr[49432]= 618347408;
assign addr[49433]= 470399716;
assign addr[49434]= 320065829;
assign addr[49435]= 168108346;
assign addr[49436]= 15298099;
assign addr[49437]= -137589750;
assign addr[49438]= -289779648;
assign addr[49439]= -440499581;
assign addr[49440]= -588984994;
assign addr[49441]= -734482665;
assign addr[49442]= -876254528;
assign addr[49443]= -1013581418;
assign addr[49444]= -1145766716;
assign addr[49445]= -1272139887;
assign addr[49446]= -1392059879;
assign addr[49447]= -1504918373;
assign addr[49448]= -1610142873;
assign addr[49449]= -1707199606;
assign addr[49450]= -1795596234;
assign addr[49451]= -1874884346;
assign addr[49452]= -1944661739;
assign addr[49453]= -2004574453;
assign addr[49454]= -2054318569;
assign addr[49455]= -2093641749;
assign addr[49456]= -2122344521;
assign addr[49457]= -2140281282;
assign addr[49458]= -2147361045;
assign addr[49459]= -2143547897;
assign addr[49460]= -2128861181;
assign addr[49461]= -2103375398;
assign addr[49462]= -2067219829;
assign addr[49463]= -2020577882;
assign addr[49464]= -1963686155;
assign addr[49465]= -1896833245;
assign addr[49466]= -1820358275;
assign addr[49467]= -1734649179;
assign addr[49468]= -1640140734;
assign addr[49469]= -1537312353;
assign addr[49470]= -1426685652;
assign addr[49471]= -1308821808;
assign addr[49472]= -1184318708;
assign addr[49473]= -1053807919;
assign addr[49474]= -917951481;
assign addr[49475]= -777438554;
assign addr[49476]= -632981917;
assign addr[49477]= -485314355;
assign addr[49478]= -335184940;
assign addr[49479]= -183355234;
assign addr[49480]= -30595422;
assign addr[49481]= 122319591;
assign addr[49482]= 274614114;
assign addr[49483]= 425515602;
assign addr[49484]= 574258580;
assign addr[49485]= 720088517;
assign addr[49486]= 862265664;
assign addr[49487]= 1000068799;
assign addr[49488]= 1132798888;
assign addr[49489]= 1259782632;
assign addr[49490]= 1380375881;
assign addr[49491]= 1493966902;
assign addr[49492]= 1599979481;
assign addr[49493]= 1697875851;
assign addr[49494]= 1787159411;
assign addr[49495]= 1867377253;
assign addr[49496]= 1938122457;
assign addr[49497]= 1999036154;
assign addr[49498]= 2049809346;
assign addr[49499]= 2090184478;
assign addr[49500]= 2119956737;
assign addr[49501]= 2138975100;
assign addr[49502]= 2147143090;
assign addr[49503]= 2144419275;
assign addr[49504]= 2130817471;
assign addr[49505]= 2106406677;
assign addr[49506]= 2071310720;
assign addr[49507]= 2025707632;
assign addr[49508]= 1969828744;
assign addr[49509]= 1903957513;
assign addr[49510]= 1828428082;
assign addr[49511]= 1743623590;
assign addr[49512]= 1649974225;
assign addr[49513]= 1547955041;
assign addr[49514]= 1438083551;
assign addr[49515]= 1320917099;
assign addr[49516]= 1197050035;
assign addr[49517]= 1067110699;
assign addr[49518]= 931758235;
assign addr[49519]= 791679244;
assign addr[49520]= 647584304;
assign addr[49521]= 500204365;
assign addr[49522]= 350287041;
assign addr[49523]= 198592817;
assign addr[49524]= 45891193;
assign addr[49525]= -107043224;
assign addr[49526]= -259434643;
assign addr[49527]= -410510029;
assign addr[49528]= -559503022;
assign addr[49529]= -705657826;
assign addr[49530]= -848233042;
assign addr[49531]= -986505429;
assign addr[49532]= -1119773573;
assign addr[49533]= -1247361445;
assign addr[49534]= -1368621831;
assign addr[49535]= -1482939614;
assign addr[49536]= -1589734894;
assign addr[49537]= -1688465931;
assign addr[49538]= -1778631892;
assign addr[49539]= -1859775393;
assign addr[49540]= -1931484818;
assign addr[49541]= -1993396407;
assign addr[49542]= -2045196100;
assign addr[49543]= -2086621133;
assign addr[49544]= -2117461370;
assign addr[49545]= -2137560369;
assign addr[49546]= -2146816171;
assign addr[49547]= -2145181827;
assign addr[49548]= -2132665626;
assign addr[49549]= -2109331059;
assign addr[49550]= -2075296495;
assign addr[49551]= -2030734582;
assign addr[49552]= -1975871368;
assign addr[49553]= -1910985158;
assign addr[49554]= -1836405100;
assign addr[49555]= -1752509516;
assign addr[49556]= -1659723983;
assign addr[49557]= -1558519173;
assign addr[49558]= -1449408469;
assign addr[49559]= -1332945355;
assign addr[49560]= -1209720613;
assign addr[49561]= -1080359326;
assign addr[49562]= -945517704;
assign addr[49563]= -805879757;
assign addr[49564]= -662153826;
assign addr[49565]= -515068990;
assign addr[49566]= -365371365;
assign addr[49567]= -213820322;
assign addr[49568]= -61184634;
assign addr[49569]= 91761426;
assign addr[49570]= 244242007;
assign addr[49571]= 395483624;
assign addr[49572]= 544719071;
assign addr[49573]= 691191324;
assign addr[49574]= 834157373;
assign addr[49575]= 972891995;
assign addr[49576]= 1106691431;
assign addr[49577]= 1234876957;
assign addr[49578]= 1356798326;
assign addr[49579]= 1471837070;
assign addr[49580]= 1579409630;
assign addr[49581]= 1678970324;
assign addr[49582]= 1770014111;
assign addr[49583]= 1852079154;
assign addr[49584]= 1924749160;
assign addr[49585]= 1987655498;
assign addr[49586]= 2040479063;
assign addr[49587]= 2082951896;
assign addr[49588]= 2114858546;
assign addr[49589]= 2136037160;
assign addr[49590]= 2146380306;
assign addr[49591]= 2145835515;
assign addr[49592]= 2134405552;
assign addr[49593]= 2112148396;
assign addr[49594]= 2079176953;
assign addr[49595]= 2035658475;
assign addr[49596]= 1981813720;
assign addr[49597]= 1917915825;
assign addr[49598]= 1844288924;
assign addr[49599]= 1761306505;
assign addr[49600]= 1669389513;
assign addr[49601]= 1569004214;
assign addr[49602]= 1460659832;
assign addr[49603]= 1344905966;
assign addr[49604]= 1222329801;
assign addr[49605]= 1093553126;
assign addr[49606]= 959229189;
assign addr[49607]= 820039373;
assign addr[49608]= 676689746;
assign addr[49609]= 529907477;
assign addr[49610]= 380437148;
assign addr[49611]= 229036977;
assign addr[49612]= 76474970;
assign addr[49613]= -76474970;
assign addr[49614]= -229036977;
assign addr[49615]= -380437148;
assign addr[49616]= -529907477;
assign addr[49617]= -676689746;
assign addr[49618]= -820039373;
assign addr[49619]= -959229189;
assign addr[49620]= -1093553126;
assign addr[49621]= -1222329801;
assign addr[49622]= -1344905966;
assign addr[49623]= -1460659832;
assign addr[49624]= -1569004214;
assign addr[49625]= -1669389513;
assign addr[49626]= -1761306505;
assign addr[49627]= -1844288924;
assign addr[49628]= -1917915825;
assign addr[49629]= -1981813720;
assign addr[49630]= -2035658475;
assign addr[49631]= -2079176953;
assign addr[49632]= -2112148396;
assign addr[49633]= -2134405552;
assign addr[49634]= -2145835515;
assign addr[49635]= -2146380306;
assign addr[49636]= -2136037160;
assign addr[49637]= -2114858546;
assign addr[49638]= -2082951896;
assign addr[49639]= -2040479063;
assign addr[49640]= -1987655498;
assign addr[49641]= -1924749160;
assign addr[49642]= -1852079154;
assign addr[49643]= -1770014111;
assign addr[49644]= -1678970324;
assign addr[49645]= -1579409630;
assign addr[49646]= -1471837070;
assign addr[49647]= -1356798326;
assign addr[49648]= -1234876957;
assign addr[49649]= -1106691431;
assign addr[49650]= -972891995;
assign addr[49651]= -834157373;
assign addr[49652]= -691191324;
assign addr[49653]= -544719071;
assign addr[49654]= -395483624;
assign addr[49655]= -244242007;
assign addr[49656]= -91761426;
assign addr[49657]= 61184634;
assign addr[49658]= 213820322;
assign addr[49659]= 365371365;
assign addr[49660]= 515068990;
assign addr[49661]= 662153826;
assign addr[49662]= 805879757;
assign addr[49663]= 945517704;
assign addr[49664]= 1080359326;
assign addr[49665]= 1209720613;
assign addr[49666]= 1332945355;
assign addr[49667]= 1449408469;
assign addr[49668]= 1558519173;
assign addr[49669]= 1659723983;
assign addr[49670]= 1752509516;
assign addr[49671]= 1836405100;
assign addr[49672]= 1910985158;
assign addr[49673]= 1975871368;
assign addr[49674]= 2030734582;
assign addr[49675]= 2075296495;
assign addr[49676]= 2109331059;
assign addr[49677]= 2132665626;
assign addr[49678]= 2145181827;
assign addr[49679]= 2146816171;
assign addr[49680]= 2137560369;
assign addr[49681]= 2117461370;
assign addr[49682]= 2086621133;
assign addr[49683]= 2045196100;
assign addr[49684]= 1993396407;
assign addr[49685]= 1931484818;
assign addr[49686]= 1859775393;
assign addr[49687]= 1778631892;
assign addr[49688]= 1688465931;
assign addr[49689]= 1589734894;
assign addr[49690]= 1482939614;
assign addr[49691]= 1368621831;
assign addr[49692]= 1247361445;
assign addr[49693]= 1119773573;
assign addr[49694]= 986505429;
assign addr[49695]= 848233042;
assign addr[49696]= 705657826;
assign addr[49697]= 559503022;
assign addr[49698]= 410510029;
assign addr[49699]= 259434643;
assign addr[49700]= 107043224;
assign addr[49701]= -45891193;
assign addr[49702]= -198592817;
assign addr[49703]= -350287041;
assign addr[49704]= -500204365;
assign addr[49705]= -647584304;
assign addr[49706]= -791679244;
assign addr[49707]= -931758235;
assign addr[49708]= -1067110699;
assign addr[49709]= -1197050035;
assign addr[49710]= -1320917099;
assign addr[49711]= -1438083551;
assign addr[49712]= -1547955041;
assign addr[49713]= -1649974225;
assign addr[49714]= -1743623590;
assign addr[49715]= -1828428082;
assign addr[49716]= -1903957513;
assign addr[49717]= -1969828744;
assign addr[49718]= -2025707632;
assign addr[49719]= -2071310720;
assign addr[49720]= -2106406677;
assign addr[49721]= -2130817471;
assign addr[49722]= -2144419275;
assign addr[49723]= -2147143090;
assign addr[49724]= -2138975100;
assign addr[49725]= -2119956737;
assign addr[49726]= -2090184478;
assign addr[49727]= -2049809346;
assign addr[49728]= -1999036154;
assign addr[49729]= -1938122457;
assign addr[49730]= -1867377253;
assign addr[49731]= -1787159411;
assign addr[49732]= -1697875851;
assign addr[49733]= -1599979481;
assign addr[49734]= -1493966902;
assign addr[49735]= -1380375881;
assign addr[49736]= -1259782632;
assign addr[49737]= -1132798888;
assign addr[49738]= -1000068799;
assign addr[49739]= -862265664;
assign addr[49740]= -720088517;
assign addr[49741]= -574258580;
assign addr[49742]= -425515602;
assign addr[49743]= -274614114;
assign addr[49744]= -122319591;
assign addr[49745]= 30595422;
assign addr[49746]= 183355234;
assign addr[49747]= 335184940;
assign addr[49748]= 485314355;
assign addr[49749]= 632981917;
assign addr[49750]= 777438554;
assign addr[49751]= 917951481;
assign addr[49752]= 1053807919;
assign addr[49753]= 1184318708;
assign addr[49754]= 1308821808;
assign addr[49755]= 1426685652;
assign addr[49756]= 1537312353;
assign addr[49757]= 1640140734;
assign addr[49758]= 1734649179;
assign addr[49759]= 1820358275;
assign addr[49760]= 1896833245;
assign addr[49761]= 1963686155;
assign addr[49762]= 2020577882;
assign addr[49763]= 2067219829;
assign addr[49764]= 2103375398;
assign addr[49765]= 2128861181;
assign addr[49766]= 2143547897;
assign addr[49767]= 2147361045;
assign addr[49768]= 2140281282;
assign addr[49769]= 2122344521;
assign addr[49770]= 2093641749;
assign addr[49771]= 2054318569;
assign addr[49772]= 2004574453;
assign addr[49773]= 1944661739;
assign addr[49774]= 1874884346;
assign addr[49775]= 1795596234;
assign addr[49776]= 1707199606;
assign addr[49777]= 1610142873;
assign addr[49778]= 1504918373;
assign addr[49779]= 1392059879;
assign addr[49780]= 1272139887;
assign addr[49781]= 1145766716;
assign addr[49782]= 1013581418;
assign addr[49783]= 876254528;
assign addr[49784]= 734482665;
assign addr[49785]= 588984994;
assign addr[49786]= 440499581;
assign addr[49787]= 289779648;
assign addr[49788]= 137589750;
assign addr[49789]= -15298099;
assign addr[49790]= -168108346;
assign addr[49791]= -320065829;
assign addr[49792]= -470399716;
assign addr[49793]= -618347408;
assign addr[49794]= -763158411;
assign addr[49795]= -904098143;
assign addr[49796]= -1040451659;
assign addr[49797]= -1171527280;
assign addr[49798]= -1296660098;
assign addr[49799]= -1415215352;
assign addr[49800]= -1526591649;
assign addr[49801]= -1630224009;
assign addr[49802]= -1725586737;
assign addr[49803]= -1812196087;
assign addr[49804]= -1889612716;
assign addr[49805]= -1957443913;
assign addr[49806]= -2015345591;
assign addr[49807]= -2063024031;
assign addr[49808]= -2100237377;
assign addr[49809]= -2126796855;
assign addr[49810]= -2142567738;
assign addr[49811]= -2147470025;
assign addr[49812]= -2141478848;
assign addr[49813]= -2124624598;
assign addr[49814]= -2096992772;
assign addr[49815]= -2058723538;
assign addr[49816]= -2010011024;
assign addr[49817]= -1951102334;
assign addr[49818]= -1882296293;
assign addr[49819]= -1803941934;
assign addr[49820]= -1716436725;
assign addr[49821]= -1620224553;
assign addr[49822]= -1515793473;
assign addr[49823]= -1403673233;
assign addr[49824]= -1284432584;
assign addr[49825]= -1158676398;
assign addr[49826]= -1027042599;
assign addr[49827]= -890198924;
assign addr[49828]= -748839539;
assign addr[49829]= -603681519;
assign addr[49830]= -455461206;
assign addr[49831]= -304930476;
assign addr[49832]= -152852926;
assign addr[49833]= 0;
assign addr[49834]= 152852926;
assign addr[49835]= 304930476;
assign addr[49836]= 455461206;
assign addr[49837]= 603681519;
assign addr[49838]= 748839539;
assign addr[49839]= 890198924;
assign addr[49840]= 1027042599;
assign addr[49841]= 1158676398;
assign addr[49842]= 1284432584;
assign addr[49843]= 1403673233;
assign addr[49844]= 1515793473;
assign addr[49845]= 1620224553;
assign addr[49846]= 1716436725;
assign addr[49847]= 1803941934;
assign addr[49848]= 1882296293;
assign addr[49849]= 1951102334;
assign addr[49850]= 2010011024;
assign addr[49851]= 2058723538;
assign addr[49852]= 2096992772;
assign addr[49853]= 2124624598;
assign addr[49854]= 2141478848;
assign addr[49855]= 2147470025;
assign addr[49856]= 2142567738;
assign addr[49857]= 2126796855;
assign addr[49858]= 2100237377;
assign addr[49859]= 2063024031;
assign addr[49860]= 2015345591;
assign addr[49861]= 1957443913;
assign addr[49862]= 1889612716;
assign addr[49863]= 1812196087;
assign addr[49864]= 1725586737;
assign addr[49865]= 1630224009;
assign addr[49866]= 1526591649;
assign addr[49867]= 1415215352;
assign addr[49868]= 1296660098;
assign addr[49869]= 1171527280;
assign addr[49870]= 1040451659;
assign addr[49871]= 904098143;
assign addr[49872]= 763158411;
assign addr[49873]= 618347408;
assign addr[49874]= 470399716;
assign addr[49875]= 320065829;
assign addr[49876]= 168108346;
assign addr[49877]= 15298099;
assign addr[49878]= -137589750;
assign addr[49879]= -289779648;
assign addr[49880]= -440499581;
assign addr[49881]= -588984994;
assign addr[49882]= -734482665;
assign addr[49883]= -876254528;
assign addr[49884]= -1013581418;
assign addr[49885]= -1145766716;
assign addr[49886]= -1272139887;
assign addr[49887]= -1392059879;
assign addr[49888]= -1504918373;
assign addr[49889]= -1610142873;
assign addr[49890]= -1707199606;
assign addr[49891]= -1795596234;
assign addr[49892]= -1874884346;
assign addr[49893]= -1944661739;
assign addr[49894]= -2004574453;
assign addr[49895]= -2054318569;
assign addr[49896]= -2093641749;
assign addr[49897]= -2122344521;
assign addr[49898]= -2140281282;
assign addr[49899]= -2147361045;
assign addr[49900]= -2143547897;
assign addr[49901]= -2128861181;
assign addr[49902]= -2103375398;
assign addr[49903]= -2067219829;
assign addr[49904]= -2020577882;
assign addr[49905]= -1963686155;
assign addr[49906]= -1896833245;
assign addr[49907]= -1820358275;
assign addr[49908]= -1734649179;
assign addr[49909]= -1640140734;
assign addr[49910]= -1537312353;
assign addr[49911]= -1426685652;
assign addr[49912]= -1308821808;
assign addr[49913]= -1184318708;
assign addr[49914]= -1053807919;
assign addr[49915]= -917951481;
assign addr[49916]= -777438554;
assign addr[49917]= -632981917;
assign addr[49918]= -485314355;
assign addr[49919]= -335184940;
assign addr[49920]= -183355234;
assign addr[49921]= -30595422;
assign addr[49922]= 122319591;
assign addr[49923]= 274614114;
assign addr[49924]= 425515602;
assign addr[49925]= 574258580;
assign addr[49926]= 720088517;
assign addr[49927]= 862265664;
assign addr[49928]= 1000068799;
assign addr[49929]= 1132798888;
assign addr[49930]= 1259782632;
assign addr[49931]= 1380375881;
assign addr[49932]= 1493966902;
assign addr[49933]= 1599979481;
assign addr[49934]= 1697875851;
assign addr[49935]= 1787159411;
assign addr[49936]= 1867377253;
assign addr[49937]= 1938122457;
assign addr[49938]= 1999036154;
assign addr[49939]= 2049809346;
assign addr[49940]= 2090184478;
assign addr[49941]= 2119956737;
assign addr[49942]= 2138975100;
assign addr[49943]= 2147143090;
assign addr[49944]= 2144419275;
assign addr[49945]= 2130817471;
assign addr[49946]= 2106406677;
assign addr[49947]= 2071310720;
assign addr[49948]= 2025707632;
assign addr[49949]= 1969828744;
assign addr[49950]= 1903957513;
assign addr[49951]= 1828428082;
assign addr[49952]= 1743623590;
assign addr[49953]= 1649974225;
assign addr[49954]= 1547955041;
assign addr[49955]= 1438083551;
assign addr[49956]= 1320917099;
assign addr[49957]= 1197050035;
assign addr[49958]= 1067110699;
assign addr[49959]= 931758235;
assign addr[49960]= 791679244;
assign addr[49961]= 647584304;
assign addr[49962]= 500204365;
assign addr[49963]= 350287041;
assign addr[49964]= 198592817;
assign addr[49965]= 45891193;
assign addr[49966]= -107043224;
assign addr[49967]= -259434643;
assign addr[49968]= -410510029;
assign addr[49969]= -559503022;
assign addr[49970]= -705657826;
assign addr[49971]= -848233042;
assign addr[49972]= -986505429;
assign addr[49973]= -1119773573;
assign addr[49974]= -1247361445;
assign addr[49975]= -1368621831;
assign addr[49976]= -1482939614;
assign addr[49977]= -1589734894;
assign addr[49978]= -1688465931;
assign addr[49979]= -1778631892;
assign addr[49980]= -1859775393;
assign addr[49981]= -1931484818;
assign addr[49982]= -1993396407;
assign addr[49983]= -2045196100;
assign addr[49984]= -2086621133;
assign addr[49985]= -2117461370;
assign addr[49986]= -2137560369;
assign addr[49987]= -2146816171;
assign addr[49988]= -2145181827;
assign addr[49989]= -2132665626;
assign addr[49990]= -2109331059;
assign addr[49991]= -2075296495;
assign addr[49992]= -2030734582;
assign addr[49993]= -1975871368;
assign addr[49994]= -1910985158;
assign addr[49995]= -1836405100;
assign addr[49996]= -1752509516;
assign addr[49997]= -1659723983;
assign addr[49998]= -1558519173;
assign addr[49999]= -1449408469;
assign addr[50000]= -1332945355;
assign addr[50001]= -1209720613;
assign addr[50002]= -1080359326;
assign addr[50003]= -945517704;
assign addr[50004]= -805879757;
assign addr[50005]= -662153826;
assign addr[50006]= -515068990;
assign addr[50007]= -365371365;
assign addr[50008]= -213820322;
assign addr[50009]= -61184634;
assign addr[50010]= 91761426;
assign addr[50011]= 244242007;
assign addr[50012]= 395483624;
assign addr[50013]= 544719071;
assign addr[50014]= 691191324;
assign addr[50015]= 834157373;
assign addr[50016]= 972891995;
assign addr[50017]= 1106691431;
assign addr[50018]= 1234876957;
assign addr[50019]= 1356798326;
assign addr[50020]= 1471837070;
assign addr[50021]= 1579409630;
assign addr[50022]= 1678970324;
assign addr[50023]= 1770014111;
assign addr[50024]= 1852079154;
assign addr[50025]= 1924749160;
assign addr[50026]= 1987655498;
assign addr[50027]= 2040479063;
assign addr[50028]= 2082951896;
assign addr[50029]= 2114858546;
assign addr[50030]= 2136037160;
assign addr[50031]= 2146380306;
assign addr[50032]= 2145835515;
assign addr[50033]= 2134405552;
assign addr[50034]= 2112148396;
assign addr[50035]= 2079176953;
assign addr[50036]= 2035658475;
assign addr[50037]= 1981813720;
assign addr[50038]= 1917915825;
assign addr[50039]= 1844288924;
assign addr[50040]= 1761306505;
assign addr[50041]= 1669389513;
assign addr[50042]= 1569004214;
assign addr[50043]= 1460659832;
assign addr[50044]= 1344905966;
assign addr[50045]= 1222329801;
assign addr[50046]= 1093553126;
assign addr[50047]= 959229189;
assign addr[50048]= 820039373;
assign addr[50049]= 676689746;
assign addr[50050]= 529907477;
assign addr[50051]= 380437148;
assign addr[50052]= 229036977;
assign addr[50053]= 76474970;
assign addr[50054]= -76474970;
assign addr[50055]= -229036977;
assign addr[50056]= -380437148;
assign addr[50057]= -529907477;
assign addr[50058]= -676689746;
assign addr[50059]= -820039373;
assign addr[50060]= -959229189;
assign addr[50061]= -1093553126;
assign addr[50062]= -1222329801;
assign addr[50063]= -1344905966;
assign addr[50064]= -1460659832;
assign addr[50065]= -1569004214;
assign addr[50066]= -1669389513;
assign addr[50067]= -1761306505;
assign addr[50068]= -1844288924;
assign addr[50069]= -1917915825;
assign addr[50070]= -1981813720;
assign addr[50071]= -2035658475;
assign addr[50072]= -2079176953;
assign addr[50073]= -2112148396;
assign addr[50074]= -2134405552;
assign addr[50075]= -2145835515;
assign addr[50076]= -2146380306;
assign addr[50077]= -2136037160;
assign addr[50078]= -2114858546;
assign addr[50079]= -2082951896;
assign addr[50080]= -2040479063;
assign addr[50081]= -1987655498;
assign addr[50082]= -1924749160;
assign addr[50083]= -1852079154;
assign addr[50084]= -1770014111;
assign addr[50085]= -1678970324;
assign addr[50086]= -1579409630;
assign addr[50087]= -1471837070;
assign addr[50088]= -1356798326;
assign addr[50089]= -1234876957;
assign addr[50090]= -1106691431;
assign addr[50091]= -972891995;
assign addr[50092]= -834157373;
assign addr[50093]= -691191324;
assign addr[50094]= -544719071;
assign addr[50095]= -395483624;
assign addr[50096]= -244242007;
assign addr[50097]= -91761426;
assign addr[50098]= 61184634;
assign addr[50099]= 213820322;
assign addr[50100]= 365371365;
assign addr[50101]= 515068990;
assign addr[50102]= 662153826;
assign addr[50103]= 805879757;
assign addr[50104]= 945517704;
assign addr[50105]= 1080359326;
assign addr[50106]= 1209720613;
assign addr[50107]= 1332945355;
assign addr[50108]= 1449408469;
assign addr[50109]= 1558519173;
assign addr[50110]= 1659723983;
assign addr[50111]= 1752509516;
assign addr[50112]= 1836405100;
assign addr[50113]= 1910985158;
assign addr[50114]= 1975871368;
assign addr[50115]= 2030734582;
assign addr[50116]= 2075296495;
assign addr[50117]= 2109331059;
assign addr[50118]= 2132665626;
assign addr[50119]= 2145181827;
assign addr[50120]= 2146816171;
assign addr[50121]= 2137560369;
assign addr[50122]= 2117461370;
assign addr[50123]= 2086621133;
assign addr[50124]= 2045196100;
assign addr[50125]= 1993396407;
assign addr[50126]= 1931484818;
assign addr[50127]= 1859775393;
assign addr[50128]= 1778631892;
assign addr[50129]= 1688465931;
assign addr[50130]= 1589734894;
assign addr[50131]= 1482939614;
assign addr[50132]= 1368621831;
assign addr[50133]= 1247361445;
assign addr[50134]= 1119773573;
assign addr[50135]= 986505429;
assign addr[50136]= 848233042;
assign addr[50137]= 705657826;
assign addr[50138]= 559503022;
assign addr[50139]= 410510029;
assign addr[50140]= 259434643;
assign addr[50141]= 107043224;
assign addr[50142]= -45891193;
assign addr[50143]= -198592817;
assign addr[50144]= -350287041;
assign addr[50145]= -500204365;
assign addr[50146]= -647584304;
assign addr[50147]= -791679244;
assign addr[50148]= -931758235;
assign addr[50149]= -1067110699;
assign addr[50150]= -1197050035;
assign addr[50151]= -1320917099;
assign addr[50152]= -1438083551;
assign addr[50153]= -1547955041;
assign addr[50154]= -1649974225;
assign addr[50155]= -1743623590;
assign addr[50156]= -1828428082;
assign addr[50157]= -1903957513;
assign addr[50158]= -1969828744;
assign addr[50159]= -2025707632;
assign addr[50160]= -2071310720;
assign addr[50161]= -2106406677;
assign addr[50162]= -2130817471;
assign addr[50163]= -2144419275;
assign addr[50164]= -2147143090;
assign addr[50165]= -2138975100;
assign addr[50166]= -2119956737;
assign addr[50167]= -2090184478;
assign addr[50168]= -2049809346;
assign addr[50169]= -1999036154;
assign addr[50170]= -1938122457;
assign addr[50171]= -1867377253;
assign addr[50172]= -1787159411;
assign addr[50173]= -1697875851;
assign addr[50174]= -1599979481;
assign addr[50175]= -1493966902;
assign addr[50176]= -1380375881;
assign addr[50177]= -1259782632;
assign addr[50178]= -1132798888;
assign addr[50179]= -1000068799;
assign addr[50180]= -862265664;
assign addr[50181]= -720088517;
assign addr[50182]= -574258580;
assign addr[50183]= -425515602;
assign addr[50184]= -274614114;
assign addr[50185]= -122319591;
assign addr[50186]= 30595422;
assign addr[50187]= 183355234;
assign addr[50188]= 335184940;
assign addr[50189]= 485314355;
assign addr[50190]= 632981917;
assign addr[50191]= 777438554;
assign addr[50192]= 917951481;
assign addr[50193]= 1053807919;
assign addr[50194]= 1184318708;
assign addr[50195]= 1308821808;
assign addr[50196]= 1426685652;
assign addr[50197]= 1537312353;
assign addr[50198]= 1640140734;
assign addr[50199]= 1734649179;
assign addr[50200]= 1820358275;
assign addr[50201]= 1896833245;
assign addr[50202]= 1963686155;
assign addr[50203]= 2020577882;
assign addr[50204]= 2067219829;
assign addr[50205]= 2103375398;
assign addr[50206]= 2128861181;
assign addr[50207]= 2143547897;
assign addr[50208]= 2147361045;
assign addr[50209]= 2140281282;
assign addr[50210]= 2122344521;
assign addr[50211]= 2093641749;
assign addr[50212]= 2054318569;
assign addr[50213]= 2004574453;
assign addr[50214]= 1944661739;
assign addr[50215]= 1874884346;
assign addr[50216]= 1795596234;
assign addr[50217]= 1707199606;
assign addr[50218]= 1610142873;
assign addr[50219]= 1504918373;
assign addr[50220]= 1392059879;
assign addr[50221]= 1272139887;
assign addr[50222]= 1145766716;
assign addr[50223]= 1013581418;
assign addr[50224]= 876254528;
assign addr[50225]= 734482665;
assign addr[50226]= 588984994;
assign addr[50227]= 440499581;
assign addr[50228]= 289779648;
assign addr[50229]= 137589750;
assign addr[50230]= -15298099;
assign addr[50231]= -168108346;
assign addr[50232]= -320065829;
assign addr[50233]= -470399716;
assign addr[50234]= -618347408;
assign addr[50235]= -763158411;
assign addr[50236]= -904098143;
assign addr[50237]= -1040451659;
assign addr[50238]= -1171527280;
assign addr[50239]= -1296660098;
assign addr[50240]= -1415215352;
assign addr[50241]= -1526591649;
assign addr[50242]= -1630224009;
assign addr[50243]= -1725586737;
assign addr[50244]= -1812196087;
assign addr[50245]= -1889612716;
assign addr[50246]= -1957443913;
assign addr[50247]= -2015345591;
assign addr[50248]= -2063024031;
assign addr[50249]= -2100237377;
assign addr[50250]= -2126796855;
assign addr[50251]= -2142567738;
assign addr[50252]= -2147470025;
assign addr[50253]= -2141478848;
assign addr[50254]= -2124624598;
assign addr[50255]= -2096992772;
assign addr[50256]= -2058723538;
assign addr[50257]= -2010011024;
assign addr[50258]= -1951102334;
assign addr[50259]= -1882296293;
assign addr[50260]= -1803941934;
assign addr[50261]= -1716436725;
assign addr[50262]= -1620224553;
assign addr[50263]= -1515793473;
assign addr[50264]= -1403673233;
assign addr[50265]= -1284432584;
assign addr[50266]= -1158676398;
assign addr[50267]= -1027042599;
assign addr[50268]= -890198924;
assign addr[50269]= -748839539;
assign addr[50270]= -603681519;
assign addr[50271]= -455461206;
assign addr[50272]= -304930476;
assign addr[50273]= -152852926;
assign addr[50274]= 0;
assign addr[50275]= 152852926;
assign addr[50276]= 304930476;
assign addr[50277]= 455461206;
assign addr[50278]= 603681519;
assign addr[50279]= 748839539;
assign addr[50280]= 890198924;
assign addr[50281]= 1027042599;
assign addr[50282]= 1158676398;
assign addr[50283]= 1284432584;
assign addr[50284]= 1403673233;
assign addr[50285]= 1515793473;
assign addr[50286]= 1620224553;
assign addr[50287]= 1716436725;
assign addr[50288]= 1803941934;
assign addr[50289]= 1882296293;
assign addr[50290]= 1951102334;
assign addr[50291]= 2010011024;
assign addr[50292]= 2058723538;
assign addr[50293]= 2096992772;
assign addr[50294]= 2124624598;
assign addr[50295]= 2141478848;
assign addr[50296]= 2147470025;
assign addr[50297]= 2142567738;
assign addr[50298]= 2126796855;
assign addr[50299]= 2100237377;
assign addr[50300]= 2063024031;
assign addr[50301]= 2015345591;
assign addr[50302]= 1957443913;
assign addr[50303]= 1889612716;
assign addr[50304]= 1812196087;
assign addr[50305]= 1725586737;
assign addr[50306]= 1630224009;
assign addr[50307]= 1526591649;
assign addr[50308]= 1415215352;
assign addr[50309]= 1296660098;
assign addr[50310]= 1171527280;
assign addr[50311]= 1040451659;
assign addr[50312]= 904098143;
assign addr[50313]= 763158411;
assign addr[50314]= 618347408;
assign addr[50315]= 470399716;
assign addr[50316]= 320065829;
assign addr[50317]= 168108346;
assign addr[50318]= 15298099;
assign addr[50319]= -137589750;
assign addr[50320]= -289779648;
assign addr[50321]= -440499581;
assign addr[50322]= -588984994;
assign addr[50323]= -734482665;
assign addr[50324]= -876254528;
assign addr[50325]= -1013581418;
assign addr[50326]= -1145766716;
assign addr[50327]= -1272139887;
assign addr[50328]= -1392059879;
assign addr[50329]= -1504918373;
assign addr[50330]= -1610142873;
assign addr[50331]= -1707199606;
assign addr[50332]= -1795596234;
assign addr[50333]= -1874884346;
assign addr[50334]= -1944661739;
assign addr[50335]= -2004574453;
assign addr[50336]= -2054318569;
assign addr[50337]= -2093641749;
assign addr[50338]= -2122344521;
assign addr[50339]= -2140281282;
assign addr[50340]= -2147361045;
assign addr[50341]= -2143547897;
assign addr[50342]= -2128861181;
assign addr[50343]= -2103375398;
assign addr[50344]= -2067219829;
assign addr[50345]= -2020577882;
assign addr[50346]= -1963686155;
assign addr[50347]= -1896833245;
assign addr[50348]= -1820358275;
assign addr[50349]= -1734649179;
assign addr[50350]= -1640140734;
assign addr[50351]= -1537312353;
assign addr[50352]= -1426685652;
assign addr[50353]= -1308821808;
assign addr[50354]= -1184318708;
assign addr[50355]= -1053807919;
assign addr[50356]= -917951481;
assign addr[50357]= -777438554;
assign addr[50358]= -632981917;
assign addr[50359]= -485314355;
assign addr[50360]= -335184940;
assign addr[50361]= -183355234;
assign addr[50362]= -30595422;
assign addr[50363]= 122319591;
assign addr[50364]= 274614114;
assign addr[50365]= 425515602;
assign addr[50366]= 574258580;
assign addr[50367]= 720088517;
assign addr[50368]= 862265664;
assign addr[50369]= 1000068799;
assign addr[50370]= 1132798888;
assign addr[50371]= 1259782632;
assign addr[50372]= 1380375881;
assign addr[50373]= 1493966902;
assign addr[50374]= 1599979481;
assign addr[50375]= 1697875851;
assign addr[50376]= 1787159411;
assign addr[50377]= 1867377253;
assign addr[50378]= 1938122457;
assign addr[50379]= 1999036154;
assign addr[50380]= 2049809346;
assign addr[50381]= 2090184478;
assign addr[50382]= 2119956737;
assign addr[50383]= 2138975100;
assign addr[50384]= 2147143090;
assign addr[50385]= 2144419275;
assign addr[50386]= 2130817471;
assign addr[50387]= 2106406677;
assign addr[50388]= 2071310720;
assign addr[50389]= 2025707632;
assign addr[50390]= 1969828744;
assign addr[50391]= 1903957513;
assign addr[50392]= 1828428082;
assign addr[50393]= 1743623590;
assign addr[50394]= 1649974225;
assign addr[50395]= 1547955041;
assign addr[50396]= 1438083551;
assign addr[50397]= 1320917099;
assign addr[50398]= 1197050035;
assign addr[50399]= 1067110699;
assign addr[50400]= 931758235;
assign addr[50401]= 791679244;
assign addr[50402]= 647584304;
assign addr[50403]= 500204365;
assign addr[50404]= 350287041;
assign addr[50405]= 198592817;
assign addr[50406]= 45891193;
assign addr[50407]= -107043224;
assign addr[50408]= -259434643;
assign addr[50409]= -410510029;
assign addr[50410]= -559503022;
assign addr[50411]= -705657826;
assign addr[50412]= -848233042;
assign addr[50413]= -986505429;
assign addr[50414]= -1119773573;
assign addr[50415]= -1247361445;
assign addr[50416]= -1368621831;
assign addr[50417]= -1482939614;
assign addr[50418]= -1589734894;
assign addr[50419]= -1688465931;
assign addr[50420]= -1778631892;
assign addr[50421]= -1859775393;
assign addr[50422]= -1931484818;
assign addr[50423]= -1993396407;
assign addr[50424]= -2045196100;
assign addr[50425]= -2086621133;
assign addr[50426]= -2117461370;
assign addr[50427]= -2137560369;
assign addr[50428]= -2146816171;
assign addr[50429]= -2145181827;
assign addr[50430]= -2132665626;
assign addr[50431]= -2109331059;
assign addr[50432]= -2075296495;
assign addr[50433]= -2030734582;
assign addr[50434]= -1975871368;
assign addr[50435]= -1910985158;
assign addr[50436]= -1836405100;
assign addr[50437]= -1752509516;
assign addr[50438]= -1659723983;
assign addr[50439]= -1558519173;
assign addr[50440]= -1449408469;
assign addr[50441]= -1332945355;
assign addr[50442]= -1209720613;
assign addr[50443]= -1080359326;
assign addr[50444]= -945517704;
assign addr[50445]= -805879757;
assign addr[50446]= -662153826;
assign addr[50447]= -515068990;
assign addr[50448]= -365371365;
assign addr[50449]= -213820322;
assign addr[50450]= -61184634;
assign addr[50451]= 91761426;
assign addr[50452]= 244242007;
assign addr[50453]= 395483624;
assign addr[50454]= 544719071;
assign addr[50455]= 691191324;
assign addr[50456]= 834157373;
assign addr[50457]= 972891995;
assign addr[50458]= 1106691431;
assign addr[50459]= 1234876957;
assign addr[50460]= 1356798326;
assign addr[50461]= 1471837070;
assign addr[50462]= 1579409630;
assign addr[50463]= 1678970324;
assign addr[50464]= 1770014111;
assign addr[50465]= 1852079154;
assign addr[50466]= 1924749160;
assign addr[50467]= 1987655498;
assign addr[50468]= 2040479063;
assign addr[50469]= 2082951896;
assign addr[50470]= 2114858546;
assign addr[50471]= 2136037160;
assign addr[50472]= 2146380306;
assign addr[50473]= 2145835515;
assign addr[50474]= 2134405552;
assign addr[50475]= 2112148396;
assign addr[50476]= 2079176953;
assign addr[50477]= 2035658475;
assign addr[50478]= 1981813720;
assign addr[50479]= 1917915825;
assign addr[50480]= 1844288924;
assign addr[50481]= 1761306505;
assign addr[50482]= 1669389513;
assign addr[50483]= 1569004214;
assign addr[50484]= 1460659832;
assign addr[50485]= 1344905966;
assign addr[50486]= 1222329801;
assign addr[50487]= 1093553126;
assign addr[50488]= 959229189;
assign addr[50489]= 820039373;
assign addr[50490]= 676689746;
assign addr[50491]= 529907477;
assign addr[50492]= 380437148;
assign addr[50493]= 229036977;
assign addr[50494]= 76474970;
assign addr[50495]= -76474970;
assign addr[50496]= -229036977;
assign addr[50497]= -380437148;
assign addr[50498]= -529907477;
assign addr[50499]= -676689746;
assign addr[50500]= -820039373;
assign addr[50501]= -959229189;
assign addr[50502]= -1093553126;
assign addr[50503]= -1222329801;
assign addr[50504]= -1344905966;
assign addr[50505]= -1460659832;
assign addr[50506]= -1569004214;
assign addr[50507]= -1669389513;
assign addr[50508]= -1761306505;
assign addr[50509]= -1844288924;
assign addr[50510]= -1917915825;
assign addr[50511]= -1981813720;
assign addr[50512]= -2035658475;
assign addr[50513]= -2079176953;
assign addr[50514]= -2112148396;
assign addr[50515]= -2134405552;
assign addr[50516]= -2145835515;
assign addr[50517]= -2146380306;
assign addr[50518]= -2136037160;
assign addr[50519]= -2114858546;
assign addr[50520]= -2082951896;
assign addr[50521]= -2040479063;
assign addr[50522]= -1987655498;
assign addr[50523]= -1924749160;
assign addr[50524]= -1852079154;
assign addr[50525]= -1770014111;
assign addr[50526]= -1678970324;
assign addr[50527]= -1579409630;
assign addr[50528]= -1471837070;
assign addr[50529]= -1356798326;
assign addr[50530]= -1234876957;
assign addr[50531]= -1106691431;
assign addr[50532]= -972891995;
assign addr[50533]= -834157373;
assign addr[50534]= -691191324;
assign addr[50535]= -544719071;
assign addr[50536]= -395483624;
assign addr[50537]= -244242007;
assign addr[50538]= -91761426;
assign addr[50539]= 61184634;
assign addr[50540]= 213820322;
assign addr[50541]= 365371365;
assign addr[50542]= 515068990;
assign addr[50543]= 662153826;
assign addr[50544]= 805879757;
assign addr[50545]= 945517704;
assign addr[50546]= 1080359326;
assign addr[50547]= 1209720613;
assign addr[50548]= 1332945355;
assign addr[50549]= 1449408469;
assign addr[50550]= 1558519173;
assign addr[50551]= 1659723983;
assign addr[50552]= 1752509516;
assign addr[50553]= 1836405100;
assign addr[50554]= 1910985158;
assign addr[50555]= 1975871368;
assign addr[50556]= 2030734582;
assign addr[50557]= 2075296495;
assign addr[50558]= 2109331059;
assign addr[50559]= 2132665626;
assign addr[50560]= 2145181827;
assign addr[50561]= 2146816171;
assign addr[50562]= 2137560369;
assign addr[50563]= 2117461370;
assign addr[50564]= 2086621133;
assign addr[50565]= 2045196100;
assign addr[50566]= 1993396407;
assign addr[50567]= 1931484818;
assign addr[50568]= 1859775393;
assign addr[50569]= 1778631892;
assign addr[50570]= 1688465931;
assign addr[50571]= 1589734894;
assign addr[50572]= 1482939614;
assign addr[50573]= 1368621831;
assign addr[50574]= 1247361445;
assign addr[50575]= 1119773573;
assign addr[50576]= 986505429;
assign addr[50577]= 848233042;
assign addr[50578]= 705657826;
assign addr[50579]= 559503022;
assign addr[50580]= 410510029;
assign addr[50581]= 259434643;
assign addr[50582]= 107043224;
assign addr[50583]= -45891193;
assign addr[50584]= -198592817;
assign addr[50585]= -350287041;
assign addr[50586]= -500204365;
assign addr[50587]= -647584304;
assign addr[50588]= -791679244;
assign addr[50589]= -931758235;
assign addr[50590]= -1067110699;
assign addr[50591]= -1197050035;
assign addr[50592]= -1320917099;
assign addr[50593]= -1438083551;
assign addr[50594]= -1547955041;
assign addr[50595]= -1649974225;
assign addr[50596]= -1743623590;
assign addr[50597]= -1828428082;
assign addr[50598]= -1903957513;
assign addr[50599]= -1969828744;
assign addr[50600]= -2025707632;
assign addr[50601]= -2071310720;
assign addr[50602]= -2106406677;
assign addr[50603]= -2130817471;
assign addr[50604]= -2144419275;
assign addr[50605]= -2147143090;
assign addr[50606]= -2138975100;
assign addr[50607]= -2119956737;
assign addr[50608]= -2090184478;
assign addr[50609]= -2049809346;
assign addr[50610]= -1999036154;
assign addr[50611]= -1938122457;
assign addr[50612]= -1867377253;
assign addr[50613]= -1787159411;
assign addr[50614]= -1697875851;
assign addr[50615]= -1599979481;
assign addr[50616]= -1493966902;
assign addr[50617]= -1380375881;
assign addr[50618]= -1259782632;
assign addr[50619]= -1132798888;
assign addr[50620]= -1000068799;
assign addr[50621]= -862265664;
assign addr[50622]= -720088517;
assign addr[50623]= -574258580;
assign addr[50624]= -425515602;
assign addr[50625]= -274614114;
assign addr[50626]= -122319591;
assign addr[50627]= 30595422;
assign addr[50628]= 183355234;
assign addr[50629]= 335184940;
assign addr[50630]= 485314355;
assign addr[50631]= 632981917;
assign addr[50632]= 777438554;
assign addr[50633]= 917951481;
assign addr[50634]= 1053807919;
assign addr[50635]= 1184318708;
assign addr[50636]= 1308821808;
assign addr[50637]= 1426685652;
assign addr[50638]= 1537312353;
assign addr[50639]= 1640140734;
assign addr[50640]= 1734649179;
assign addr[50641]= 1820358275;
assign addr[50642]= 1896833245;
assign addr[50643]= 1963686155;
assign addr[50644]= 2020577882;
assign addr[50645]= 2067219829;
assign addr[50646]= 2103375398;
assign addr[50647]= 2128861181;
assign addr[50648]= 2143547897;
assign addr[50649]= 2147361045;
assign addr[50650]= 2140281282;
assign addr[50651]= 2122344521;
assign addr[50652]= 2093641749;
assign addr[50653]= 2054318569;
assign addr[50654]= 2004574453;
assign addr[50655]= 1944661739;
assign addr[50656]= 1874884346;
assign addr[50657]= 1795596234;
assign addr[50658]= 1707199606;
assign addr[50659]= 1610142873;
assign addr[50660]= 1504918373;
assign addr[50661]= 1392059879;
assign addr[50662]= 1272139887;
assign addr[50663]= 1145766716;
assign addr[50664]= 1013581418;
assign addr[50665]= 876254528;
assign addr[50666]= 734482665;
assign addr[50667]= 588984994;
assign addr[50668]= 440499581;
assign addr[50669]= 289779648;
assign addr[50670]= 137589750;
assign addr[50671]= -15298099;
assign addr[50672]= -168108346;
assign addr[50673]= -320065829;
assign addr[50674]= -470399716;
assign addr[50675]= -618347408;
assign addr[50676]= -763158411;
assign addr[50677]= -904098143;
assign addr[50678]= -1040451659;
assign addr[50679]= -1171527280;
assign addr[50680]= -1296660098;
assign addr[50681]= -1415215352;
assign addr[50682]= -1526591649;
assign addr[50683]= -1630224009;
assign addr[50684]= -1725586737;
assign addr[50685]= -1812196087;
assign addr[50686]= -1889612716;
assign addr[50687]= -1957443913;
assign addr[50688]= -2015345591;
assign addr[50689]= -2063024031;
assign addr[50690]= -2100237377;
assign addr[50691]= -2126796855;
assign addr[50692]= -2142567738;
assign addr[50693]= -2147470025;
assign addr[50694]= -2141478848;
assign addr[50695]= -2124624598;
assign addr[50696]= -2096992772;
assign addr[50697]= -2058723538;
assign addr[50698]= -2010011024;
assign addr[50699]= -1951102334;
assign addr[50700]= -1882296293;
assign addr[50701]= -1803941934;
assign addr[50702]= -1716436725;
assign addr[50703]= -1620224553;
assign addr[50704]= -1515793473;
assign addr[50705]= -1403673233;
assign addr[50706]= -1284432584;
assign addr[50707]= -1158676398;
assign addr[50708]= -1027042599;
assign addr[50709]= -890198924;
assign addr[50710]= -748839539;
assign addr[50711]= -603681519;
assign addr[50712]= -455461206;
assign addr[50713]= -304930476;
assign addr[50714]= -152852926;
assign addr[50715]= 0;
assign addr[50716]= 152852926;
assign addr[50717]= 304930476;
assign addr[50718]= 455461206;
assign addr[50719]= 603681519;
assign addr[50720]= 748839539;
assign addr[50721]= 890198924;
assign addr[50722]= 1027042599;
assign addr[50723]= 1158676398;
assign addr[50724]= 1284432584;
assign addr[50725]= 1403673233;
assign addr[50726]= 1515793473;
assign addr[50727]= 1620224553;
assign addr[50728]= 1716436725;
assign addr[50729]= 1803941934;
assign addr[50730]= 1882296293;
assign addr[50731]= 1951102334;
assign addr[50732]= 2010011024;
assign addr[50733]= 2058723538;
assign addr[50734]= 2096992772;
assign addr[50735]= 2124624598;
assign addr[50736]= 2141478848;
assign addr[50737]= 2147470025;
assign addr[50738]= 2142567738;
assign addr[50739]= 2126796855;
assign addr[50740]= 2100237377;
assign addr[50741]= 2063024031;
assign addr[50742]= 2015345591;
assign addr[50743]= 1957443913;
assign addr[50744]= 1889612716;
assign addr[50745]= 1812196087;
assign addr[50746]= 1725586737;
assign addr[50747]= 1630224009;
assign addr[50748]= 1526591649;
assign addr[50749]= 1415215352;
assign addr[50750]= 1296660098;
assign addr[50751]= 1171527280;
assign addr[50752]= 1040451659;
assign addr[50753]= 904098143;
assign addr[50754]= 763158411;
assign addr[50755]= 618347408;
assign addr[50756]= 470399716;
assign addr[50757]= 320065829;
assign addr[50758]= 168108346;
assign addr[50759]= 15298099;
assign addr[50760]= -137589750;
assign addr[50761]= -289779648;
assign addr[50762]= -440499581;
assign addr[50763]= -588984994;
assign addr[50764]= -734482665;
assign addr[50765]= -876254528;
assign addr[50766]= -1013581418;
assign addr[50767]= -1145766716;
assign addr[50768]= -1272139887;
assign addr[50769]= -1392059879;
assign addr[50770]= -1504918373;
assign addr[50771]= -1610142873;
assign addr[50772]= -1707199606;
assign addr[50773]= -1795596234;
assign addr[50774]= -1874884346;
assign addr[50775]= -1944661739;
assign addr[50776]= -2004574453;
assign addr[50777]= -2054318569;
assign addr[50778]= -2093641749;
assign addr[50779]= -2122344521;
assign addr[50780]= -2140281282;
assign addr[50781]= -2147361045;
assign addr[50782]= -2143547897;
assign addr[50783]= -2128861181;
assign addr[50784]= -2103375398;
assign addr[50785]= -2067219829;
assign addr[50786]= -2020577882;
assign addr[50787]= -1963686155;
assign addr[50788]= -1896833245;
assign addr[50789]= -1820358275;
assign addr[50790]= -1734649179;
assign addr[50791]= -1640140734;
assign addr[50792]= -1537312353;
assign addr[50793]= -1426685652;
assign addr[50794]= -1308821808;
assign addr[50795]= -1184318708;
assign addr[50796]= -1053807919;
assign addr[50797]= -917951481;
assign addr[50798]= -777438554;
assign addr[50799]= -632981917;
assign addr[50800]= -485314355;
assign addr[50801]= -335184940;
assign addr[50802]= -183355234;
assign addr[50803]= -30595422;
assign addr[50804]= 122319591;
assign addr[50805]= 274614114;
assign addr[50806]= 425515602;
assign addr[50807]= 574258580;
assign addr[50808]= 720088517;
assign addr[50809]= 862265664;
assign addr[50810]= 1000068799;
assign addr[50811]= 1132798888;
assign addr[50812]= 1259782632;
assign addr[50813]= 1380375881;
assign addr[50814]= 1493966902;
assign addr[50815]= 1599979481;
assign addr[50816]= 1697875851;
assign addr[50817]= 1787159411;
assign addr[50818]= 1867377253;
assign addr[50819]= 1938122457;
assign addr[50820]= 1999036154;
assign addr[50821]= 2049809346;
assign addr[50822]= 2090184478;
assign addr[50823]= 2119956737;
assign addr[50824]= 2138975100;
assign addr[50825]= 2147143090;
assign addr[50826]= 2144419275;
assign addr[50827]= 2130817471;
assign addr[50828]= 2106406677;
assign addr[50829]= 2071310720;
assign addr[50830]= 2025707632;
assign addr[50831]= 1969828744;
assign addr[50832]= 1903957513;
assign addr[50833]= 1828428082;
assign addr[50834]= 1743623590;
assign addr[50835]= 1649974225;
assign addr[50836]= 1547955041;
assign addr[50837]= 1438083551;
assign addr[50838]= 1320917099;
assign addr[50839]= 1197050035;
assign addr[50840]= 1067110699;
assign addr[50841]= 931758235;
assign addr[50842]= 791679244;
assign addr[50843]= 647584304;
assign addr[50844]= 500204365;
assign addr[50845]= 350287041;
assign addr[50846]= 198592817;
assign addr[50847]= 45891193;
assign addr[50848]= -107043224;
assign addr[50849]= -259434643;
assign addr[50850]= -410510029;
assign addr[50851]= -559503022;
assign addr[50852]= -705657826;
assign addr[50853]= -848233042;
assign addr[50854]= -986505429;
assign addr[50855]= -1119773573;
assign addr[50856]= -1247361445;
assign addr[50857]= -1368621831;
assign addr[50858]= -1482939614;
assign addr[50859]= -1589734894;
assign addr[50860]= -1688465931;
assign addr[50861]= -1778631892;
assign addr[50862]= -1859775393;
assign addr[50863]= -1931484818;
assign addr[50864]= -1993396407;
assign addr[50865]= -2045196100;
assign addr[50866]= -2086621133;
assign addr[50867]= -2117461370;
assign addr[50868]= -2137560369;
assign addr[50869]= -2146816171;
assign addr[50870]= -2145181827;
assign addr[50871]= -2132665626;
assign addr[50872]= -2109331059;
assign addr[50873]= -2075296495;
assign addr[50874]= -2030734582;
assign addr[50875]= -1975871368;
assign addr[50876]= -1910985158;
assign addr[50877]= -1836405100;
assign addr[50878]= -1752509516;
assign addr[50879]= -1659723983;
assign addr[50880]= -1558519173;
assign addr[50881]= -1449408469;
assign addr[50882]= -1332945355;
assign addr[50883]= -1209720613;
assign addr[50884]= -1080359326;
assign addr[50885]= -945517704;
assign addr[50886]= -805879757;
assign addr[50887]= -662153826;
assign addr[50888]= -515068990;
assign addr[50889]= -365371365;
assign addr[50890]= -213820322;
assign addr[50891]= -61184634;
assign addr[50892]= 91761426;
assign addr[50893]= 244242007;
assign addr[50894]= 395483624;
assign addr[50895]= 544719071;
assign addr[50896]= 691191324;
assign addr[50897]= 834157373;
assign addr[50898]= 972891995;
assign addr[50899]= 1106691431;
assign addr[50900]= 1234876957;
assign addr[50901]= 1356798326;
assign addr[50902]= 1471837070;
assign addr[50903]= 1579409630;
assign addr[50904]= 1678970324;
assign addr[50905]= 1770014111;
assign addr[50906]= 1852079154;
assign addr[50907]= 1924749160;
assign addr[50908]= 1987655498;
assign addr[50909]= 2040479063;
assign addr[50910]= 2082951896;
assign addr[50911]= 2114858546;
assign addr[50912]= 2136037160;
assign addr[50913]= 2146380306;
assign addr[50914]= 2145835515;
assign addr[50915]= 2134405552;
assign addr[50916]= 2112148396;
assign addr[50917]= 2079176953;
assign addr[50918]= 2035658475;
assign addr[50919]= 1981813720;
assign addr[50920]= 1917915825;
assign addr[50921]= 1844288924;
assign addr[50922]= 1761306505;
assign addr[50923]= 1669389513;
assign addr[50924]= 1569004214;
assign addr[50925]= 1460659832;
assign addr[50926]= 1344905966;
assign addr[50927]= 1222329801;
assign addr[50928]= 1093553126;
assign addr[50929]= 959229189;
assign addr[50930]= 820039373;
assign addr[50931]= 676689746;
assign addr[50932]= 529907477;
assign addr[50933]= 380437148;
assign addr[50934]= 229036977;
assign addr[50935]= 76474970;
assign addr[50936]= -76474970;
assign addr[50937]= -229036977;
assign addr[50938]= -380437148;
assign addr[50939]= -529907477;
assign addr[50940]= -676689746;
assign addr[50941]= -820039373;
assign addr[50942]= -959229189;
assign addr[50943]= -1093553126;
assign addr[50944]= -1222329801;
assign addr[50945]= -1344905966;
assign addr[50946]= -1460659832;
assign addr[50947]= -1569004214;
assign addr[50948]= -1669389513;
assign addr[50949]= -1761306505;
assign addr[50950]= -1844288924;
assign addr[50951]= -1917915825;
assign addr[50952]= -1981813720;
assign addr[50953]= -2035658475;
assign addr[50954]= -2079176953;
assign addr[50955]= -2112148396;
assign addr[50956]= -2134405552;
assign addr[50957]= -2145835515;
assign addr[50958]= -2146380306;
assign addr[50959]= -2136037160;
assign addr[50960]= -2114858546;
assign addr[50961]= -2082951896;
assign addr[50962]= -2040479063;
assign addr[50963]= -1987655498;
assign addr[50964]= -1924749160;
assign addr[50965]= -1852079154;
assign addr[50966]= -1770014111;
assign addr[50967]= -1678970324;
assign addr[50968]= -1579409630;
assign addr[50969]= -1471837070;
assign addr[50970]= -1356798326;
assign addr[50971]= -1234876957;
assign addr[50972]= -1106691431;
assign addr[50973]= -972891995;
assign addr[50974]= -834157373;
assign addr[50975]= -691191324;
assign addr[50976]= -544719071;
assign addr[50977]= -395483624;
assign addr[50978]= -244242007;
assign addr[50979]= -91761426;
assign addr[50980]= 61184634;
assign addr[50981]= 213820322;
assign addr[50982]= 365371365;
assign addr[50983]= 515068990;
assign addr[50984]= 662153826;
assign addr[50985]= 805879757;
assign addr[50986]= 945517704;
assign addr[50987]= 1080359326;
assign addr[50988]= 1209720613;
assign addr[50989]= 1332945355;
assign addr[50990]= 1449408469;
assign addr[50991]= 1558519173;
assign addr[50992]= 1659723983;
assign addr[50993]= 1752509516;
assign addr[50994]= 1836405100;
assign addr[50995]= 1910985158;
assign addr[50996]= 1975871368;
assign addr[50997]= 2030734582;
assign addr[50998]= 2075296495;
assign addr[50999]= 2109331059;
assign addr[51000]= 2132665626;
assign addr[51001]= 2145181827;
assign addr[51002]= 2146816171;
assign addr[51003]= 2137560369;
assign addr[51004]= 2117461370;
assign addr[51005]= 2086621133;
assign addr[51006]= 2045196100;
assign addr[51007]= 1993396407;
assign addr[51008]= 1931484818;
assign addr[51009]= 1859775393;
assign addr[51010]= 1778631892;
assign addr[51011]= 1688465931;
assign addr[51012]= 1589734894;
assign addr[51013]= 1482939614;
assign addr[51014]= 1368621831;
assign addr[51015]= 1247361445;
assign addr[51016]= 1119773573;
assign addr[51017]= 986505429;
assign addr[51018]= 848233042;
assign addr[51019]= 705657826;
assign addr[51020]= 559503022;
assign addr[51021]= 410510029;
assign addr[51022]= 259434643;
assign addr[51023]= 107043224;
assign addr[51024]= -45891193;
assign addr[51025]= -198592817;
assign addr[51026]= -350287041;
assign addr[51027]= -500204365;
assign addr[51028]= -647584304;
assign addr[51029]= -791679244;
assign addr[51030]= -931758235;
assign addr[51031]= -1067110699;
assign addr[51032]= -1197050035;
assign addr[51033]= -1320917099;
assign addr[51034]= -1438083551;
assign addr[51035]= -1547955041;
assign addr[51036]= -1649974225;
assign addr[51037]= -1743623590;
assign addr[51038]= -1828428082;
assign addr[51039]= -1903957513;
assign addr[51040]= -1969828744;
assign addr[51041]= -2025707632;
assign addr[51042]= -2071310720;
assign addr[51043]= -2106406677;
assign addr[51044]= -2130817471;
assign addr[51045]= -2144419275;
assign addr[51046]= -2147143090;
assign addr[51047]= -2138975100;
assign addr[51048]= -2119956737;
assign addr[51049]= -2090184478;
assign addr[51050]= -2049809346;
assign addr[51051]= -1999036154;
assign addr[51052]= -1938122457;
assign addr[51053]= -1867377253;
assign addr[51054]= -1787159411;
assign addr[51055]= -1697875851;
assign addr[51056]= -1599979481;
assign addr[51057]= -1493966902;
assign addr[51058]= -1380375881;
assign addr[51059]= -1259782632;
assign addr[51060]= -1132798888;
assign addr[51061]= -1000068799;
assign addr[51062]= -862265664;
assign addr[51063]= -720088517;
assign addr[51064]= -574258580;
assign addr[51065]= -425515602;
assign addr[51066]= -274614114;
assign addr[51067]= -122319591;
assign addr[51068]= 30595422;
assign addr[51069]= 183355234;
assign addr[51070]= 335184940;
assign addr[51071]= 485314355;
assign addr[51072]= 632981917;
assign addr[51073]= 777438554;
assign addr[51074]= 917951481;
assign addr[51075]= 1053807919;
assign addr[51076]= 1184318708;
assign addr[51077]= 1308821808;
assign addr[51078]= 1426685652;
assign addr[51079]= 1537312353;
assign addr[51080]= 1640140734;
assign addr[51081]= 1734649179;
assign addr[51082]= 1820358275;
assign addr[51083]= 1896833245;
assign addr[51084]= 1963686155;
assign addr[51085]= 2020577882;
assign addr[51086]= 2067219829;
assign addr[51087]= 2103375398;
assign addr[51088]= 2128861181;
assign addr[51089]= 2143547897;
assign addr[51090]= 2147361045;
assign addr[51091]= 2140281282;
assign addr[51092]= 2122344521;
assign addr[51093]= 2093641749;
assign addr[51094]= 2054318569;
assign addr[51095]= 2004574453;
assign addr[51096]= 1944661739;
assign addr[51097]= 1874884346;
assign addr[51098]= 1795596234;
assign addr[51099]= 1707199606;
assign addr[51100]= 1610142873;
assign addr[51101]= 1504918373;
assign addr[51102]= 1392059879;
assign addr[51103]= 1272139887;
assign addr[51104]= 1145766716;
assign addr[51105]= 1013581418;
assign addr[51106]= 876254528;
assign addr[51107]= 734482665;
assign addr[51108]= 588984994;
assign addr[51109]= 440499581;
assign addr[51110]= 289779648;
assign addr[51111]= 137589750;
assign addr[51112]= -15298099;
assign addr[51113]= -168108346;
assign addr[51114]= -320065829;
assign addr[51115]= -470399716;
assign addr[51116]= -618347408;
assign addr[51117]= -763158411;
assign addr[51118]= -904098143;
assign addr[51119]= -1040451659;
assign addr[51120]= -1171527280;
assign addr[51121]= -1296660098;
assign addr[51122]= -1415215352;
assign addr[51123]= -1526591649;
assign addr[51124]= -1630224009;
assign addr[51125]= -1725586737;
assign addr[51126]= -1812196087;
assign addr[51127]= -1889612716;
assign addr[51128]= -1957443913;
assign addr[51129]= -2015345591;
assign addr[51130]= -2063024031;
assign addr[51131]= -2100237377;
assign addr[51132]= -2126796855;
assign addr[51133]= -2142567738;
assign addr[51134]= -2147470025;
assign addr[51135]= -2141478848;
assign addr[51136]= -2124624598;
assign addr[51137]= -2096992772;
assign addr[51138]= -2058723538;
assign addr[51139]= -2010011024;
assign addr[51140]= -1951102334;
assign addr[51141]= -1882296293;
assign addr[51142]= -1803941934;
assign addr[51143]= -1716436725;
assign addr[51144]= -1620224553;
assign addr[51145]= -1515793473;
assign addr[51146]= -1403673233;
assign addr[51147]= -1284432584;
assign addr[51148]= -1158676398;
assign addr[51149]= -1027042599;
assign addr[51150]= -890198924;
assign addr[51151]= -748839539;
assign addr[51152]= -603681519;
assign addr[51153]= -455461206;
assign addr[51154]= -304930476;
assign addr[51155]= -152852926;
assign addr[51156]= 0;
assign addr[51157]= 152852926;
assign addr[51158]= 304930476;
assign addr[51159]= 455461206;
assign addr[51160]= 603681519;
assign addr[51161]= 748839539;
assign addr[51162]= 890198924;
assign addr[51163]= 1027042599;
assign addr[51164]= 1158676398;
assign addr[51165]= 1284432584;
assign addr[51166]= 1403673233;
assign addr[51167]= 1515793473;
assign addr[51168]= 1620224553;
assign addr[51169]= 1716436725;
assign addr[51170]= 1803941934;
assign addr[51171]= 1882296293;
assign addr[51172]= 1951102334;
assign addr[51173]= 2010011024;
assign addr[51174]= 2058723538;
assign addr[51175]= 2096992772;
assign addr[51176]= 2124624598;
assign addr[51177]= 2141478848;
assign addr[51178]= 2147470025;
assign addr[51179]= 2142567738;
assign addr[51180]= 2126796855;
assign addr[51181]= 2100237377;
assign addr[51182]= 2063024031;
assign addr[51183]= 2015345591;
assign addr[51184]= 1957443913;
assign addr[51185]= 1889612716;
assign addr[51186]= 1812196087;
assign addr[51187]= 1725586737;
assign addr[51188]= 1630224009;
assign addr[51189]= 1526591649;
assign addr[51190]= 1415215352;
assign addr[51191]= 1296660098;
assign addr[51192]= 1171527280;
assign addr[51193]= 1040451659;
assign addr[51194]= 904098143;
assign addr[51195]= 763158411;
assign addr[51196]= 618347408;
assign addr[51197]= 470399716;
assign addr[51198]= 320065829;
assign addr[51199]= 168108346;
assign addr[51200]= 15298099;
assign addr[51201]= -137589750;
assign addr[51202]= -289779648;
assign addr[51203]= -440499581;
assign addr[51204]= -588984994;
assign addr[51205]= -734482665;
assign addr[51206]= -876254528;
assign addr[51207]= -1013581418;
assign addr[51208]= -1145766716;
assign addr[51209]= -1272139887;
assign addr[51210]= -1392059879;
assign addr[51211]= -1504918373;
assign addr[51212]= -1610142873;
assign addr[51213]= -1707199606;
assign addr[51214]= -1795596234;
assign addr[51215]= -1874884346;
assign addr[51216]= -1944661739;
assign addr[51217]= -2004574453;
assign addr[51218]= -2054318569;
assign addr[51219]= -2093641749;
assign addr[51220]= -2122344521;
assign addr[51221]= -2140281282;
assign addr[51222]= -2147361045;
assign addr[51223]= -2143547897;
assign addr[51224]= -2128861181;
assign addr[51225]= -2103375398;
assign addr[51226]= -2067219829;
assign addr[51227]= -2020577882;
assign addr[51228]= -1963686155;
assign addr[51229]= -1896833245;
assign addr[51230]= -1820358275;
assign addr[51231]= -1734649179;
assign addr[51232]= -1640140734;
assign addr[51233]= -1537312353;
assign addr[51234]= -1426685652;
assign addr[51235]= -1308821808;
assign addr[51236]= -1184318708;
assign addr[51237]= -1053807919;
assign addr[51238]= -917951481;
assign addr[51239]= -777438554;
assign addr[51240]= -632981917;
assign addr[51241]= -485314355;
assign addr[51242]= -335184940;
assign addr[51243]= -183355234;
assign addr[51244]= -30595422;
assign addr[51245]= 122319591;
assign addr[51246]= 274614114;
assign addr[51247]= 425515602;
assign addr[51248]= 574258580;
assign addr[51249]= 720088517;
assign addr[51250]= 862265664;
assign addr[51251]= 1000068799;
assign addr[51252]= 1132798888;
assign addr[51253]= 1259782632;
assign addr[51254]= 1380375881;
assign addr[51255]= 1493966902;
assign addr[51256]= 1599979481;
assign addr[51257]= 1697875851;
assign addr[51258]= 1787159411;
assign addr[51259]= 1867377253;
assign addr[51260]= 1938122457;
assign addr[51261]= 1999036154;
assign addr[51262]= 2049809346;
assign addr[51263]= 2090184478;
assign addr[51264]= 2119956737;
assign addr[51265]= 2138975100;
assign addr[51266]= 2147143090;
assign addr[51267]= 2144419275;
assign addr[51268]= 2130817471;
assign addr[51269]= 2106406677;
assign addr[51270]= 2071310720;
assign addr[51271]= 2025707632;
assign addr[51272]= 1969828744;
assign addr[51273]= 1903957513;
assign addr[51274]= 1828428082;
assign addr[51275]= 1743623590;
assign addr[51276]= 1649974225;
assign addr[51277]= 1547955041;
assign addr[51278]= 1438083551;
assign addr[51279]= 1320917099;
assign addr[51280]= 1197050035;
assign addr[51281]= 1067110699;
assign addr[51282]= 931758235;
assign addr[51283]= 791679244;
assign addr[51284]= 647584304;
assign addr[51285]= 500204365;
assign addr[51286]= 350287041;
assign addr[51287]= 198592817;
assign addr[51288]= 45891193;
assign addr[51289]= -107043224;
assign addr[51290]= -259434643;
assign addr[51291]= -410510029;
assign addr[51292]= -559503022;
assign addr[51293]= -705657826;
assign addr[51294]= -848233042;
assign addr[51295]= -986505429;
assign addr[51296]= -1119773573;
assign addr[51297]= -1247361445;
assign addr[51298]= -1368621831;
assign addr[51299]= -1482939614;
assign addr[51300]= -1589734894;
assign addr[51301]= -1688465931;
assign addr[51302]= -1778631892;
assign addr[51303]= -1859775393;
assign addr[51304]= -1931484818;
assign addr[51305]= -1993396407;
assign addr[51306]= -2045196100;
assign addr[51307]= -2086621133;
assign addr[51308]= -2117461370;
assign addr[51309]= -2137560369;
assign addr[51310]= -2146816171;
assign addr[51311]= -2145181827;
assign addr[51312]= -2132665626;
assign addr[51313]= -2109331059;
assign addr[51314]= -2075296495;
assign addr[51315]= -2030734582;
assign addr[51316]= -1975871368;
assign addr[51317]= -1910985158;
assign addr[51318]= -1836405100;
assign addr[51319]= -1752509516;
assign addr[51320]= -1659723983;
assign addr[51321]= -1558519173;
assign addr[51322]= -1449408469;
assign addr[51323]= -1332945355;
assign addr[51324]= -1209720613;
assign addr[51325]= -1080359326;
assign addr[51326]= -945517704;
assign addr[51327]= -805879757;
assign addr[51328]= -662153826;
assign addr[51329]= -515068990;
assign addr[51330]= -365371365;
assign addr[51331]= -213820322;
assign addr[51332]= -61184634;
assign addr[51333]= 91761426;
assign addr[51334]= 244242007;
assign addr[51335]= 395483624;
assign addr[51336]= 544719071;
assign addr[51337]= 691191324;
assign addr[51338]= 834157373;
assign addr[51339]= 972891995;
assign addr[51340]= 1106691431;
assign addr[51341]= 1234876957;
assign addr[51342]= 1356798326;
assign addr[51343]= 1471837070;
assign addr[51344]= 1579409630;
assign addr[51345]= 1678970324;
assign addr[51346]= 1770014111;
assign addr[51347]= 1852079154;
assign addr[51348]= 1924749160;
assign addr[51349]= 1987655498;
assign addr[51350]= 2040479063;
assign addr[51351]= 2082951896;
assign addr[51352]= 2114858546;
assign addr[51353]= 2136037160;
assign addr[51354]= 2146380306;
assign addr[51355]= 2145835515;
assign addr[51356]= 2134405552;
assign addr[51357]= 2112148396;
assign addr[51358]= 2079176953;
assign addr[51359]= 2035658475;
assign addr[51360]= 1981813720;
assign addr[51361]= 1917915825;
assign addr[51362]= 1844288924;
assign addr[51363]= 1761306505;
assign addr[51364]= 1669389513;
assign addr[51365]= 1569004214;
assign addr[51366]= 1460659832;
assign addr[51367]= 1344905966;
assign addr[51368]= 1222329801;
assign addr[51369]= 1093553126;
assign addr[51370]= 959229189;
assign addr[51371]= 820039373;
assign addr[51372]= 676689746;
assign addr[51373]= 529907477;
assign addr[51374]= 380437148;
assign addr[51375]= 229036977;
assign addr[51376]= 76474970;
assign addr[51377]= -76474970;
assign addr[51378]= -229036977;
assign addr[51379]= -380437148;
assign addr[51380]= -529907477;
assign addr[51381]= -676689746;
assign addr[51382]= -820039373;
assign addr[51383]= -959229189;
assign addr[51384]= -1093553126;
assign addr[51385]= -1222329801;
assign addr[51386]= -1344905966;
assign addr[51387]= -1460659832;
assign addr[51388]= -1569004214;
assign addr[51389]= -1669389513;
assign addr[51390]= -1761306505;
assign addr[51391]= -1844288924;
assign addr[51392]= -1917915825;
assign addr[51393]= -1981813720;
assign addr[51394]= -2035658475;
assign addr[51395]= -2079176953;
assign addr[51396]= -2112148396;
assign addr[51397]= -2134405552;
assign addr[51398]= -2145835515;
assign addr[51399]= -2146380306;
assign addr[51400]= -2136037160;
assign addr[51401]= -2114858546;
assign addr[51402]= -2082951896;
assign addr[51403]= -2040479063;
assign addr[51404]= -1987655498;
assign addr[51405]= -1924749160;
assign addr[51406]= -1852079154;
assign addr[51407]= -1770014111;
assign addr[51408]= -1678970324;
assign addr[51409]= -1579409630;
assign addr[51410]= -1471837070;
assign addr[51411]= -1356798326;
assign addr[51412]= -1234876957;
assign addr[51413]= -1106691431;
assign addr[51414]= -972891995;
assign addr[51415]= -834157373;
assign addr[51416]= -691191324;
assign addr[51417]= -544719071;
assign addr[51418]= -395483624;
assign addr[51419]= -244242007;
assign addr[51420]= -91761426;
assign addr[51421]= 61184634;
assign addr[51422]= 213820322;
assign addr[51423]= 365371365;
assign addr[51424]= 515068990;
assign addr[51425]= 662153826;
assign addr[51426]= 805879757;
assign addr[51427]= 945517704;
assign addr[51428]= 1080359326;
assign addr[51429]= 1209720613;
assign addr[51430]= 1332945355;
assign addr[51431]= 1449408469;
assign addr[51432]= 1558519173;
assign addr[51433]= 1659723983;
assign addr[51434]= 1752509516;
assign addr[51435]= 1836405100;
assign addr[51436]= 1910985158;
assign addr[51437]= 1975871368;
assign addr[51438]= 2030734582;
assign addr[51439]= 2075296495;
assign addr[51440]= 2109331059;
assign addr[51441]= 2132665626;
assign addr[51442]= 2145181827;
assign addr[51443]= 2146816171;
assign addr[51444]= 2137560369;
assign addr[51445]= 2117461370;
assign addr[51446]= 2086621133;
assign addr[51447]= 2045196100;
assign addr[51448]= 1993396407;
assign addr[51449]= 1931484818;
assign addr[51450]= 1859775393;
assign addr[51451]= 1778631892;
assign addr[51452]= 1688465931;
assign addr[51453]= 1589734894;
assign addr[51454]= 1482939614;
assign addr[51455]= 1368621831;
assign addr[51456]= 1247361445;
assign addr[51457]= 1119773573;
assign addr[51458]= 986505429;
assign addr[51459]= 848233042;
assign addr[51460]= 705657826;
assign addr[51461]= 559503022;
assign addr[51462]= 410510029;
assign addr[51463]= 259434643;
assign addr[51464]= 107043224;
assign addr[51465]= -45891193;
assign addr[51466]= -198592817;
assign addr[51467]= -350287041;
assign addr[51468]= -500204365;
assign addr[51469]= -647584304;
assign addr[51470]= -791679244;
assign addr[51471]= -931758235;
assign addr[51472]= -1067110699;
assign addr[51473]= -1197050035;
assign addr[51474]= -1320917099;
assign addr[51475]= -1438083551;
assign addr[51476]= -1547955041;
assign addr[51477]= -1649974225;
assign addr[51478]= -1743623590;
assign addr[51479]= -1828428082;
assign addr[51480]= -1903957513;
assign addr[51481]= -1969828744;
assign addr[51482]= -2025707632;
assign addr[51483]= -2071310720;
assign addr[51484]= -2106406677;
assign addr[51485]= -2130817471;
assign addr[51486]= -2144419275;
assign addr[51487]= -2147143090;
assign addr[51488]= -2138975100;
assign addr[51489]= -2119956737;
assign addr[51490]= -2090184478;
assign addr[51491]= -2049809346;
assign addr[51492]= -1999036154;
assign addr[51493]= -1938122457;
assign addr[51494]= -1867377253;
assign addr[51495]= -1787159411;
assign addr[51496]= -1697875851;
assign addr[51497]= -1599979481;
assign addr[51498]= -1493966902;
assign addr[51499]= -1380375881;
assign addr[51500]= -1259782632;
assign addr[51501]= -1132798888;
assign addr[51502]= -1000068799;
assign addr[51503]= -862265664;
assign addr[51504]= -720088517;
assign addr[51505]= -574258580;
assign addr[51506]= -425515602;
assign addr[51507]= -274614114;
assign addr[51508]= -122319591;
assign addr[51509]= 30595422;
assign addr[51510]= 183355234;
assign addr[51511]= 335184940;
assign addr[51512]= 485314355;
assign addr[51513]= 632981917;
assign addr[51514]= 777438554;
assign addr[51515]= 917951481;
assign addr[51516]= 1053807919;
assign addr[51517]= 1184318708;
assign addr[51518]= 1308821808;
assign addr[51519]= 1426685652;
assign addr[51520]= 1537312353;
assign addr[51521]= 1640140734;
assign addr[51522]= 1734649179;
assign addr[51523]= 1820358275;
assign addr[51524]= 1896833245;
assign addr[51525]= 1963686155;
assign addr[51526]= 2020577882;
assign addr[51527]= 2067219829;
assign addr[51528]= 2103375398;
assign addr[51529]= 2128861181;
assign addr[51530]= 2143547897;
assign addr[51531]= 2147361045;
assign addr[51532]= 2140281282;
assign addr[51533]= 2122344521;
assign addr[51534]= 2093641749;
assign addr[51535]= 2054318569;
assign addr[51536]= 2004574453;
assign addr[51537]= 1944661739;
assign addr[51538]= 1874884346;
assign addr[51539]= 1795596234;
assign addr[51540]= 1707199606;
assign addr[51541]= 1610142873;
assign addr[51542]= 1504918373;
assign addr[51543]= 1392059879;
assign addr[51544]= 1272139887;
assign addr[51545]= 1145766716;
assign addr[51546]= 1013581418;
assign addr[51547]= 876254528;
assign addr[51548]= 734482665;
assign addr[51549]= 588984994;
assign addr[51550]= 440499581;
assign addr[51551]= 289779648;
assign addr[51552]= 137589750;
assign addr[51553]= -15298099;
assign addr[51554]= -168108346;
assign addr[51555]= -320065829;
assign addr[51556]= -470399716;
assign addr[51557]= -618347408;
assign addr[51558]= -763158411;
assign addr[51559]= -904098143;
assign addr[51560]= -1040451659;
assign addr[51561]= -1171527280;
assign addr[51562]= -1296660098;
assign addr[51563]= -1415215352;
assign addr[51564]= -1526591649;
assign addr[51565]= -1630224009;
assign addr[51566]= -1725586737;
assign addr[51567]= -1812196087;
assign addr[51568]= -1889612716;
assign addr[51569]= -1957443913;
assign addr[51570]= -2015345591;
assign addr[51571]= -2063024031;
assign addr[51572]= -2100237377;
assign addr[51573]= -2126796855;
assign addr[51574]= -2142567738;
assign addr[51575]= -2147470025;
assign addr[51576]= -2141478848;
assign addr[51577]= -2124624598;
assign addr[51578]= -2096992772;
assign addr[51579]= -2058723538;
assign addr[51580]= -2010011024;
assign addr[51581]= -1951102334;
assign addr[51582]= -1882296293;
assign addr[51583]= -1803941934;
assign addr[51584]= -1716436725;
assign addr[51585]= -1620224553;
assign addr[51586]= -1515793473;
assign addr[51587]= -1403673233;
assign addr[51588]= -1284432584;
assign addr[51589]= -1158676398;
assign addr[51590]= -1027042599;
assign addr[51591]= -890198924;
assign addr[51592]= -748839539;
assign addr[51593]= -603681519;
assign addr[51594]= -455461206;
assign addr[51595]= -304930476;
assign addr[51596]= -152852926;
assign addr[51597]= 0;
assign addr[51598]= 152852926;
assign addr[51599]= 304930476;
assign addr[51600]= 455461206;
assign addr[51601]= 603681519;
assign addr[51602]= 748839539;
assign addr[51603]= 890198924;
assign addr[51604]= 1027042599;
assign addr[51605]= 1158676398;
assign addr[51606]= 1284432584;
assign addr[51607]= 1403673233;
assign addr[51608]= 1515793473;
assign addr[51609]= 1620224553;
assign addr[51610]= 1716436725;
assign addr[51611]= 1803941934;
assign addr[51612]= 1882296293;
assign addr[51613]= 1951102334;
assign addr[51614]= 2010011024;
assign addr[51615]= 2058723538;
assign addr[51616]= 2096992772;
assign addr[51617]= 2124624598;
assign addr[51618]= 2141478848;
assign addr[51619]= 2147470025;
assign addr[51620]= 2142567738;
assign addr[51621]= 2126796855;
assign addr[51622]= 2100237377;
assign addr[51623]= 2063024031;
assign addr[51624]= 2015345591;
assign addr[51625]= 1957443913;
assign addr[51626]= 1889612716;
assign addr[51627]= 1812196087;
assign addr[51628]= 1725586737;
assign addr[51629]= 1630224009;
assign addr[51630]= 1526591649;
assign addr[51631]= 1415215352;
assign addr[51632]= 1296660098;
assign addr[51633]= 1171527280;
assign addr[51634]= 1040451659;
assign addr[51635]= 904098143;
assign addr[51636]= 763158411;
assign addr[51637]= 618347408;
assign addr[51638]= 470399716;
assign addr[51639]= 320065829;
assign addr[51640]= 168108346;
assign addr[51641]= 15298099;
assign addr[51642]= -137589750;
assign addr[51643]= -289779648;
assign addr[51644]= -440499581;
assign addr[51645]= -588984994;
assign addr[51646]= -734482665;
assign addr[51647]= -876254528;
assign addr[51648]= -1013581418;
assign addr[51649]= -1145766716;
assign addr[51650]= -1272139887;
assign addr[51651]= -1392059879;
assign addr[51652]= -1504918373;
assign addr[51653]= -1610142873;
assign addr[51654]= -1707199606;
assign addr[51655]= -1795596234;
assign addr[51656]= -1874884346;
assign addr[51657]= -1944661739;
assign addr[51658]= -2004574453;
assign addr[51659]= -2054318569;
assign addr[51660]= -2093641749;
assign addr[51661]= -2122344521;
assign addr[51662]= -2140281282;
assign addr[51663]= -2147361045;
assign addr[51664]= -2143547897;
assign addr[51665]= -2128861181;
assign addr[51666]= -2103375398;
assign addr[51667]= -2067219829;
assign addr[51668]= -2020577882;
assign addr[51669]= -1963686155;
assign addr[51670]= -1896833245;
assign addr[51671]= -1820358275;
assign addr[51672]= -1734649179;
assign addr[51673]= -1640140734;
assign addr[51674]= -1537312353;
assign addr[51675]= -1426685652;
assign addr[51676]= -1308821808;
assign addr[51677]= -1184318708;
assign addr[51678]= -1053807919;
assign addr[51679]= -917951481;
assign addr[51680]= -777438554;
assign addr[51681]= -632981917;
assign addr[51682]= -485314355;
assign addr[51683]= -335184940;
assign addr[51684]= -183355234;
assign addr[51685]= -30595422;
assign addr[51686]= 122319591;
assign addr[51687]= 274614114;
assign addr[51688]= 425515602;
assign addr[51689]= 574258580;
assign addr[51690]= 720088517;
assign addr[51691]= 862265664;
assign addr[51692]= 1000068799;
assign addr[51693]= 1132798888;
assign addr[51694]= 1259782632;
assign addr[51695]= 1380375881;
assign addr[51696]= 1493966902;
assign addr[51697]= 1599979481;
assign addr[51698]= 1697875851;
assign addr[51699]= 1787159411;
assign addr[51700]= 1867377253;
assign addr[51701]= 1938122457;
assign addr[51702]= 1999036154;
assign addr[51703]= 2049809346;
assign addr[51704]= 2090184478;
assign addr[51705]= 2119956737;
assign addr[51706]= 2138975100;
assign addr[51707]= 2147143090;
assign addr[51708]= 2144419275;
assign addr[51709]= 2130817471;
assign addr[51710]= 2106406677;
assign addr[51711]= 2071310720;
assign addr[51712]= 2025707632;
assign addr[51713]= 1969828744;
assign addr[51714]= 1903957513;
assign addr[51715]= 1828428082;
assign addr[51716]= 1743623590;
assign addr[51717]= 1649974225;
assign addr[51718]= 1547955041;
assign addr[51719]= 1438083551;
assign addr[51720]= 1320917099;
assign addr[51721]= 1197050035;
assign addr[51722]= 1067110699;
assign addr[51723]= 931758235;
assign addr[51724]= 791679244;
assign addr[51725]= 647584304;
assign addr[51726]= 500204365;
assign addr[51727]= 350287041;
assign addr[51728]= 198592817;
assign addr[51729]= 45891193;
assign addr[51730]= -107043224;
assign addr[51731]= -259434643;
assign addr[51732]= -410510029;
assign addr[51733]= -559503022;
assign addr[51734]= -705657826;
assign addr[51735]= -848233042;
assign addr[51736]= -986505429;
assign addr[51737]= -1119773573;
assign addr[51738]= -1247361445;
assign addr[51739]= -1368621831;
assign addr[51740]= -1482939614;
assign addr[51741]= -1589734894;
assign addr[51742]= -1688465931;
assign addr[51743]= -1778631892;
assign addr[51744]= -1859775393;
assign addr[51745]= -1931484818;
assign addr[51746]= -1993396407;
assign addr[51747]= -2045196100;
assign addr[51748]= -2086621133;
assign addr[51749]= -2117461370;
assign addr[51750]= -2137560369;
assign addr[51751]= -2146816171;
assign addr[51752]= -2145181827;
assign addr[51753]= -2132665626;
assign addr[51754]= -2109331059;
assign addr[51755]= -2075296495;
assign addr[51756]= -2030734582;
assign addr[51757]= -1975871368;
assign addr[51758]= -1910985158;
assign addr[51759]= -1836405100;
assign addr[51760]= -1752509516;
assign addr[51761]= -1659723983;
assign addr[51762]= -1558519173;
assign addr[51763]= -1449408469;
assign addr[51764]= -1332945355;
assign addr[51765]= -1209720613;
assign addr[51766]= -1080359326;
assign addr[51767]= -945517704;
assign addr[51768]= -805879757;
assign addr[51769]= -662153826;
assign addr[51770]= -515068990;
assign addr[51771]= -365371365;
assign addr[51772]= -213820322;
assign addr[51773]= -61184634;
assign addr[51774]= 91761426;
assign addr[51775]= 244242007;
assign addr[51776]= 395483624;
assign addr[51777]= 544719071;
assign addr[51778]= 691191324;
assign addr[51779]= 834157373;
assign addr[51780]= 972891995;
assign addr[51781]= 1106691431;
assign addr[51782]= 1234876957;
assign addr[51783]= 1356798326;
assign addr[51784]= 1471837070;
assign addr[51785]= 1579409630;
assign addr[51786]= 1678970324;
assign addr[51787]= 1770014111;
assign addr[51788]= 1852079154;
assign addr[51789]= 1924749160;
assign addr[51790]= 1987655498;
assign addr[51791]= 2040479063;
assign addr[51792]= 2082951896;
assign addr[51793]= 2114858546;
assign addr[51794]= 2136037160;
assign addr[51795]= 2146380306;
assign addr[51796]= 2145835515;
assign addr[51797]= 2134405552;
assign addr[51798]= 2112148396;
assign addr[51799]= 2079176953;
assign addr[51800]= 2035658475;
assign addr[51801]= 1981813720;
assign addr[51802]= 1917915825;
assign addr[51803]= 1844288924;
assign addr[51804]= 1761306505;
assign addr[51805]= 1669389513;
assign addr[51806]= 1569004214;
assign addr[51807]= 1460659832;
assign addr[51808]= 1344905966;
assign addr[51809]= 1222329801;
assign addr[51810]= 1093553126;
assign addr[51811]= 959229189;
assign addr[51812]= 820039373;
assign addr[51813]= 676689746;
assign addr[51814]= 529907477;
assign addr[51815]= 380437148;
assign addr[51816]= 229036977;
assign addr[51817]= 76474970;
assign addr[51818]= -76474970;
assign addr[51819]= -229036977;
assign addr[51820]= -380437148;
assign addr[51821]= -529907477;
assign addr[51822]= -676689746;
assign addr[51823]= -820039373;
assign addr[51824]= -959229189;
assign addr[51825]= -1093553126;
assign addr[51826]= -1222329801;
assign addr[51827]= -1344905966;
assign addr[51828]= -1460659832;
assign addr[51829]= -1569004214;
assign addr[51830]= -1669389513;
assign addr[51831]= -1761306505;
assign addr[51832]= -1844288924;
assign addr[51833]= -1917915825;
assign addr[51834]= -1981813720;
assign addr[51835]= -2035658475;
assign addr[51836]= -2079176953;
assign addr[51837]= -2112148396;
assign addr[51838]= -2134405552;
assign addr[51839]= -2145835515;
assign addr[51840]= -2146380306;
assign addr[51841]= -2136037160;
assign addr[51842]= -2114858546;
assign addr[51843]= -2082951896;
assign addr[51844]= -2040479063;
assign addr[51845]= -1987655498;
assign addr[51846]= -1924749160;
assign addr[51847]= -1852079154;
assign addr[51848]= -1770014111;
assign addr[51849]= -1678970324;
assign addr[51850]= -1579409630;
assign addr[51851]= -1471837070;
assign addr[51852]= -1356798326;
assign addr[51853]= -1234876957;
assign addr[51854]= -1106691431;
assign addr[51855]= -972891995;
assign addr[51856]= -834157373;
assign addr[51857]= -691191324;
assign addr[51858]= -544719071;
assign addr[51859]= -395483624;
assign addr[51860]= -244242007;
assign addr[51861]= -91761426;
assign addr[51862]= 61184634;
assign addr[51863]= 213820322;
assign addr[51864]= 365371365;
assign addr[51865]= 515068990;
assign addr[51866]= 662153826;
assign addr[51867]= 805879757;
assign addr[51868]= 945517704;
assign addr[51869]= 1080359326;
assign addr[51870]= 1209720613;
assign addr[51871]= 1332945355;
assign addr[51872]= 1449408469;
assign addr[51873]= 1558519173;
assign addr[51874]= 1659723983;
assign addr[51875]= 1752509516;
assign addr[51876]= 1836405100;
assign addr[51877]= 1910985158;
assign addr[51878]= 1975871368;
assign addr[51879]= 2030734582;
assign addr[51880]= 2075296495;
assign addr[51881]= 2109331059;
assign addr[51882]= 2132665626;
assign addr[51883]= 2145181827;
assign addr[51884]= 2146816171;
assign addr[51885]= 2137560369;
assign addr[51886]= 2117461370;
assign addr[51887]= 2086621133;
assign addr[51888]= 2045196100;
assign addr[51889]= 1993396407;
assign addr[51890]= 1931484818;
assign addr[51891]= 1859775393;
assign addr[51892]= 1778631892;
assign addr[51893]= 1688465931;
assign addr[51894]= 1589734894;
assign addr[51895]= 1482939614;
assign addr[51896]= 1368621831;
assign addr[51897]= 1247361445;
assign addr[51898]= 1119773573;
assign addr[51899]= 986505429;
assign addr[51900]= 848233042;
assign addr[51901]= 705657826;
assign addr[51902]= 559503022;
assign addr[51903]= 410510029;
assign addr[51904]= 259434643;
assign addr[51905]= 107043224;
assign addr[51906]= -45891193;
assign addr[51907]= -198592817;
assign addr[51908]= -350287041;
assign addr[51909]= -500204365;
assign addr[51910]= -647584304;
assign addr[51911]= -791679244;
assign addr[51912]= -931758235;
assign addr[51913]= -1067110699;
assign addr[51914]= -1197050035;
assign addr[51915]= -1320917099;
assign addr[51916]= -1438083551;
assign addr[51917]= -1547955041;
assign addr[51918]= -1649974225;
assign addr[51919]= -1743623590;
assign addr[51920]= -1828428082;
assign addr[51921]= -1903957513;
assign addr[51922]= -1969828744;
assign addr[51923]= -2025707632;
assign addr[51924]= -2071310720;
assign addr[51925]= -2106406677;
assign addr[51926]= -2130817471;
assign addr[51927]= -2144419275;
assign addr[51928]= -2147143090;
assign addr[51929]= -2138975100;
assign addr[51930]= -2119956737;
assign addr[51931]= -2090184478;
assign addr[51932]= -2049809346;
assign addr[51933]= -1999036154;
assign addr[51934]= -1938122457;
assign addr[51935]= -1867377253;
assign addr[51936]= -1787159411;
assign addr[51937]= -1697875851;
assign addr[51938]= -1599979481;
assign addr[51939]= -1493966902;
assign addr[51940]= -1380375881;
assign addr[51941]= -1259782632;
assign addr[51942]= -1132798888;
assign addr[51943]= -1000068799;
assign addr[51944]= -862265664;
assign addr[51945]= -720088517;
assign addr[51946]= -574258580;
assign addr[51947]= -425515602;
assign addr[51948]= -274614114;
assign addr[51949]= -122319591;
assign addr[51950]= 30595422;
assign addr[51951]= 183355234;
assign addr[51952]= 335184940;
assign addr[51953]= 485314355;
assign addr[51954]= 632981917;
assign addr[51955]= 777438554;
assign addr[51956]= 917951481;
assign addr[51957]= 1053807919;
assign addr[51958]= 1184318708;
assign addr[51959]= 1308821808;
assign addr[51960]= 1426685652;
assign addr[51961]= 1537312353;
assign addr[51962]= 1640140734;
assign addr[51963]= 1734649179;
assign addr[51964]= 1820358275;
assign addr[51965]= 1896833245;
assign addr[51966]= 1963686155;
assign addr[51967]= 2020577882;
assign addr[51968]= 2067219829;
assign addr[51969]= 2103375398;
assign addr[51970]= 2128861181;
assign addr[51971]= 2143547897;
assign addr[51972]= 2147361045;
assign addr[51973]= 2140281282;
assign addr[51974]= 2122344521;
assign addr[51975]= 2093641749;
assign addr[51976]= 2054318569;
assign addr[51977]= 2004574453;
assign addr[51978]= 1944661739;
assign addr[51979]= 1874884346;
assign addr[51980]= 1795596234;
assign addr[51981]= 1707199606;
assign addr[51982]= 1610142873;
assign addr[51983]= 1504918373;
assign addr[51984]= 1392059879;
assign addr[51985]= 1272139887;
assign addr[51986]= 1145766716;
assign addr[51987]= 1013581418;
assign addr[51988]= 876254528;
assign addr[51989]= 734482665;
assign addr[51990]= 588984994;
assign addr[51991]= 440499581;
assign addr[51992]= 289779648;
assign addr[51993]= 137589750;
assign addr[51994]= -15298099;
assign addr[51995]= -168108346;
assign addr[51996]= -320065829;
assign addr[51997]= -470399716;
assign addr[51998]= -618347408;
assign addr[51999]= -763158411;
assign addr[52000]= -904098143;
assign addr[52001]= -1040451659;
assign addr[52002]= -1171527280;
assign addr[52003]= -1296660098;
assign addr[52004]= -1415215352;
assign addr[52005]= -1526591649;
assign addr[52006]= -1630224009;
assign addr[52007]= -1725586737;
assign addr[52008]= -1812196087;
assign addr[52009]= -1889612716;
assign addr[52010]= -1957443913;
assign addr[52011]= -2015345591;
assign addr[52012]= -2063024031;
assign addr[52013]= -2100237377;
assign addr[52014]= -2126796855;
assign addr[52015]= -2142567738;
assign addr[52016]= -2147470025;
assign addr[52017]= -2141478848;
assign addr[52018]= -2124624598;
assign addr[52019]= -2096992772;
assign addr[52020]= -2058723538;
assign addr[52021]= -2010011024;
assign addr[52022]= -1951102334;
assign addr[52023]= -1882296293;
assign addr[52024]= -1803941934;
assign addr[52025]= -1716436725;
assign addr[52026]= -1620224553;
assign addr[52027]= -1515793473;
assign addr[52028]= -1403673233;
assign addr[52029]= -1284432584;
assign addr[52030]= -1158676398;
assign addr[52031]= -1027042599;
assign addr[52032]= -890198924;
assign addr[52033]= -748839539;
assign addr[52034]= -603681519;
assign addr[52035]= -455461206;
assign addr[52036]= -304930476;
assign addr[52037]= -152852926;
assign addr[52038]= 0;
assign addr[52039]= 152852926;
assign addr[52040]= 304930476;
assign addr[52041]= 455461206;
assign addr[52042]= 603681519;
assign addr[52043]= 748839539;
assign addr[52044]= 890198924;
assign addr[52045]= 1027042599;
assign addr[52046]= 1158676398;
assign addr[52047]= 1284432584;
assign addr[52048]= 1403673233;
assign addr[52049]= 1515793473;
assign addr[52050]= 1620224553;
assign addr[52051]= 1716436725;
assign addr[52052]= 1803941934;
assign addr[52053]= 1882296293;
assign addr[52054]= 1951102334;
assign addr[52055]= 2010011024;
assign addr[52056]= 2058723538;
assign addr[52057]= 2096992772;
assign addr[52058]= 2124624598;
assign addr[52059]= 2141478848;
assign addr[52060]= 2147470025;
assign addr[52061]= 2142567738;
assign addr[52062]= 2126796855;
assign addr[52063]= 2100237377;
assign addr[52064]= 2063024031;
assign addr[52065]= 2015345591;
assign addr[52066]= 1957443913;
assign addr[52067]= 1889612716;
assign addr[52068]= 1812196087;
assign addr[52069]= 1725586737;
assign addr[52070]= 1630224009;
assign addr[52071]= 1526591649;
assign addr[52072]= 1415215352;
assign addr[52073]= 1296660098;
assign addr[52074]= 1171527280;
assign addr[52075]= 1040451659;
assign addr[52076]= 904098143;
assign addr[52077]= 763158411;
assign addr[52078]= 618347408;
assign addr[52079]= 470399716;
assign addr[52080]= 320065829;
assign addr[52081]= 168108346;
assign addr[52082]= 15298099;
assign addr[52083]= -137589750;
assign addr[52084]= -289779648;
assign addr[52085]= -440499581;
assign addr[52086]= -588984994;
assign addr[52087]= -734482665;
assign addr[52088]= -876254528;
assign addr[52089]= -1013581418;
assign addr[52090]= -1145766716;
assign addr[52091]= -1272139887;
assign addr[52092]= -1392059879;
assign addr[52093]= -1504918373;
assign addr[52094]= -1610142873;
assign addr[52095]= -1707199606;
assign addr[52096]= -1795596234;
assign addr[52097]= -1874884346;
assign addr[52098]= -1944661739;
assign addr[52099]= -2004574453;
assign addr[52100]= -2054318569;
assign addr[52101]= -2093641749;
assign addr[52102]= -2122344521;
assign addr[52103]= -2140281282;
assign addr[52104]= -2147361045;
assign addr[52105]= -2143547897;
assign addr[52106]= -2128861181;
assign addr[52107]= -2103375398;
assign addr[52108]= -2067219829;
assign addr[52109]= -2020577882;
assign addr[52110]= -1963686155;
assign addr[52111]= -1896833245;
assign addr[52112]= -1820358275;
assign addr[52113]= -1734649179;
assign addr[52114]= -1640140734;
assign addr[52115]= -1537312353;
assign addr[52116]= -1426685652;
assign addr[52117]= -1308821808;
assign addr[52118]= -1184318708;
assign addr[52119]= -1053807919;
assign addr[52120]= -917951481;
assign addr[52121]= -777438554;
assign addr[52122]= -632981917;
assign addr[52123]= -485314355;
assign addr[52124]= -335184940;
assign addr[52125]= -183355234;
assign addr[52126]= -30595422;
assign addr[52127]= 122319591;
assign addr[52128]= 274614114;
assign addr[52129]= 425515602;
assign addr[52130]= 574258580;
assign addr[52131]= 720088517;
assign addr[52132]= 862265664;
assign addr[52133]= 1000068799;
assign addr[52134]= 1132798888;
assign addr[52135]= 1259782632;
assign addr[52136]= 1380375881;
assign addr[52137]= 1493966902;
assign addr[52138]= 1599979481;
assign addr[52139]= 1697875851;
assign addr[52140]= 1787159411;
assign addr[52141]= 1867377253;
assign addr[52142]= 1938122457;
assign addr[52143]= 1999036154;
assign addr[52144]= 2049809346;
assign addr[52145]= 2090184478;
assign addr[52146]= 2119956737;
assign addr[52147]= 2138975100;
assign addr[52148]= 2147143090;
assign addr[52149]= 2144419275;
assign addr[52150]= 2130817471;
assign addr[52151]= 2106406677;
assign addr[52152]= 2071310720;
assign addr[52153]= 2025707632;
assign addr[52154]= 1969828744;
assign addr[52155]= 1903957513;
assign addr[52156]= 1828428082;
assign addr[52157]= 1743623590;
assign addr[52158]= 1649974225;
assign addr[52159]= 1547955041;
assign addr[52160]= 1438083551;
assign addr[52161]= 1320917099;
assign addr[52162]= 1197050035;
assign addr[52163]= 1067110699;
assign addr[52164]= 931758235;
assign addr[52165]= 791679244;
assign addr[52166]= 647584304;
assign addr[52167]= 500204365;
assign addr[52168]= 350287041;
assign addr[52169]= 198592817;
assign addr[52170]= 45891193;
assign addr[52171]= -107043224;
assign addr[52172]= -259434643;
assign addr[52173]= -410510029;
assign addr[52174]= -559503022;
assign addr[52175]= -705657826;
assign addr[52176]= -848233042;
assign addr[52177]= -986505429;
assign addr[52178]= -1119773573;
assign addr[52179]= -1247361445;
assign addr[52180]= -1368621831;
assign addr[52181]= -1482939614;
assign addr[52182]= -1589734894;
assign addr[52183]= -1688465931;
assign addr[52184]= -1778631892;
assign addr[52185]= -1859775393;
assign addr[52186]= -1931484818;
assign addr[52187]= -1993396407;
assign addr[52188]= -2045196100;
assign addr[52189]= -2086621133;
assign addr[52190]= -2117461370;
assign addr[52191]= -2137560369;
assign addr[52192]= -2146816171;
assign addr[52193]= -2145181827;
assign addr[52194]= -2132665626;
assign addr[52195]= -2109331059;
assign addr[52196]= -2075296495;
assign addr[52197]= -2030734582;
assign addr[52198]= -1975871368;
assign addr[52199]= -1910985158;
assign addr[52200]= -1836405100;
assign addr[52201]= -1752509516;
assign addr[52202]= -1659723983;
assign addr[52203]= -1558519173;
assign addr[52204]= -1449408469;
assign addr[52205]= -1332945355;
assign addr[52206]= -1209720613;
assign addr[52207]= -1080359326;
assign addr[52208]= -945517704;
assign addr[52209]= -805879757;
assign addr[52210]= -662153826;
assign addr[52211]= -515068990;
assign addr[52212]= -365371365;
assign addr[52213]= -213820322;
assign addr[52214]= -61184634;
assign addr[52215]= 91761426;
assign addr[52216]= 244242007;
assign addr[52217]= 395483624;
assign addr[52218]= 544719071;
assign addr[52219]= 691191324;
assign addr[52220]= 834157373;
assign addr[52221]= 972891995;
assign addr[52222]= 1106691431;
assign addr[52223]= 1234876957;
assign addr[52224]= 1356798326;
assign addr[52225]= 1471837070;
assign addr[52226]= 1579409630;
assign addr[52227]= 1678970324;
assign addr[52228]= 1770014111;
assign addr[52229]= 1852079154;
assign addr[52230]= 1924749160;
assign addr[52231]= 1987655498;
assign addr[52232]= 2040479063;
assign addr[52233]= 2082951896;
assign addr[52234]= 2114858546;
assign addr[52235]= 2136037160;
assign addr[52236]= 2146380306;
assign addr[52237]= 2145835515;
assign addr[52238]= 2134405552;
assign addr[52239]= 2112148396;
assign addr[52240]= 2079176953;
assign addr[52241]= 2035658475;
assign addr[52242]= 1981813720;
assign addr[52243]= 1917915825;
assign addr[52244]= 1844288924;
assign addr[52245]= 1761306505;
assign addr[52246]= 1669389513;
assign addr[52247]= 1569004214;
assign addr[52248]= 1460659832;
assign addr[52249]= 1344905966;
assign addr[52250]= 1222329801;
assign addr[52251]= 1093553126;
assign addr[52252]= 959229189;
assign addr[52253]= 820039373;
assign addr[52254]= 676689746;
assign addr[52255]= 529907477;
assign addr[52256]= 380437148;
assign addr[52257]= 229036977;
assign addr[52258]= 76474970;
assign addr[52259]= -76474970;
assign addr[52260]= -229036977;
assign addr[52261]= -380437148;
assign addr[52262]= -529907477;
assign addr[52263]= -676689746;
assign addr[52264]= -820039373;
assign addr[52265]= -959229189;
assign addr[52266]= -1093553126;
assign addr[52267]= -1222329801;
assign addr[52268]= -1344905966;
assign addr[52269]= -1460659832;
assign addr[52270]= -1569004214;
assign addr[52271]= -1669389513;
assign addr[52272]= -1761306505;
assign addr[52273]= -1844288924;
assign addr[52274]= -1917915825;
assign addr[52275]= -1981813720;
assign addr[52276]= -2035658475;
assign addr[52277]= -2079176953;
assign addr[52278]= -2112148396;
assign addr[52279]= -2134405552;
assign addr[52280]= -2145835515;
assign addr[52281]= -2146380306;
assign addr[52282]= -2136037160;
assign addr[52283]= -2114858546;
assign addr[52284]= -2082951896;
assign addr[52285]= -2040479063;
assign addr[52286]= -1987655498;
assign addr[52287]= -1924749160;
assign addr[52288]= -1852079154;
assign addr[52289]= -1770014111;
assign addr[52290]= -1678970324;
assign addr[52291]= -1579409630;
assign addr[52292]= -1471837070;
assign addr[52293]= -1356798326;
assign addr[52294]= -1234876957;
assign addr[52295]= -1106691431;
assign addr[52296]= -972891995;
assign addr[52297]= -834157373;
assign addr[52298]= -691191324;
assign addr[52299]= -544719071;
assign addr[52300]= -395483624;
assign addr[52301]= -244242007;
assign addr[52302]= -91761426;
assign addr[52303]= 61184634;
assign addr[52304]= 213820322;
assign addr[52305]= 365371365;
assign addr[52306]= 515068990;
assign addr[52307]= 662153826;
assign addr[52308]= 805879757;
assign addr[52309]= 945517704;
assign addr[52310]= 1080359326;
assign addr[52311]= 1209720613;
assign addr[52312]= 1332945355;
assign addr[52313]= 1449408469;
assign addr[52314]= 1558519173;
assign addr[52315]= 1659723983;
assign addr[52316]= 1752509516;
assign addr[52317]= 1836405100;
assign addr[52318]= 1910985158;
assign addr[52319]= 1975871368;
assign addr[52320]= 2030734582;
assign addr[52321]= 2075296495;
assign addr[52322]= 2109331059;
assign addr[52323]= 2132665626;
assign addr[52324]= 2145181827;
assign addr[52325]= 2146816171;
assign addr[52326]= 2137560369;
assign addr[52327]= 2117461370;
assign addr[52328]= 2086621133;
assign addr[52329]= 2045196100;
assign addr[52330]= 1993396407;
assign addr[52331]= 1931484818;
assign addr[52332]= 1859775393;
assign addr[52333]= 1778631892;
assign addr[52334]= 1688465931;
assign addr[52335]= 1589734894;
assign addr[52336]= 1482939614;
assign addr[52337]= 1368621831;
assign addr[52338]= 1247361445;
assign addr[52339]= 1119773573;
assign addr[52340]= 986505429;
assign addr[52341]= 848233042;
assign addr[52342]= 705657826;
assign addr[52343]= 559503022;
assign addr[52344]= 410510029;
assign addr[52345]= 259434643;
assign addr[52346]= 107043224;
assign addr[52347]= -45891193;
assign addr[52348]= -198592817;
assign addr[52349]= -350287041;
assign addr[52350]= -500204365;
assign addr[52351]= -647584304;
assign addr[52352]= -791679244;
assign addr[52353]= -931758235;
assign addr[52354]= -1067110699;
assign addr[52355]= -1197050035;
assign addr[52356]= -1320917099;
assign addr[52357]= -1438083551;
assign addr[52358]= -1547955041;
assign addr[52359]= -1649974225;
assign addr[52360]= -1743623590;
assign addr[52361]= -1828428082;
assign addr[52362]= -1903957513;
assign addr[52363]= -1969828744;
assign addr[52364]= -2025707632;
assign addr[52365]= -2071310720;
assign addr[52366]= -2106406677;
assign addr[52367]= -2130817471;
assign addr[52368]= -2144419275;
assign addr[52369]= -2147143090;
assign addr[52370]= -2138975100;
assign addr[52371]= -2119956737;
assign addr[52372]= -2090184478;
assign addr[52373]= -2049809346;
assign addr[52374]= -1999036154;
assign addr[52375]= -1938122457;
assign addr[52376]= -1867377253;
assign addr[52377]= -1787159411;
assign addr[52378]= -1697875851;
assign addr[52379]= -1599979481;
assign addr[52380]= -1493966902;
assign addr[52381]= -1380375881;
assign addr[52382]= -1259782632;
assign addr[52383]= -1132798888;
assign addr[52384]= -1000068799;
assign addr[52385]= -862265664;
assign addr[52386]= -720088517;
assign addr[52387]= -574258580;
assign addr[52388]= -425515602;
assign addr[52389]= -274614114;
assign addr[52390]= -122319591;
assign addr[52391]= 30595422;
assign addr[52392]= 183355234;
assign addr[52393]= 335184940;
assign addr[52394]= 485314355;
assign addr[52395]= 632981917;
assign addr[52396]= 777438554;
assign addr[52397]= 917951481;
assign addr[52398]= 1053807919;
assign addr[52399]= 1184318708;
assign addr[52400]= 1308821808;
assign addr[52401]= 1426685652;
assign addr[52402]= 1537312353;
assign addr[52403]= 1640140734;
assign addr[52404]= 1734649179;
assign addr[52405]= 1820358275;
assign addr[52406]= 1896833245;
assign addr[52407]= 1963686155;
assign addr[52408]= 2020577882;
assign addr[52409]= 2067219829;
assign addr[52410]= 2103375398;
assign addr[52411]= 2128861181;
assign addr[52412]= 2143547897;
assign addr[52413]= 2147361045;
assign addr[52414]= 2140281282;
assign addr[52415]= 2122344521;
assign addr[52416]= 2093641749;
assign addr[52417]= 2054318569;
assign addr[52418]= 2004574453;
assign addr[52419]= 1944661739;
assign addr[52420]= 1874884346;
assign addr[52421]= 1795596234;
assign addr[52422]= 1707199606;
assign addr[52423]= 1610142873;
assign addr[52424]= 1504918373;
assign addr[52425]= 1392059879;
assign addr[52426]= 1272139887;
assign addr[52427]= 1145766716;
assign addr[52428]= 1013581418;
assign addr[52429]= 876254528;
assign addr[52430]= 734482665;
assign addr[52431]= 588984994;
assign addr[52432]= 440499581;
assign addr[52433]= 289779648;
assign addr[52434]= 137589750;
assign addr[52435]= -15298099;
assign addr[52436]= -168108346;
assign addr[52437]= -320065829;
assign addr[52438]= -470399716;
assign addr[52439]= -618347408;
assign addr[52440]= -763158411;
assign addr[52441]= -904098143;
assign addr[52442]= -1040451659;
assign addr[52443]= -1171527280;
assign addr[52444]= -1296660098;
assign addr[52445]= -1415215352;
assign addr[52446]= -1526591649;
assign addr[52447]= -1630224009;
assign addr[52448]= -1725586737;
assign addr[52449]= -1812196087;
assign addr[52450]= -1889612716;
assign addr[52451]= -1957443913;
assign addr[52452]= -2015345591;
assign addr[52453]= -2063024031;
assign addr[52454]= -2100237377;
assign addr[52455]= -2126796855;
assign addr[52456]= -2142567738;
assign addr[52457]= -2147470025;
assign addr[52458]= -2141478848;
assign addr[52459]= -2124624598;
assign addr[52460]= -2096992772;
assign addr[52461]= -2058723538;
assign addr[52462]= -2010011024;
assign addr[52463]= -1951102334;
assign addr[52464]= -1882296293;
assign addr[52465]= -1803941934;
assign addr[52466]= -1716436725;
assign addr[52467]= -1620224553;
assign addr[52468]= -1515793473;
assign addr[52469]= -1403673233;
assign addr[52470]= -1284432584;
assign addr[52471]= -1158676398;
assign addr[52472]= -1027042599;
assign addr[52473]= -890198924;
assign addr[52474]= -748839539;
assign addr[52475]= -603681519;
assign addr[52476]= -455461206;
assign addr[52477]= -304930476;
assign addr[52478]= -152852926;
assign addr[52479]= 0;
assign addr[52480]= 152852926;
assign addr[52481]= 304930476;
assign addr[52482]= 455461206;
assign addr[52483]= 603681519;
assign addr[52484]= 748839539;
assign addr[52485]= 890198924;
assign addr[52486]= 1027042599;
assign addr[52487]= 1158676398;
assign addr[52488]= 1284432584;
assign addr[52489]= 1403673233;
assign addr[52490]= 1515793473;
assign addr[52491]= 1620224553;
assign addr[52492]= 1716436725;
assign addr[52493]= 1803941934;
assign addr[52494]= 1882296293;
assign addr[52495]= 1951102334;
assign addr[52496]= 2010011024;
assign addr[52497]= 2058723538;
assign addr[52498]= 2096992772;
assign addr[52499]= 2124624598;
assign addr[52500]= 2141478848;
assign addr[52501]= 2147470025;
assign addr[52502]= 2142567738;
assign addr[52503]= 2126796855;
assign addr[52504]= 2100237377;
assign addr[52505]= 2063024031;
assign addr[52506]= 2015345591;
assign addr[52507]= 1957443913;
assign addr[52508]= 1889612716;
assign addr[52509]= 1812196087;
assign addr[52510]= 1725586737;
assign addr[52511]= 1630224009;
assign addr[52512]= 1526591649;
assign addr[52513]= 1415215352;
assign addr[52514]= 1296660098;
assign addr[52515]= 1171527280;
assign addr[52516]= 1040451659;
assign addr[52517]= 904098143;
assign addr[52518]= 763158411;
assign addr[52519]= 618347408;
assign addr[52520]= 470399716;
assign addr[52521]= 320065829;
assign addr[52522]= 168108346;
assign addr[52523]= 15298099;
assign addr[52524]= -137589750;
assign addr[52525]= -289779648;
assign addr[52526]= -440499581;
assign addr[52527]= -588984994;
assign addr[52528]= -734482665;
assign addr[52529]= -876254528;
assign addr[52530]= -1013581418;
assign addr[52531]= -1145766716;
assign addr[52532]= -1272139887;
assign addr[52533]= -1392059879;
assign addr[52534]= -1504918373;
assign addr[52535]= -1610142873;
assign addr[52536]= -1707199606;
assign addr[52537]= -1795596234;
assign addr[52538]= -1874884346;
assign addr[52539]= -1944661739;
assign addr[52540]= -2004574453;
assign addr[52541]= -2054318569;
assign addr[52542]= -2093641749;
assign addr[52543]= -2122344521;
assign addr[52544]= -2140281282;
assign addr[52545]= -2147361045;
assign addr[52546]= -2143547897;
assign addr[52547]= -2128861181;
assign addr[52548]= -2103375398;
assign addr[52549]= -2067219829;
assign addr[52550]= -2020577882;
assign addr[52551]= -1963686155;
assign addr[52552]= -1896833245;
assign addr[52553]= -1820358275;
assign addr[52554]= -1734649179;
assign addr[52555]= -1640140734;
assign addr[52556]= -1537312353;
assign addr[52557]= -1426685652;
assign addr[52558]= -1308821808;
assign addr[52559]= -1184318708;
assign addr[52560]= -1053807919;
assign addr[52561]= -917951481;
assign addr[52562]= -777438554;
assign addr[52563]= -632981917;
assign addr[52564]= -485314355;
assign addr[52565]= -335184940;
assign addr[52566]= -183355234;
assign addr[52567]= -30595422;
assign addr[52568]= 122319591;
assign addr[52569]= 274614114;
assign addr[52570]= 425515602;
assign addr[52571]= 574258580;
assign addr[52572]= 720088517;
assign addr[52573]= 862265664;
assign addr[52574]= 1000068799;
assign addr[52575]= 1132798888;
assign addr[52576]= 1259782632;
assign addr[52577]= 1380375881;
assign addr[52578]= 1493966902;
assign addr[52579]= 1599979481;
assign addr[52580]= 1697875851;
assign addr[52581]= 1787159411;
assign addr[52582]= 1867377253;
assign addr[52583]= 1938122457;
assign addr[52584]= 1999036154;
assign addr[52585]= 2049809346;
assign addr[52586]= 2090184478;
assign addr[52587]= 2119956737;
assign addr[52588]= 2138975100;
assign addr[52589]= 2147143090;
assign addr[52590]= 2144419275;
assign addr[52591]= 2130817471;
assign addr[52592]= 2106406677;
assign addr[52593]= 2071310720;
assign addr[52594]= 2025707632;
assign addr[52595]= 1969828744;
assign addr[52596]= 1903957513;
assign addr[52597]= 1828428082;
assign addr[52598]= 1743623590;
assign addr[52599]= 1649974225;
assign addr[52600]= 1547955041;
assign addr[52601]= 1438083551;
assign addr[52602]= 1320917099;
assign addr[52603]= 1197050035;
assign addr[52604]= 1067110699;
assign addr[52605]= 931758235;
assign addr[52606]= 791679244;
assign addr[52607]= 647584304;
assign addr[52608]= 500204365;
assign addr[52609]= 350287041;
assign addr[52610]= 198592817;
assign addr[52611]= 45891193;
assign addr[52612]= -107043224;
assign addr[52613]= -259434643;
assign addr[52614]= -410510029;
assign addr[52615]= -559503022;
assign addr[52616]= -705657826;
assign addr[52617]= -848233042;
assign addr[52618]= -986505429;
assign addr[52619]= -1119773573;
assign addr[52620]= -1247361445;
assign addr[52621]= -1368621831;
assign addr[52622]= -1482939614;
assign addr[52623]= -1589734894;
assign addr[52624]= -1688465931;
assign addr[52625]= -1778631892;
assign addr[52626]= -1859775393;
assign addr[52627]= -1931484818;
assign addr[52628]= -1993396407;
assign addr[52629]= -2045196100;
assign addr[52630]= -2086621133;
assign addr[52631]= -2117461370;
assign addr[52632]= -2137560369;
assign addr[52633]= -2146816171;
assign addr[52634]= -2145181827;
assign addr[52635]= -2132665626;
assign addr[52636]= -2109331059;
assign addr[52637]= -2075296495;
assign addr[52638]= -2030734582;
assign addr[52639]= -1975871368;
assign addr[52640]= -1910985158;
assign addr[52641]= -1836405100;
assign addr[52642]= -1752509516;
assign addr[52643]= -1659723983;
assign addr[52644]= -1558519173;
assign addr[52645]= -1449408469;
assign addr[52646]= -1332945355;
assign addr[52647]= -1209720613;
assign addr[52648]= -1080359326;
assign addr[52649]= -945517704;
assign addr[52650]= -805879757;
assign addr[52651]= -662153826;
assign addr[52652]= -515068990;
assign addr[52653]= -365371365;
assign addr[52654]= -213820322;
assign addr[52655]= -61184634;
assign addr[52656]= 91761426;
assign addr[52657]= 244242007;
assign addr[52658]= 395483624;
assign addr[52659]= 544719071;
assign addr[52660]= 691191324;
assign addr[52661]= 834157373;
assign addr[52662]= 972891995;
assign addr[52663]= 1106691431;
assign addr[52664]= 1234876957;
assign addr[52665]= 1356798326;
assign addr[52666]= 1471837070;
assign addr[52667]= 1579409630;
assign addr[52668]= 1678970324;
assign addr[52669]= 1770014111;
assign addr[52670]= 1852079154;
assign addr[52671]= 1924749160;
assign addr[52672]= 1987655498;
assign addr[52673]= 2040479063;
assign addr[52674]= 2082951896;
assign addr[52675]= 2114858546;
assign addr[52676]= 2136037160;
assign addr[52677]= 2146380306;
assign addr[52678]= 2145835515;
assign addr[52679]= 2134405552;
assign addr[52680]= 2112148396;
assign addr[52681]= 2079176953;
assign addr[52682]= 2035658475;
assign addr[52683]= 1981813720;
assign addr[52684]= 1917915825;
assign addr[52685]= 1844288924;
assign addr[52686]= 1761306505;
assign addr[52687]= 1669389513;
assign addr[52688]= 1569004214;
assign addr[52689]= 1460659832;
assign addr[52690]= 1344905966;
assign addr[52691]= 1222329801;
assign addr[52692]= 1093553126;
assign addr[52693]= 959229189;
assign addr[52694]= 820039373;
assign addr[52695]= 676689746;
assign addr[52696]= 529907477;
assign addr[52697]= 380437148;
assign addr[52698]= 229036977;
assign addr[52699]= 76474970;
assign addr[52700]= -76474970;
assign addr[52701]= -229036977;
assign addr[52702]= -380437148;
assign addr[52703]= -529907477;
assign addr[52704]= -676689746;
assign addr[52705]= -820039373;
assign addr[52706]= -959229189;
assign addr[52707]= -1093553126;
assign addr[52708]= -1222329801;
assign addr[52709]= -1344905966;
assign addr[52710]= -1460659832;
assign addr[52711]= -1569004214;
assign addr[52712]= -1669389513;
assign addr[52713]= -1761306505;
assign addr[52714]= -1844288924;
assign addr[52715]= -1917915825;
assign addr[52716]= -1981813720;
assign addr[52717]= -2035658475;
assign addr[52718]= -2079176953;
assign addr[52719]= -2112148396;
assign addr[52720]= -2134405552;
assign addr[52721]= -2145835515;
assign addr[52722]= -2146380306;
assign addr[52723]= -2136037160;
assign addr[52724]= -2114858546;
assign addr[52725]= -2082951896;
assign addr[52726]= -2040479063;
assign addr[52727]= -1987655498;
assign addr[52728]= -1924749160;
assign addr[52729]= -1852079154;
assign addr[52730]= -1770014111;
assign addr[52731]= -1678970324;
assign addr[52732]= -1579409630;
assign addr[52733]= -1471837070;
assign addr[52734]= -1356798326;
assign addr[52735]= -1234876957;
assign addr[52736]= -1106691431;
assign addr[52737]= -972891995;
assign addr[52738]= -834157373;
assign addr[52739]= -691191324;
assign addr[52740]= -544719071;
assign addr[52741]= -395483624;
assign addr[52742]= -244242007;
assign addr[52743]= -91761426;
assign addr[52744]= 61184634;
assign addr[52745]= 213820322;
assign addr[52746]= 365371365;
assign addr[52747]= 515068990;
assign addr[52748]= 662153826;
assign addr[52749]= 805879757;
assign addr[52750]= 945517704;
assign addr[52751]= 1080359326;
assign addr[52752]= 1209720613;
assign addr[52753]= 1332945355;
assign addr[52754]= 1449408469;
assign addr[52755]= 1558519173;
assign addr[52756]= 1659723983;
assign addr[52757]= 1752509516;
assign addr[52758]= 1836405100;
assign addr[52759]= 1910985158;
assign addr[52760]= 1975871368;
assign addr[52761]= 2030734582;
assign addr[52762]= 2075296495;
assign addr[52763]= 2109331059;
assign addr[52764]= 2132665626;
assign addr[52765]= 2145181827;
assign addr[52766]= 2146816171;
assign addr[52767]= 2137560369;
assign addr[52768]= 2117461370;
assign addr[52769]= 2086621133;
assign addr[52770]= 2045196100;
assign addr[52771]= 1993396407;
assign addr[52772]= 1931484818;
assign addr[52773]= 1859775393;
assign addr[52774]= 1778631892;
assign addr[52775]= 1688465931;
assign addr[52776]= 1589734894;
assign addr[52777]= 1482939614;
assign addr[52778]= 1368621831;
assign addr[52779]= 1247361445;
assign addr[52780]= 1119773573;
assign addr[52781]= 986505429;
assign addr[52782]= 848233042;
assign addr[52783]= 705657826;
assign addr[52784]= 559503022;
assign addr[52785]= 410510029;
assign addr[52786]= 259434643;
assign addr[52787]= 107043224;
assign addr[52788]= -45891193;
assign addr[52789]= -198592817;
assign addr[52790]= -350287041;
assign addr[52791]= -500204365;
assign addr[52792]= -647584304;
assign addr[52793]= -791679244;
assign addr[52794]= -931758235;
assign addr[52795]= -1067110699;
assign addr[52796]= -1197050035;
assign addr[52797]= -1320917099;
assign addr[52798]= -1438083551;
assign addr[52799]= -1547955041;
assign addr[52800]= -1649974225;
assign addr[52801]= -1743623590;
assign addr[52802]= -1828428082;
assign addr[52803]= -1903957513;
assign addr[52804]= -1969828744;
assign addr[52805]= -2025707632;
assign addr[52806]= -2071310720;
assign addr[52807]= -2106406677;
assign addr[52808]= -2130817471;
assign addr[52809]= -2144419275;
assign addr[52810]= -2147143090;
assign addr[52811]= -2138975100;
assign addr[52812]= -2119956737;
assign addr[52813]= -2090184478;
assign addr[52814]= -2049809346;
assign addr[52815]= -1999036154;
assign addr[52816]= -1938122457;
assign addr[52817]= -1867377253;
assign addr[52818]= -1787159411;
assign addr[52819]= -1697875851;
assign addr[52820]= -1599979481;
assign addr[52821]= -1493966902;
assign addr[52822]= -1380375881;
assign addr[52823]= -1259782632;
assign addr[52824]= -1132798888;
assign addr[52825]= -1000068799;
assign addr[52826]= -862265664;
assign addr[52827]= -720088517;
assign addr[52828]= -574258580;
assign addr[52829]= -425515602;
assign addr[52830]= -274614114;
assign addr[52831]= -122319591;
assign addr[52832]= 30595422;
assign addr[52833]= 183355234;
assign addr[52834]= 335184940;
assign addr[52835]= 485314355;
assign addr[52836]= 632981917;
assign addr[52837]= 777438554;
assign addr[52838]= 917951481;
assign addr[52839]= 1053807919;
assign addr[52840]= 1184318708;
assign addr[52841]= 1308821808;
assign addr[52842]= 1426685652;
assign addr[52843]= 1537312353;
assign addr[52844]= 1640140734;
assign addr[52845]= 1734649179;
assign addr[52846]= 1820358275;
assign addr[52847]= 1896833245;
assign addr[52848]= 1963686155;
assign addr[52849]= 2020577882;
assign addr[52850]= 2067219829;
assign addr[52851]= 2103375398;
assign addr[52852]= 2128861181;
assign addr[52853]= 2143547897;
assign addr[52854]= 2147361045;
assign addr[52855]= 2140281282;
assign addr[52856]= 2122344521;
assign addr[52857]= 2093641749;
assign addr[52858]= 2054318569;
assign addr[52859]= 2004574453;
assign addr[52860]= 1944661739;
assign addr[52861]= 1874884346;
assign addr[52862]= 1795596234;
assign addr[52863]= 1707199606;
assign addr[52864]= 1610142873;
assign addr[52865]= 1504918373;
assign addr[52866]= 1392059879;
assign addr[52867]= 1272139887;
assign addr[52868]= 1145766716;
assign addr[52869]= 1013581418;
assign addr[52870]= 876254528;
assign addr[52871]= 734482665;
assign addr[52872]= 588984994;
assign addr[52873]= 440499581;
assign addr[52874]= 289779648;
assign addr[52875]= 137589750;
assign addr[52876]= -15298099;
assign addr[52877]= -168108346;
assign addr[52878]= -320065829;
assign addr[52879]= -470399716;
assign addr[52880]= -618347408;
assign addr[52881]= -763158411;
assign addr[52882]= -904098143;
assign addr[52883]= -1040451659;
assign addr[52884]= -1171527280;
assign addr[52885]= -1296660098;
assign addr[52886]= -1415215352;
assign addr[52887]= -1526591649;
assign addr[52888]= -1630224009;
assign addr[52889]= -1725586737;
assign addr[52890]= -1812196087;
assign addr[52891]= -1889612716;
assign addr[52892]= -1957443913;
assign addr[52893]= -2015345591;
assign addr[52894]= -2063024031;
assign addr[52895]= -2100237377;
assign addr[52896]= -2126796855;
assign addr[52897]= -2142567738;
assign addr[52898]= -2147470025;
assign addr[52899]= -2141478848;
assign addr[52900]= -2124624598;
assign addr[52901]= -2096992772;
assign addr[52902]= -2058723538;
assign addr[52903]= -2010011024;
assign addr[52904]= -1951102334;
assign addr[52905]= -1882296293;
assign addr[52906]= -1803941934;
assign addr[52907]= -1716436725;
assign addr[52908]= -1620224553;
assign addr[52909]= -1515793473;
assign addr[52910]= -1403673233;
assign addr[52911]= -1284432584;
assign addr[52912]= -1158676398;
assign addr[52913]= -1027042599;
assign addr[52914]= -890198924;
assign addr[52915]= -748839539;
assign addr[52916]= -603681519;
assign addr[52917]= -455461206;
assign addr[52918]= -304930476;
assign addr[52919]= -152852926;
assign addr[52920]= 0;
assign addr[52921]= 152852926;
assign addr[52922]= 304930476;
assign addr[52923]= 455461206;
assign addr[52924]= 603681519;
assign addr[52925]= 748839539;
assign addr[52926]= 890198924;
assign addr[52927]= 1027042599;
assign addr[52928]= 1158676398;
assign addr[52929]= 1284432584;
assign addr[52930]= 1403673233;
assign addr[52931]= 1515793473;
assign addr[52932]= 1620224553;
assign addr[52933]= 1716436725;
assign addr[52934]= 1803941934;
assign addr[52935]= 1882296293;
assign addr[52936]= 1951102334;
assign addr[52937]= 2010011024;
assign addr[52938]= 2058723538;
assign addr[52939]= 2096992772;
assign addr[52940]= 2124624598;
assign addr[52941]= 2141478848;
assign addr[52942]= 2147470025;
assign addr[52943]= 2142567738;
assign addr[52944]= 2126796855;
assign addr[52945]= 2100237377;
assign addr[52946]= 2063024031;
assign addr[52947]= 2015345591;
assign addr[52948]= 1957443913;
assign addr[52949]= 1889612716;
assign addr[52950]= 1812196087;
assign addr[52951]= 1725586737;
assign addr[52952]= 1630224009;
assign addr[52953]= 1526591649;
assign addr[52954]= 1415215352;
assign addr[52955]= 1296660098;
assign addr[52956]= 1171527280;
assign addr[52957]= 1040451659;
assign addr[52958]= 904098143;
assign addr[52959]= 763158411;
assign addr[52960]= 618347408;
assign addr[52961]= 470399716;
assign addr[52962]= 320065829;
assign addr[52963]= 168108346;
assign addr[52964]= 15298099;
assign addr[52965]= -137589750;
assign addr[52966]= -289779648;
assign addr[52967]= -440499581;
assign addr[52968]= -588984994;
assign addr[52969]= -734482665;
assign addr[52970]= -876254528;
assign addr[52971]= -1013581418;
assign addr[52972]= -1145766716;
assign addr[52973]= -1272139887;
assign addr[52974]= -1392059879;
assign addr[52975]= -1504918373;
assign addr[52976]= -1610142873;
assign addr[52977]= -1707199606;
assign addr[52978]= -1795596234;
assign addr[52979]= -1874884346;
assign addr[52980]= -1944661739;
assign addr[52981]= -2004574453;
assign addr[52982]= -2054318569;
assign addr[52983]= -2093641749;
assign addr[52984]= -2122344521;
assign addr[52985]= -2140281282;
assign addr[52986]= -2147361045;
assign addr[52987]= -2143547897;
assign addr[52988]= -2128861181;
assign addr[52989]= -2103375398;
assign addr[52990]= -2067219829;
assign addr[52991]= -2020577882;
assign addr[52992]= -1963686155;
assign addr[52993]= -1896833245;
assign addr[52994]= -1820358275;
assign addr[52995]= -1734649179;
assign addr[52996]= -1640140734;
assign addr[52997]= -1537312353;
assign addr[52998]= -1426685652;
assign addr[52999]= -1308821808;
assign addr[53000]= -1184318708;
assign addr[53001]= -1053807919;
assign addr[53002]= -917951481;
assign addr[53003]= -777438554;
assign addr[53004]= -632981917;
assign addr[53005]= -485314355;
assign addr[53006]= -335184940;
assign addr[53007]= -183355234;
assign addr[53008]= -30595422;
assign addr[53009]= 122319591;
assign addr[53010]= 274614114;
assign addr[53011]= 425515602;
assign addr[53012]= 574258580;
assign addr[53013]= 720088517;
assign addr[53014]= 862265664;
assign addr[53015]= 1000068799;
assign addr[53016]= 1132798888;
assign addr[53017]= 1259782632;
assign addr[53018]= 1380375881;
assign addr[53019]= 1493966902;
assign addr[53020]= 1599979481;
assign addr[53021]= 1697875851;
assign addr[53022]= 1787159411;
assign addr[53023]= 1867377253;
assign addr[53024]= 1938122457;
assign addr[53025]= 1999036154;
assign addr[53026]= 2049809346;
assign addr[53027]= 2090184478;
assign addr[53028]= 2119956737;
assign addr[53029]= 2138975100;
assign addr[53030]= 2147143090;
assign addr[53031]= 2144419275;
assign addr[53032]= 2130817471;
assign addr[53033]= 2106406677;
assign addr[53034]= 2071310720;
assign addr[53035]= 2025707632;
assign addr[53036]= 1969828744;
assign addr[53037]= 1903957513;
assign addr[53038]= 1828428082;
assign addr[53039]= 1743623590;
assign addr[53040]= 1649974225;
assign addr[53041]= 1547955041;
assign addr[53042]= 1438083551;
assign addr[53043]= 1320917099;
assign addr[53044]= 1197050035;
assign addr[53045]= 1067110699;
assign addr[53046]= 931758235;
assign addr[53047]= 791679244;
assign addr[53048]= 647584304;
assign addr[53049]= 500204365;
assign addr[53050]= 350287041;
assign addr[53051]= 198592817;
assign addr[53052]= 45891193;
assign addr[53053]= -107043224;
assign addr[53054]= -259434643;
assign addr[53055]= -410510029;
assign addr[53056]= -559503022;
assign addr[53057]= -705657826;
assign addr[53058]= -848233042;
assign addr[53059]= -986505429;
assign addr[53060]= -1119773573;
assign addr[53061]= -1247361445;
assign addr[53062]= -1368621831;
assign addr[53063]= -1482939614;
assign addr[53064]= -1589734894;
assign addr[53065]= -1688465931;
assign addr[53066]= -1778631892;
assign addr[53067]= -1859775393;
assign addr[53068]= -1931484818;
assign addr[53069]= -1993396407;
assign addr[53070]= -2045196100;
assign addr[53071]= -2086621133;
assign addr[53072]= -2117461370;
assign addr[53073]= -2137560369;
assign addr[53074]= -2146816171;
assign addr[53075]= -2145181827;
assign addr[53076]= -2132665626;
assign addr[53077]= -2109331059;
assign addr[53078]= -2075296495;
assign addr[53079]= -2030734582;
assign addr[53080]= -1975871368;
assign addr[53081]= -1910985158;
assign addr[53082]= -1836405100;
assign addr[53083]= -1752509516;
assign addr[53084]= -1659723983;
assign addr[53085]= -1558519173;
assign addr[53086]= -1449408469;
assign addr[53087]= -1332945355;
assign addr[53088]= -1209720613;
assign addr[53089]= -1080359326;
assign addr[53090]= -945517704;
assign addr[53091]= -805879757;
assign addr[53092]= -662153826;
assign addr[53093]= -515068990;
assign addr[53094]= -365371365;
assign addr[53095]= -213820322;
assign addr[53096]= -61184634;
assign addr[53097]= 91761426;
assign addr[53098]= 244242007;
assign addr[53099]= 395483624;
assign addr[53100]= 544719071;
assign addr[53101]= 691191324;
assign addr[53102]= 834157373;
assign addr[53103]= 972891995;
assign addr[53104]= 1106691431;
assign addr[53105]= 1234876957;
assign addr[53106]= 1356798326;
assign addr[53107]= 1471837070;
assign addr[53108]= 1579409630;
assign addr[53109]= 1678970324;
assign addr[53110]= 1770014111;
assign addr[53111]= 1852079154;
assign addr[53112]= 1924749160;
assign addr[53113]= 1987655498;
assign addr[53114]= 2040479063;
assign addr[53115]= 2082951896;
assign addr[53116]= 2114858546;
assign addr[53117]= 2136037160;
assign addr[53118]= 2146380306;
assign addr[53119]= 2145835515;
assign addr[53120]= 2134405552;
assign addr[53121]= 2112148396;
assign addr[53122]= 2079176953;
assign addr[53123]= 2035658475;
assign addr[53124]= 1981813720;
assign addr[53125]= 1917915825;
assign addr[53126]= 1844288924;
assign addr[53127]= 1761306505;
assign addr[53128]= 1669389513;
assign addr[53129]= 1569004214;
assign addr[53130]= 1460659832;
assign addr[53131]= 1344905966;
assign addr[53132]= 1222329801;
assign addr[53133]= 1093553126;
assign addr[53134]= 959229189;
assign addr[53135]= 820039373;
assign addr[53136]= 676689746;
assign addr[53137]= 529907477;
assign addr[53138]= 380437148;
assign addr[53139]= 229036977;
assign addr[53140]= 76474970;
assign addr[53141]= -76474970;
assign addr[53142]= -229036977;
assign addr[53143]= -380437148;
assign addr[53144]= -529907477;
assign addr[53145]= -676689746;
assign addr[53146]= -820039373;
assign addr[53147]= -959229189;
assign addr[53148]= -1093553126;
assign addr[53149]= -1222329801;
assign addr[53150]= -1344905966;
assign addr[53151]= -1460659832;
assign addr[53152]= -1569004214;
assign addr[53153]= -1669389513;
assign addr[53154]= -1761306505;
assign addr[53155]= -1844288924;
assign addr[53156]= -1917915825;
assign addr[53157]= -1981813720;
assign addr[53158]= -2035658475;
assign addr[53159]= -2079176953;
assign addr[53160]= -2112148396;
assign addr[53161]= -2134405552;
assign addr[53162]= -2145835515;
assign addr[53163]= -2146380306;
assign addr[53164]= -2136037160;
assign addr[53165]= -2114858546;
assign addr[53166]= -2082951896;
assign addr[53167]= -2040479063;
assign addr[53168]= -1987655498;
assign addr[53169]= -1924749160;
assign addr[53170]= -1852079154;
assign addr[53171]= -1770014111;
assign addr[53172]= -1678970324;
assign addr[53173]= -1579409630;
assign addr[53174]= -1471837070;
assign addr[53175]= -1356798326;
assign addr[53176]= -1234876957;
assign addr[53177]= -1106691431;
assign addr[53178]= -972891995;
assign addr[53179]= -834157373;
assign addr[53180]= -691191324;
assign addr[53181]= -544719071;
assign addr[53182]= -395483624;
assign addr[53183]= -244242007;
assign addr[53184]= -91761426;
assign addr[53185]= 61184634;
assign addr[53186]= 213820322;
assign addr[53187]= 365371365;
assign addr[53188]= 515068990;
assign addr[53189]= 662153826;
assign addr[53190]= 805879757;
assign addr[53191]= 945517704;
assign addr[53192]= 1080359326;
assign addr[53193]= 1209720613;
assign addr[53194]= 1332945355;
assign addr[53195]= 1449408469;
assign addr[53196]= 1558519173;
assign addr[53197]= 1659723983;
assign addr[53198]= 1752509516;
assign addr[53199]= 1836405100;
assign addr[53200]= 1910985158;
assign addr[53201]= 1975871368;
assign addr[53202]= 2030734582;
assign addr[53203]= 2075296495;
assign addr[53204]= 2109331059;
assign addr[53205]= 2132665626;
assign addr[53206]= 2145181827;
assign addr[53207]= 2146816171;
assign addr[53208]= 2137560369;
assign addr[53209]= 2117461370;
assign addr[53210]= 2086621133;
assign addr[53211]= 2045196100;
assign addr[53212]= 1993396407;
assign addr[53213]= 1931484818;
assign addr[53214]= 1859775393;
assign addr[53215]= 1778631892;
assign addr[53216]= 1688465931;
assign addr[53217]= 1589734894;
assign addr[53218]= 1482939614;
assign addr[53219]= 1368621831;
assign addr[53220]= 1247361445;
assign addr[53221]= 1119773573;
assign addr[53222]= 986505429;
assign addr[53223]= 848233042;
assign addr[53224]= 705657826;
assign addr[53225]= 559503022;
assign addr[53226]= 410510029;
assign addr[53227]= 259434643;
assign addr[53228]= 107043224;
assign addr[53229]= -45891193;
assign addr[53230]= -198592817;
assign addr[53231]= -350287041;
assign addr[53232]= -500204365;
assign addr[53233]= -647584304;
assign addr[53234]= -791679244;
assign addr[53235]= -931758235;
assign addr[53236]= -1067110699;
assign addr[53237]= -1197050035;
assign addr[53238]= -1320917099;
assign addr[53239]= -1438083551;
assign addr[53240]= -1547955041;
assign addr[53241]= -1649974225;
assign addr[53242]= -1743623590;
assign addr[53243]= -1828428082;
assign addr[53244]= -1903957513;
assign addr[53245]= -1969828744;
assign addr[53246]= -2025707632;
assign addr[53247]= -2071310720;
assign addr[53248]= -2106406677;
assign addr[53249]= -2130817471;
assign addr[53250]= -2144419275;
assign addr[53251]= -2147143090;
assign addr[53252]= -2138975100;
assign addr[53253]= -2119956737;
assign addr[53254]= -2090184478;
assign addr[53255]= -2049809346;
assign addr[53256]= -1999036154;
assign addr[53257]= -1938122457;
assign addr[53258]= -1867377253;
assign addr[53259]= -1787159411;
assign addr[53260]= -1697875851;
assign addr[53261]= -1599979481;
assign addr[53262]= -1493966902;
assign addr[53263]= -1380375881;
assign addr[53264]= -1259782632;
assign addr[53265]= -1132798888;
assign addr[53266]= -1000068799;
assign addr[53267]= -862265664;
assign addr[53268]= -720088517;
assign addr[53269]= -574258580;
assign addr[53270]= -425515602;
assign addr[53271]= -274614114;
assign addr[53272]= -122319591;
assign addr[53273]= 30595422;
assign addr[53274]= 183355234;
assign addr[53275]= 335184940;
assign addr[53276]= 485314355;
assign addr[53277]= 632981917;
assign addr[53278]= 777438554;
assign addr[53279]= 917951481;
assign addr[53280]= 1053807919;
assign addr[53281]= 1184318708;
assign addr[53282]= 1308821808;
assign addr[53283]= 1426685652;
assign addr[53284]= 1537312353;
assign addr[53285]= 1640140734;
assign addr[53286]= 1734649179;
assign addr[53287]= 1820358275;
assign addr[53288]= 1896833245;
assign addr[53289]= 1963686155;
assign addr[53290]= 2020577882;
assign addr[53291]= 2067219829;
assign addr[53292]= 2103375398;
assign addr[53293]= 2128861181;
assign addr[53294]= 2143547897;
assign addr[53295]= 2147361045;
assign addr[53296]= 2140281282;
assign addr[53297]= 2122344521;
assign addr[53298]= 2093641749;
assign addr[53299]= 2054318569;
assign addr[53300]= 2004574453;
assign addr[53301]= 1944661739;
assign addr[53302]= 1874884346;
assign addr[53303]= 1795596234;
assign addr[53304]= 1707199606;
assign addr[53305]= 1610142873;
assign addr[53306]= 1504918373;
assign addr[53307]= 1392059879;
assign addr[53308]= 1272139887;
assign addr[53309]= 1145766716;
assign addr[53310]= 1013581418;
assign addr[53311]= 876254528;
assign addr[53312]= 734482665;
assign addr[53313]= 588984994;
assign addr[53314]= 440499581;
assign addr[53315]= 289779648;
assign addr[53316]= 137589750;
assign addr[53317]= -15298099;
assign addr[53318]= -168108346;
assign addr[53319]= -320065829;
assign addr[53320]= -470399716;
assign addr[53321]= -618347408;
assign addr[53322]= -763158411;
assign addr[53323]= -904098143;
assign addr[53324]= -1040451659;
assign addr[53325]= -1171527280;
assign addr[53326]= -1296660098;
assign addr[53327]= -1415215352;
assign addr[53328]= -1526591649;
assign addr[53329]= -1630224009;
assign addr[53330]= -1725586737;
assign addr[53331]= -1812196087;
assign addr[53332]= -1889612716;
assign addr[53333]= -1957443913;
assign addr[53334]= -2015345591;
assign addr[53335]= -2063024031;
assign addr[53336]= -2100237377;
assign addr[53337]= -2126796855;
assign addr[53338]= -2142567738;
assign addr[53339]= -2147470025;
assign addr[53340]= -2141478848;
assign addr[53341]= -2124624598;
assign addr[53342]= -2096992772;
assign addr[53343]= -2058723538;
assign addr[53344]= -2010011024;
assign addr[53345]= -1951102334;
assign addr[53346]= -1882296293;
assign addr[53347]= -1803941934;
assign addr[53348]= -1716436725;
assign addr[53349]= -1620224553;
assign addr[53350]= -1515793473;
assign addr[53351]= -1403673233;
assign addr[53352]= -1284432584;
assign addr[53353]= -1158676398;
assign addr[53354]= -1027042599;
assign addr[53355]= -890198924;
assign addr[53356]= -748839539;
assign addr[53357]= -603681519;
assign addr[53358]= -455461206;
assign addr[53359]= -304930476;
assign addr[53360]= -152852926;
assign addr[53361]= 0;
assign addr[53362]= 152852926;
assign addr[53363]= 304930476;
assign addr[53364]= 455461206;
assign addr[53365]= 603681519;
assign addr[53366]= 748839539;
assign addr[53367]= 890198924;
assign addr[53368]= 1027042599;
assign addr[53369]= 1158676398;
assign addr[53370]= 1284432584;
assign addr[53371]= 1403673233;
assign addr[53372]= 1515793473;
assign addr[53373]= 1620224553;
assign addr[53374]= 1716436725;
assign addr[53375]= 1803941934;
assign addr[53376]= 1882296293;
assign addr[53377]= 1951102334;
assign addr[53378]= 2010011024;
assign addr[53379]= 2058723538;
assign addr[53380]= 2096992772;
assign addr[53381]= 2124624598;
assign addr[53382]= 2141478848;
assign addr[53383]= 2147470025;
assign addr[53384]= 2142567738;
assign addr[53385]= 2126796855;
assign addr[53386]= 2100237377;
assign addr[53387]= 2063024031;
assign addr[53388]= 2015345591;
assign addr[53389]= 1957443913;
assign addr[53390]= 1889612716;
assign addr[53391]= 1812196087;
assign addr[53392]= 1725586737;
assign addr[53393]= 1630224009;
assign addr[53394]= 1526591649;
assign addr[53395]= 1415215352;
assign addr[53396]= 1296660098;
assign addr[53397]= 1171527280;
assign addr[53398]= 1040451659;
assign addr[53399]= 904098143;
assign addr[53400]= 763158411;
assign addr[53401]= 618347408;
assign addr[53402]= 470399716;
assign addr[53403]= 320065829;
assign addr[53404]= 168108346;
assign addr[53405]= 15298099;
assign addr[53406]= -137589750;
assign addr[53407]= -289779648;
assign addr[53408]= -440499581;
assign addr[53409]= -588984994;
assign addr[53410]= -734482665;
assign addr[53411]= -876254528;
assign addr[53412]= -1013581418;
assign addr[53413]= -1145766716;
assign addr[53414]= -1272139887;
assign addr[53415]= -1392059879;
assign addr[53416]= -1504918373;
assign addr[53417]= -1610142873;
assign addr[53418]= -1707199606;
assign addr[53419]= -1795596234;
assign addr[53420]= -1874884346;
assign addr[53421]= -1944661739;
assign addr[53422]= -2004574453;
assign addr[53423]= -2054318569;
assign addr[53424]= -2093641749;
assign addr[53425]= -2122344521;
assign addr[53426]= -2140281282;
assign addr[53427]= -2147361045;
assign addr[53428]= -2143547897;
assign addr[53429]= -2128861181;
assign addr[53430]= -2103375398;
assign addr[53431]= -2067219829;
assign addr[53432]= -2020577882;
assign addr[53433]= -1963686155;
assign addr[53434]= -1896833245;
assign addr[53435]= -1820358275;
assign addr[53436]= -1734649179;
assign addr[53437]= -1640140734;
assign addr[53438]= -1537312353;
assign addr[53439]= -1426685652;
assign addr[53440]= -1308821808;
assign addr[53441]= -1184318708;
assign addr[53442]= -1053807919;
assign addr[53443]= -917951481;
assign addr[53444]= -777438554;
assign addr[53445]= -632981917;
assign addr[53446]= -485314355;
assign addr[53447]= -335184940;
assign addr[53448]= -183355234;
assign addr[53449]= -30595422;
assign addr[53450]= 122319591;
assign addr[53451]= 274614114;
assign addr[53452]= 425515602;
assign addr[53453]= 574258580;
assign addr[53454]= 720088517;
assign addr[53455]= 862265664;
assign addr[53456]= 1000068799;
assign addr[53457]= 1132798888;
assign addr[53458]= 1259782632;
assign addr[53459]= 1380375881;
assign addr[53460]= 1493966902;
assign addr[53461]= 1599979481;
assign addr[53462]= 1697875851;
assign addr[53463]= 1787159411;
assign addr[53464]= 1867377253;
assign addr[53465]= 1938122457;
assign addr[53466]= 1999036154;
assign addr[53467]= 2049809346;
assign addr[53468]= 2090184478;
assign addr[53469]= 2119956737;
assign addr[53470]= 2138975100;
assign addr[53471]= 2147143090;
assign addr[53472]= 2144419275;
assign addr[53473]= 2130817471;
assign addr[53474]= 2106406677;
assign addr[53475]= 2071310720;
assign addr[53476]= 2025707632;
assign addr[53477]= 1969828744;
assign addr[53478]= 1903957513;
assign addr[53479]= 1828428082;
assign addr[53480]= 1743623590;
assign addr[53481]= 1649974225;
assign addr[53482]= 1547955041;
assign addr[53483]= 1438083551;
assign addr[53484]= 1320917099;
assign addr[53485]= 1197050035;
assign addr[53486]= 1067110699;
assign addr[53487]= 931758235;
assign addr[53488]= 791679244;
assign addr[53489]= 647584304;
assign addr[53490]= 500204365;
assign addr[53491]= 350287041;
assign addr[53492]= 198592817;
assign addr[53493]= 45891193;
assign addr[53494]= -107043224;
assign addr[53495]= -259434643;
assign addr[53496]= -410510029;
assign addr[53497]= -559503022;
assign addr[53498]= -705657826;
assign addr[53499]= -848233042;
assign addr[53500]= -986505429;
assign addr[53501]= -1119773573;
assign addr[53502]= -1247361445;
assign addr[53503]= -1368621831;
assign addr[53504]= -1482939614;
assign addr[53505]= -1589734894;
assign addr[53506]= -1688465931;
assign addr[53507]= -1778631892;
assign addr[53508]= -1859775393;
assign addr[53509]= -1931484818;
assign addr[53510]= -1993396407;
assign addr[53511]= -2045196100;
assign addr[53512]= -2086621133;
assign addr[53513]= -2117461370;
assign addr[53514]= -2137560369;
assign addr[53515]= -2146816171;
assign addr[53516]= -2145181827;
assign addr[53517]= -2132665626;
assign addr[53518]= -2109331059;
assign addr[53519]= -2075296495;
assign addr[53520]= -2030734582;
assign addr[53521]= -1975871368;
assign addr[53522]= -1910985158;
assign addr[53523]= -1836405100;
assign addr[53524]= -1752509516;
assign addr[53525]= -1659723983;
assign addr[53526]= -1558519173;
assign addr[53527]= -1449408469;
assign addr[53528]= -1332945355;
assign addr[53529]= -1209720613;
assign addr[53530]= -1080359326;
assign addr[53531]= -945517704;
assign addr[53532]= -805879757;
assign addr[53533]= -662153826;
assign addr[53534]= -515068990;
assign addr[53535]= -365371365;
assign addr[53536]= -213820322;
assign addr[53537]= -61184634;
assign addr[53538]= 91761426;
assign addr[53539]= 244242007;
assign addr[53540]= 395483624;
assign addr[53541]= 544719071;
assign addr[53542]= 691191324;
assign addr[53543]= 834157373;
assign addr[53544]= 972891995;
assign addr[53545]= 1106691431;
assign addr[53546]= 1234876957;
assign addr[53547]= 1356798326;
assign addr[53548]= 1471837070;
assign addr[53549]= 1579409630;
assign addr[53550]= 1678970324;
assign addr[53551]= 1770014111;
assign addr[53552]= 1852079154;
assign addr[53553]= 1924749160;
assign addr[53554]= 1987655498;
assign addr[53555]= 2040479063;
assign addr[53556]= 2082951896;
assign addr[53557]= 2114858546;
assign addr[53558]= 2136037160;
assign addr[53559]= 2146380306;
assign addr[53560]= 2145835515;
assign addr[53561]= 2134405552;
assign addr[53562]= 2112148396;
assign addr[53563]= 2079176953;
assign addr[53564]= 2035658475;
assign addr[53565]= 1981813720;
assign addr[53566]= 1917915825;
assign addr[53567]= 1844288924;
assign addr[53568]= 1761306505;
assign addr[53569]= 1669389513;
assign addr[53570]= 1569004214;
assign addr[53571]= 1460659832;
assign addr[53572]= 1344905966;
assign addr[53573]= 1222329801;
assign addr[53574]= 1093553126;
assign addr[53575]= 959229189;
assign addr[53576]= 820039373;
assign addr[53577]= 676689746;
assign addr[53578]= 529907477;
assign addr[53579]= 380437148;
assign addr[53580]= 229036977;
assign addr[53581]= 76474970;
assign addr[53582]= -76474970;
assign addr[53583]= -229036977;
assign addr[53584]= -380437148;
assign addr[53585]= -529907477;
assign addr[53586]= -676689746;
assign addr[53587]= -820039373;
assign addr[53588]= -959229189;
assign addr[53589]= -1093553126;
assign addr[53590]= -1222329801;
assign addr[53591]= -1344905966;
assign addr[53592]= -1460659832;
assign addr[53593]= -1569004214;
assign addr[53594]= -1669389513;
assign addr[53595]= -1761306505;
assign addr[53596]= -1844288924;
assign addr[53597]= -1917915825;
assign addr[53598]= -1981813720;
assign addr[53599]= -2035658475;
assign addr[53600]= -2079176953;
assign addr[53601]= -2112148396;
assign addr[53602]= -2134405552;
assign addr[53603]= -2145835515;
assign addr[53604]= -2146380306;
assign addr[53605]= -2136037160;
assign addr[53606]= -2114858546;
assign addr[53607]= -2082951896;
assign addr[53608]= -2040479063;
assign addr[53609]= -1987655498;
assign addr[53610]= -1924749160;
assign addr[53611]= -1852079154;
assign addr[53612]= -1770014111;
assign addr[53613]= -1678970324;
assign addr[53614]= -1579409630;
assign addr[53615]= -1471837070;
assign addr[53616]= -1356798326;
assign addr[53617]= -1234876957;
assign addr[53618]= -1106691431;
assign addr[53619]= -972891995;
assign addr[53620]= -834157373;
assign addr[53621]= -691191324;
assign addr[53622]= -544719071;
assign addr[53623]= -395483624;
assign addr[53624]= -244242007;
assign addr[53625]= -91761426;
assign addr[53626]= 61184634;
assign addr[53627]= 213820322;
assign addr[53628]= 365371365;
assign addr[53629]= 515068990;
assign addr[53630]= 662153826;
assign addr[53631]= 805879757;
assign addr[53632]= 945517704;
assign addr[53633]= 1080359326;
assign addr[53634]= 1209720613;
assign addr[53635]= 1332945355;
assign addr[53636]= 1449408469;
assign addr[53637]= 1558519173;
assign addr[53638]= 1659723983;
assign addr[53639]= 1752509516;
assign addr[53640]= 1836405100;
assign addr[53641]= 1910985158;
assign addr[53642]= 1975871368;
assign addr[53643]= 2030734582;
assign addr[53644]= 2075296495;
assign addr[53645]= 2109331059;
assign addr[53646]= 2132665626;
assign addr[53647]= 2145181827;
assign addr[53648]= 2146816171;
assign addr[53649]= 2137560369;
assign addr[53650]= 2117461370;
assign addr[53651]= 2086621133;
assign addr[53652]= 2045196100;
assign addr[53653]= 1993396407;
assign addr[53654]= 1931484818;
assign addr[53655]= 1859775393;
assign addr[53656]= 1778631892;
assign addr[53657]= 1688465931;
assign addr[53658]= 1589734894;
assign addr[53659]= 1482939614;
assign addr[53660]= 1368621831;
assign addr[53661]= 1247361445;
assign addr[53662]= 1119773573;
assign addr[53663]= 986505429;
assign addr[53664]= 848233042;
assign addr[53665]= 705657826;
assign addr[53666]= 559503022;
assign addr[53667]= 410510029;
assign addr[53668]= 259434643;
assign addr[53669]= 107043224;
assign addr[53670]= -45891193;
assign addr[53671]= -198592817;
assign addr[53672]= -350287041;
assign addr[53673]= -500204365;
assign addr[53674]= -647584304;
assign addr[53675]= -791679244;
assign addr[53676]= -931758235;
assign addr[53677]= -1067110699;
assign addr[53678]= -1197050035;
assign addr[53679]= -1320917099;
assign addr[53680]= -1438083551;
assign addr[53681]= -1547955041;
assign addr[53682]= -1649974225;
assign addr[53683]= -1743623590;
assign addr[53684]= -1828428082;
assign addr[53685]= -1903957513;
assign addr[53686]= -1969828744;
assign addr[53687]= -2025707632;
assign addr[53688]= -2071310720;
assign addr[53689]= -2106406677;
assign addr[53690]= -2130817471;
assign addr[53691]= -2144419275;
assign addr[53692]= -2147143090;
assign addr[53693]= -2138975100;
assign addr[53694]= -2119956737;
assign addr[53695]= -2090184478;
assign addr[53696]= -2049809346;
assign addr[53697]= -1999036154;
assign addr[53698]= -1938122457;
assign addr[53699]= -1867377253;
assign addr[53700]= -1787159411;
assign addr[53701]= -1697875851;
assign addr[53702]= -1599979481;
assign addr[53703]= -1493966902;
assign addr[53704]= -1380375881;
assign addr[53705]= -1259782632;
assign addr[53706]= -1132798888;
assign addr[53707]= -1000068799;
assign addr[53708]= -862265664;
assign addr[53709]= -720088517;
assign addr[53710]= -574258580;
assign addr[53711]= -425515602;
assign addr[53712]= -274614114;
assign addr[53713]= -122319591;
assign addr[53714]= 30595422;
assign addr[53715]= 183355234;
assign addr[53716]= 335184940;
assign addr[53717]= 485314355;
assign addr[53718]= 632981917;
assign addr[53719]= 777438554;
assign addr[53720]= 917951481;
assign addr[53721]= 1053807919;
assign addr[53722]= 1184318708;
assign addr[53723]= 1308821808;
assign addr[53724]= 1426685652;
assign addr[53725]= 1537312353;
assign addr[53726]= 1640140734;
assign addr[53727]= 1734649179;
assign addr[53728]= 1820358275;
assign addr[53729]= 1896833245;
assign addr[53730]= 1963686155;
assign addr[53731]= 2020577882;
assign addr[53732]= 2067219829;
assign addr[53733]= 2103375398;
assign addr[53734]= 2128861181;
assign addr[53735]= 2143547897;
assign addr[53736]= 2147361045;
assign addr[53737]= 2140281282;
assign addr[53738]= 2122344521;
assign addr[53739]= 2093641749;
assign addr[53740]= 2054318569;
assign addr[53741]= 2004574453;
assign addr[53742]= 1944661739;
assign addr[53743]= 1874884346;
assign addr[53744]= 1795596234;
assign addr[53745]= 1707199606;
assign addr[53746]= 1610142873;
assign addr[53747]= 1504918373;
assign addr[53748]= 1392059879;
assign addr[53749]= 1272139887;
assign addr[53750]= 1145766716;
assign addr[53751]= 1013581418;
assign addr[53752]= 876254528;
assign addr[53753]= 734482665;
assign addr[53754]= 588984994;
assign addr[53755]= 440499581;
assign addr[53756]= 289779648;
assign addr[53757]= 137589750;
assign addr[53758]= -15298099;
assign addr[53759]= -168108346;
assign addr[53760]= -320065829;
assign addr[53761]= -470399716;
assign addr[53762]= -618347408;
assign addr[53763]= -763158411;
assign addr[53764]= -904098143;
assign addr[53765]= -1040451659;
assign addr[53766]= -1171527280;
assign addr[53767]= -1296660098;
assign addr[53768]= -1415215352;
assign addr[53769]= -1526591649;
assign addr[53770]= -1630224009;
assign addr[53771]= -1725586737;
assign addr[53772]= -1812196087;
assign addr[53773]= -1889612716;
assign addr[53774]= -1957443913;
assign addr[53775]= -2015345591;
assign addr[53776]= -2063024031;
assign addr[53777]= -2100237377;
assign addr[53778]= -2126796855;
assign addr[53779]= -2142567738;
assign addr[53780]= -2147470025;
assign addr[53781]= -2141478848;
assign addr[53782]= -2124624598;
assign addr[53783]= -2096992772;
assign addr[53784]= -2058723538;
assign addr[53785]= -2010011024;
assign addr[53786]= -1951102334;
assign addr[53787]= -1882296293;
assign addr[53788]= -1803941934;
assign addr[53789]= -1716436725;
assign addr[53790]= -1620224553;
assign addr[53791]= -1515793473;
assign addr[53792]= -1403673233;
assign addr[53793]= -1284432584;
assign addr[53794]= -1158676398;
assign addr[53795]= -1027042599;
assign addr[53796]= -890198924;
assign addr[53797]= -748839539;
assign addr[53798]= -603681519;
assign addr[53799]= -455461206;
assign addr[53800]= -304930476;
assign addr[53801]= -152852926;
assign addr[53802]= 0;
assign addr[53803]= 152852926;
assign addr[53804]= 304930476;
assign addr[53805]= 455461206;
assign addr[53806]= 603681519;
assign addr[53807]= 748839539;
assign addr[53808]= 890198924;
assign addr[53809]= 1027042599;
assign addr[53810]= 1158676398;
assign addr[53811]= 1284432584;
assign addr[53812]= 1403673233;
assign addr[53813]= 1515793473;
assign addr[53814]= 1620224553;
assign addr[53815]= 1716436725;
assign addr[53816]= 1803941934;
assign addr[53817]= 1882296293;
assign addr[53818]= 1951102334;
assign addr[53819]= 2010011024;
assign addr[53820]= 2058723538;
assign addr[53821]= 2096992772;
assign addr[53822]= 2124624598;
assign addr[53823]= 2141478848;
assign addr[53824]= 2147470025;
assign addr[53825]= 2142567738;
assign addr[53826]= 2126796855;
assign addr[53827]= 2100237377;
assign addr[53828]= 2063024031;
assign addr[53829]= 2015345591;
assign addr[53830]= 1957443913;
assign addr[53831]= 1889612716;
assign addr[53832]= 1812196087;
assign addr[53833]= 1725586737;
assign addr[53834]= 1630224009;
assign addr[53835]= 1526591649;
assign addr[53836]= 1415215352;
assign addr[53837]= 1296660098;
assign addr[53838]= 1171527280;
assign addr[53839]= 1040451659;
assign addr[53840]= 904098143;
assign addr[53841]= 763158411;
assign addr[53842]= 618347408;
assign addr[53843]= 470399716;
assign addr[53844]= 320065829;
assign addr[53845]= 168108346;
assign addr[53846]= 15298099;
assign addr[53847]= -137589750;
assign addr[53848]= -289779648;
assign addr[53849]= -440499581;
assign addr[53850]= -588984994;
assign addr[53851]= -734482665;
assign addr[53852]= -876254528;
assign addr[53853]= -1013581418;
assign addr[53854]= -1145766716;
assign addr[53855]= -1272139887;
assign addr[53856]= -1392059879;
assign addr[53857]= -1504918373;
assign addr[53858]= -1610142873;
assign addr[53859]= -1707199606;
assign addr[53860]= -1795596234;
assign addr[53861]= -1874884346;
assign addr[53862]= -1944661739;
assign addr[53863]= -2004574453;
assign addr[53864]= -2054318569;
assign addr[53865]= -2093641749;
assign addr[53866]= -2122344521;
assign addr[53867]= -2140281282;
assign addr[53868]= -2147361045;
assign addr[53869]= -2143547897;
assign addr[53870]= -2128861181;
assign addr[53871]= -2103375398;
assign addr[53872]= -2067219829;
assign addr[53873]= -2020577882;
assign addr[53874]= -1963686155;
assign addr[53875]= -1896833245;
assign addr[53876]= -1820358275;
assign addr[53877]= -1734649179;
assign addr[53878]= -1640140734;
assign addr[53879]= -1537312353;
assign addr[53880]= -1426685652;
assign addr[53881]= -1308821808;
assign addr[53882]= -1184318708;
assign addr[53883]= -1053807919;
assign addr[53884]= -917951481;
assign addr[53885]= -777438554;
assign addr[53886]= -632981917;
assign addr[53887]= -485314355;
assign addr[53888]= -335184940;
assign addr[53889]= -183355234;
assign addr[53890]= -30595422;
assign addr[53891]= 122319591;
assign addr[53892]= 274614114;
assign addr[53893]= 425515602;
assign addr[53894]= 574258580;
assign addr[53895]= 720088517;
assign addr[53896]= 862265664;
assign addr[53897]= 1000068799;
assign addr[53898]= 1132798888;
assign addr[53899]= 1259782632;
assign addr[53900]= 1380375881;
assign addr[53901]= 1493966902;
assign addr[53902]= 1599979481;
assign addr[53903]= 1697875851;
assign addr[53904]= 1787159411;
assign addr[53905]= 1867377253;
assign addr[53906]= 1938122457;
assign addr[53907]= 1999036154;
assign addr[53908]= 2049809346;
assign addr[53909]= 2090184478;
assign addr[53910]= 2119956737;
assign addr[53911]= 2138975100;
assign addr[53912]= 2147143090;
assign addr[53913]= 2144419275;
assign addr[53914]= 2130817471;
assign addr[53915]= 2106406677;
assign addr[53916]= 2071310720;
assign addr[53917]= 2025707632;
assign addr[53918]= 1969828744;
assign addr[53919]= 1903957513;
assign addr[53920]= 1828428082;
assign addr[53921]= 1743623590;
assign addr[53922]= 1649974225;
assign addr[53923]= 1547955041;
assign addr[53924]= 1438083551;
assign addr[53925]= 1320917099;
assign addr[53926]= 1197050035;
assign addr[53927]= 1067110699;
assign addr[53928]= 931758235;
assign addr[53929]= 791679244;
assign addr[53930]= 647584304;
assign addr[53931]= 500204365;
assign addr[53932]= 350287041;
assign addr[53933]= 198592817;
assign addr[53934]= 45891193;
assign addr[53935]= -107043224;
assign addr[53936]= -259434643;
assign addr[53937]= -410510029;
assign addr[53938]= -559503022;
assign addr[53939]= -705657826;
assign addr[53940]= -848233042;
assign addr[53941]= -986505429;
assign addr[53942]= -1119773573;
assign addr[53943]= -1247361445;
assign addr[53944]= -1368621831;
assign addr[53945]= -1482939614;
assign addr[53946]= -1589734894;
assign addr[53947]= -1688465931;
assign addr[53948]= -1778631892;
assign addr[53949]= -1859775393;
assign addr[53950]= -1931484818;
assign addr[53951]= -1993396407;
assign addr[53952]= -2045196100;
assign addr[53953]= -2086621133;
assign addr[53954]= -2117461370;
assign addr[53955]= -2137560369;
assign addr[53956]= -2146816171;
assign addr[53957]= -2145181827;
assign addr[53958]= -2132665626;
assign addr[53959]= -2109331059;
assign addr[53960]= -2075296495;
assign addr[53961]= -2030734582;
assign addr[53962]= -1975871368;
assign addr[53963]= -1910985158;
assign addr[53964]= -1836405100;
assign addr[53965]= -1752509516;
assign addr[53966]= -1659723983;
assign addr[53967]= -1558519173;
assign addr[53968]= -1449408469;
assign addr[53969]= -1332945355;
assign addr[53970]= -1209720613;
assign addr[53971]= -1080359326;
assign addr[53972]= -945517704;
assign addr[53973]= -805879757;
assign addr[53974]= -662153826;
assign addr[53975]= -515068990;
assign addr[53976]= -365371365;
assign addr[53977]= -213820322;
assign addr[53978]= -61184634;
assign addr[53979]= 91761426;
assign addr[53980]= 244242007;
assign addr[53981]= 395483624;
assign addr[53982]= 544719071;
assign addr[53983]= 691191324;
assign addr[53984]= 834157373;
assign addr[53985]= 972891995;
assign addr[53986]= 1106691431;
assign addr[53987]= 1234876957;
assign addr[53988]= 1356798326;
assign addr[53989]= 1471837070;
assign addr[53990]= 1579409630;
assign addr[53991]= 1678970324;
assign addr[53992]= 1770014111;
assign addr[53993]= 1852079154;
assign addr[53994]= 1924749160;
assign addr[53995]= 1987655498;
assign addr[53996]= 2040479063;
assign addr[53997]= 2082951896;
assign addr[53998]= 2114858546;
assign addr[53999]= 2136037160;
assign addr[54000]= 2146380306;
assign addr[54001]= 2145835515;
assign addr[54002]= 2134405552;
assign addr[54003]= 2112148396;
assign addr[54004]= 2079176953;
assign addr[54005]= 2035658475;
assign addr[54006]= 1981813720;
assign addr[54007]= 1917915825;
assign addr[54008]= 1844288924;
assign addr[54009]= 1761306505;
assign addr[54010]= 1669389513;
assign addr[54011]= 1569004214;
assign addr[54012]= 1460659832;
assign addr[54013]= 1344905966;
assign addr[54014]= 1222329801;
assign addr[54015]= 1093553126;
assign addr[54016]= 959229189;
assign addr[54017]= 820039373;
assign addr[54018]= 676689746;
assign addr[54019]= 529907477;
assign addr[54020]= 380437148;
assign addr[54021]= 229036977;
assign addr[54022]= 76474970;
assign addr[54023]= -76474970;
assign addr[54024]= -229036977;
assign addr[54025]= -380437148;
assign addr[54026]= -529907477;
assign addr[54027]= -676689746;
assign addr[54028]= -820039373;
assign addr[54029]= -959229189;
assign addr[54030]= -1093553126;
assign addr[54031]= -1222329801;
assign addr[54032]= -1344905966;
assign addr[54033]= -1460659832;
assign addr[54034]= -1569004214;
assign addr[54035]= -1669389513;
assign addr[54036]= -1761306505;
assign addr[54037]= -1844288924;
assign addr[54038]= -1917915825;
assign addr[54039]= -1981813720;
assign addr[54040]= -2035658475;
assign addr[54041]= -2079176953;
assign addr[54042]= -2112148396;
assign addr[54043]= -2134405552;
assign addr[54044]= -2145835515;
assign addr[54045]= -2146380306;
assign addr[54046]= -2136037160;
assign addr[54047]= -2114858546;
assign addr[54048]= -2082951896;
assign addr[54049]= -2040479063;
assign addr[54050]= -1987655498;
assign addr[54051]= -1924749160;
assign addr[54052]= -1852079154;
assign addr[54053]= -1770014111;
assign addr[54054]= -1678970324;
assign addr[54055]= -1579409630;
assign addr[54056]= -1471837070;
assign addr[54057]= -1356798326;
assign addr[54058]= -1234876957;
assign addr[54059]= -1106691431;
assign addr[54060]= -972891995;
assign addr[54061]= -834157373;
assign addr[54062]= -691191324;
assign addr[54063]= -544719071;
assign addr[54064]= -395483624;
assign addr[54065]= -244242007;
assign addr[54066]= -91761426;
assign addr[54067]= 61184634;
assign addr[54068]= 213820322;
assign addr[54069]= 365371365;
assign addr[54070]= 515068990;
assign addr[54071]= 662153826;
assign addr[54072]= 805879757;
assign addr[54073]= 945517704;
assign addr[54074]= 1080359326;
assign addr[54075]= 1209720613;
assign addr[54076]= 1332945355;
assign addr[54077]= 1449408469;
assign addr[54078]= 1558519173;
assign addr[54079]= 1659723983;
assign addr[54080]= 1752509516;
assign addr[54081]= 1836405100;
assign addr[54082]= 1910985158;
assign addr[54083]= 1975871368;
assign addr[54084]= 2030734582;
assign addr[54085]= 2075296495;
assign addr[54086]= 2109331059;
assign addr[54087]= 2132665626;
assign addr[54088]= 2145181827;
assign addr[54089]= 2146816171;
assign addr[54090]= 2137560369;
assign addr[54091]= 2117461370;
assign addr[54092]= 2086621133;
assign addr[54093]= 2045196100;
assign addr[54094]= 1993396407;
assign addr[54095]= 1931484818;
assign addr[54096]= 1859775393;
assign addr[54097]= 1778631892;
assign addr[54098]= 1688465931;
assign addr[54099]= 1589734894;
assign addr[54100]= 1482939614;
assign addr[54101]= 1368621831;
assign addr[54102]= 1247361445;
assign addr[54103]= 1119773573;
assign addr[54104]= 986505429;
assign addr[54105]= 848233042;
assign addr[54106]= 705657826;
assign addr[54107]= 559503022;
assign addr[54108]= 410510029;
assign addr[54109]= 259434643;
assign addr[54110]= 107043224;
assign addr[54111]= -45891193;
assign addr[54112]= -198592817;
assign addr[54113]= -350287041;
assign addr[54114]= -500204365;
assign addr[54115]= -647584304;
assign addr[54116]= -791679244;
assign addr[54117]= -931758235;
assign addr[54118]= -1067110699;
assign addr[54119]= -1197050035;
assign addr[54120]= -1320917099;
assign addr[54121]= -1438083551;
assign addr[54122]= -1547955041;
assign addr[54123]= -1649974225;
assign addr[54124]= -1743623590;
assign addr[54125]= -1828428082;
assign addr[54126]= -1903957513;
assign addr[54127]= -1969828744;
assign addr[54128]= -2025707632;
assign addr[54129]= -2071310720;
assign addr[54130]= -2106406677;
assign addr[54131]= -2130817471;
assign addr[54132]= -2144419275;
assign addr[54133]= -2147143090;
assign addr[54134]= -2138975100;
assign addr[54135]= -2119956737;
assign addr[54136]= -2090184478;
assign addr[54137]= -2049809346;
assign addr[54138]= -1999036154;
assign addr[54139]= -1938122457;
assign addr[54140]= -1867377253;
assign addr[54141]= -1787159411;
assign addr[54142]= -1697875851;
assign addr[54143]= -1599979481;
assign addr[54144]= -1493966902;
assign addr[54145]= -1380375881;
assign addr[54146]= -1259782632;
assign addr[54147]= -1132798888;
assign addr[54148]= -1000068799;
assign addr[54149]= -862265664;
assign addr[54150]= -720088517;
assign addr[54151]= -574258580;
assign addr[54152]= -425515602;
assign addr[54153]= -274614114;
assign addr[54154]= -122319591;
assign addr[54155]= 30595422;
assign addr[54156]= 183355234;
assign addr[54157]= 335184940;
assign addr[54158]= 485314355;
assign addr[54159]= 632981917;
assign addr[54160]= 777438554;
assign addr[54161]= 917951481;
assign addr[54162]= 1053807919;
assign addr[54163]= 1184318708;
assign addr[54164]= 1308821808;
assign addr[54165]= 1426685652;
assign addr[54166]= 1537312353;
assign addr[54167]= 1640140734;
assign addr[54168]= 1734649179;
assign addr[54169]= 1820358275;
assign addr[54170]= 1896833245;
assign addr[54171]= 1963686155;
assign addr[54172]= 2020577882;
assign addr[54173]= 2067219829;
assign addr[54174]= 2103375398;
assign addr[54175]= 2128861181;
assign addr[54176]= 2143547897;
assign addr[54177]= 2147361045;
assign addr[54178]= 2140281282;
assign addr[54179]= 2122344521;
assign addr[54180]= 2093641749;
assign addr[54181]= 2054318569;
assign addr[54182]= 2004574453;
assign addr[54183]= 1944661739;
assign addr[54184]= 1874884346;
assign addr[54185]= 1795596234;
assign addr[54186]= 1707199606;
assign addr[54187]= 1610142873;
assign addr[54188]= 1504918373;
assign addr[54189]= 1392059879;
assign addr[54190]= 1272139887;
assign addr[54191]= 1145766716;
assign addr[54192]= 1013581418;
assign addr[54193]= 876254528;
assign addr[54194]= 734482665;
assign addr[54195]= 588984994;
assign addr[54196]= 440499581;
assign addr[54197]= 289779648;
assign addr[54198]= 137589750;
assign addr[54199]= -15298099;
assign addr[54200]= -168108346;
assign addr[54201]= -320065829;
assign addr[54202]= -470399716;
assign addr[54203]= -618347408;
assign addr[54204]= -763158411;
assign addr[54205]= -904098143;
assign addr[54206]= -1040451659;
assign addr[54207]= -1171527280;
assign addr[54208]= -1296660098;
assign addr[54209]= -1415215352;
assign addr[54210]= -1526591649;
assign addr[54211]= -1630224009;
assign addr[54212]= -1725586737;
assign addr[54213]= -1812196087;
assign addr[54214]= -1889612716;
assign addr[54215]= -1957443913;
assign addr[54216]= -2015345591;
assign addr[54217]= -2063024031;
assign addr[54218]= -2100237377;
assign addr[54219]= -2126796855;
assign addr[54220]= -2142567738;
assign addr[54221]= -2147470025;
assign addr[54222]= -2141478848;
assign addr[54223]= -2124624598;
assign addr[54224]= -2096992772;
assign addr[54225]= -2058723538;
assign addr[54226]= -2010011024;
assign addr[54227]= -1951102334;
assign addr[54228]= -1882296293;
assign addr[54229]= -1803941934;
assign addr[54230]= -1716436725;
assign addr[54231]= -1620224553;
assign addr[54232]= -1515793473;
assign addr[54233]= -1403673233;
assign addr[54234]= -1284432584;
assign addr[54235]= -1158676398;
assign addr[54236]= -1027042599;
assign addr[54237]= -890198924;
assign addr[54238]= -748839539;
assign addr[54239]= -603681519;
assign addr[54240]= -455461206;
assign addr[54241]= -304930476;
assign addr[54242]= -152852926;
assign addr[54243]= 0;
assign addr[54244]= 152852926;
assign addr[54245]= 304930476;
assign addr[54246]= 455461206;
assign addr[54247]= 603681519;
assign addr[54248]= 748839539;
assign addr[54249]= 890198924;
assign addr[54250]= 1027042599;
assign addr[54251]= 1158676398;
assign addr[54252]= 1284432584;
assign addr[54253]= 1403673233;
assign addr[54254]= 1515793473;
assign addr[54255]= 1620224553;
assign addr[54256]= 1716436725;
assign addr[54257]= 1803941934;
assign addr[54258]= 1882296293;
assign addr[54259]= 1951102334;
assign addr[54260]= 2010011024;
assign addr[54261]= 2058723538;
assign addr[54262]= 2096992772;
assign addr[54263]= 2124624598;
assign addr[54264]= 2141478848;
assign addr[54265]= 2147470025;
assign addr[54266]= 2142567738;
assign addr[54267]= 2126796855;
assign addr[54268]= 2100237377;
assign addr[54269]= 2063024031;
assign addr[54270]= 2015345591;
assign addr[54271]= 1957443913;
assign addr[54272]= 1889612716;
assign addr[54273]= 1812196087;
assign addr[54274]= 1725586737;
assign addr[54275]= 1630224009;
assign addr[54276]= 1526591649;
assign addr[54277]= 1415215352;
assign addr[54278]= 1296660098;
assign addr[54279]= 1171527280;
assign addr[54280]= 1040451659;
assign addr[54281]= 904098143;
assign addr[54282]= 763158411;
assign addr[54283]= 618347408;
assign addr[54284]= 470399716;
assign addr[54285]= 320065829;
assign addr[54286]= 168108346;
assign addr[54287]= 15298099;
assign addr[54288]= -137589750;
assign addr[54289]= -289779648;
assign addr[54290]= -440499581;
assign addr[54291]= -588984994;
assign addr[54292]= -734482665;
assign addr[54293]= -876254528;
assign addr[54294]= -1013581418;
assign addr[54295]= -1145766716;
assign addr[54296]= -1272139887;
assign addr[54297]= -1392059879;
assign addr[54298]= -1504918373;
assign addr[54299]= -1610142873;
assign addr[54300]= -1707199606;
assign addr[54301]= -1795596234;
assign addr[54302]= -1874884346;
assign addr[54303]= -1944661739;
assign addr[54304]= -2004574453;
assign addr[54305]= -2054318569;
assign addr[54306]= -2093641749;
assign addr[54307]= -2122344521;
assign addr[54308]= -2140281282;
assign addr[54309]= -2147361045;
assign addr[54310]= -2143547897;
assign addr[54311]= -2128861181;
assign addr[54312]= -2103375398;
assign addr[54313]= -2067219829;
assign addr[54314]= -2020577882;
assign addr[54315]= -1963686155;
assign addr[54316]= -1896833245;
assign addr[54317]= -1820358275;
assign addr[54318]= -1734649179;
assign addr[54319]= -1640140734;
assign addr[54320]= -1537312353;
assign addr[54321]= -1426685652;
assign addr[54322]= -1308821808;
assign addr[54323]= -1184318708;
assign addr[54324]= -1053807919;
assign addr[54325]= -917951481;
assign addr[54326]= -777438554;
assign addr[54327]= -632981917;
assign addr[54328]= -485314355;
assign addr[54329]= -335184940;
assign addr[54330]= -183355234;
assign addr[54331]= -30595422;
assign addr[54332]= 122319591;
assign addr[54333]= 274614114;
assign addr[54334]= 425515602;
assign addr[54335]= 574258580;
assign addr[54336]= 720088517;
assign addr[54337]= 862265664;
assign addr[54338]= 1000068799;
assign addr[54339]= 1132798888;
assign addr[54340]= 1259782632;
assign addr[54341]= 1380375881;
assign addr[54342]= 1493966902;
assign addr[54343]= 1599979481;
assign addr[54344]= 1697875851;
assign addr[54345]= 1787159411;
assign addr[54346]= 1867377253;
assign addr[54347]= 1938122457;
assign addr[54348]= 1999036154;
assign addr[54349]= 2049809346;
assign addr[54350]= 2090184478;
assign addr[54351]= 2119956737;
assign addr[54352]= 2138975100;
assign addr[54353]= 2147143090;
assign addr[54354]= 2144419275;
assign addr[54355]= 2130817471;
assign addr[54356]= 2106406677;
assign addr[54357]= 2071310720;
assign addr[54358]= 2025707632;
assign addr[54359]= 1969828744;
assign addr[54360]= 1903957513;
assign addr[54361]= 1828428082;
assign addr[54362]= 1743623590;
assign addr[54363]= 1649974225;
assign addr[54364]= 1547955041;
assign addr[54365]= 1438083551;
assign addr[54366]= 1320917099;
assign addr[54367]= 1197050035;
assign addr[54368]= 1067110699;
assign addr[54369]= 931758235;
assign addr[54370]= 791679244;
assign addr[54371]= 647584304;
assign addr[54372]= 500204365;
assign addr[54373]= 350287041;
assign addr[54374]= 198592817;
assign addr[54375]= 45891193;
assign addr[54376]= -107043224;
assign addr[54377]= -259434643;
assign addr[54378]= -410510029;
assign addr[54379]= -559503022;
assign addr[54380]= -705657826;
assign addr[54381]= -848233042;
assign addr[54382]= -986505429;
assign addr[54383]= -1119773573;
assign addr[54384]= -1247361445;
assign addr[54385]= -1368621831;
assign addr[54386]= -1482939614;
assign addr[54387]= -1589734894;
assign addr[54388]= -1688465931;
assign addr[54389]= -1778631892;
assign addr[54390]= -1859775393;
assign addr[54391]= -1931484818;
assign addr[54392]= -1993396407;
assign addr[54393]= -2045196100;
assign addr[54394]= -2086621133;
assign addr[54395]= -2117461370;
assign addr[54396]= -2137560369;
assign addr[54397]= -2146816171;
assign addr[54398]= -2145181827;
assign addr[54399]= -2132665626;
assign addr[54400]= -2109331059;
assign addr[54401]= -2075296495;
assign addr[54402]= -2030734582;
assign addr[54403]= -1975871368;
assign addr[54404]= -1910985158;
assign addr[54405]= -1836405100;
assign addr[54406]= -1752509516;
assign addr[54407]= -1659723983;
assign addr[54408]= -1558519173;
assign addr[54409]= -1449408469;
assign addr[54410]= -1332945355;
assign addr[54411]= -1209720613;
assign addr[54412]= -1080359326;
assign addr[54413]= -945517704;
assign addr[54414]= -805879757;
assign addr[54415]= -662153826;
assign addr[54416]= -515068990;
assign addr[54417]= -365371365;
assign addr[54418]= -213820322;
assign addr[54419]= -61184634;
assign addr[54420]= 91761426;
assign addr[54421]= 244242007;
assign addr[54422]= 395483624;
assign addr[54423]= 544719071;
assign addr[54424]= 691191324;
assign addr[54425]= 834157373;
assign addr[54426]= 972891995;
assign addr[54427]= 1106691431;
assign addr[54428]= 1234876957;
assign addr[54429]= 1356798326;
assign addr[54430]= 1471837070;
assign addr[54431]= 1579409630;
assign addr[54432]= 1678970324;
assign addr[54433]= 1770014111;
assign addr[54434]= 1852079154;
assign addr[54435]= 1924749160;
assign addr[54436]= 1987655498;
assign addr[54437]= 2040479063;
assign addr[54438]= 2082951896;
assign addr[54439]= 2114858546;
assign addr[54440]= 2136037160;
assign addr[54441]= 2146380306;
assign addr[54442]= 2145835515;
assign addr[54443]= 2134405552;
assign addr[54444]= 2112148396;
assign addr[54445]= 2079176953;
assign addr[54446]= 2035658475;
assign addr[54447]= 1981813720;
assign addr[54448]= 1917915825;
assign addr[54449]= 1844288924;
assign addr[54450]= 1761306505;
assign addr[54451]= 1669389513;
assign addr[54452]= 1569004214;
assign addr[54453]= 1460659832;
assign addr[54454]= 1344905966;
assign addr[54455]= 1222329801;
assign addr[54456]= 1093553126;
assign addr[54457]= 959229189;
assign addr[54458]= 820039373;
assign addr[54459]= 676689746;
assign addr[54460]= 529907477;
assign addr[54461]= 380437148;
assign addr[54462]= 229036977;
assign addr[54463]= 76474970;
assign addr[54464]= -76474970;
assign addr[54465]= -229036977;
assign addr[54466]= -380437148;
assign addr[54467]= -529907477;
assign addr[54468]= -676689746;
assign addr[54469]= -820039373;
assign addr[54470]= -959229189;
assign addr[54471]= -1093553126;
assign addr[54472]= -1222329801;
assign addr[54473]= -1344905966;
assign addr[54474]= -1460659832;
assign addr[54475]= -1569004214;
assign addr[54476]= -1669389513;
assign addr[54477]= -1761306505;
assign addr[54478]= -1844288924;
assign addr[54479]= -1917915825;
assign addr[54480]= -1981813720;
assign addr[54481]= -2035658475;
assign addr[54482]= -2079176953;
assign addr[54483]= -2112148396;
assign addr[54484]= -2134405552;
assign addr[54485]= -2145835515;
assign addr[54486]= -2146380306;
assign addr[54487]= -2136037160;
assign addr[54488]= -2114858546;
assign addr[54489]= -2082951896;
assign addr[54490]= -2040479063;
assign addr[54491]= -1987655498;
assign addr[54492]= -1924749160;
assign addr[54493]= -1852079154;
assign addr[54494]= -1770014111;
assign addr[54495]= -1678970324;
assign addr[54496]= -1579409630;
assign addr[54497]= -1471837070;
assign addr[54498]= -1356798326;
assign addr[54499]= -1234876957;
assign addr[54500]= -1106691431;
assign addr[54501]= -972891995;
assign addr[54502]= -834157373;
assign addr[54503]= -691191324;
assign addr[54504]= -544719071;
assign addr[54505]= -395483624;
assign addr[54506]= -244242007;
assign addr[54507]= -91761426;
assign addr[54508]= 61184634;
assign addr[54509]= 213820322;
assign addr[54510]= 365371365;
assign addr[54511]= 515068990;
assign addr[54512]= 662153826;
assign addr[54513]= 805879757;
assign addr[54514]= 945517704;
assign addr[54515]= 1080359326;
assign addr[54516]= 1209720613;
assign addr[54517]= 1332945355;
assign addr[54518]= 1449408469;
assign addr[54519]= 1558519173;
assign addr[54520]= 1659723983;
assign addr[54521]= 1752509516;
assign addr[54522]= 1836405100;
assign addr[54523]= 1910985158;
assign addr[54524]= 1975871368;
assign addr[54525]= 2030734582;
assign addr[54526]= 2075296495;
assign addr[54527]= 2109331059;
assign addr[54528]= 2132665626;
assign addr[54529]= 2145181827;
assign addr[54530]= 2146816171;
assign addr[54531]= 2137560369;
assign addr[54532]= 2117461370;
assign addr[54533]= 2086621133;
assign addr[54534]= 2045196100;
assign addr[54535]= 1993396407;
assign addr[54536]= 1931484818;
assign addr[54537]= 1859775393;
assign addr[54538]= 1778631892;
assign addr[54539]= 1688465931;
assign addr[54540]= 1589734894;
assign addr[54541]= 1482939614;
assign addr[54542]= 1368621831;
assign addr[54543]= 1247361445;
assign addr[54544]= 1119773573;
assign addr[54545]= 986505429;
assign addr[54546]= 848233042;
assign addr[54547]= 705657826;
assign addr[54548]= 559503022;
assign addr[54549]= 410510029;
assign addr[54550]= 259434643;
assign addr[54551]= 107043224;
assign addr[54552]= -45891193;
assign addr[54553]= -198592817;
assign addr[54554]= -350287041;
assign addr[54555]= -500204365;
assign addr[54556]= -647584304;
assign addr[54557]= -791679244;
assign addr[54558]= -931758235;
assign addr[54559]= -1067110699;
assign addr[54560]= -1197050035;
assign addr[54561]= -1320917099;
assign addr[54562]= -1438083551;
assign addr[54563]= -1547955041;
assign addr[54564]= -1649974225;
assign addr[54565]= -1743623590;
assign addr[54566]= -1828428082;
assign addr[54567]= -1903957513;
assign addr[54568]= -1969828744;
assign addr[54569]= -2025707632;
assign addr[54570]= -2071310720;
assign addr[54571]= -2106406677;
assign addr[54572]= -2130817471;
assign addr[54573]= -2144419275;
assign addr[54574]= -2147143090;
assign addr[54575]= -2138975100;
assign addr[54576]= -2119956737;
assign addr[54577]= -2090184478;
assign addr[54578]= -2049809346;
assign addr[54579]= -1999036154;
assign addr[54580]= -1938122457;
assign addr[54581]= -1867377253;
assign addr[54582]= -1787159411;
assign addr[54583]= -1697875851;
assign addr[54584]= -1599979481;
assign addr[54585]= -1493966902;
assign addr[54586]= -1380375881;
assign addr[54587]= -1259782632;
assign addr[54588]= -1132798888;
assign addr[54589]= -1000068799;
assign addr[54590]= -862265664;
assign addr[54591]= -720088517;
assign addr[54592]= -574258580;
assign addr[54593]= -425515602;
assign addr[54594]= -274614114;
assign addr[54595]= -122319591;
assign addr[54596]= 30595422;
assign addr[54597]= 183355234;
assign addr[54598]= 335184940;
assign addr[54599]= 485314355;
assign addr[54600]= 632981917;
assign addr[54601]= 777438554;
assign addr[54602]= 917951481;
assign addr[54603]= 1053807919;
assign addr[54604]= 1184318708;
assign addr[54605]= 1308821808;
assign addr[54606]= 1426685652;
assign addr[54607]= 1537312353;
assign addr[54608]= 1640140734;
assign addr[54609]= 1734649179;
assign addr[54610]= 1820358275;
assign addr[54611]= 1896833245;
assign addr[54612]= 1963686155;
assign addr[54613]= 2020577882;
assign addr[54614]= 2067219829;
assign addr[54615]= 2103375398;
assign addr[54616]= 2128861181;
assign addr[54617]= 2143547897;
assign addr[54618]= 2147361045;
assign addr[54619]= 2140281282;
assign addr[54620]= 2122344521;
assign addr[54621]= 2093641749;
assign addr[54622]= 2054318569;
assign addr[54623]= 2004574453;
assign addr[54624]= 1944661739;
assign addr[54625]= 1874884346;
assign addr[54626]= 1795596234;
assign addr[54627]= 1707199606;
assign addr[54628]= 1610142873;
assign addr[54629]= 1504918373;
assign addr[54630]= 1392059879;
assign addr[54631]= 1272139887;
assign addr[54632]= 1145766716;
assign addr[54633]= 1013581418;
assign addr[54634]= 876254528;
assign addr[54635]= 734482665;
assign addr[54636]= 588984994;
assign addr[54637]= 440499581;
assign addr[54638]= 289779648;
assign addr[54639]= 137589750;
assign addr[54640]= -15298099;
assign addr[54641]= -168108346;
assign addr[54642]= -320065829;
assign addr[54643]= -470399716;
assign addr[54644]= -618347408;
assign addr[54645]= -763158411;
assign addr[54646]= -904098143;
assign addr[54647]= -1040451659;
assign addr[54648]= -1171527280;
assign addr[54649]= -1296660098;
assign addr[54650]= -1415215352;
assign addr[54651]= -1526591649;
assign addr[54652]= -1630224009;
assign addr[54653]= -1725586737;
assign addr[54654]= -1812196087;
assign addr[54655]= -1889612716;
assign addr[54656]= -1957443913;
assign addr[54657]= -2015345591;
assign addr[54658]= -2063024031;
assign addr[54659]= -2100237377;
assign addr[54660]= -2126796855;
assign addr[54661]= -2142567738;
assign addr[54662]= -2147470025;
assign addr[54663]= -2141478848;
assign addr[54664]= -2124624598;
assign addr[54665]= -2096992772;
assign addr[54666]= -2058723538;
assign addr[54667]= -2010011024;
assign addr[54668]= -1951102334;
assign addr[54669]= -1882296293;
assign addr[54670]= -1803941934;
assign addr[54671]= -1716436725;
assign addr[54672]= -1620224553;
assign addr[54673]= -1515793473;
assign addr[54674]= -1403673233;
assign addr[54675]= -1284432584;
assign addr[54676]= -1158676398;
assign addr[54677]= -1027042599;
assign addr[54678]= -890198924;
assign addr[54679]= -748839539;
assign addr[54680]= -603681519;
assign addr[54681]= -455461206;
assign addr[54682]= -304930476;
assign addr[54683]= -152852926;
assign addr[54684]= 0;
assign addr[54685]= 152852926;
assign addr[54686]= 304930476;
assign addr[54687]= 455461206;
assign addr[54688]= 603681519;
assign addr[54689]= 748839539;
assign addr[54690]= 890198924;
assign addr[54691]= 1027042599;
assign addr[54692]= 1158676398;
assign addr[54693]= 1284432584;
assign addr[54694]= 1403673233;
assign addr[54695]= 1515793473;
assign addr[54696]= 1620224553;
assign addr[54697]= 1716436725;
assign addr[54698]= 1803941934;
assign addr[54699]= 1882296293;
assign addr[54700]= 1951102334;
assign addr[54701]= 2010011024;
assign addr[54702]= 2058723538;
assign addr[54703]= 2096992772;
assign addr[54704]= 2124624598;
assign addr[54705]= 2141478848;
assign addr[54706]= 2147470025;
assign addr[54707]= 2142567738;
assign addr[54708]= 2126796855;
assign addr[54709]= 2100237377;
assign addr[54710]= 2063024031;
assign addr[54711]= 2015345591;
assign addr[54712]= 1957443913;
assign addr[54713]= 1889612716;
assign addr[54714]= 1812196087;
assign addr[54715]= 1725586737;
assign addr[54716]= 1630224009;
assign addr[54717]= 1526591649;
assign addr[54718]= 1415215352;
assign addr[54719]= 1296660098;
assign addr[54720]= 1171527280;
assign addr[54721]= 1040451659;
assign addr[54722]= 904098143;
assign addr[54723]= 763158411;
assign addr[54724]= 618347408;
assign addr[54725]= 470399716;
assign addr[54726]= 320065829;
assign addr[54727]= 168108346;
assign addr[54728]= 15298099;
assign addr[54729]= -137589750;
assign addr[54730]= -289779648;
assign addr[54731]= -440499581;
assign addr[54732]= -588984994;
assign addr[54733]= -734482665;
assign addr[54734]= -876254528;
assign addr[54735]= -1013581418;
assign addr[54736]= -1145766716;
assign addr[54737]= -1272139887;
assign addr[54738]= -1392059879;
assign addr[54739]= -1504918373;
assign addr[54740]= -1610142873;
assign addr[54741]= -1707199606;
assign addr[54742]= -1795596234;
assign addr[54743]= -1874884346;
assign addr[54744]= -1944661739;
assign addr[54745]= -2004574453;
assign addr[54746]= -2054318569;
assign addr[54747]= -2093641749;
assign addr[54748]= -2122344521;
assign addr[54749]= -2140281282;
assign addr[54750]= -2147361045;
assign addr[54751]= -2143547897;
assign addr[54752]= -2128861181;
assign addr[54753]= -2103375398;
assign addr[54754]= -2067219829;
assign addr[54755]= -2020577882;
assign addr[54756]= -1963686155;
assign addr[54757]= -1896833245;
assign addr[54758]= -1820358275;
assign addr[54759]= -1734649179;
assign addr[54760]= -1640140734;
assign addr[54761]= -1537312353;
assign addr[54762]= -1426685652;
assign addr[54763]= -1308821808;
assign addr[54764]= -1184318708;
assign addr[54765]= -1053807919;
assign addr[54766]= -917951481;
assign addr[54767]= -777438554;
assign addr[54768]= -632981917;
assign addr[54769]= -485314355;
assign addr[54770]= -335184940;
assign addr[54771]= -183355234;
assign addr[54772]= -30595422;
assign addr[54773]= 122319591;
assign addr[54774]= 274614114;
assign addr[54775]= 425515602;
assign addr[54776]= 574258580;
assign addr[54777]= 720088517;
assign addr[54778]= 862265664;
assign addr[54779]= 1000068799;
assign addr[54780]= 1132798888;
assign addr[54781]= 1259782632;
assign addr[54782]= 1380375881;
assign addr[54783]= 1493966902;
assign addr[54784]= 1599979481;
assign addr[54785]= 1697875851;
assign addr[54786]= 1787159411;
assign addr[54787]= 1867377253;
assign addr[54788]= 1938122457;
assign addr[54789]= 1999036154;
assign addr[54790]= 2049809346;
assign addr[54791]= 2090184478;
assign addr[54792]= 2119956737;
assign addr[54793]= 2138975100;
assign addr[54794]= 2147143090;
assign addr[54795]= 2144419275;
assign addr[54796]= 2130817471;
assign addr[54797]= 2106406677;
assign addr[54798]= 2071310720;
assign addr[54799]= 2025707632;
assign addr[54800]= 1969828744;
assign addr[54801]= 1903957513;
assign addr[54802]= 1828428082;
assign addr[54803]= 1743623590;
assign addr[54804]= 1649974225;
assign addr[54805]= 1547955041;
assign addr[54806]= 1438083551;
assign addr[54807]= 1320917099;
assign addr[54808]= 1197050035;
assign addr[54809]= 1067110699;
assign addr[54810]= 931758235;
assign addr[54811]= 791679244;
assign addr[54812]= 647584304;
assign addr[54813]= 500204365;
assign addr[54814]= 350287041;
assign addr[54815]= 198592817;
assign addr[54816]= 45891193;
assign addr[54817]= -107043224;
assign addr[54818]= -259434643;
assign addr[54819]= -410510029;
assign addr[54820]= -559503022;
assign addr[54821]= -705657826;
assign addr[54822]= -848233042;
assign addr[54823]= -986505429;
assign addr[54824]= -1119773573;
assign addr[54825]= -1247361445;
assign addr[54826]= -1368621831;
assign addr[54827]= -1482939614;
assign addr[54828]= -1589734894;
assign addr[54829]= -1688465931;
assign addr[54830]= -1778631892;
assign addr[54831]= -1859775393;
assign addr[54832]= -1931484818;
assign addr[54833]= -1993396407;
assign addr[54834]= -2045196100;
assign addr[54835]= -2086621133;
assign addr[54836]= -2117461370;
assign addr[54837]= -2137560369;
assign addr[54838]= -2146816171;
assign addr[54839]= -2145181827;
assign addr[54840]= -2132665626;
assign addr[54841]= -2109331059;
assign addr[54842]= -2075296495;
assign addr[54843]= -2030734582;
assign addr[54844]= -1975871368;
assign addr[54845]= -1910985158;
assign addr[54846]= -1836405100;
assign addr[54847]= -1752509516;
assign addr[54848]= -1659723983;
assign addr[54849]= -1558519173;
assign addr[54850]= -1449408469;
assign addr[54851]= -1332945355;
assign addr[54852]= -1209720613;
assign addr[54853]= -1080359326;
assign addr[54854]= -945517704;
assign addr[54855]= -805879757;
assign addr[54856]= -662153826;
assign addr[54857]= -515068990;
assign addr[54858]= -365371365;
assign addr[54859]= -213820322;
assign addr[54860]= -61184634;
assign addr[54861]= 91761426;
assign addr[54862]= 244242007;
assign addr[54863]= 395483624;
assign addr[54864]= 544719071;
assign addr[54865]= 691191324;
assign addr[54866]= 834157373;
assign addr[54867]= 972891995;
assign addr[54868]= 1106691431;
assign addr[54869]= 1234876957;
assign addr[54870]= 1356798326;
assign addr[54871]= 1471837070;
assign addr[54872]= 1579409630;
assign addr[54873]= 1678970324;
assign addr[54874]= 1770014111;
assign addr[54875]= 1852079154;
assign addr[54876]= 1924749160;
assign addr[54877]= 1987655498;
assign addr[54878]= 2040479063;
assign addr[54879]= 2082951896;
assign addr[54880]= 2114858546;
assign addr[54881]= 2136037160;
assign addr[54882]= 2146380306;
assign addr[54883]= 2145835515;
assign addr[54884]= 2134405552;
assign addr[54885]= 2112148396;
assign addr[54886]= 2079176953;
assign addr[54887]= 2035658475;
assign addr[54888]= 1981813720;
assign addr[54889]= 1917915825;
assign addr[54890]= 1844288924;
assign addr[54891]= 1761306505;
assign addr[54892]= 1669389513;
assign addr[54893]= 1569004214;
assign addr[54894]= 1460659832;
assign addr[54895]= 1344905966;
assign addr[54896]= 1222329801;
assign addr[54897]= 1093553126;
assign addr[54898]= 959229189;
assign addr[54899]= 820039373;
assign addr[54900]= 676689746;
assign addr[54901]= 529907477;
assign addr[54902]= 380437148;
assign addr[54903]= 229036977;
assign addr[54904]= 76474970;
assign addr[54905]= -76474970;
assign addr[54906]= -229036977;
assign addr[54907]= -380437148;
assign addr[54908]= -529907477;
assign addr[54909]= -676689746;
assign addr[54910]= -820039373;
assign addr[54911]= -959229189;
assign addr[54912]= -1093553126;
assign addr[54913]= -1222329801;
assign addr[54914]= -1344905966;
assign addr[54915]= -1460659832;
assign addr[54916]= -1569004214;
assign addr[54917]= -1669389513;
assign addr[54918]= -1761306505;
assign addr[54919]= -1844288924;
assign addr[54920]= -1917915825;
assign addr[54921]= -1981813720;
assign addr[54922]= -2035658475;
assign addr[54923]= -2079176953;
assign addr[54924]= -2112148396;
assign addr[54925]= -2134405552;
assign addr[54926]= -2145835515;
assign addr[54927]= -2146380306;
assign addr[54928]= -2136037160;
assign addr[54929]= -2114858546;
assign addr[54930]= -2082951896;
assign addr[54931]= -2040479063;
assign addr[54932]= -1987655498;
assign addr[54933]= -1924749160;
assign addr[54934]= -1852079154;
assign addr[54935]= -1770014111;
assign addr[54936]= -1678970324;
assign addr[54937]= -1579409630;
assign addr[54938]= -1471837070;
assign addr[54939]= -1356798326;
assign addr[54940]= -1234876957;
assign addr[54941]= -1106691431;
assign addr[54942]= -972891995;
assign addr[54943]= -834157373;
assign addr[54944]= -691191324;
assign addr[54945]= -544719071;
assign addr[54946]= -395483624;
assign addr[54947]= -244242007;
assign addr[54948]= -91761426;
assign addr[54949]= 61184634;
assign addr[54950]= 213820322;
assign addr[54951]= 365371365;
assign addr[54952]= 515068990;
assign addr[54953]= 662153826;
assign addr[54954]= 805879757;
assign addr[54955]= 945517704;
assign addr[54956]= 1080359326;
assign addr[54957]= 1209720613;
assign addr[54958]= 1332945355;
assign addr[54959]= 1449408469;
assign addr[54960]= 1558519173;
assign addr[54961]= 1659723983;
assign addr[54962]= 1752509516;
assign addr[54963]= 1836405100;
assign addr[54964]= 1910985158;
assign addr[54965]= 1975871368;
assign addr[54966]= 2030734582;
assign addr[54967]= 2075296495;
assign addr[54968]= 2109331059;
assign addr[54969]= 2132665626;
assign addr[54970]= 2145181827;
assign addr[54971]= 2146816171;
assign addr[54972]= 2137560369;
assign addr[54973]= 2117461370;
assign addr[54974]= 2086621133;
assign addr[54975]= 2045196100;
assign addr[54976]= 1993396407;
assign addr[54977]= 1931484818;
assign addr[54978]= 1859775393;
assign addr[54979]= 1778631892;
assign addr[54980]= 1688465931;
assign addr[54981]= 1589734894;
assign addr[54982]= 1482939614;
assign addr[54983]= 1368621831;
assign addr[54984]= 1247361445;
assign addr[54985]= 1119773573;
assign addr[54986]= 986505429;
assign addr[54987]= 848233042;
assign addr[54988]= 705657826;
assign addr[54989]= 559503022;
assign addr[54990]= 410510029;
assign addr[54991]= 259434643;
assign addr[54992]= 107043224;
assign addr[54993]= -45891193;
assign addr[54994]= -198592817;
assign addr[54995]= -350287041;
assign addr[54996]= -500204365;
assign addr[54997]= -647584304;
assign addr[54998]= -791679244;
assign addr[54999]= -931758235;
assign addr[55000]= -1067110699;
assign addr[55001]= -1197050035;
assign addr[55002]= -1320917099;
assign addr[55003]= -1438083551;
assign addr[55004]= -1547955041;
assign addr[55005]= -1649974225;
assign addr[55006]= -1743623590;
assign addr[55007]= -1828428082;
assign addr[55008]= -1903957513;
assign addr[55009]= -1969828744;
assign addr[55010]= -2025707632;
assign addr[55011]= -2071310720;
assign addr[55012]= -2106406677;
assign addr[55013]= -2130817471;
assign addr[55014]= -2144419275;
assign addr[55015]= -2147143090;
assign addr[55016]= -2138975100;
assign addr[55017]= -2119956737;
assign addr[55018]= -2090184478;
assign addr[55019]= -2049809346;
assign addr[55020]= -1999036154;
assign addr[55021]= -1938122457;
assign addr[55022]= -1867377253;
assign addr[55023]= -1787159411;
assign addr[55024]= -1697875851;
assign addr[55025]= -1599979481;
assign addr[55026]= -1493966902;
assign addr[55027]= -1380375881;
assign addr[55028]= -1259782632;
assign addr[55029]= -1132798888;
assign addr[55030]= -1000068799;
assign addr[55031]= -862265664;
assign addr[55032]= -720088517;
assign addr[55033]= -574258580;
assign addr[55034]= -425515602;
assign addr[55035]= -274614114;
assign addr[55036]= -122319591;
assign addr[55037]= 30595422;
assign addr[55038]= 183355234;
assign addr[55039]= 335184940;
assign addr[55040]= 485314355;
assign addr[55041]= 632981917;
assign addr[55042]= 777438554;
assign addr[55043]= 917951481;
assign addr[55044]= 1053807919;
assign addr[55045]= 1184318708;
assign addr[55046]= 1308821808;
assign addr[55047]= 1426685652;
assign addr[55048]= 1537312353;
assign addr[55049]= 1640140734;
assign addr[55050]= 1734649179;
assign addr[55051]= 1820358275;
assign addr[55052]= 1896833245;
assign addr[55053]= 1963686155;
assign addr[55054]= 2020577882;
assign addr[55055]= 2067219829;
assign addr[55056]= 2103375398;
assign addr[55057]= 2128861181;
assign addr[55058]= 2143547897;
assign addr[55059]= 2147361045;
assign addr[55060]= 2140281282;
assign addr[55061]= 2122344521;
assign addr[55062]= 2093641749;
assign addr[55063]= 2054318569;
assign addr[55064]= 2004574453;
assign addr[55065]= 1944661739;
assign addr[55066]= 1874884346;
assign addr[55067]= 1795596234;
assign addr[55068]= 1707199606;
assign addr[55069]= 1610142873;
assign addr[55070]= 1504918373;
assign addr[55071]= 1392059879;
assign addr[55072]= 1272139887;
assign addr[55073]= 1145766716;
assign addr[55074]= 1013581418;
assign addr[55075]= 876254528;
assign addr[55076]= 734482665;
assign addr[55077]= 588984994;
assign addr[55078]= 440499581;
assign addr[55079]= 289779648;
assign addr[55080]= 137589750;
assign addr[55081]= -15298099;
assign addr[55082]= -168108346;
assign addr[55083]= -320065829;
assign addr[55084]= -470399716;
assign addr[55085]= -618347408;
assign addr[55086]= -763158411;
assign addr[55087]= -904098143;
assign addr[55088]= -1040451659;
assign addr[55089]= -1171527280;
assign addr[55090]= -1296660098;
assign addr[55091]= -1415215352;
assign addr[55092]= -1526591649;
assign addr[55093]= -1630224009;
assign addr[55094]= -1725586737;
assign addr[55095]= -1812196087;
assign addr[55096]= -1889612716;
assign addr[55097]= -1957443913;
assign addr[55098]= -2015345591;
assign addr[55099]= -2063024031;
assign addr[55100]= -2100237377;
assign addr[55101]= -2126796855;
assign addr[55102]= -2142567738;
assign addr[55103]= -2147470025;
assign addr[55104]= -2141478848;
assign addr[55105]= -2124624598;
assign addr[55106]= -2096992772;
assign addr[55107]= -2058723538;
assign addr[55108]= -2010011024;
assign addr[55109]= -1951102334;
assign addr[55110]= -1882296293;
assign addr[55111]= -1803941934;
assign addr[55112]= -1716436725;
assign addr[55113]= -1620224553;
assign addr[55114]= -1515793473;
assign addr[55115]= -1403673233;
assign addr[55116]= -1284432584;
assign addr[55117]= -1158676398;
assign addr[55118]= -1027042599;
assign addr[55119]= -890198924;
assign addr[55120]= -748839539;
assign addr[55121]= -603681519;
assign addr[55122]= -455461206;
assign addr[55123]= -304930476;
assign addr[55124]= -152852926;
assign addr[55125]= 0;
assign addr[55126]= 152852926;
assign addr[55127]= 304930476;
assign addr[55128]= 455461206;
assign addr[55129]= 603681519;
assign addr[55130]= 748839539;
assign addr[55131]= 890198924;
assign addr[55132]= 1027042599;
assign addr[55133]= 1158676398;
assign addr[55134]= 1284432584;
assign addr[55135]= 1403673233;
assign addr[55136]= 1515793473;
assign addr[55137]= 1620224553;
assign addr[55138]= 1716436725;
assign addr[55139]= 1803941934;
assign addr[55140]= 1882296293;
assign addr[55141]= 1951102334;
assign addr[55142]= 2010011024;
assign addr[55143]= 2058723538;
assign addr[55144]= 2096992772;
assign addr[55145]= 2124624598;
assign addr[55146]= 2141478848;
assign addr[55147]= 2147470025;
assign addr[55148]= 2142567738;
assign addr[55149]= 2126796855;
assign addr[55150]= 2100237377;
assign addr[55151]= 2063024031;
assign addr[55152]= 2015345591;
assign addr[55153]= 1957443913;
assign addr[55154]= 1889612716;
assign addr[55155]= 1812196087;
assign addr[55156]= 1725586737;
assign addr[55157]= 1630224009;
assign addr[55158]= 1526591649;
assign addr[55159]= 1415215352;
assign addr[55160]= 1296660098;
assign addr[55161]= 1171527280;
assign addr[55162]= 1040451659;
assign addr[55163]= 904098143;
assign addr[55164]= 763158411;
assign addr[55165]= 618347408;
assign addr[55166]= 470399716;
assign addr[55167]= 320065829;
assign addr[55168]= 168108346;
assign addr[55169]= 15298099;
assign addr[55170]= -137589750;
assign addr[55171]= -289779648;
assign addr[55172]= -440499581;
assign addr[55173]= -588984994;
assign addr[55174]= -734482665;
assign addr[55175]= -876254528;
assign addr[55176]= -1013581418;
assign addr[55177]= -1145766716;
assign addr[55178]= -1272139887;
assign addr[55179]= -1392059879;
assign addr[55180]= -1504918373;
assign addr[55181]= -1610142873;
assign addr[55182]= -1707199606;
assign addr[55183]= -1795596234;
assign addr[55184]= -1874884346;
assign addr[55185]= -1944661739;
assign addr[55186]= -2004574453;
assign addr[55187]= -2054318569;
assign addr[55188]= -2093641749;
assign addr[55189]= -2122344521;
assign addr[55190]= -2140281282;
assign addr[55191]= -2147361045;
assign addr[55192]= -2143547897;
assign addr[55193]= -2128861181;
assign addr[55194]= -2103375398;
assign addr[55195]= -2067219829;
assign addr[55196]= -2020577882;
assign addr[55197]= -1963686155;
assign addr[55198]= -1896833245;
assign addr[55199]= -1820358275;
assign addr[55200]= -1734649179;
assign addr[55201]= -1640140734;
assign addr[55202]= -1537312353;
assign addr[55203]= -1426685652;
assign addr[55204]= -1308821808;
assign addr[55205]= -1184318708;
assign addr[55206]= -1053807919;
assign addr[55207]= -917951481;
assign addr[55208]= -777438554;
assign addr[55209]= -632981917;
assign addr[55210]= -485314355;
assign addr[55211]= -335184940;
assign addr[55212]= -183355234;
assign addr[55213]= -30595422;
assign addr[55214]= 122319591;
assign addr[55215]= 274614114;
assign addr[55216]= 425515602;
assign addr[55217]= 574258580;
assign addr[55218]= 720088517;
assign addr[55219]= 862265664;
assign addr[55220]= 1000068799;
assign addr[55221]= 1132798888;
assign addr[55222]= 1259782632;
assign addr[55223]= 1380375881;
assign addr[55224]= 1493966902;
assign addr[55225]= 1599979481;
assign addr[55226]= 1697875851;
assign addr[55227]= 1787159411;
assign addr[55228]= 1867377253;
assign addr[55229]= 1938122457;
assign addr[55230]= 1999036154;
assign addr[55231]= 2049809346;
assign addr[55232]= 2090184478;
assign addr[55233]= 2119956737;
assign addr[55234]= 2138975100;
assign addr[55235]= 2147143090;
assign addr[55236]= 2144419275;
assign addr[55237]= 2130817471;
assign addr[55238]= 2106406677;
assign addr[55239]= 2071310720;
assign addr[55240]= 2025707632;
assign addr[55241]= 1969828744;
assign addr[55242]= 1903957513;
assign addr[55243]= 1828428082;
assign addr[55244]= 1743623590;
assign addr[55245]= 1649974225;
assign addr[55246]= 1547955041;
assign addr[55247]= 1438083551;
assign addr[55248]= 1320917099;
assign addr[55249]= 1197050035;
assign addr[55250]= 1067110699;
assign addr[55251]= 931758235;
assign addr[55252]= 791679244;
assign addr[55253]= 647584304;
assign addr[55254]= 500204365;
assign addr[55255]= 350287041;
assign addr[55256]= 198592817;
assign addr[55257]= 45891193;
assign addr[55258]= -107043224;
assign addr[55259]= -259434643;
assign addr[55260]= -410510029;
assign addr[55261]= -559503022;
assign addr[55262]= -705657826;
assign addr[55263]= -848233042;
assign addr[55264]= -986505429;
assign addr[55265]= -1119773573;
assign addr[55266]= -1247361445;
assign addr[55267]= -1368621831;
assign addr[55268]= -1482939614;
assign addr[55269]= -1589734894;
assign addr[55270]= -1688465931;
assign addr[55271]= -1778631892;
assign addr[55272]= -1859775393;
assign addr[55273]= -1931484818;
assign addr[55274]= -1993396407;
assign addr[55275]= -2045196100;
assign addr[55276]= -2086621133;
assign addr[55277]= -2117461370;
assign addr[55278]= -2137560369;
assign addr[55279]= -2146816171;
assign addr[55280]= -2145181827;
assign addr[55281]= -2132665626;
assign addr[55282]= -2109331059;
assign addr[55283]= -2075296495;
assign addr[55284]= -2030734582;
assign addr[55285]= -1975871368;
assign addr[55286]= -1910985158;
assign addr[55287]= -1836405100;
assign addr[55288]= -1752509516;
assign addr[55289]= -1659723983;
assign addr[55290]= -1558519173;
assign addr[55291]= -1449408469;
assign addr[55292]= -1332945355;
assign addr[55293]= -1209720613;
assign addr[55294]= -1080359326;
assign addr[55295]= -945517704;
assign addr[55296]= -805879757;
assign addr[55297]= -662153826;
assign addr[55298]= -515068990;
assign addr[55299]= -365371365;
assign addr[55300]= -213820322;
assign addr[55301]= -61184634;
assign addr[55302]= 91761426;
assign addr[55303]= 244242007;
assign addr[55304]= 395483624;
assign addr[55305]= 544719071;
assign addr[55306]= 691191324;
assign addr[55307]= 834157373;
assign addr[55308]= 972891995;
assign addr[55309]= 1106691431;
assign addr[55310]= 1234876957;
assign addr[55311]= 1356798326;
assign addr[55312]= 1471837070;
assign addr[55313]= 1579409630;
assign addr[55314]= 1678970324;
assign addr[55315]= 1770014111;
assign addr[55316]= 1852079154;
assign addr[55317]= 1924749160;
assign addr[55318]= 1987655498;
assign addr[55319]= 2040479063;
assign addr[55320]= 2082951896;
assign addr[55321]= 2114858546;
assign addr[55322]= 2136037160;
assign addr[55323]= 2146380306;
assign addr[55324]= 2145835515;
assign addr[55325]= 2134405552;
assign addr[55326]= 2112148396;
assign addr[55327]= 2079176953;
assign addr[55328]= 2035658475;
assign addr[55329]= 1981813720;
assign addr[55330]= 1917915825;
assign addr[55331]= 1844288924;
assign addr[55332]= 1761306505;
assign addr[55333]= 1669389513;
assign addr[55334]= 1569004214;
assign addr[55335]= 1460659832;
assign addr[55336]= 1344905966;
assign addr[55337]= 1222329801;
assign addr[55338]= 1093553126;
assign addr[55339]= 959229189;
assign addr[55340]= 820039373;
assign addr[55341]= 676689746;
assign addr[55342]= 529907477;
assign addr[55343]= 380437148;
assign addr[55344]= 229036977;
assign addr[55345]= 76474970;
assign addr[55346]= -76474970;
assign addr[55347]= -229036977;
assign addr[55348]= -380437148;
assign addr[55349]= -529907477;
assign addr[55350]= -676689746;
assign addr[55351]= -820039373;
assign addr[55352]= -959229189;
assign addr[55353]= -1093553126;
assign addr[55354]= -1222329801;
assign addr[55355]= -1344905966;
assign addr[55356]= -1460659832;
assign addr[55357]= -1569004214;
assign addr[55358]= -1669389513;
assign addr[55359]= -1761306505;
assign addr[55360]= -1844288924;
assign addr[55361]= -1917915825;
assign addr[55362]= -1981813720;
assign addr[55363]= -2035658475;
assign addr[55364]= -2079176953;
assign addr[55365]= -2112148396;
assign addr[55366]= -2134405552;
assign addr[55367]= -2145835515;
assign addr[55368]= -2146380306;
assign addr[55369]= -2136037160;
assign addr[55370]= -2114858546;
assign addr[55371]= -2082951896;
assign addr[55372]= -2040479063;
assign addr[55373]= -1987655498;
assign addr[55374]= -1924749160;
assign addr[55375]= -1852079154;
assign addr[55376]= -1770014111;
assign addr[55377]= -1678970324;
assign addr[55378]= -1579409630;
assign addr[55379]= -1471837070;
assign addr[55380]= -1356798326;
assign addr[55381]= -1234876957;
assign addr[55382]= -1106691431;
assign addr[55383]= -972891995;
assign addr[55384]= -834157373;
assign addr[55385]= -691191324;
assign addr[55386]= -544719071;
assign addr[55387]= -395483624;
assign addr[55388]= -244242007;
assign addr[55389]= -91761426;
assign addr[55390]= 61184634;
assign addr[55391]= 213820322;
assign addr[55392]= 365371365;
assign addr[55393]= 515068990;
assign addr[55394]= 662153826;
assign addr[55395]= 805879757;
assign addr[55396]= 945517704;
assign addr[55397]= 1080359326;
assign addr[55398]= 1209720613;
assign addr[55399]= 1332945355;
assign addr[55400]= 1449408469;
assign addr[55401]= 1558519173;
assign addr[55402]= 1659723983;
assign addr[55403]= 1752509516;
assign addr[55404]= 1836405100;
assign addr[55405]= 1910985158;
assign addr[55406]= 1975871368;
assign addr[55407]= 2030734582;
assign addr[55408]= 2075296495;
assign addr[55409]= 2109331059;
assign addr[55410]= 2132665626;
assign addr[55411]= 2145181827;
assign addr[55412]= 2146816171;
assign addr[55413]= 2137560369;
assign addr[55414]= 2117461370;
assign addr[55415]= 2086621133;
assign addr[55416]= 2045196100;
assign addr[55417]= 1993396407;
assign addr[55418]= 1931484818;
assign addr[55419]= 1859775393;
assign addr[55420]= 1778631892;
assign addr[55421]= 1688465931;
assign addr[55422]= 1589734894;
assign addr[55423]= 1482939614;
assign addr[55424]= 1368621831;
assign addr[55425]= 1247361445;
assign addr[55426]= 1119773573;
assign addr[55427]= 986505429;
assign addr[55428]= 848233042;
assign addr[55429]= 705657826;
assign addr[55430]= 559503022;
assign addr[55431]= 410510029;
assign addr[55432]= 259434643;
assign addr[55433]= 107043224;
assign addr[55434]= -45891193;
assign addr[55435]= -198592817;
assign addr[55436]= -350287041;
assign addr[55437]= -500204365;
assign addr[55438]= -647584304;
assign addr[55439]= -791679244;
assign addr[55440]= -931758235;
assign addr[55441]= -1067110699;
assign addr[55442]= -1197050035;
assign addr[55443]= -1320917099;
assign addr[55444]= -1438083551;
assign addr[55445]= -1547955041;
assign addr[55446]= -1649974225;
assign addr[55447]= -1743623590;
assign addr[55448]= -1828428082;
assign addr[55449]= -1903957513;
assign addr[55450]= -1969828744;
assign addr[55451]= -2025707632;
assign addr[55452]= -2071310720;
assign addr[55453]= -2106406677;
assign addr[55454]= -2130817471;
assign addr[55455]= -2144419275;
assign addr[55456]= -2147143090;
assign addr[55457]= -2138975100;
assign addr[55458]= -2119956737;
assign addr[55459]= -2090184478;
assign addr[55460]= -2049809346;
assign addr[55461]= -1999036154;
assign addr[55462]= -1938122457;
assign addr[55463]= -1867377253;
assign addr[55464]= -1787159411;
assign addr[55465]= -1697875851;
assign addr[55466]= -1599979481;
assign addr[55467]= -1493966902;
assign addr[55468]= -1380375881;
assign addr[55469]= -1259782632;
assign addr[55470]= -1132798888;
assign addr[55471]= -1000068799;
assign addr[55472]= -862265664;
assign addr[55473]= -720088517;
assign addr[55474]= -574258580;
assign addr[55475]= -425515602;
assign addr[55476]= -274614114;
assign addr[55477]= -122319591;
assign addr[55478]= 30595422;
assign addr[55479]= 183355234;
assign addr[55480]= 335184940;
assign addr[55481]= 485314355;
assign addr[55482]= 632981917;
assign addr[55483]= 777438554;
assign addr[55484]= 917951481;
assign addr[55485]= 1053807919;
assign addr[55486]= 1184318708;
assign addr[55487]= 1308821808;
assign addr[55488]= 1426685652;
assign addr[55489]= 1537312353;
assign addr[55490]= 1640140734;
assign addr[55491]= 1734649179;
assign addr[55492]= 1820358275;
assign addr[55493]= 1896833245;
assign addr[55494]= 1963686155;
assign addr[55495]= 2020577882;
assign addr[55496]= 2067219829;
assign addr[55497]= 2103375398;
assign addr[55498]= 2128861181;
assign addr[55499]= 2143547897;
assign addr[55500]= 2147361045;
assign addr[55501]= 2140281282;
assign addr[55502]= 2122344521;
assign addr[55503]= 2093641749;
assign addr[55504]= 2054318569;
assign addr[55505]= 2004574453;
assign addr[55506]= 1944661739;
assign addr[55507]= 1874884346;
assign addr[55508]= 1795596234;
assign addr[55509]= 1707199606;
assign addr[55510]= 1610142873;
assign addr[55511]= 1504918373;
assign addr[55512]= 1392059879;
assign addr[55513]= 1272139887;
assign addr[55514]= 1145766716;
assign addr[55515]= 1013581418;
assign addr[55516]= 876254528;
assign addr[55517]= 734482665;
assign addr[55518]= 588984994;
assign addr[55519]= 440499581;
assign addr[55520]= 289779648;
assign addr[55521]= 137589750;
assign addr[55522]= -15298099;
assign addr[55523]= -168108346;
assign addr[55524]= -320065829;
assign addr[55525]= -470399716;
assign addr[55526]= -618347408;
assign addr[55527]= -763158411;
assign addr[55528]= -904098143;
assign addr[55529]= -1040451659;
assign addr[55530]= -1171527280;
assign addr[55531]= -1296660098;
assign addr[55532]= -1415215352;
assign addr[55533]= -1526591649;
assign addr[55534]= -1630224009;
assign addr[55535]= -1725586737;
assign addr[55536]= -1812196087;
assign addr[55537]= -1889612716;
assign addr[55538]= -1957443913;
assign addr[55539]= -2015345591;
assign addr[55540]= -2063024031;
assign addr[55541]= -2100237377;
assign addr[55542]= -2126796855;
assign addr[55543]= -2142567738;
assign addr[55544]= -2147470025;
assign addr[55545]= -2141478848;
assign addr[55546]= -2124624598;
assign addr[55547]= -2096992772;
assign addr[55548]= -2058723538;
assign addr[55549]= -2010011024;
assign addr[55550]= -1951102334;
assign addr[55551]= -1882296293;
assign addr[55552]= -1803941934;
assign addr[55553]= -1716436725;
assign addr[55554]= -1620224553;
assign addr[55555]= -1515793473;
assign addr[55556]= -1403673233;
assign addr[55557]= -1284432584;
assign addr[55558]= -1158676398;
assign addr[55559]= -1027042599;
assign addr[55560]= -890198924;
assign addr[55561]= -748839539;
assign addr[55562]= -603681519;
assign addr[55563]= -455461206;
assign addr[55564]= -304930476;
assign addr[55565]= -152852926;
assign addr[55566]= 0;
assign addr[55567]= 152852926;
assign addr[55568]= 304930476;
assign addr[55569]= 455461206;
assign addr[55570]= 603681519;
assign addr[55571]= 748839539;
assign addr[55572]= 890198924;
assign addr[55573]= 1027042599;
assign addr[55574]= 1158676398;
assign addr[55575]= 1284432584;
assign addr[55576]= 1403673233;
assign addr[55577]= 1515793473;
assign addr[55578]= 1620224553;
assign addr[55579]= 1716436725;
assign addr[55580]= 1803941934;
assign addr[55581]= 1882296293;
assign addr[55582]= 1951102334;
assign addr[55583]= 2010011024;
assign addr[55584]= 2058723538;
assign addr[55585]= 2096992772;
assign addr[55586]= 2124624598;
assign addr[55587]= 2141478848;
assign addr[55588]= 2147470025;
assign addr[55589]= 2142567738;
assign addr[55590]= 2126796855;
assign addr[55591]= 2100237377;
assign addr[55592]= 2063024031;
assign addr[55593]= 2015345591;
assign addr[55594]= 1957443913;
assign addr[55595]= 1889612716;
assign addr[55596]= 1812196087;
assign addr[55597]= 1725586737;
assign addr[55598]= 1630224009;
assign addr[55599]= 1526591649;
assign addr[55600]= 1415215352;
assign addr[55601]= 1296660098;
assign addr[55602]= 1171527280;
assign addr[55603]= 1040451659;
assign addr[55604]= 904098143;
assign addr[55605]= 763158411;
assign addr[55606]= 618347408;
assign addr[55607]= 470399716;
assign addr[55608]= 320065829;
assign addr[55609]= 168108346;
assign addr[55610]= 15298099;
assign addr[55611]= -137589750;
assign addr[55612]= -289779648;
assign addr[55613]= -440499581;
assign addr[55614]= -588984994;
assign addr[55615]= -734482665;
assign addr[55616]= -876254528;
assign addr[55617]= -1013581418;
assign addr[55618]= -1145766716;
assign addr[55619]= -1272139887;
assign addr[55620]= -1392059879;
assign addr[55621]= -1504918373;
assign addr[55622]= -1610142873;
assign addr[55623]= -1707199606;
assign addr[55624]= -1795596234;
assign addr[55625]= -1874884346;
assign addr[55626]= -1944661739;
assign addr[55627]= -2004574453;
assign addr[55628]= -2054318569;
assign addr[55629]= -2093641749;
assign addr[55630]= -2122344521;
assign addr[55631]= -2140281282;
assign addr[55632]= -2147361045;
assign addr[55633]= -2143547897;
assign addr[55634]= -2128861181;
assign addr[55635]= -2103375398;
assign addr[55636]= -2067219829;
assign addr[55637]= -2020577882;
assign addr[55638]= -1963686155;
assign addr[55639]= -1896833245;
assign addr[55640]= -1820358275;
assign addr[55641]= -1734649179;
assign addr[55642]= -1640140734;
assign addr[55643]= -1537312353;
assign addr[55644]= -1426685652;
assign addr[55645]= -1308821808;
assign addr[55646]= -1184318708;
assign addr[55647]= -1053807919;
assign addr[55648]= -917951481;
assign addr[55649]= -777438554;
assign addr[55650]= -632981917;
assign addr[55651]= -485314355;
assign addr[55652]= -335184940;
assign addr[55653]= -183355234;
assign addr[55654]= -30595422;
assign addr[55655]= 122319591;
assign addr[55656]= 274614114;
assign addr[55657]= 425515602;
assign addr[55658]= 574258580;
assign addr[55659]= 720088517;
assign addr[55660]= 862265664;
assign addr[55661]= 1000068799;
assign addr[55662]= 1132798888;
assign addr[55663]= 1259782632;
assign addr[55664]= 1380375881;
assign addr[55665]= 1493966902;
assign addr[55666]= 1599979481;
assign addr[55667]= 1697875851;
assign addr[55668]= 1787159411;
assign addr[55669]= 1867377253;
assign addr[55670]= 1938122457;
assign addr[55671]= 1999036154;
assign addr[55672]= 2049809346;
assign addr[55673]= 2090184478;
assign addr[55674]= 2119956737;
assign addr[55675]= 2138975100;
assign addr[55676]= 2147143090;
assign addr[55677]= 2144419275;
assign addr[55678]= 2130817471;
assign addr[55679]= 2106406677;
assign addr[55680]= 2071310720;
assign addr[55681]= 2025707632;
assign addr[55682]= 1969828744;
assign addr[55683]= 1903957513;
assign addr[55684]= 1828428082;
assign addr[55685]= 1743623590;
assign addr[55686]= 1649974225;
assign addr[55687]= 1547955041;
assign addr[55688]= 1438083551;
assign addr[55689]= 1320917099;
assign addr[55690]= 1197050035;
assign addr[55691]= 1067110699;
assign addr[55692]= 931758235;
assign addr[55693]= 791679244;
assign addr[55694]= 647584304;
assign addr[55695]= 500204365;
assign addr[55696]= 350287041;
assign addr[55697]= 198592817;
assign addr[55698]= 45891193;
assign addr[55699]= -107043224;
assign addr[55700]= -259434643;
assign addr[55701]= -410510029;
assign addr[55702]= -559503022;
assign addr[55703]= -705657826;
assign addr[55704]= -848233042;
assign addr[55705]= -986505429;
assign addr[55706]= -1119773573;
assign addr[55707]= -1247361445;
assign addr[55708]= -1368621831;
assign addr[55709]= -1482939614;
assign addr[55710]= -1589734894;
assign addr[55711]= -1688465931;
assign addr[55712]= -1778631892;
assign addr[55713]= -1859775393;
assign addr[55714]= -1931484818;
assign addr[55715]= -1993396407;
assign addr[55716]= -2045196100;
assign addr[55717]= -2086621133;
assign addr[55718]= -2117461370;
assign addr[55719]= -2137560369;
assign addr[55720]= -2146816171;
assign addr[55721]= -2145181827;
assign addr[55722]= -2132665626;
assign addr[55723]= -2109331059;
assign addr[55724]= -2075296495;
assign addr[55725]= -2030734582;
assign addr[55726]= -1975871368;
assign addr[55727]= -1910985158;
assign addr[55728]= -1836405100;
assign addr[55729]= -1752509516;
assign addr[55730]= -1659723983;
assign addr[55731]= -1558519173;
assign addr[55732]= -1449408469;
assign addr[55733]= -1332945355;
assign addr[55734]= -1209720613;
assign addr[55735]= -1080359326;
assign addr[55736]= -945517704;
assign addr[55737]= -805879757;
assign addr[55738]= -662153826;
assign addr[55739]= -515068990;
assign addr[55740]= -365371365;
assign addr[55741]= -213820322;
assign addr[55742]= -61184634;
assign addr[55743]= 91761426;
assign addr[55744]= 244242007;
assign addr[55745]= 395483624;
assign addr[55746]= 544719071;
assign addr[55747]= 691191324;
assign addr[55748]= 834157373;
assign addr[55749]= 972891995;
assign addr[55750]= 1106691431;
assign addr[55751]= 1234876957;
assign addr[55752]= 1356798326;
assign addr[55753]= 1471837070;
assign addr[55754]= 1579409630;
assign addr[55755]= 1678970324;
assign addr[55756]= 1770014111;
assign addr[55757]= 1852079154;
assign addr[55758]= 1924749160;
assign addr[55759]= 1987655498;
assign addr[55760]= 2040479063;
assign addr[55761]= 2082951896;
assign addr[55762]= 2114858546;
assign addr[55763]= 2136037160;
assign addr[55764]= 2146380306;
assign addr[55765]= 2145835515;
assign addr[55766]= 2134405552;
assign addr[55767]= 2112148396;
assign addr[55768]= 2079176953;
assign addr[55769]= 2035658475;
assign addr[55770]= 1981813720;
assign addr[55771]= 1917915825;
assign addr[55772]= 1844288924;
assign addr[55773]= 1761306505;
assign addr[55774]= 1669389513;
assign addr[55775]= 1569004214;
assign addr[55776]= 1460659832;
assign addr[55777]= 1344905966;
assign addr[55778]= 1222329801;
assign addr[55779]= 1093553126;
assign addr[55780]= 959229189;
assign addr[55781]= 820039373;
assign addr[55782]= 676689746;
assign addr[55783]= 529907477;
assign addr[55784]= 380437148;
assign addr[55785]= 229036977;
assign addr[55786]= 76474970;
assign addr[55787]= -76474970;
assign addr[55788]= -229036977;
assign addr[55789]= -380437148;
assign addr[55790]= -529907477;
assign addr[55791]= -676689746;
assign addr[55792]= -820039373;
assign addr[55793]= -959229189;
assign addr[55794]= -1093553126;
assign addr[55795]= -1222329801;
assign addr[55796]= -1344905966;
assign addr[55797]= -1460659832;
assign addr[55798]= -1569004214;
assign addr[55799]= -1669389513;
assign addr[55800]= -1761306505;
assign addr[55801]= -1844288924;
assign addr[55802]= -1917915825;
assign addr[55803]= -1981813720;
assign addr[55804]= -2035658475;
assign addr[55805]= -2079176953;
assign addr[55806]= -2112148396;
assign addr[55807]= -2134405552;
assign addr[55808]= -2145835515;
assign addr[55809]= -2146380306;
assign addr[55810]= -2136037160;
assign addr[55811]= -2114858546;
assign addr[55812]= -2082951896;
assign addr[55813]= -2040479063;
assign addr[55814]= -1987655498;
assign addr[55815]= -1924749160;
assign addr[55816]= -1852079154;
assign addr[55817]= -1770014111;
assign addr[55818]= -1678970324;
assign addr[55819]= -1579409630;
assign addr[55820]= -1471837070;
assign addr[55821]= -1356798326;
assign addr[55822]= -1234876957;
assign addr[55823]= -1106691431;
assign addr[55824]= -972891995;
assign addr[55825]= -834157373;
assign addr[55826]= -691191324;
assign addr[55827]= -544719071;
assign addr[55828]= -395483624;
assign addr[55829]= -244242007;
assign addr[55830]= -91761426;
assign addr[55831]= 61184634;
assign addr[55832]= 213820322;
assign addr[55833]= 365371365;
assign addr[55834]= 515068990;
assign addr[55835]= 662153826;
assign addr[55836]= 805879757;
assign addr[55837]= 945517704;
assign addr[55838]= 1080359326;
assign addr[55839]= 1209720613;
assign addr[55840]= 1332945355;
assign addr[55841]= 1449408469;
assign addr[55842]= 1558519173;
assign addr[55843]= 1659723983;
assign addr[55844]= 1752509516;
assign addr[55845]= 1836405100;
assign addr[55846]= 1910985158;
assign addr[55847]= 1975871368;
assign addr[55848]= 2030734582;
assign addr[55849]= 2075296495;
assign addr[55850]= 2109331059;
assign addr[55851]= 2132665626;
assign addr[55852]= 2145181827;
assign addr[55853]= 2146816171;
assign addr[55854]= 2137560369;
assign addr[55855]= 2117461370;
assign addr[55856]= 2086621133;
assign addr[55857]= 2045196100;
assign addr[55858]= 1993396407;
assign addr[55859]= 1931484818;
assign addr[55860]= 1859775393;
assign addr[55861]= 1778631892;
assign addr[55862]= 1688465931;
assign addr[55863]= 1589734894;
assign addr[55864]= 1482939614;
assign addr[55865]= 1368621831;
assign addr[55866]= 1247361445;
assign addr[55867]= 1119773573;
assign addr[55868]= 986505429;
assign addr[55869]= 848233042;
assign addr[55870]= 705657826;
assign addr[55871]= 559503022;
assign addr[55872]= 410510029;
assign addr[55873]= 259434643;
assign addr[55874]= 107043224;
assign addr[55875]= -45891193;
assign addr[55876]= -198592817;
assign addr[55877]= -350287041;
assign addr[55878]= -500204365;
assign addr[55879]= -647584304;
assign addr[55880]= -791679244;
assign addr[55881]= -931758235;
assign addr[55882]= -1067110699;
assign addr[55883]= -1197050035;
assign addr[55884]= -1320917099;
assign addr[55885]= -1438083551;
assign addr[55886]= -1547955041;
assign addr[55887]= -1649974225;
assign addr[55888]= -1743623590;
assign addr[55889]= -1828428082;
assign addr[55890]= -1903957513;
assign addr[55891]= -1969828744;
assign addr[55892]= -2025707632;
assign addr[55893]= -2071310720;
assign addr[55894]= -2106406677;
assign addr[55895]= -2130817471;
assign addr[55896]= -2144419275;
assign addr[55897]= -2147143090;
assign addr[55898]= -2138975100;
assign addr[55899]= -2119956737;
assign addr[55900]= -2090184478;
assign addr[55901]= -2049809346;
assign addr[55902]= -1999036154;
assign addr[55903]= -1938122457;
assign addr[55904]= -1867377253;
assign addr[55905]= -1787159411;
assign addr[55906]= -1697875851;
assign addr[55907]= -1599979481;
assign addr[55908]= -1493966902;
assign addr[55909]= -1380375881;
assign addr[55910]= -1259782632;
assign addr[55911]= -1132798888;
assign addr[55912]= -1000068799;
assign addr[55913]= -862265664;
assign addr[55914]= -720088517;
assign addr[55915]= -574258580;
assign addr[55916]= -425515602;
assign addr[55917]= -274614114;
assign addr[55918]= -122319591;
assign addr[55919]= 30595422;
assign addr[55920]= 183355234;
assign addr[55921]= 335184940;
assign addr[55922]= 485314355;
assign addr[55923]= 632981917;
assign addr[55924]= 777438554;
assign addr[55925]= 917951481;
assign addr[55926]= 1053807919;
assign addr[55927]= 1184318708;
assign addr[55928]= 1308821808;
assign addr[55929]= 1426685652;
assign addr[55930]= 1537312353;
assign addr[55931]= 1640140734;
assign addr[55932]= 1734649179;
assign addr[55933]= 1820358275;
assign addr[55934]= 1896833245;
assign addr[55935]= 1963686155;
assign addr[55936]= 2020577882;
assign addr[55937]= 2067219829;
assign addr[55938]= 2103375398;
assign addr[55939]= 2128861181;
assign addr[55940]= 2143547897;
assign addr[55941]= 2147361045;
assign addr[55942]= 2140281282;
assign addr[55943]= 2122344521;
assign addr[55944]= 2093641749;
assign addr[55945]= 2054318569;
assign addr[55946]= 2004574453;
assign addr[55947]= 1944661739;
assign addr[55948]= 1874884346;
assign addr[55949]= 1795596234;
assign addr[55950]= 1707199606;
assign addr[55951]= 1610142873;
assign addr[55952]= 1504918373;
assign addr[55953]= 1392059879;
assign addr[55954]= 1272139887;
assign addr[55955]= 1145766716;
assign addr[55956]= 1013581418;
assign addr[55957]= 876254528;
assign addr[55958]= 734482665;
assign addr[55959]= 588984994;
assign addr[55960]= 440499581;
assign addr[55961]= 289779648;
assign addr[55962]= 137589750;
assign addr[55963]= -15298099;
assign addr[55964]= -168108346;
assign addr[55965]= -320065829;
assign addr[55966]= -470399716;
assign addr[55967]= -618347408;
assign addr[55968]= -763158411;
assign addr[55969]= -904098143;
assign addr[55970]= -1040451659;
assign addr[55971]= -1171527280;
assign addr[55972]= -1296660098;
assign addr[55973]= -1415215352;
assign addr[55974]= -1526591649;
assign addr[55975]= -1630224009;
assign addr[55976]= -1725586737;
assign addr[55977]= -1812196087;
assign addr[55978]= -1889612716;
assign addr[55979]= -1957443913;
assign addr[55980]= -2015345591;
assign addr[55981]= -2063024031;
assign addr[55982]= -2100237377;
assign addr[55983]= -2126796855;
assign addr[55984]= -2142567738;
assign addr[55985]= -2147470025;
assign addr[55986]= -2141478848;
assign addr[55987]= -2124624598;
assign addr[55988]= -2096992772;
assign addr[55989]= -2058723538;
assign addr[55990]= -2010011024;
assign addr[55991]= -1951102334;
assign addr[55992]= -1882296293;
assign addr[55993]= -1803941934;
assign addr[55994]= -1716436725;
assign addr[55995]= -1620224553;
assign addr[55996]= -1515793473;
assign addr[55997]= -1403673233;
assign addr[55998]= -1284432584;
assign addr[55999]= -1158676398;
assign addr[56000]= -1027042599;
assign addr[56001]= -890198924;
assign addr[56002]= -748839539;
assign addr[56003]= -603681519;
assign addr[56004]= -455461206;
assign addr[56005]= -304930476;
assign addr[56006]= -152852926;
assign addr[56007]= 0;
assign addr[56008]= 152852926;
assign addr[56009]= 304930476;
assign addr[56010]= 455461206;
assign addr[56011]= 603681519;
assign addr[56012]= 748839539;
assign addr[56013]= 890198924;
assign addr[56014]= 1027042599;
assign addr[56015]= 1158676398;
assign addr[56016]= 1284432584;
assign addr[56017]= 1403673233;
assign addr[56018]= 1515793473;
assign addr[56019]= 1620224553;
assign addr[56020]= 1716436725;
assign addr[56021]= 1803941934;
assign addr[56022]= 1882296293;
assign addr[56023]= 1951102334;
assign addr[56024]= 2010011024;
assign addr[56025]= 2058723538;
assign addr[56026]= 2096992772;
assign addr[56027]= 2124624598;
assign addr[56028]= 2141478848;
assign addr[56029]= 2147470025;
assign addr[56030]= 2142567738;
assign addr[56031]= 2126796855;
assign addr[56032]= 2100237377;
assign addr[56033]= 2063024031;
assign addr[56034]= 2015345591;
assign addr[56035]= 1957443913;
assign addr[56036]= 1889612716;
assign addr[56037]= 1812196087;
assign addr[56038]= 1725586737;
assign addr[56039]= 1630224009;
assign addr[56040]= 1526591649;
assign addr[56041]= 1415215352;
assign addr[56042]= 1296660098;
assign addr[56043]= 1171527280;
assign addr[56044]= 1040451659;
assign addr[56045]= 904098143;
assign addr[56046]= 763158411;
assign addr[56047]= 618347408;
assign addr[56048]= 470399716;
assign addr[56049]= 320065829;
assign addr[56050]= 168108346;
assign addr[56051]= 15298099;
assign addr[56052]= -137589750;
assign addr[56053]= -289779648;
assign addr[56054]= -440499581;
assign addr[56055]= -588984994;
assign addr[56056]= -734482665;
assign addr[56057]= -876254528;
assign addr[56058]= -1013581418;
assign addr[56059]= -1145766716;
assign addr[56060]= -1272139887;
assign addr[56061]= -1392059879;
assign addr[56062]= -1504918373;
assign addr[56063]= -1610142873;
assign addr[56064]= -1707199606;
assign addr[56065]= -1795596234;
assign addr[56066]= -1874884346;
assign addr[56067]= -1944661739;
assign addr[56068]= -2004574453;
assign addr[56069]= -2054318569;
assign addr[56070]= -2093641749;
assign addr[56071]= -2122344521;
assign addr[56072]= -2140281282;
assign addr[56073]= -2147361045;
assign addr[56074]= -2143547897;
assign addr[56075]= -2128861181;
assign addr[56076]= -2103375398;
assign addr[56077]= -2067219829;
assign addr[56078]= -2020577882;
assign addr[56079]= -1963686155;
assign addr[56080]= -1896833245;
assign addr[56081]= -1820358275;
assign addr[56082]= -1734649179;
assign addr[56083]= -1640140734;
assign addr[56084]= -1537312353;
assign addr[56085]= -1426685652;
assign addr[56086]= -1308821808;
assign addr[56087]= -1184318708;
assign addr[56088]= -1053807919;
assign addr[56089]= -917951481;
assign addr[56090]= -777438554;
assign addr[56091]= -632981917;
assign addr[56092]= -485314355;
assign addr[56093]= -335184940;
assign addr[56094]= -183355234;
assign addr[56095]= -30595422;
assign addr[56096]= 122319591;
assign addr[56097]= 274614114;
assign addr[56098]= 425515602;
assign addr[56099]= 574258580;
assign addr[56100]= 720088517;
assign addr[56101]= 862265664;
assign addr[56102]= 1000068799;
assign addr[56103]= 1132798888;
assign addr[56104]= 1259782632;
assign addr[56105]= 1380375881;
assign addr[56106]= 1493966902;
assign addr[56107]= 1599979481;
assign addr[56108]= 1697875851;
assign addr[56109]= 1787159411;
assign addr[56110]= 1867377253;
assign addr[56111]= 1938122457;
assign addr[56112]= 1999036154;
assign addr[56113]= 2049809346;
assign addr[56114]= 2090184478;
assign addr[56115]= 2119956737;
assign addr[56116]= 2138975100;
assign addr[56117]= 2147143090;
assign addr[56118]= 2144419275;
assign addr[56119]= 2130817471;
assign addr[56120]= 2106406677;
assign addr[56121]= 2071310720;
assign addr[56122]= 2025707632;
assign addr[56123]= 1969828744;
assign addr[56124]= 1903957513;
assign addr[56125]= 1828428082;
assign addr[56126]= 1743623590;
assign addr[56127]= 1649974225;
assign addr[56128]= 1547955041;
assign addr[56129]= 1438083551;
assign addr[56130]= 1320917099;
assign addr[56131]= 1197050035;
assign addr[56132]= 1067110699;
assign addr[56133]= 931758235;
assign addr[56134]= 791679244;
assign addr[56135]= 647584304;
assign addr[56136]= 500204365;
assign addr[56137]= 350287041;
assign addr[56138]= 198592817;
assign addr[56139]= 45891193;
assign addr[56140]= -107043224;
assign addr[56141]= -259434643;
assign addr[56142]= -410510029;
assign addr[56143]= -559503022;
assign addr[56144]= -705657826;
assign addr[56145]= -848233042;
assign addr[56146]= -986505429;
assign addr[56147]= -1119773573;
assign addr[56148]= -1247361445;
assign addr[56149]= -1368621831;
assign addr[56150]= -1482939614;
assign addr[56151]= -1589734894;
assign addr[56152]= -1688465931;
assign addr[56153]= -1778631892;
assign addr[56154]= -1859775393;
assign addr[56155]= -1931484818;
assign addr[56156]= -1993396407;
assign addr[56157]= -2045196100;
assign addr[56158]= -2086621133;
assign addr[56159]= -2117461370;
assign addr[56160]= -2137560369;
assign addr[56161]= -2146816171;
assign addr[56162]= -2145181827;
assign addr[56163]= -2132665626;
assign addr[56164]= -2109331059;
assign addr[56165]= -2075296495;
assign addr[56166]= -2030734582;
assign addr[56167]= -1975871368;
assign addr[56168]= -1910985158;
assign addr[56169]= -1836405100;
assign addr[56170]= -1752509516;
assign addr[56171]= -1659723983;
assign addr[56172]= -1558519173;
assign addr[56173]= -1449408469;
assign addr[56174]= -1332945355;
assign addr[56175]= -1209720613;
assign addr[56176]= -1080359326;
assign addr[56177]= -945517704;
assign addr[56178]= -805879757;
assign addr[56179]= -662153826;
assign addr[56180]= -515068990;
assign addr[56181]= -365371365;
assign addr[56182]= -213820322;
assign addr[56183]= -61184634;
assign addr[56184]= 91761426;
assign addr[56185]= 244242007;
assign addr[56186]= 395483624;
assign addr[56187]= 544719071;
assign addr[56188]= 691191324;
assign addr[56189]= 834157373;
assign addr[56190]= 972891995;
assign addr[56191]= 1106691431;
assign addr[56192]= 1234876957;
assign addr[56193]= 1356798326;
assign addr[56194]= 1471837070;
assign addr[56195]= 1579409630;
assign addr[56196]= 1678970324;
assign addr[56197]= 1770014111;
assign addr[56198]= 1852079154;
assign addr[56199]= 1924749160;
assign addr[56200]= 1987655498;
assign addr[56201]= 2040479063;
assign addr[56202]= 2082951896;
assign addr[56203]= 2114858546;
assign addr[56204]= 2136037160;
assign addr[56205]= 2146380306;
assign addr[56206]= 2145835515;
assign addr[56207]= 2134405552;
assign addr[56208]= 2112148396;
assign addr[56209]= 2079176953;
assign addr[56210]= 2035658475;
assign addr[56211]= 1981813720;
assign addr[56212]= 1917915825;
assign addr[56213]= 1844288924;
assign addr[56214]= 1761306505;
assign addr[56215]= 1669389513;
assign addr[56216]= 1569004214;
assign addr[56217]= 1460659832;
assign addr[56218]= 1344905966;
assign addr[56219]= 1222329801;
assign addr[56220]= 1093553126;
assign addr[56221]= 959229189;
assign addr[56222]= 820039373;
assign addr[56223]= 676689746;
assign addr[56224]= 529907477;
assign addr[56225]= 380437148;
assign addr[56226]= 229036977;
assign addr[56227]= 76474970;
assign addr[56228]= -76474970;
assign addr[56229]= -229036977;
assign addr[56230]= -380437148;
assign addr[56231]= -529907477;
assign addr[56232]= -676689746;
assign addr[56233]= -820039373;
assign addr[56234]= -959229189;
assign addr[56235]= -1093553126;
assign addr[56236]= -1222329801;
assign addr[56237]= -1344905966;
assign addr[56238]= -1460659832;
assign addr[56239]= -1569004214;
assign addr[56240]= -1669389513;
assign addr[56241]= -1761306505;
assign addr[56242]= -1844288924;
assign addr[56243]= -1917915825;
assign addr[56244]= -1981813720;
assign addr[56245]= -2035658475;
assign addr[56246]= -2079176953;
assign addr[56247]= -2112148396;
assign addr[56248]= -2134405552;
assign addr[56249]= -2145835515;
assign addr[56250]= -2146380306;
assign addr[56251]= -2136037160;
assign addr[56252]= -2114858546;
assign addr[56253]= -2082951896;
assign addr[56254]= -2040479063;
assign addr[56255]= -1987655498;
assign addr[56256]= -1924749160;
assign addr[56257]= -1852079154;
assign addr[56258]= -1770014111;
assign addr[56259]= -1678970324;
assign addr[56260]= -1579409630;
assign addr[56261]= -1471837070;
assign addr[56262]= -1356798326;
assign addr[56263]= -1234876957;
assign addr[56264]= -1106691431;
assign addr[56265]= -972891995;
assign addr[56266]= -834157373;
assign addr[56267]= -691191324;
assign addr[56268]= -544719071;
assign addr[56269]= -395483624;
assign addr[56270]= -244242007;
assign addr[56271]= -91761426;
assign addr[56272]= 61184634;
assign addr[56273]= 213820322;
assign addr[56274]= 365371365;
assign addr[56275]= 515068990;
assign addr[56276]= 662153826;
assign addr[56277]= 805879757;
assign addr[56278]= 945517704;
assign addr[56279]= 1080359326;
assign addr[56280]= 1209720613;
assign addr[56281]= 1332945355;
assign addr[56282]= 1449408469;
assign addr[56283]= 1558519173;
assign addr[56284]= 1659723983;
assign addr[56285]= 1752509516;
assign addr[56286]= 1836405100;
assign addr[56287]= 1910985158;
assign addr[56288]= 1975871368;
assign addr[56289]= 2030734582;
assign addr[56290]= 2075296495;
assign addr[56291]= 2109331059;
assign addr[56292]= 2132665626;
assign addr[56293]= 2145181827;
assign addr[56294]= 2146816171;
assign addr[56295]= 2137560369;
assign addr[56296]= 2117461370;
assign addr[56297]= 2086621133;
assign addr[56298]= 2045196100;
assign addr[56299]= 1993396407;
assign addr[56300]= 1931484818;
assign addr[56301]= 1859775393;
assign addr[56302]= 1778631892;
assign addr[56303]= 1688465931;
assign addr[56304]= 1589734894;
assign addr[56305]= 1482939614;
assign addr[56306]= 1368621831;
assign addr[56307]= 1247361445;
assign addr[56308]= 1119773573;
assign addr[56309]= 986505429;
assign addr[56310]= 848233042;
assign addr[56311]= 705657826;
assign addr[56312]= 559503022;
assign addr[56313]= 410510029;
assign addr[56314]= 259434643;
assign addr[56315]= 107043224;
assign addr[56316]= -45891193;
assign addr[56317]= -198592817;
assign addr[56318]= -350287041;
assign addr[56319]= -500204365;
assign addr[56320]= -647584304;
assign addr[56321]= -791679244;
assign addr[56322]= -931758235;
assign addr[56323]= -1067110699;
assign addr[56324]= -1197050035;
assign addr[56325]= -1320917099;
assign addr[56326]= -1438083551;
assign addr[56327]= -1547955041;
assign addr[56328]= -1649974225;
assign addr[56329]= -1743623590;
assign addr[56330]= -1828428082;
assign addr[56331]= -1903957513;
assign addr[56332]= -1969828744;
assign addr[56333]= -2025707632;
assign addr[56334]= -2071310720;
assign addr[56335]= -2106406677;
assign addr[56336]= -2130817471;
assign addr[56337]= -2144419275;
assign addr[56338]= -2147143090;
assign addr[56339]= -2138975100;
assign addr[56340]= -2119956737;
assign addr[56341]= -2090184478;
assign addr[56342]= -2049809346;
assign addr[56343]= -1999036154;
assign addr[56344]= -1938122457;
assign addr[56345]= -1867377253;
assign addr[56346]= -1787159411;
assign addr[56347]= -1697875851;
assign addr[56348]= -1599979481;
assign addr[56349]= -1493966902;
assign addr[56350]= -1380375881;
assign addr[56351]= -1259782632;
assign addr[56352]= -1132798888;
assign addr[56353]= -1000068799;
assign addr[56354]= -862265664;
assign addr[56355]= -720088517;
assign addr[56356]= -574258580;
assign addr[56357]= -425515602;
assign addr[56358]= -274614114;
assign addr[56359]= -122319591;
assign addr[56360]= 30595422;
assign addr[56361]= 183355234;
assign addr[56362]= 335184940;
assign addr[56363]= 485314355;
assign addr[56364]= 632981917;
assign addr[56365]= 777438554;
assign addr[56366]= 917951481;
assign addr[56367]= 1053807919;
assign addr[56368]= 1184318708;
assign addr[56369]= 1308821808;
assign addr[56370]= 1426685652;
assign addr[56371]= 1537312353;
assign addr[56372]= 1640140734;
assign addr[56373]= 1734649179;
assign addr[56374]= 1820358275;
assign addr[56375]= 1896833245;
assign addr[56376]= 1963686155;
assign addr[56377]= 2020577882;
assign addr[56378]= 2067219829;
assign addr[56379]= 2103375398;
assign addr[56380]= 2128861181;
assign addr[56381]= 2143547897;
assign addr[56382]= 2147361045;
assign addr[56383]= 2140281282;
assign addr[56384]= 2122344521;
assign addr[56385]= 2093641749;
assign addr[56386]= 2054318569;
assign addr[56387]= 2004574453;
assign addr[56388]= 1944661739;
assign addr[56389]= 1874884346;
assign addr[56390]= 1795596234;
assign addr[56391]= 1707199606;
assign addr[56392]= 1610142873;
assign addr[56393]= 1504918373;
assign addr[56394]= 1392059879;
assign addr[56395]= 1272139887;
assign addr[56396]= 1145766716;
assign addr[56397]= 1013581418;
assign addr[56398]= 876254528;
assign addr[56399]= 734482665;
assign addr[56400]= 588984994;
assign addr[56401]= 440499581;
assign addr[56402]= 289779648;
assign addr[56403]= 137589750;
assign addr[56404]= -15298099;
assign addr[56405]= -168108346;
assign addr[56406]= -320065829;
assign addr[56407]= -470399716;
assign addr[56408]= -618347408;
assign addr[56409]= -763158411;
assign addr[56410]= -904098143;
assign addr[56411]= -1040451659;
assign addr[56412]= -1171527280;
assign addr[56413]= -1296660098;
assign addr[56414]= -1415215352;
assign addr[56415]= -1526591649;
assign addr[56416]= -1630224009;
assign addr[56417]= -1725586737;
assign addr[56418]= -1812196087;
assign addr[56419]= -1889612716;
assign addr[56420]= -1957443913;
assign addr[56421]= -2015345591;
assign addr[56422]= -2063024031;
assign addr[56423]= -2100237377;
assign addr[56424]= -2126796855;
assign addr[56425]= -2142567738;
assign addr[56426]= -2147470025;
assign addr[56427]= -2141478848;
assign addr[56428]= -2124624598;
assign addr[56429]= -2096992772;
assign addr[56430]= -2058723538;
assign addr[56431]= -2010011024;
assign addr[56432]= -1951102334;
assign addr[56433]= -1882296293;
assign addr[56434]= -1803941934;
assign addr[56435]= -1716436725;
assign addr[56436]= -1620224553;
assign addr[56437]= -1515793473;
assign addr[56438]= -1403673233;
assign addr[56439]= -1284432584;
assign addr[56440]= -1158676398;
assign addr[56441]= -1027042599;
assign addr[56442]= -890198924;
assign addr[56443]= -748839539;
assign addr[56444]= -603681519;
assign addr[56445]= -455461206;
assign addr[56446]= -304930476;
assign addr[56447]= -152852926;
assign addr[56448]= 0;
assign addr[56449]= 152852926;
assign addr[56450]= 304930476;
assign addr[56451]= 455461206;
assign addr[56452]= 603681519;
assign addr[56453]= 748839539;
assign addr[56454]= 890198924;
assign addr[56455]= 1027042599;
assign addr[56456]= 1158676398;
assign addr[56457]= 1284432584;
assign addr[56458]= 1403673233;
assign addr[56459]= 1515793473;
assign addr[56460]= 1620224553;
assign addr[56461]= 1716436725;
assign addr[56462]= 1803941934;
assign addr[56463]= 1882296293;
assign addr[56464]= 1951102334;
assign addr[56465]= 2010011024;
assign addr[56466]= 2058723538;
assign addr[56467]= 2096992772;
assign addr[56468]= 2124624598;
assign addr[56469]= 2141478848;
assign addr[56470]= 2147470025;
assign addr[56471]= 2142567738;
assign addr[56472]= 2126796855;
assign addr[56473]= 2100237377;
assign addr[56474]= 2063024031;
assign addr[56475]= 2015345591;
assign addr[56476]= 1957443913;
assign addr[56477]= 1889612716;
assign addr[56478]= 1812196087;
assign addr[56479]= 1725586737;
assign addr[56480]= 1630224009;
assign addr[56481]= 1526591649;
assign addr[56482]= 1415215352;
assign addr[56483]= 1296660098;
assign addr[56484]= 1171527280;
assign addr[56485]= 1040451659;
assign addr[56486]= 904098143;
assign addr[56487]= 763158411;
assign addr[56488]= 618347408;
assign addr[56489]= 470399716;
assign addr[56490]= 320065829;
assign addr[56491]= 168108346;
assign addr[56492]= 15298099;
assign addr[56493]= -137589750;
assign addr[56494]= -289779648;
assign addr[56495]= -440499581;
assign addr[56496]= -588984994;
assign addr[56497]= -734482665;
assign addr[56498]= -876254528;
assign addr[56499]= -1013581418;
assign addr[56500]= -1145766716;
assign addr[56501]= -1272139887;
assign addr[56502]= -1392059879;
assign addr[56503]= -1504918373;
assign addr[56504]= -1610142873;
assign addr[56505]= -1707199606;
assign addr[56506]= -1795596234;
assign addr[56507]= -1874884346;
assign addr[56508]= -1944661739;
assign addr[56509]= -2004574453;
assign addr[56510]= -2054318569;
assign addr[56511]= -2093641749;
assign addr[56512]= -2122344521;
assign addr[56513]= -2140281282;
assign addr[56514]= -2147361045;
assign addr[56515]= -2143547897;
assign addr[56516]= -2128861181;
assign addr[56517]= -2103375398;
assign addr[56518]= -2067219829;
assign addr[56519]= -2020577882;
assign addr[56520]= -1963686155;
assign addr[56521]= -1896833245;
assign addr[56522]= -1820358275;
assign addr[56523]= -1734649179;
assign addr[56524]= -1640140734;
assign addr[56525]= -1537312353;
assign addr[56526]= -1426685652;
assign addr[56527]= -1308821808;
assign addr[56528]= -1184318708;
assign addr[56529]= -1053807919;
assign addr[56530]= -917951481;
assign addr[56531]= -777438554;
assign addr[56532]= -632981917;
assign addr[56533]= -485314355;
assign addr[56534]= -335184940;
assign addr[56535]= -183355234;
assign addr[56536]= -30595422;
assign addr[56537]= 122319591;
assign addr[56538]= 274614114;
assign addr[56539]= 425515602;
assign addr[56540]= 574258580;
assign addr[56541]= 720088517;
assign addr[56542]= 862265664;
assign addr[56543]= 1000068799;
assign addr[56544]= 1132798888;
assign addr[56545]= 1259782632;
assign addr[56546]= 1380375881;
assign addr[56547]= 1493966902;
assign addr[56548]= 1599979481;
assign addr[56549]= 1697875851;
assign addr[56550]= 1787159411;
assign addr[56551]= 1867377253;
assign addr[56552]= 1938122457;
assign addr[56553]= 1999036154;
assign addr[56554]= 2049809346;
assign addr[56555]= 2090184478;
assign addr[56556]= 2119956737;
assign addr[56557]= 2138975100;
assign addr[56558]= 2147143090;
assign addr[56559]= 2144419275;
assign addr[56560]= 2130817471;
assign addr[56561]= 2106406677;
assign addr[56562]= 2071310720;
assign addr[56563]= 2025707632;
assign addr[56564]= 1969828744;
assign addr[56565]= 1903957513;
assign addr[56566]= 1828428082;
assign addr[56567]= 1743623590;
assign addr[56568]= 1649974225;
assign addr[56569]= 1547955041;
assign addr[56570]= 1438083551;
assign addr[56571]= 1320917099;
assign addr[56572]= 1197050035;
assign addr[56573]= 1067110699;
assign addr[56574]= 931758235;
assign addr[56575]= 791679244;
assign addr[56576]= 647584304;
assign addr[56577]= 500204365;
assign addr[56578]= 350287041;
assign addr[56579]= 198592817;
assign addr[56580]= 45891193;
assign addr[56581]= -107043224;
assign addr[56582]= -259434643;
assign addr[56583]= -410510029;
assign addr[56584]= -559503022;
assign addr[56585]= -705657826;
assign addr[56586]= -848233042;
assign addr[56587]= -986505429;
assign addr[56588]= -1119773573;
assign addr[56589]= -1247361445;
assign addr[56590]= -1368621831;
assign addr[56591]= -1482939614;
assign addr[56592]= -1589734894;
assign addr[56593]= -1688465931;
assign addr[56594]= -1778631892;
assign addr[56595]= -1859775393;
assign addr[56596]= -1931484818;
assign addr[56597]= -1993396407;
assign addr[56598]= -2045196100;
assign addr[56599]= -2086621133;
assign addr[56600]= -2117461370;
assign addr[56601]= -2137560369;
assign addr[56602]= -2146816171;
assign addr[56603]= -2145181827;
assign addr[56604]= -2132665626;
assign addr[56605]= -2109331059;
assign addr[56606]= -2075296495;
assign addr[56607]= -2030734582;
assign addr[56608]= -1975871368;
assign addr[56609]= -1910985158;
assign addr[56610]= -1836405100;
assign addr[56611]= -1752509516;
assign addr[56612]= -1659723983;
assign addr[56613]= -1558519173;
assign addr[56614]= -1449408469;
assign addr[56615]= -1332945355;
assign addr[56616]= -1209720613;
assign addr[56617]= -1080359326;
assign addr[56618]= -945517704;
assign addr[56619]= -805879757;
assign addr[56620]= -662153826;
assign addr[56621]= -515068990;
assign addr[56622]= -365371365;
assign addr[56623]= -213820322;
assign addr[56624]= -61184634;
assign addr[56625]= 91761426;
assign addr[56626]= 244242007;
assign addr[56627]= 395483624;
assign addr[56628]= 544719071;
assign addr[56629]= 691191324;
assign addr[56630]= 834157373;
assign addr[56631]= 972891995;
assign addr[56632]= 1106691431;
assign addr[56633]= 1234876957;
assign addr[56634]= 1356798326;
assign addr[56635]= 1471837070;
assign addr[56636]= 1579409630;
assign addr[56637]= 1678970324;
assign addr[56638]= 1770014111;
assign addr[56639]= 1852079154;
assign addr[56640]= 1924749160;
assign addr[56641]= 1987655498;
assign addr[56642]= 2040479063;
assign addr[56643]= 2082951896;
assign addr[56644]= 2114858546;
assign addr[56645]= 2136037160;
assign addr[56646]= 2146380306;
assign addr[56647]= 2145835515;
assign addr[56648]= 2134405552;
assign addr[56649]= 2112148396;
assign addr[56650]= 2079176953;
assign addr[56651]= 2035658475;
assign addr[56652]= 1981813720;
assign addr[56653]= 1917915825;
assign addr[56654]= 1844288924;
assign addr[56655]= 1761306505;
assign addr[56656]= 1669389513;
assign addr[56657]= 1569004214;
assign addr[56658]= 1460659832;
assign addr[56659]= 1344905966;
assign addr[56660]= 1222329801;
assign addr[56661]= 1093553126;
assign addr[56662]= 959229189;
assign addr[56663]= 820039373;
assign addr[56664]= 676689746;
assign addr[56665]= 529907477;
assign addr[56666]= 380437148;
assign addr[56667]= 229036977;
assign addr[56668]= 76474970;
assign addr[56669]= -76474970;
assign addr[56670]= -229036977;
assign addr[56671]= -380437148;
assign addr[56672]= -529907477;
assign addr[56673]= -676689746;
assign addr[56674]= -820039373;
assign addr[56675]= -959229189;
assign addr[56676]= -1093553126;
assign addr[56677]= -1222329801;
assign addr[56678]= -1344905966;
assign addr[56679]= -1460659832;
assign addr[56680]= -1569004214;
assign addr[56681]= -1669389513;
assign addr[56682]= -1761306505;
assign addr[56683]= -1844288924;
assign addr[56684]= -1917915825;
assign addr[56685]= -1981813720;
assign addr[56686]= -2035658475;
assign addr[56687]= -2079176953;
assign addr[56688]= -2112148396;
assign addr[56689]= -2134405552;
assign addr[56690]= -2145835515;
assign addr[56691]= -2146380306;
assign addr[56692]= -2136037160;
assign addr[56693]= -2114858546;
assign addr[56694]= -2082951896;
assign addr[56695]= -2040479063;
assign addr[56696]= -1987655498;
assign addr[56697]= -1924749160;
assign addr[56698]= -1852079154;
assign addr[56699]= -1770014111;
assign addr[56700]= -1678970324;
assign addr[56701]= -1579409630;
assign addr[56702]= -1471837070;
assign addr[56703]= -1356798326;
assign addr[56704]= -1234876957;
assign addr[56705]= -1106691431;
assign addr[56706]= -972891995;
assign addr[56707]= -834157373;
assign addr[56708]= -691191324;
assign addr[56709]= -544719071;
assign addr[56710]= -395483624;
assign addr[56711]= -244242007;
assign addr[56712]= -91761426;
assign addr[56713]= 61184634;
assign addr[56714]= 213820322;
assign addr[56715]= 365371365;
assign addr[56716]= 515068990;
assign addr[56717]= 662153826;
assign addr[56718]= 805879757;
assign addr[56719]= 945517704;
assign addr[56720]= 1080359326;
assign addr[56721]= 1209720613;
assign addr[56722]= 1332945355;
assign addr[56723]= 1449408469;
assign addr[56724]= 1558519173;
assign addr[56725]= 1659723983;
assign addr[56726]= 1752509516;
assign addr[56727]= 1836405100;
assign addr[56728]= 1910985158;
assign addr[56729]= 1975871368;
assign addr[56730]= 2030734582;
assign addr[56731]= 2075296495;
assign addr[56732]= 2109331059;
assign addr[56733]= 2132665626;
assign addr[56734]= 2145181827;
assign addr[56735]= 2146816171;
assign addr[56736]= 2137560369;
assign addr[56737]= 2117461370;
assign addr[56738]= 2086621133;
assign addr[56739]= 2045196100;
assign addr[56740]= 1993396407;
assign addr[56741]= 1931484818;
assign addr[56742]= 1859775393;
assign addr[56743]= 1778631892;
assign addr[56744]= 1688465931;
assign addr[56745]= 1589734894;
assign addr[56746]= 1482939614;
assign addr[56747]= 1368621831;
assign addr[56748]= 1247361445;
assign addr[56749]= 1119773573;
assign addr[56750]= 986505429;
assign addr[56751]= 848233042;
assign addr[56752]= 705657826;
assign addr[56753]= 559503022;
assign addr[56754]= 410510029;
assign addr[56755]= 259434643;
assign addr[56756]= 107043224;
assign addr[56757]= -45891193;
assign addr[56758]= -198592817;
assign addr[56759]= -350287041;
assign addr[56760]= -500204365;
assign addr[56761]= -647584304;
assign addr[56762]= -791679244;
assign addr[56763]= -931758235;
assign addr[56764]= -1067110699;
assign addr[56765]= -1197050035;
assign addr[56766]= -1320917099;
assign addr[56767]= -1438083551;
assign addr[56768]= -1547955041;
assign addr[56769]= -1649974225;
assign addr[56770]= -1743623590;
assign addr[56771]= -1828428082;
assign addr[56772]= -1903957513;
assign addr[56773]= -1969828744;
assign addr[56774]= -2025707632;
assign addr[56775]= -2071310720;
assign addr[56776]= -2106406677;
assign addr[56777]= -2130817471;
assign addr[56778]= -2144419275;
assign addr[56779]= -2147143090;
assign addr[56780]= -2138975100;
assign addr[56781]= -2119956737;
assign addr[56782]= -2090184478;
assign addr[56783]= -2049809346;
assign addr[56784]= -1999036154;
assign addr[56785]= -1938122457;
assign addr[56786]= -1867377253;
assign addr[56787]= -1787159411;
assign addr[56788]= -1697875851;
assign addr[56789]= -1599979481;
assign addr[56790]= -1493966902;
assign addr[56791]= -1380375881;
assign addr[56792]= -1259782632;
assign addr[56793]= -1132798888;
assign addr[56794]= -1000068799;
assign addr[56795]= -862265664;
assign addr[56796]= -720088517;
assign addr[56797]= -574258580;
assign addr[56798]= -425515602;
assign addr[56799]= -274614114;
assign addr[56800]= -122319591;
assign addr[56801]= 30595422;
assign addr[56802]= 183355234;
assign addr[56803]= 335184940;
assign addr[56804]= 485314355;
assign addr[56805]= 632981917;
assign addr[56806]= 777438554;
assign addr[56807]= 917951481;
assign addr[56808]= 1053807919;
assign addr[56809]= 1184318708;
assign addr[56810]= 1308821808;
assign addr[56811]= 1426685652;
assign addr[56812]= 1537312353;
assign addr[56813]= 1640140734;
assign addr[56814]= 1734649179;
assign addr[56815]= 1820358275;
assign addr[56816]= 1896833245;
assign addr[56817]= 1963686155;
assign addr[56818]= 2020577882;
assign addr[56819]= 2067219829;
assign addr[56820]= 2103375398;
assign addr[56821]= 2128861181;
assign addr[56822]= 2143547897;
assign addr[56823]= 2147361045;
assign addr[56824]= 2140281282;
assign addr[56825]= 2122344521;
assign addr[56826]= 2093641749;
assign addr[56827]= 2054318569;
assign addr[56828]= 2004574453;
assign addr[56829]= 1944661739;
assign addr[56830]= 1874884346;
assign addr[56831]= 1795596234;
assign addr[56832]= 1707199606;
assign addr[56833]= 1610142873;
assign addr[56834]= 1504918373;
assign addr[56835]= 1392059879;
assign addr[56836]= 1272139887;
assign addr[56837]= 1145766716;
assign addr[56838]= 1013581418;
assign addr[56839]= 876254528;
assign addr[56840]= 734482665;
assign addr[56841]= 588984994;
assign addr[56842]= 440499581;
assign addr[56843]= 289779648;
assign addr[56844]= 137589750;
assign addr[56845]= -15298099;
assign addr[56846]= -168108346;
assign addr[56847]= -320065829;
assign addr[56848]= -470399716;
assign addr[56849]= -618347408;
assign addr[56850]= -763158411;
assign addr[56851]= -904098143;
assign addr[56852]= -1040451659;
assign addr[56853]= -1171527280;
assign addr[56854]= -1296660098;
assign addr[56855]= -1415215352;
assign addr[56856]= -1526591649;
assign addr[56857]= -1630224009;
assign addr[56858]= -1725586737;
assign addr[56859]= -1812196087;
assign addr[56860]= -1889612716;
assign addr[56861]= -1957443913;
assign addr[56862]= -2015345591;
assign addr[56863]= -2063024031;
assign addr[56864]= -2100237377;
assign addr[56865]= -2126796855;
assign addr[56866]= -2142567738;
assign addr[56867]= -2147470025;
assign addr[56868]= -2141478848;
assign addr[56869]= -2124624598;
assign addr[56870]= -2096992772;
assign addr[56871]= -2058723538;
assign addr[56872]= -2010011024;
assign addr[56873]= -1951102334;
assign addr[56874]= -1882296293;
assign addr[56875]= -1803941934;
assign addr[56876]= -1716436725;
assign addr[56877]= -1620224553;
assign addr[56878]= -1515793473;
assign addr[56879]= -1403673233;
assign addr[56880]= -1284432584;
assign addr[56881]= -1158676398;
assign addr[56882]= -1027042599;
assign addr[56883]= -890198924;
assign addr[56884]= -748839539;
assign addr[56885]= -603681519;
assign addr[56886]= -455461206;
assign addr[56887]= -304930476;
assign addr[56888]= -152852926;
assign addr[56889]= 0;
assign addr[56890]= 152852926;
assign addr[56891]= 304930476;
assign addr[56892]= 455461206;
assign addr[56893]= 603681519;
assign addr[56894]= 748839539;
assign addr[56895]= 890198924;
assign addr[56896]= 1027042599;
assign addr[56897]= 1158676398;
assign addr[56898]= 1284432584;
assign addr[56899]= 1403673233;
assign addr[56900]= 1515793473;
assign addr[56901]= 1620224553;
assign addr[56902]= 1716436725;
assign addr[56903]= 1803941934;
assign addr[56904]= 1882296293;
assign addr[56905]= 1951102334;
assign addr[56906]= 2010011024;
assign addr[56907]= 2058723538;
assign addr[56908]= 2096992772;
assign addr[56909]= 2124624598;
assign addr[56910]= 2141478848;
assign addr[56911]= 2147470025;
assign addr[56912]= 2142567738;
assign addr[56913]= 2126796855;
assign addr[56914]= 2100237377;
assign addr[56915]= 2063024031;
assign addr[56916]= 2015345591;
assign addr[56917]= 1957443913;
assign addr[56918]= 1889612716;
assign addr[56919]= 1812196087;
assign addr[56920]= 1725586737;
assign addr[56921]= 1630224009;
assign addr[56922]= 1526591649;
assign addr[56923]= 1415215352;
assign addr[56924]= 1296660098;
assign addr[56925]= 1171527280;
assign addr[56926]= 1040451659;
assign addr[56927]= 904098143;
assign addr[56928]= 763158411;
assign addr[56929]= 618347408;
assign addr[56930]= 470399716;
assign addr[56931]= 320065829;
assign addr[56932]= 168108346;
assign addr[56933]= 15298099;
assign addr[56934]= -137589750;
assign addr[56935]= -289779648;
assign addr[56936]= -440499581;
assign addr[56937]= -588984994;
assign addr[56938]= -734482665;
assign addr[56939]= -876254528;
assign addr[56940]= -1013581418;
assign addr[56941]= -1145766716;
assign addr[56942]= -1272139887;
assign addr[56943]= -1392059879;
assign addr[56944]= -1504918373;
assign addr[56945]= -1610142873;
assign addr[56946]= -1707199606;
assign addr[56947]= -1795596234;
assign addr[56948]= -1874884346;
assign addr[56949]= -1944661739;
assign addr[56950]= -2004574453;
assign addr[56951]= -2054318569;
assign addr[56952]= -2093641749;
assign addr[56953]= -2122344521;
assign addr[56954]= -2140281282;
assign addr[56955]= -2147361045;
assign addr[56956]= -2143547897;
assign addr[56957]= -2128861181;
assign addr[56958]= -2103375398;
assign addr[56959]= -2067219829;
assign addr[56960]= -2020577882;
assign addr[56961]= -1963686155;
assign addr[56962]= -1896833245;
assign addr[56963]= -1820358275;
assign addr[56964]= -1734649179;
assign addr[56965]= -1640140734;
assign addr[56966]= -1537312353;
assign addr[56967]= -1426685652;
assign addr[56968]= -1308821808;
assign addr[56969]= -1184318708;
assign addr[56970]= -1053807919;
assign addr[56971]= -917951481;
assign addr[56972]= -777438554;
assign addr[56973]= -632981917;
assign addr[56974]= -485314355;
assign addr[56975]= -335184940;
assign addr[56976]= -183355234;
assign addr[56977]= -30595422;
assign addr[56978]= 122319591;
assign addr[56979]= 274614114;
assign addr[56980]= 425515602;
assign addr[56981]= 574258580;
assign addr[56982]= 720088517;
assign addr[56983]= 862265664;
assign addr[56984]= 1000068799;
assign addr[56985]= 1132798888;
assign addr[56986]= 1259782632;
assign addr[56987]= 1380375881;
assign addr[56988]= 1493966902;
assign addr[56989]= 1599979481;
assign addr[56990]= 1697875851;
assign addr[56991]= 1787159411;
assign addr[56992]= 1867377253;
assign addr[56993]= 1938122457;
assign addr[56994]= 1999036154;
assign addr[56995]= 2049809346;
assign addr[56996]= 2090184478;
assign addr[56997]= 2119956737;
assign addr[56998]= 2138975100;
assign addr[56999]= 2147143090;
assign addr[57000]= 2144419275;
assign addr[57001]= 2130817471;
assign addr[57002]= 2106406677;
assign addr[57003]= 2071310720;
assign addr[57004]= 2025707632;
assign addr[57005]= 1969828744;
assign addr[57006]= 1903957513;
assign addr[57007]= 1828428082;
assign addr[57008]= 1743623590;
assign addr[57009]= 1649974225;
assign addr[57010]= 1547955041;
assign addr[57011]= 1438083551;
assign addr[57012]= 1320917099;
assign addr[57013]= 1197050035;
assign addr[57014]= 1067110699;
assign addr[57015]= 931758235;
assign addr[57016]= 791679244;
assign addr[57017]= 647584304;
assign addr[57018]= 500204365;
assign addr[57019]= 350287041;
assign addr[57020]= 198592817;
assign addr[57021]= 45891193;
assign addr[57022]= -107043224;
assign addr[57023]= -259434643;
assign addr[57024]= -410510029;
assign addr[57025]= -559503022;
assign addr[57026]= -705657826;
assign addr[57027]= -848233042;
assign addr[57028]= -986505429;
assign addr[57029]= -1119773573;
assign addr[57030]= -1247361445;
assign addr[57031]= -1368621831;
assign addr[57032]= -1482939614;
assign addr[57033]= -1589734894;
assign addr[57034]= -1688465931;
assign addr[57035]= -1778631892;
assign addr[57036]= -1859775393;
assign addr[57037]= -1931484818;
assign addr[57038]= -1993396407;
assign addr[57039]= -2045196100;
assign addr[57040]= -2086621133;
assign addr[57041]= -2117461370;
assign addr[57042]= -2137560369;
assign addr[57043]= -2146816171;
assign addr[57044]= -2145181827;
assign addr[57045]= -2132665626;
assign addr[57046]= -2109331059;
assign addr[57047]= -2075296495;
assign addr[57048]= -2030734582;
assign addr[57049]= -1975871368;
assign addr[57050]= -1910985158;
assign addr[57051]= -1836405100;
assign addr[57052]= -1752509516;
assign addr[57053]= -1659723983;
assign addr[57054]= -1558519173;
assign addr[57055]= -1449408469;
assign addr[57056]= -1332945355;
assign addr[57057]= -1209720613;
assign addr[57058]= -1080359326;
assign addr[57059]= -945517704;
assign addr[57060]= -805879757;
assign addr[57061]= -662153826;
assign addr[57062]= -515068990;
assign addr[57063]= -365371365;
assign addr[57064]= -213820322;
assign addr[57065]= -61184634;
assign addr[57066]= 91761426;
assign addr[57067]= 244242007;
assign addr[57068]= 395483624;
assign addr[57069]= 544719071;
assign addr[57070]= 691191324;
assign addr[57071]= 834157373;
assign addr[57072]= 972891995;
assign addr[57073]= 1106691431;
assign addr[57074]= 1234876957;
assign addr[57075]= 1356798326;
assign addr[57076]= 1471837070;
assign addr[57077]= 1579409630;
assign addr[57078]= 1678970324;
assign addr[57079]= 1770014111;
assign addr[57080]= 1852079154;
assign addr[57081]= 1924749160;
assign addr[57082]= 1987655498;
assign addr[57083]= 2040479063;
assign addr[57084]= 2082951896;
assign addr[57085]= 2114858546;
assign addr[57086]= 2136037160;
assign addr[57087]= 2146380306;
assign addr[57088]= 2145835515;
assign addr[57089]= 2134405552;
assign addr[57090]= 2112148396;
assign addr[57091]= 2079176953;
assign addr[57092]= 2035658475;
assign addr[57093]= 1981813720;
assign addr[57094]= 1917915825;
assign addr[57095]= 1844288924;
assign addr[57096]= 1761306505;
assign addr[57097]= 1669389513;
assign addr[57098]= 1569004214;
assign addr[57099]= 1460659832;
assign addr[57100]= 1344905966;
assign addr[57101]= 1222329801;
assign addr[57102]= 1093553126;
assign addr[57103]= 959229189;
assign addr[57104]= 820039373;
assign addr[57105]= 676689746;
assign addr[57106]= 529907477;
assign addr[57107]= 380437148;
assign addr[57108]= 229036977;
assign addr[57109]= 76474970;
assign addr[57110]= -76474970;
assign addr[57111]= -229036977;
assign addr[57112]= -380437148;
assign addr[57113]= -529907477;
assign addr[57114]= -676689746;
assign addr[57115]= -820039373;
assign addr[57116]= -959229189;
assign addr[57117]= -1093553126;
assign addr[57118]= -1222329801;
assign addr[57119]= -1344905966;
assign addr[57120]= -1460659832;
assign addr[57121]= -1569004214;
assign addr[57122]= -1669389513;
assign addr[57123]= -1761306505;
assign addr[57124]= -1844288924;
assign addr[57125]= -1917915825;
assign addr[57126]= -1981813720;
assign addr[57127]= -2035658475;
assign addr[57128]= -2079176953;
assign addr[57129]= -2112148396;
assign addr[57130]= -2134405552;
assign addr[57131]= -2145835515;
assign addr[57132]= -2146380306;
assign addr[57133]= -2136037160;
assign addr[57134]= -2114858546;
assign addr[57135]= -2082951896;
assign addr[57136]= -2040479063;
assign addr[57137]= -1987655498;
assign addr[57138]= -1924749160;
assign addr[57139]= -1852079154;
assign addr[57140]= -1770014111;
assign addr[57141]= -1678970324;
assign addr[57142]= -1579409630;
assign addr[57143]= -1471837070;
assign addr[57144]= -1356798326;
assign addr[57145]= -1234876957;
assign addr[57146]= -1106691431;
assign addr[57147]= -972891995;
assign addr[57148]= -834157373;
assign addr[57149]= -691191324;
assign addr[57150]= -544719071;
assign addr[57151]= -395483624;
assign addr[57152]= -244242007;
assign addr[57153]= -91761426;
assign addr[57154]= 61184634;
assign addr[57155]= 213820322;
assign addr[57156]= 365371365;
assign addr[57157]= 515068990;
assign addr[57158]= 662153826;
assign addr[57159]= 805879757;
assign addr[57160]= 945517704;
assign addr[57161]= 1080359326;
assign addr[57162]= 1209720613;
assign addr[57163]= 1332945355;
assign addr[57164]= 1449408469;
assign addr[57165]= 1558519173;
assign addr[57166]= 1659723983;
assign addr[57167]= 1752509516;
assign addr[57168]= 1836405100;
assign addr[57169]= 1910985158;
assign addr[57170]= 1975871368;
assign addr[57171]= 2030734582;
assign addr[57172]= 2075296495;
assign addr[57173]= 2109331059;
assign addr[57174]= 2132665626;
assign addr[57175]= 2145181827;
assign addr[57176]= 2146816171;
assign addr[57177]= 2137560369;
assign addr[57178]= 2117461370;
assign addr[57179]= 2086621133;
assign addr[57180]= 2045196100;
assign addr[57181]= 1993396407;
assign addr[57182]= 1931484818;
assign addr[57183]= 1859775393;
assign addr[57184]= 1778631892;
assign addr[57185]= 1688465931;
assign addr[57186]= 1589734894;
assign addr[57187]= 1482939614;
assign addr[57188]= 1368621831;
assign addr[57189]= 1247361445;
assign addr[57190]= 1119773573;
assign addr[57191]= 986505429;
assign addr[57192]= 848233042;
assign addr[57193]= 705657826;
assign addr[57194]= 559503022;
assign addr[57195]= 410510029;
assign addr[57196]= 259434643;
assign addr[57197]= 107043224;
assign addr[57198]= -45891193;
assign addr[57199]= -198592817;
assign addr[57200]= -350287041;
assign addr[57201]= -500204365;
assign addr[57202]= -647584304;
assign addr[57203]= -791679244;
assign addr[57204]= -931758235;
assign addr[57205]= -1067110699;
assign addr[57206]= -1197050035;
assign addr[57207]= -1320917099;
assign addr[57208]= -1438083551;
assign addr[57209]= -1547955041;
assign addr[57210]= -1649974225;
assign addr[57211]= -1743623590;
assign addr[57212]= -1828428082;
assign addr[57213]= -1903957513;
assign addr[57214]= -1969828744;
assign addr[57215]= -2025707632;
assign addr[57216]= -2071310720;
assign addr[57217]= -2106406677;
assign addr[57218]= -2130817471;
assign addr[57219]= -2144419275;
assign addr[57220]= -2147143090;
assign addr[57221]= -2138975100;
assign addr[57222]= -2119956737;
assign addr[57223]= -2090184478;
assign addr[57224]= -2049809346;
assign addr[57225]= -1999036154;
assign addr[57226]= -1938122457;
assign addr[57227]= -1867377253;
assign addr[57228]= -1787159411;
assign addr[57229]= -1697875851;
assign addr[57230]= -1599979481;
assign addr[57231]= -1493966902;
assign addr[57232]= -1380375881;
assign addr[57233]= -1259782632;
assign addr[57234]= -1132798888;
assign addr[57235]= -1000068799;
assign addr[57236]= -862265664;
assign addr[57237]= -720088517;
assign addr[57238]= -574258580;
assign addr[57239]= -425515602;
assign addr[57240]= -274614114;
assign addr[57241]= -122319591;
assign addr[57242]= 30595422;
assign addr[57243]= 183355234;
assign addr[57244]= 335184940;
assign addr[57245]= 485314355;
assign addr[57246]= 632981917;
assign addr[57247]= 777438554;
assign addr[57248]= 917951481;
assign addr[57249]= 1053807919;
assign addr[57250]= 1184318708;
assign addr[57251]= 1308821808;
assign addr[57252]= 1426685652;
assign addr[57253]= 1537312353;
assign addr[57254]= 1640140734;
assign addr[57255]= 1734649179;
assign addr[57256]= 1820358275;
assign addr[57257]= 1896833245;
assign addr[57258]= 1963686155;
assign addr[57259]= 2020577882;
assign addr[57260]= 2067219829;
assign addr[57261]= 2103375398;
assign addr[57262]= 2128861181;
assign addr[57263]= 2143547897;
assign addr[57264]= 2147361045;
assign addr[57265]= 2140281282;
assign addr[57266]= 2122344521;
assign addr[57267]= 2093641749;
assign addr[57268]= 2054318569;
assign addr[57269]= 2004574453;
assign addr[57270]= 1944661739;
assign addr[57271]= 1874884346;
assign addr[57272]= 1795596234;
assign addr[57273]= 1707199606;
assign addr[57274]= 1610142873;
assign addr[57275]= 1504918373;
assign addr[57276]= 1392059879;
assign addr[57277]= 1272139887;
assign addr[57278]= 1145766716;
assign addr[57279]= 1013581418;
assign addr[57280]= 876254528;
assign addr[57281]= 734482665;
assign addr[57282]= 588984994;
assign addr[57283]= 440499581;
assign addr[57284]= 289779648;
assign addr[57285]= 137589750;
assign addr[57286]= -15298099;
assign addr[57287]= -168108346;
assign addr[57288]= -320065829;
assign addr[57289]= -470399716;
assign addr[57290]= -618347408;
assign addr[57291]= -763158411;
assign addr[57292]= -904098143;
assign addr[57293]= -1040451659;
assign addr[57294]= -1171527280;
assign addr[57295]= -1296660098;
assign addr[57296]= -1415215352;
assign addr[57297]= -1526591649;
assign addr[57298]= -1630224009;
assign addr[57299]= -1725586737;
assign addr[57300]= -1812196087;
assign addr[57301]= -1889612716;
assign addr[57302]= -1957443913;
assign addr[57303]= -2015345591;
assign addr[57304]= -2063024031;
assign addr[57305]= -2100237377;
assign addr[57306]= -2126796855;
assign addr[57307]= -2142567738;
assign addr[57308]= -2147470025;
assign addr[57309]= -2141478848;
assign addr[57310]= -2124624598;
assign addr[57311]= -2096992772;
assign addr[57312]= -2058723538;
assign addr[57313]= -2010011024;
assign addr[57314]= -1951102334;
assign addr[57315]= -1882296293;
assign addr[57316]= -1803941934;
assign addr[57317]= -1716436725;
assign addr[57318]= -1620224553;
assign addr[57319]= -1515793473;
assign addr[57320]= -1403673233;
assign addr[57321]= -1284432584;
assign addr[57322]= -1158676398;
assign addr[57323]= -1027042599;
assign addr[57324]= -890198924;
assign addr[57325]= -748839539;
assign addr[57326]= -603681519;
assign addr[57327]= -455461206;
assign addr[57328]= -304930476;
assign addr[57329]= -152852926;
assign addr[57330]= 0;
assign addr[57331]= 152852926;
assign addr[57332]= 304930476;
assign addr[57333]= 455461206;
assign addr[57334]= 603681519;
assign addr[57335]= 748839539;
assign addr[57336]= 890198924;
assign addr[57337]= 1027042599;
assign addr[57338]= 1158676398;
assign addr[57339]= 1284432584;
assign addr[57340]= 1403673233;
assign addr[57341]= 1515793473;
assign addr[57342]= 1620224553;
assign addr[57343]= 1716436725;
assign addr[57344]= 1803941934;
assign addr[57345]= 1882296293;
assign addr[57346]= 1951102334;
assign addr[57347]= 2010011024;
assign addr[57348]= 2058723538;
assign addr[57349]= 2096992772;
assign addr[57350]= 2124624598;
assign addr[57351]= 2141478848;
assign addr[57352]= 2147470025;
assign addr[57353]= 2142567738;
assign addr[57354]= 2126796855;
assign addr[57355]= 2100237377;
assign addr[57356]= 2063024031;
assign addr[57357]= 2015345591;
assign addr[57358]= 1957443913;
assign addr[57359]= 1889612716;
assign addr[57360]= 1812196087;
assign addr[57361]= 1725586737;
assign addr[57362]= 1630224009;
assign addr[57363]= 1526591649;
assign addr[57364]= 1415215352;
assign addr[57365]= 1296660098;
assign addr[57366]= 1171527280;
assign addr[57367]= 1040451659;
assign addr[57368]= 904098143;
assign addr[57369]= 763158411;
assign addr[57370]= 618347408;
assign addr[57371]= 470399716;
assign addr[57372]= 320065829;
assign addr[57373]= 168108346;
assign addr[57374]= 15298099;
assign addr[57375]= -137589750;
assign addr[57376]= -289779648;
assign addr[57377]= -440499581;
assign addr[57378]= -588984994;
assign addr[57379]= -734482665;
assign addr[57380]= -876254528;
assign addr[57381]= -1013581418;
assign addr[57382]= -1145766716;
assign addr[57383]= -1272139887;
assign addr[57384]= -1392059879;
assign addr[57385]= -1504918373;
assign addr[57386]= -1610142873;
assign addr[57387]= -1707199606;
assign addr[57388]= -1795596234;
assign addr[57389]= -1874884346;
assign addr[57390]= -1944661739;
assign addr[57391]= -2004574453;
assign addr[57392]= -2054318569;
assign addr[57393]= -2093641749;
assign addr[57394]= -2122344521;
assign addr[57395]= -2140281282;
assign addr[57396]= -2147361045;
assign addr[57397]= -2143547897;
assign addr[57398]= -2128861181;
assign addr[57399]= -2103375398;
assign addr[57400]= -2067219829;
assign addr[57401]= -2020577882;
assign addr[57402]= -1963686155;
assign addr[57403]= -1896833245;
assign addr[57404]= -1820358275;
assign addr[57405]= -1734649179;
assign addr[57406]= -1640140734;
assign addr[57407]= -1537312353;
assign addr[57408]= -1426685652;
assign addr[57409]= -1308821808;
assign addr[57410]= -1184318708;
assign addr[57411]= -1053807919;
assign addr[57412]= -917951481;
assign addr[57413]= -777438554;
assign addr[57414]= -632981917;
assign addr[57415]= -485314355;
assign addr[57416]= -335184940;
assign addr[57417]= -183355234;
assign addr[57418]= -30595422;
assign addr[57419]= 122319591;
assign addr[57420]= 274614114;
assign addr[57421]= 425515602;
assign addr[57422]= 574258580;
assign addr[57423]= 720088517;
assign addr[57424]= 862265664;
assign addr[57425]= 1000068799;
assign addr[57426]= 1132798888;
assign addr[57427]= 1259782632;
assign addr[57428]= 1380375881;
assign addr[57429]= 1493966902;
assign addr[57430]= 1599979481;
assign addr[57431]= 1697875851;
assign addr[57432]= 1787159411;
assign addr[57433]= 1867377253;
assign addr[57434]= 1938122457;
assign addr[57435]= 1999036154;
assign addr[57436]= 2049809346;
assign addr[57437]= 2090184478;
assign addr[57438]= 2119956737;
assign addr[57439]= 2138975100;
assign addr[57440]= 2147143090;
assign addr[57441]= 2144419275;
assign addr[57442]= 2130817471;
assign addr[57443]= 2106406677;
assign addr[57444]= 2071310720;
assign addr[57445]= 2025707632;
assign addr[57446]= 1969828744;
assign addr[57447]= 1903957513;
assign addr[57448]= 1828428082;
assign addr[57449]= 1743623590;
assign addr[57450]= 1649974225;
assign addr[57451]= 1547955041;
assign addr[57452]= 1438083551;
assign addr[57453]= 1320917099;
assign addr[57454]= 1197050035;
assign addr[57455]= 1067110699;
assign addr[57456]= 931758235;
assign addr[57457]= 791679244;
assign addr[57458]= 647584304;
assign addr[57459]= 500204365;
assign addr[57460]= 350287041;
assign addr[57461]= 198592817;
assign addr[57462]= 45891193;
assign addr[57463]= -107043224;
assign addr[57464]= -259434643;
assign addr[57465]= -410510029;
assign addr[57466]= -559503022;
assign addr[57467]= -705657826;
assign addr[57468]= -848233042;
assign addr[57469]= -986505429;
assign addr[57470]= -1119773573;
assign addr[57471]= -1247361445;
assign addr[57472]= -1368621831;
assign addr[57473]= -1482939614;
assign addr[57474]= -1589734894;
assign addr[57475]= -1688465931;
assign addr[57476]= -1778631892;
assign addr[57477]= -1859775393;
assign addr[57478]= -1931484818;
assign addr[57479]= -1993396407;
assign addr[57480]= -2045196100;
assign addr[57481]= -2086621133;
assign addr[57482]= -2117461370;
assign addr[57483]= -2137560369;
assign addr[57484]= -2146816171;
assign addr[57485]= -2145181827;
assign addr[57486]= -2132665626;
assign addr[57487]= -2109331059;
assign addr[57488]= -2075296495;
assign addr[57489]= -2030734582;
assign addr[57490]= -1975871368;
assign addr[57491]= -1910985158;
assign addr[57492]= -1836405100;
assign addr[57493]= -1752509516;
assign addr[57494]= -1659723983;
assign addr[57495]= -1558519173;
assign addr[57496]= -1449408469;
assign addr[57497]= -1332945355;
assign addr[57498]= -1209720613;
assign addr[57499]= -1080359326;
assign addr[57500]= -945517704;
assign addr[57501]= -805879757;
assign addr[57502]= -662153826;
assign addr[57503]= -515068990;
assign addr[57504]= -365371365;
assign addr[57505]= -213820322;
assign addr[57506]= -61184634;
assign addr[57507]= 91761426;
assign addr[57508]= 244242007;
assign addr[57509]= 395483624;
assign addr[57510]= 544719071;
assign addr[57511]= 691191324;
assign addr[57512]= 834157373;
assign addr[57513]= 972891995;
assign addr[57514]= 1106691431;
assign addr[57515]= 1234876957;
assign addr[57516]= 1356798326;
assign addr[57517]= 1471837070;
assign addr[57518]= 1579409630;
assign addr[57519]= 1678970324;
assign addr[57520]= 1770014111;
assign addr[57521]= 1852079154;
assign addr[57522]= 1924749160;
assign addr[57523]= 1987655498;
assign addr[57524]= 2040479063;
assign addr[57525]= 2082951896;
assign addr[57526]= 2114858546;
assign addr[57527]= 2136037160;
assign addr[57528]= 2146380306;
assign addr[57529]= 2145835515;
assign addr[57530]= 2134405552;
assign addr[57531]= 2112148396;
assign addr[57532]= 2079176953;
assign addr[57533]= 2035658475;
assign addr[57534]= 1981813720;
assign addr[57535]= 1917915825;
assign addr[57536]= 1844288924;
assign addr[57537]= 1761306505;
assign addr[57538]= 1669389513;
assign addr[57539]= 1569004214;
assign addr[57540]= 1460659832;
assign addr[57541]= 1344905966;
assign addr[57542]= 1222329801;
assign addr[57543]= 1093553126;
assign addr[57544]= 959229189;
assign addr[57545]= 820039373;
assign addr[57546]= 676689746;
assign addr[57547]= 529907477;
assign addr[57548]= 380437148;
assign addr[57549]= 229036977;
assign addr[57550]= 76474970;
assign addr[57551]= -76474970;
assign addr[57552]= -229036977;
assign addr[57553]= -380437148;
assign addr[57554]= -529907477;
assign addr[57555]= -676689746;
assign addr[57556]= -820039373;
assign addr[57557]= -959229189;
assign addr[57558]= -1093553126;
assign addr[57559]= -1222329801;
assign addr[57560]= -1344905966;
assign addr[57561]= -1460659832;
assign addr[57562]= -1569004214;
assign addr[57563]= -1669389513;
assign addr[57564]= -1761306505;
assign addr[57565]= -1844288924;
assign addr[57566]= -1917915825;
assign addr[57567]= -1981813720;
assign addr[57568]= -2035658475;
assign addr[57569]= -2079176953;
assign addr[57570]= -2112148396;
assign addr[57571]= -2134405552;
assign addr[57572]= -2145835515;
assign addr[57573]= -2146380306;
assign addr[57574]= -2136037160;
assign addr[57575]= -2114858546;
assign addr[57576]= -2082951896;
assign addr[57577]= -2040479063;
assign addr[57578]= -1987655498;
assign addr[57579]= -1924749160;
assign addr[57580]= -1852079154;
assign addr[57581]= -1770014111;
assign addr[57582]= -1678970324;
assign addr[57583]= -1579409630;
assign addr[57584]= -1471837070;
assign addr[57585]= -1356798326;
assign addr[57586]= -1234876957;
assign addr[57587]= -1106691431;
assign addr[57588]= -972891995;
assign addr[57589]= -834157373;
assign addr[57590]= -691191324;
assign addr[57591]= -544719071;
assign addr[57592]= -395483624;
assign addr[57593]= -244242007;
assign addr[57594]= -91761426;
assign addr[57595]= 61184634;
assign addr[57596]= 213820322;
assign addr[57597]= 365371365;
assign addr[57598]= 515068990;
assign addr[57599]= 662153826;
assign addr[57600]= 805879757;
assign addr[57601]= 945517704;
assign addr[57602]= 1080359326;
assign addr[57603]= 1209720613;
assign addr[57604]= 1332945355;
assign addr[57605]= 1449408469;
assign addr[57606]= 1558519173;
assign addr[57607]= 1659723983;
assign addr[57608]= 1752509516;
assign addr[57609]= 1836405100;
assign addr[57610]= 1910985158;
assign addr[57611]= 1975871368;
assign addr[57612]= 2030734582;
assign addr[57613]= 2075296495;
assign addr[57614]= 2109331059;
assign addr[57615]= 2132665626;
assign addr[57616]= 2145181827;
assign addr[57617]= 2146816171;
assign addr[57618]= 2137560369;
assign addr[57619]= 2117461370;
assign addr[57620]= 2086621133;
assign addr[57621]= 2045196100;
assign addr[57622]= 1993396407;
assign addr[57623]= 1931484818;
assign addr[57624]= 1859775393;
assign addr[57625]= 1778631892;
assign addr[57626]= 1688465931;
assign addr[57627]= 1589734894;
assign addr[57628]= 1482939614;
assign addr[57629]= 1368621831;
assign addr[57630]= 1247361445;
assign addr[57631]= 1119773573;
assign addr[57632]= 986505429;
assign addr[57633]= 848233042;
assign addr[57634]= 705657826;
assign addr[57635]= 559503022;
assign addr[57636]= 410510029;
assign addr[57637]= 259434643;
assign addr[57638]= 107043224;
assign addr[57639]= -45891193;
assign addr[57640]= -198592817;
assign addr[57641]= -350287041;
assign addr[57642]= -500204365;
assign addr[57643]= -647584304;
assign addr[57644]= -791679244;
assign addr[57645]= -931758235;
assign addr[57646]= -1067110699;
assign addr[57647]= -1197050035;
assign addr[57648]= -1320917099;
assign addr[57649]= -1438083551;
assign addr[57650]= -1547955041;
assign addr[57651]= -1649974225;
assign addr[57652]= -1743623590;
assign addr[57653]= -1828428082;
assign addr[57654]= -1903957513;
assign addr[57655]= -1969828744;
assign addr[57656]= -2025707632;
assign addr[57657]= -2071310720;
assign addr[57658]= -2106406677;
assign addr[57659]= -2130817471;
assign addr[57660]= -2144419275;
assign addr[57661]= -2147143090;
assign addr[57662]= -2138975100;
assign addr[57663]= -2119956737;
assign addr[57664]= -2090184478;
assign addr[57665]= -2049809346;
assign addr[57666]= -1999036154;
assign addr[57667]= -1938122457;
assign addr[57668]= -1867377253;
assign addr[57669]= -1787159411;
assign addr[57670]= -1697875851;
assign addr[57671]= -1599979481;
assign addr[57672]= -1493966902;
assign addr[57673]= -1380375881;
assign addr[57674]= -1259782632;
assign addr[57675]= -1132798888;
assign addr[57676]= -1000068799;
assign addr[57677]= -862265664;
assign addr[57678]= -720088517;
assign addr[57679]= -574258580;
assign addr[57680]= -425515602;
assign addr[57681]= -274614114;
assign addr[57682]= -122319591;
assign addr[57683]= 30595422;
assign addr[57684]= 183355234;
assign addr[57685]= 335184940;
assign addr[57686]= 485314355;
assign addr[57687]= 632981917;
assign addr[57688]= 777438554;
assign addr[57689]= 917951481;
assign addr[57690]= 1053807919;
assign addr[57691]= 1184318708;
assign addr[57692]= 1308821808;
assign addr[57693]= 1426685652;
assign addr[57694]= 1537312353;
assign addr[57695]= 1640140734;
assign addr[57696]= 1734649179;
assign addr[57697]= 1820358275;
assign addr[57698]= 1896833245;
assign addr[57699]= 1963686155;
assign addr[57700]= 2020577882;
assign addr[57701]= 2067219829;
assign addr[57702]= 2103375398;
assign addr[57703]= 2128861181;
assign addr[57704]= 2143547897;
assign addr[57705]= 2147361045;
assign addr[57706]= 2140281282;
assign addr[57707]= 2122344521;
assign addr[57708]= 2093641749;
assign addr[57709]= 2054318569;
assign addr[57710]= 2004574453;
assign addr[57711]= 1944661739;
assign addr[57712]= 1874884346;
assign addr[57713]= 1795596234;
assign addr[57714]= 1707199606;
assign addr[57715]= 1610142873;
assign addr[57716]= 1504918373;
assign addr[57717]= 1392059879;
assign addr[57718]= 1272139887;
assign addr[57719]= 1145766716;
assign addr[57720]= 1013581418;
assign addr[57721]= 876254528;
assign addr[57722]= 734482665;
assign addr[57723]= 588984994;
assign addr[57724]= 440499581;
assign addr[57725]= 289779648;
assign addr[57726]= 137589750;
assign addr[57727]= -15298099;
assign addr[57728]= -168108346;
assign addr[57729]= -320065829;
assign addr[57730]= -470399716;
assign addr[57731]= -618347408;
assign addr[57732]= -763158411;
assign addr[57733]= -904098143;
assign addr[57734]= -1040451659;
assign addr[57735]= -1171527280;
assign addr[57736]= -1296660098;
assign addr[57737]= -1415215352;
assign addr[57738]= -1526591649;
assign addr[57739]= -1630224009;
assign addr[57740]= -1725586737;
assign addr[57741]= -1812196087;
assign addr[57742]= -1889612716;
assign addr[57743]= -1957443913;
assign addr[57744]= -2015345591;
assign addr[57745]= -2063024031;
assign addr[57746]= -2100237377;
assign addr[57747]= -2126796855;
assign addr[57748]= -2142567738;
assign addr[57749]= -2147470025;
assign addr[57750]= -2141478848;
assign addr[57751]= -2124624598;
assign addr[57752]= -2096992772;
assign addr[57753]= -2058723538;
assign addr[57754]= -2010011024;
assign addr[57755]= -1951102334;
assign addr[57756]= -1882296293;
assign addr[57757]= -1803941934;
assign addr[57758]= -1716436725;
assign addr[57759]= -1620224553;
assign addr[57760]= -1515793473;
assign addr[57761]= -1403673233;
assign addr[57762]= -1284432584;
assign addr[57763]= -1158676398;
assign addr[57764]= -1027042599;
assign addr[57765]= -890198924;
assign addr[57766]= -748839539;
assign addr[57767]= -603681519;
assign addr[57768]= -455461206;
assign addr[57769]= -304930476;
assign addr[57770]= -152852926;
assign addr[57771]= 0;
assign addr[57772]= 152852926;
assign addr[57773]= 304930476;
assign addr[57774]= 455461206;
assign addr[57775]= 603681519;
assign addr[57776]= 748839539;
assign addr[57777]= 890198924;
assign addr[57778]= 1027042599;
assign addr[57779]= 1158676398;
assign addr[57780]= 1284432584;
assign addr[57781]= 1403673233;
assign addr[57782]= 1515793473;
assign addr[57783]= 1620224553;
assign addr[57784]= 1716436725;
assign addr[57785]= 1803941934;
assign addr[57786]= 1882296293;
assign addr[57787]= 1951102334;
assign addr[57788]= 2010011024;
assign addr[57789]= 2058723538;
assign addr[57790]= 2096992772;
assign addr[57791]= 2124624598;
assign addr[57792]= 2141478848;
assign addr[57793]= 2147470025;
assign addr[57794]= 2142567738;
assign addr[57795]= 2126796855;
assign addr[57796]= 2100237377;
assign addr[57797]= 2063024031;
assign addr[57798]= 2015345591;
assign addr[57799]= 1957443913;
assign addr[57800]= 1889612716;
assign addr[57801]= 1812196087;
assign addr[57802]= 1725586737;
assign addr[57803]= 1630224009;
assign addr[57804]= 1526591649;
assign addr[57805]= 1415215352;
assign addr[57806]= 1296660098;
assign addr[57807]= 1171527280;
assign addr[57808]= 1040451659;
assign addr[57809]= 904098143;
assign addr[57810]= 763158411;
assign addr[57811]= 618347408;
assign addr[57812]= 470399716;
assign addr[57813]= 320065829;
assign addr[57814]= 168108346;
assign addr[57815]= 15298099;
assign addr[57816]= -137589750;
assign addr[57817]= -289779648;
assign addr[57818]= -440499581;
assign addr[57819]= -588984994;
assign addr[57820]= -734482665;
assign addr[57821]= -876254528;
assign addr[57822]= -1013581418;
assign addr[57823]= -1145766716;
assign addr[57824]= -1272139887;
assign addr[57825]= -1392059879;
assign addr[57826]= -1504918373;
assign addr[57827]= -1610142873;
assign addr[57828]= -1707199606;
assign addr[57829]= -1795596234;
assign addr[57830]= -1874884346;
assign addr[57831]= -1944661739;
assign addr[57832]= -2004574453;
assign addr[57833]= -2054318569;
assign addr[57834]= -2093641749;
assign addr[57835]= -2122344521;
assign addr[57836]= -2140281282;
assign addr[57837]= -2147361045;
assign addr[57838]= -2143547897;
assign addr[57839]= -2128861181;
assign addr[57840]= -2103375398;
assign addr[57841]= -2067219829;
assign addr[57842]= -2020577882;
assign addr[57843]= -1963686155;
assign addr[57844]= -1896833245;
assign addr[57845]= -1820358275;
assign addr[57846]= -1734649179;
assign addr[57847]= -1640140734;
assign addr[57848]= -1537312353;
assign addr[57849]= -1426685652;
assign addr[57850]= -1308821808;
assign addr[57851]= -1184318708;
assign addr[57852]= -1053807919;
assign addr[57853]= -917951481;
assign addr[57854]= -777438554;
assign addr[57855]= -632981917;
assign addr[57856]= -485314355;
assign addr[57857]= -335184940;
assign addr[57858]= -183355234;
assign addr[57859]= -30595422;
assign addr[57860]= 122319591;
assign addr[57861]= 274614114;
assign addr[57862]= 425515602;
assign addr[57863]= 574258580;
assign addr[57864]= 720088517;
assign addr[57865]= 862265664;
assign addr[57866]= 1000068799;
assign addr[57867]= 1132798888;
assign addr[57868]= 1259782632;
assign addr[57869]= 1380375881;
assign addr[57870]= 1493966902;
assign addr[57871]= 1599979481;
assign addr[57872]= 1697875851;
assign addr[57873]= 1787159411;
assign addr[57874]= 1867377253;
assign addr[57875]= 1938122457;
assign addr[57876]= 1999036154;
assign addr[57877]= 2049809346;
assign addr[57878]= 2090184478;
assign addr[57879]= 2119956737;
assign addr[57880]= 2138975100;
assign addr[57881]= 2147143090;
assign addr[57882]= 2144419275;
assign addr[57883]= 2130817471;
assign addr[57884]= 2106406677;
assign addr[57885]= 2071310720;
assign addr[57886]= 2025707632;
assign addr[57887]= 1969828744;
assign addr[57888]= 1903957513;
assign addr[57889]= 1828428082;
assign addr[57890]= 1743623590;
assign addr[57891]= 1649974225;
assign addr[57892]= 1547955041;
assign addr[57893]= 1438083551;
assign addr[57894]= 1320917099;
assign addr[57895]= 1197050035;
assign addr[57896]= 1067110699;
assign addr[57897]= 931758235;
assign addr[57898]= 791679244;
assign addr[57899]= 647584304;
assign addr[57900]= 500204365;
assign addr[57901]= 350287041;
assign addr[57902]= 198592817;
assign addr[57903]= 45891193;
assign addr[57904]= -107043224;
assign addr[57905]= -259434643;
assign addr[57906]= -410510029;
assign addr[57907]= -559503022;
assign addr[57908]= -705657826;
assign addr[57909]= -848233042;
assign addr[57910]= -986505429;
assign addr[57911]= -1119773573;
assign addr[57912]= -1247361445;
assign addr[57913]= -1368621831;
assign addr[57914]= -1482939614;
assign addr[57915]= -1589734894;
assign addr[57916]= -1688465931;
assign addr[57917]= -1778631892;
assign addr[57918]= -1859775393;
assign addr[57919]= -1931484818;
assign addr[57920]= -1993396407;
assign addr[57921]= -2045196100;
assign addr[57922]= -2086621133;
assign addr[57923]= -2117461370;
assign addr[57924]= -2137560369;
assign addr[57925]= -2146816171;
assign addr[57926]= -2145181827;
assign addr[57927]= -2132665626;
assign addr[57928]= -2109331059;
assign addr[57929]= -2075296495;
assign addr[57930]= -2030734582;
assign addr[57931]= -1975871368;
assign addr[57932]= -1910985158;
assign addr[57933]= -1836405100;
assign addr[57934]= -1752509516;
assign addr[57935]= -1659723983;
assign addr[57936]= -1558519173;
assign addr[57937]= -1449408469;
assign addr[57938]= -1332945355;
assign addr[57939]= -1209720613;
assign addr[57940]= -1080359326;
assign addr[57941]= -945517704;
assign addr[57942]= -805879757;
assign addr[57943]= -662153826;
assign addr[57944]= -515068990;
assign addr[57945]= -365371365;
assign addr[57946]= -213820322;
assign addr[57947]= -61184634;
assign addr[57948]= 91761426;
assign addr[57949]= 244242007;
assign addr[57950]= 395483624;
assign addr[57951]= 544719071;
assign addr[57952]= 691191324;
assign addr[57953]= 834157373;
assign addr[57954]= 972891995;
assign addr[57955]= 1106691431;
assign addr[57956]= 1234876957;
assign addr[57957]= 1356798326;
assign addr[57958]= 1471837070;
assign addr[57959]= 1579409630;
assign addr[57960]= 1678970324;
assign addr[57961]= 1770014111;
assign addr[57962]= 1852079154;
assign addr[57963]= 1924749160;
assign addr[57964]= 1987655498;
assign addr[57965]= 2040479063;
assign addr[57966]= 2082951896;
assign addr[57967]= 2114858546;
assign addr[57968]= 2136037160;
assign addr[57969]= 2146380306;
assign addr[57970]= 2145835515;
assign addr[57971]= 2134405552;
assign addr[57972]= 2112148396;
assign addr[57973]= 2079176953;
assign addr[57974]= 2035658475;
assign addr[57975]= 1981813720;
assign addr[57976]= 1917915825;
assign addr[57977]= 1844288924;
assign addr[57978]= 1761306505;
assign addr[57979]= 1669389513;
assign addr[57980]= 1569004214;
assign addr[57981]= 1460659832;
assign addr[57982]= 1344905966;
assign addr[57983]= 1222329801;
assign addr[57984]= 1093553126;
assign addr[57985]= 959229189;
assign addr[57986]= 820039373;
assign addr[57987]= 676689746;
assign addr[57988]= 529907477;
assign addr[57989]= 380437148;
assign addr[57990]= 229036977;
assign addr[57991]= 76474970;
assign addr[57992]= -76474970;
assign addr[57993]= -229036977;
assign addr[57994]= -380437148;
assign addr[57995]= -529907477;
assign addr[57996]= -676689746;
assign addr[57997]= -820039373;
assign addr[57998]= -959229189;
assign addr[57999]= -1093553126;
assign addr[58000]= -1222329801;
assign addr[58001]= -1344905966;
assign addr[58002]= -1460659832;
assign addr[58003]= -1569004214;
assign addr[58004]= -1669389513;
assign addr[58005]= -1761306505;
assign addr[58006]= -1844288924;
assign addr[58007]= -1917915825;
assign addr[58008]= -1981813720;
assign addr[58009]= -2035658475;
assign addr[58010]= -2079176953;
assign addr[58011]= -2112148396;
assign addr[58012]= -2134405552;
assign addr[58013]= -2145835515;
assign addr[58014]= -2146380306;
assign addr[58015]= -2136037160;
assign addr[58016]= -2114858546;
assign addr[58017]= -2082951896;
assign addr[58018]= -2040479063;
assign addr[58019]= -1987655498;
assign addr[58020]= -1924749160;
assign addr[58021]= -1852079154;
assign addr[58022]= -1770014111;
assign addr[58023]= -1678970324;
assign addr[58024]= -1579409630;
assign addr[58025]= -1471837070;
assign addr[58026]= -1356798326;
assign addr[58027]= -1234876957;
assign addr[58028]= -1106691431;
assign addr[58029]= -972891995;
assign addr[58030]= -834157373;
assign addr[58031]= -691191324;
assign addr[58032]= -544719071;
assign addr[58033]= -395483624;
assign addr[58034]= -244242007;
assign addr[58035]= -91761426;
assign addr[58036]= 61184634;
assign addr[58037]= 213820322;
assign addr[58038]= 365371365;
assign addr[58039]= 515068990;
assign addr[58040]= 662153826;
assign addr[58041]= 805879757;
assign addr[58042]= 945517704;
assign addr[58043]= 1080359326;
assign addr[58044]= 1209720613;
assign addr[58045]= 1332945355;
assign addr[58046]= 1449408469;
assign addr[58047]= 1558519173;
assign addr[58048]= 1659723983;
assign addr[58049]= 1752509516;
assign addr[58050]= 1836405100;
assign addr[58051]= 1910985158;
assign addr[58052]= 1975871368;
assign addr[58053]= 2030734582;
assign addr[58054]= 2075296495;
assign addr[58055]= 2109331059;
assign addr[58056]= 2132665626;
assign addr[58057]= 2145181827;
assign addr[58058]= 2146816171;
assign addr[58059]= 2137560369;
assign addr[58060]= 2117461370;
assign addr[58061]= 2086621133;
assign addr[58062]= 2045196100;
assign addr[58063]= 1993396407;
assign addr[58064]= 1931484818;
assign addr[58065]= 1859775393;
assign addr[58066]= 1778631892;
assign addr[58067]= 1688465931;
assign addr[58068]= 1589734894;
assign addr[58069]= 1482939614;
assign addr[58070]= 1368621831;
assign addr[58071]= 1247361445;
assign addr[58072]= 1119773573;
assign addr[58073]= 986505429;
assign addr[58074]= 848233042;
assign addr[58075]= 705657826;
assign addr[58076]= 559503022;
assign addr[58077]= 410510029;
assign addr[58078]= 259434643;
assign addr[58079]= 107043224;
assign addr[58080]= -45891193;
assign addr[58081]= -198592817;
assign addr[58082]= -350287041;
assign addr[58083]= -500204365;
assign addr[58084]= -647584304;
assign addr[58085]= -791679244;
assign addr[58086]= -931758235;
assign addr[58087]= -1067110699;
assign addr[58088]= -1197050035;
assign addr[58089]= -1320917099;
assign addr[58090]= -1438083551;
assign addr[58091]= -1547955041;
assign addr[58092]= -1649974225;
assign addr[58093]= -1743623590;
assign addr[58094]= -1828428082;
assign addr[58095]= -1903957513;
assign addr[58096]= -1969828744;
assign addr[58097]= -2025707632;
assign addr[58098]= -2071310720;
assign addr[58099]= -2106406677;
assign addr[58100]= -2130817471;
assign addr[58101]= -2144419275;
assign addr[58102]= -2147143090;
assign addr[58103]= -2138975100;
assign addr[58104]= -2119956737;
assign addr[58105]= -2090184478;
assign addr[58106]= -2049809346;
assign addr[58107]= -1999036154;
assign addr[58108]= -1938122457;
assign addr[58109]= -1867377253;
assign addr[58110]= -1787159411;
assign addr[58111]= -1697875851;
assign addr[58112]= -1599979481;
assign addr[58113]= -1493966902;
assign addr[58114]= -1380375881;
assign addr[58115]= -1259782632;
assign addr[58116]= -1132798888;
assign addr[58117]= -1000068799;
assign addr[58118]= -862265664;
assign addr[58119]= -720088517;
assign addr[58120]= -574258580;
assign addr[58121]= -425515602;
assign addr[58122]= -274614114;
assign addr[58123]= -122319591;
assign addr[58124]= 30595422;
assign addr[58125]= 183355234;
assign addr[58126]= 335184940;
assign addr[58127]= 485314355;
assign addr[58128]= 632981917;
assign addr[58129]= 777438554;
assign addr[58130]= 917951481;
assign addr[58131]= 1053807919;
assign addr[58132]= 1184318708;
assign addr[58133]= 1308821808;
assign addr[58134]= 1426685652;
assign addr[58135]= 1537312353;
assign addr[58136]= 1640140734;
assign addr[58137]= 1734649179;
assign addr[58138]= 1820358275;
assign addr[58139]= 1896833245;
assign addr[58140]= 1963686155;
assign addr[58141]= 2020577882;
assign addr[58142]= 2067219829;
assign addr[58143]= 2103375398;
assign addr[58144]= 2128861181;
assign addr[58145]= 2143547897;
assign addr[58146]= 2147361045;
assign addr[58147]= 2140281282;
assign addr[58148]= 2122344521;
assign addr[58149]= 2093641749;
assign addr[58150]= 2054318569;
assign addr[58151]= 2004574453;
assign addr[58152]= 1944661739;
assign addr[58153]= 1874884346;
assign addr[58154]= 1795596234;
assign addr[58155]= 1707199606;
assign addr[58156]= 1610142873;
assign addr[58157]= 1504918373;
assign addr[58158]= 1392059879;
assign addr[58159]= 1272139887;
assign addr[58160]= 1145766716;
assign addr[58161]= 1013581418;
assign addr[58162]= 876254528;
assign addr[58163]= 734482665;
assign addr[58164]= 588984994;
assign addr[58165]= 440499581;
assign addr[58166]= 289779648;
assign addr[58167]= 137589750;
assign addr[58168]= -15298099;
assign addr[58169]= -168108346;
assign addr[58170]= -320065829;
assign addr[58171]= -470399716;
assign addr[58172]= -618347408;
assign addr[58173]= -763158411;
assign addr[58174]= -904098143;
assign addr[58175]= -1040451659;
assign addr[58176]= -1171527280;
assign addr[58177]= -1296660098;
assign addr[58178]= -1415215352;
assign addr[58179]= -1526591649;
assign addr[58180]= -1630224009;
assign addr[58181]= -1725586737;
assign addr[58182]= -1812196087;
assign addr[58183]= -1889612716;
assign addr[58184]= -1957443913;
assign addr[58185]= -2015345591;
assign addr[58186]= -2063024031;
assign addr[58187]= -2100237377;
assign addr[58188]= -2126796855;
assign addr[58189]= -2142567738;
assign addr[58190]= -2147470025;
assign addr[58191]= -2141478848;
assign addr[58192]= -2124624598;
assign addr[58193]= -2096992772;
assign addr[58194]= -2058723538;
assign addr[58195]= -2010011024;
assign addr[58196]= -1951102334;
assign addr[58197]= -1882296293;
assign addr[58198]= -1803941934;
assign addr[58199]= -1716436725;
assign addr[58200]= -1620224553;
assign addr[58201]= -1515793473;
assign addr[58202]= -1403673233;
assign addr[58203]= -1284432584;
assign addr[58204]= -1158676398;
assign addr[58205]= -1027042599;
assign addr[58206]= -890198924;
assign addr[58207]= -748839539;
assign addr[58208]= -603681519;
assign addr[58209]= -455461206;
assign addr[58210]= -304930476;
assign addr[58211]= -152852926;
assign addr[58212]= 0;
assign addr[58213]= 152852926;
assign addr[58214]= 304930476;
assign addr[58215]= 455461206;
assign addr[58216]= 603681519;
assign addr[58217]= 748839539;
assign addr[58218]= 890198924;
assign addr[58219]= 1027042599;
assign addr[58220]= 1158676398;
assign addr[58221]= 1284432584;
assign addr[58222]= 1403673233;
assign addr[58223]= 1515793473;
assign addr[58224]= 1620224553;
assign addr[58225]= 1716436725;
assign addr[58226]= 1803941934;
assign addr[58227]= 1882296293;
assign addr[58228]= 1951102334;
assign addr[58229]= 2010011024;
assign addr[58230]= 2058723538;
assign addr[58231]= 2096992772;
assign addr[58232]= 2124624598;
assign addr[58233]= 2141478848;
assign addr[58234]= 2147470025;
assign addr[58235]= 2142567738;
assign addr[58236]= 2126796855;
assign addr[58237]= 2100237377;
assign addr[58238]= 2063024031;
assign addr[58239]= 2015345591;
assign addr[58240]= 1957443913;
assign addr[58241]= 1889612716;
assign addr[58242]= 1812196087;
assign addr[58243]= 1725586737;
assign addr[58244]= 1630224009;
assign addr[58245]= 1526591649;
assign addr[58246]= 1415215352;
assign addr[58247]= 1296660098;
assign addr[58248]= 1171527280;
assign addr[58249]= 1040451659;
assign addr[58250]= 904098143;
assign addr[58251]= 763158411;
assign addr[58252]= 618347408;
assign addr[58253]= 470399716;
assign addr[58254]= 320065829;
assign addr[58255]= 168108346;
assign addr[58256]= 15298099;
assign addr[58257]= -137589750;
assign addr[58258]= -289779648;
assign addr[58259]= -440499581;
assign addr[58260]= -588984994;
assign addr[58261]= -734482665;
assign addr[58262]= -876254528;
assign addr[58263]= -1013581418;
assign addr[58264]= -1145766716;
assign addr[58265]= -1272139887;
assign addr[58266]= -1392059879;
assign addr[58267]= -1504918373;
assign addr[58268]= -1610142873;
assign addr[58269]= -1707199606;
assign addr[58270]= -1795596234;
assign addr[58271]= -1874884346;
assign addr[58272]= -1944661739;
assign addr[58273]= -2004574453;
assign addr[58274]= -2054318569;
assign addr[58275]= -2093641749;
assign addr[58276]= -2122344521;
assign addr[58277]= -2140281282;
assign addr[58278]= -2147361045;
assign addr[58279]= -2143547897;
assign addr[58280]= -2128861181;
assign addr[58281]= -2103375398;
assign addr[58282]= -2067219829;
assign addr[58283]= -2020577882;
assign addr[58284]= -1963686155;
assign addr[58285]= -1896833245;
assign addr[58286]= -1820358275;
assign addr[58287]= -1734649179;
assign addr[58288]= -1640140734;
assign addr[58289]= -1537312353;
assign addr[58290]= -1426685652;
assign addr[58291]= -1308821808;
assign addr[58292]= -1184318708;
assign addr[58293]= -1053807919;
assign addr[58294]= -917951481;
assign addr[58295]= -777438554;
assign addr[58296]= -632981917;
assign addr[58297]= -485314355;
assign addr[58298]= -335184940;
assign addr[58299]= -183355234;
assign addr[58300]= -30595422;
assign addr[58301]= 122319591;
assign addr[58302]= 274614114;
assign addr[58303]= 425515602;
assign addr[58304]= 574258580;
assign addr[58305]= 720088517;
assign addr[58306]= 862265664;
assign addr[58307]= 1000068799;
assign addr[58308]= 1132798888;
assign addr[58309]= 1259782632;
assign addr[58310]= 1380375881;
assign addr[58311]= 1493966902;
assign addr[58312]= 1599979481;
assign addr[58313]= 1697875851;
assign addr[58314]= 1787159411;
assign addr[58315]= 1867377253;
assign addr[58316]= 1938122457;
assign addr[58317]= 1999036154;
assign addr[58318]= 2049809346;
assign addr[58319]= 2090184478;
assign addr[58320]= 2119956737;
assign addr[58321]= 2138975100;
assign addr[58322]= 2147143090;
assign addr[58323]= 2144419275;
assign addr[58324]= 2130817471;
assign addr[58325]= 2106406677;
assign addr[58326]= 2071310720;
assign addr[58327]= 2025707632;
assign addr[58328]= 1969828744;
assign addr[58329]= 1903957513;
assign addr[58330]= 1828428082;
assign addr[58331]= 1743623590;
assign addr[58332]= 1649974225;
assign addr[58333]= 1547955041;
assign addr[58334]= 1438083551;
assign addr[58335]= 1320917099;
assign addr[58336]= 1197050035;
assign addr[58337]= 1067110699;
assign addr[58338]= 931758235;
assign addr[58339]= 791679244;
assign addr[58340]= 647584304;
assign addr[58341]= 500204365;
assign addr[58342]= 350287041;
assign addr[58343]= 198592817;
assign addr[58344]= 45891193;
assign addr[58345]= -107043224;
assign addr[58346]= -259434643;
assign addr[58347]= -410510029;
assign addr[58348]= -559503022;
assign addr[58349]= -705657826;
assign addr[58350]= -848233042;
assign addr[58351]= -986505429;
assign addr[58352]= -1119773573;
assign addr[58353]= -1247361445;
assign addr[58354]= -1368621831;
assign addr[58355]= -1482939614;
assign addr[58356]= -1589734894;
assign addr[58357]= -1688465931;
assign addr[58358]= -1778631892;
assign addr[58359]= -1859775393;
assign addr[58360]= -1931484818;
assign addr[58361]= -1993396407;
assign addr[58362]= -2045196100;
assign addr[58363]= -2086621133;
assign addr[58364]= -2117461370;
assign addr[58365]= -2137560369;
assign addr[58366]= -2146816171;
assign addr[58367]= -2145181827;
assign addr[58368]= -2132665626;
assign addr[58369]= -2109331059;
assign addr[58370]= -2075296495;
assign addr[58371]= -2030734582;
assign addr[58372]= -1975871368;
assign addr[58373]= -1910985158;
assign addr[58374]= -1836405100;
assign addr[58375]= -1752509516;
assign addr[58376]= -1659723983;
assign addr[58377]= -1558519173;
assign addr[58378]= -1449408469;
assign addr[58379]= -1332945355;
assign addr[58380]= -1209720613;
assign addr[58381]= -1080359326;
assign addr[58382]= -945517704;
assign addr[58383]= -805879757;
assign addr[58384]= -662153826;
assign addr[58385]= -515068990;
assign addr[58386]= -365371365;
assign addr[58387]= -213820322;
assign addr[58388]= -61184634;
assign addr[58389]= 91761426;
assign addr[58390]= 244242007;
assign addr[58391]= 395483624;
assign addr[58392]= 544719071;
assign addr[58393]= 691191324;
assign addr[58394]= 834157373;
assign addr[58395]= 972891995;
assign addr[58396]= 1106691431;
assign addr[58397]= 1234876957;
assign addr[58398]= 1356798326;
assign addr[58399]= 1471837070;
assign addr[58400]= 1579409630;
assign addr[58401]= 1678970324;
assign addr[58402]= 1770014111;
assign addr[58403]= 1852079154;
assign addr[58404]= 1924749160;
assign addr[58405]= 1987655498;
assign addr[58406]= 2040479063;
assign addr[58407]= 2082951896;
assign addr[58408]= 2114858546;
assign addr[58409]= 2136037160;
assign addr[58410]= 2146380306;
assign addr[58411]= 2145835515;
assign addr[58412]= 2134405552;
assign addr[58413]= 2112148396;
assign addr[58414]= 2079176953;
assign addr[58415]= 2035658475;
assign addr[58416]= 1981813720;
assign addr[58417]= 1917915825;
assign addr[58418]= 1844288924;
assign addr[58419]= 1761306505;
assign addr[58420]= 1669389513;
assign addr[58421]= 1569004214;
assign addr[58422]= 1460659832;
assign addr[58423]= 1344905966;
assign addr[58424]= 1222329801;
assign addr[58425]= 1093553126;
assign addr[58426]= 959229189;
assign addr[58427]= 820039373;
assign addr[58428]= 676689746;
assign addr[58429]= 529907477;
assign addr[58430]= 380437148;
assign addr[58431]= 229036977;
assign addr[58432]= 76474970;
assign addr[58433]= -76474970;
assign addr[58434]= -229036977;
assign addr[58435]= -380437148;
assign addr[58436]= -529907477;
assign addr[58437]= -676689746;
assign addr[58438]= -820039373;
assign addr[58439]= -959229189;
assign addr[58440]= -1093553126;
assign addr[58441]= -1222329801;
assign addr[58442]= -1344905966;
assign addr[58443]= -1460659832;
assign addr[58444]= -1569004214;
assign addr[58445]= -1669389513;
assign addr[58446]= -1761306505;
assign addr[58447]= -1844288924;
assign addr[58448]= -1917915825;
assign addr[58449]= -1981813720;
assign addr[58450]= -2035658475;
assign addr[58451]= -2079176953;
assign addr[58452]= -2112148396;
assign addr[58453]= -2134405552;
assign addr[58454]= -2145835515;
assign addr[58455]= -2146380306;
assign addr[58456]= -2136037160;
assign addr[58457]= -2114858546;
assign addr[58458]= -2082951896;
assign addr[58459]= -2040479063;
assign addr[58460]= -1987655498;
assign addr[58461]= -1924749160;
assign addr[58462]= -1852079154;
assign addr[58463]= -1770014111;
assign addr[58464]= -1678970324;
assign addr[58465]= -1579409630;
assign addr[58466]= -1471837070;
assign addr[58467]= -1356798326;
assign addr[58468]= -1234876957;
assign addr[58469]= -1106691431;
assign addr[58470]= -972891995;
assign addr[58471]= -834157373;
assign addr[58472]= -691191324;
assign addr[58473]= -544719071;
assign addr[58474]= -395483624;
assign addr[58475]= -244242007;
assign addr[58476]= -91761426;
assign addr[58477]= 61184634;
assign addr[58478]= 213820322;
assign addr[58479]= 365371365;
assign addr[58480]= 515068990;
assign addr[58481]= 662153826;
assign addr[58482]= 805879757;
assign addr[58483]= 945517704;
assign addr[58484]= 1080359326;
assign addr[58485]= 1209720613;
assign addr[58486]= 1332945355;
assign addr[58487]= 1449408469;
assign addr[58488]= 1558519173;
assign addr[58489]= 1659723983;
assign addr[58490]= 1752509516;
assign addr[58491]= 1836405100;
assign addr[58492]= 1910985158;
assign addr[58493]= 1975871368;
assign addr[58494]= 2030734582;
assign addr[58495]= 2075296495;
assign addr[58496]= 2109331059;
assign addr[58497]= 2132665626;
assign addr[58498]= 2145181827;
assign addr[58499]= 2146816171;
assign addr[58500]= 2137560369;
assign addr[58501]= 2117461370;
assign addr[58502]= 2086621133;
assign addr[58503]= 2045196100;
assign addr[58504]= 1993396407;
assign addr[58505]= 1931484818;
assign addr[58506]= 1859775393;
assign addr[58507]= 1778631892;
assign addr[58508]= 1688465931;
assign addr[58509]= 1589734894;
assign addr[58510]= 1482939614;
assign addr[58511]= 1368621831;
assign addr[58512]= 1247361445;
assign addr[58513]= 1119773573;
assign addr[58514]= 986505429;
assign addr[58515]= 848233042;
assign addr[58516]= 705657826;
assign addr[58517]= 559503022;
assign addr[58518]= 410510029;
assign addr[58519]= 259434643;
assign addr[58520]= 107043224;
assign addr[58521]= -45891193;
assign addr[58522]= -198592817;
assign addr[58523]= -350287041;
assign addr[58524]= -500204365;
assign addr[58525]= -647584304;
assign addr[58526]= -791679244;
assign addr[58527]= -931758235;
assign addr[58528]= -1067110699;
assign addr[58529]= -1197050035;
assign addr[58530]= -1320917099;
assign addr[58531]= -1438083551;
assign addr[58532]= -1547955041;
assign addr[58533]= -1649974225;
assign addr[58534]= -1743623590;
assign addr[58535]= -1828428082;
assign addr[58536]= -1903957513;
assign addr[58537]= -1969828744;
assign addr[58538]= -2025707632;
assign addr[58539]= -2071310720;
assign addr[58540]= -2106406677;
assign addr[58541]= -2130817471;
assign addr[58542]= -2144419275;
assign addr[58543]= -2147143090;
assign addr[58544]= -2138975100;
assign addr[58545]= -2119956737;
assign addr[58546]= -2090184478;
assign addr[58547]= -2049809346;
assign addr[58548]= -1999036154;
assign addr[58549]= -1938122457;
assign addr[58550]= -1867377253;
assign addr[58551]= -1787159411;
assign addr[58552]= -1697875851;
assign addr[58553]= -1599979481;
assign addr[58554]= -1493966902;
assign addr[58555]= -1380375881;
assign addr[58556]= -1259782632;
assign addr[58557]= -1132798888;
assign addr[58558]= -1000068799;
assign addr[58559]= -862265664;
assign addr[58560]= -720088517;
assign addr[58561]= -574258580;
assign addr[58562]= -425515602;
assign addr[58563]= -274614114;
assign addr[58564]= -122319591;
assign addr[58565]= 30595422;
assign addr[58566]= 183355234;
assign addr[58567]= 335184940;
assign addr[58568]= 485314355;
assign addr[58569]= 632981917;
assign addr[58570]= 777438554;
assign addr[58571]= 917951481;
assign addr[58572]= 1053807919;
assign addr[58573]= 1184318708;
assign addr[58574]= 1308821808;
assign addr[58575]= 1426685652;
assign addr[58576]= 1537312353;
assign addr[58577]= 1640140734;
assign addr[58578]= 1734649179;
assign addr[58579]= 1820358275;
assign addr[58580]= 1896833245;
assign addr[58581]= 1963686155;
assign addr[58582]= 2020577882;
assign addr[58583]= 2067219829;
assign addr[58584]= 2103375398;
assign addr[58585]= 2128861181;
assign addr[58586]= 2143547897;
assign addr[58587]= 2147361045;
assign addr[58588]= 2140281282;
assign addr[58589]= 2122344521;
assign addr[58590]= 2093641749;
assign addr[58591]= 2054318569;
assign addr[58592]= 2004574453;
assign addr[58593]= 1944661739;
assign addr[58594]= 1874884346;
assign addr[58595]= 1795596234;
assign addr[58596]= 1707199606;
assign addr[58597]= 1610142873;
assign addr[58598]= 1504918373;
assign addr[58599]= 1392059879;
assign addr[58600]= 1272139887;
assign addr[58601]= 1145766716;
assign addr[58602]= 1013581418;
assign addr[58603]= 876254528;
assign addr[58604]= 734482665;
assign addr[58605]= 588984994;
assign addr[58606]= 440499581;
assign addr[58607]= 289779648;
assign addr[58608]= 137589750;
assign addr[58609]= -15298099;
assign addr[58610]= -168108346;
assign addr[58611]= -320065829;
assign addr[58612]= -470399716;
assign addr[58613]= -618347408;
assign addr[58614]= -763158411;
assign addr[58615]= -904098143;
assign addr[58616]= -1040451659;
assign addr[58617]= -1171527280;
assign addr[58618]= -1296660098;
assign addr[58619]= -1415215352;
assign addr[58620]= -1526591649;
assign addr[58621]= -1630224009;
assign addr[58622]= -1725586737;
assign addr[58623]= -1812196087;
assign addr[58624]= -1889612716;
assign addr[58625]= -1957443913;
assign addr[58626]= -2015345591;
assign addr[58627]= -2063024031;
assign addr[58628]= -2100237377;
assign addr[58629]= -2126796855;
assign addr[58630]= -2142567738;
assign addr[58631]= -2147470025;
assign addr[58632]= -2141478848;
assign addr[58633]= -2124624598;
assign addr[58634]= -2096992772;
assign addr[58635]= -2058723538;
assign addr[58636]= -2010011024;
assign addr[58637]= -1951102334;
assign addr[58638]= -1882296293;
assign addr[58639]= -1803941934;
assign addr[58640]= -1716436725;
assign addr[58641]= -1620224553;
assign addr[58642]= -1515793473;
assign addr[58643]= -1403673233;
assign addr[58644]= -1284432584;
assign addr[58645]= -1158676398;
assign addr[58646]= -1027042599;
assign addr[58647]= -890198924;
assign addr[58648]= -748839539;
assign addr[58649]= -603681519;
assign addr[58650]= -455461206;
assign addr[58651]= -304930476;
assign addr[58652]= -152852926;
assign addr[58653]= 0;
assign addr[58654]= 152852926;
assign addr[58655]= 304930476;
assign addr[58656]= 455461206;
assign addr[58657]= 603681519;
assign addr[58658]= 748839539;
assign addr[58659]= 890198924;
assign addr[58660]= 1027042599;
assign addr[58661]= 1158676398;
assign addr[58662]= 1284432584;
assign addr[58663]= 1403673233;
assign addr[58664]= 1515793473;
assign addr[58665]= 1620224553;
assign addr[58666]= 1716436725;
assign addr[58667]= 1803941934;
assign addr[58668]= 1882296293;
assign addr[58669]= 1951102334;
assign addr[58670]= 2010011024;
assign addr[58671]= 2058723538;
assign addr[58672]= 2096992772;
assign addr[58673]= 2124624598;
assign addr[58674]= 2141478848;
assign addr[58675]= 2147470025;
assign addr[58676]= 2142567738;
assign addr[58677]= 2126796855;
assign addr[58678]= 2100237377;
assign addr[58679]= 2063024031;
assign addr[58680]= 2015345591;
assign addr[58681]= 1957443913;
assign addr[58682]= 1889612716;
assign addr[58683]= 1812196087;
assign addr[58684]= 1725586737;
assign addr[58685]= 1630224009;
assign addr[58686]= 1526591649;
assign addr[58687]= 1415215352;
assign addr[58688]= 1296660098;
assign addr[58689]= 1171527280;
assign addr[58690]= 1040451659;
assign addr[58691]= 904098143;
assign addr[58692]= 763158411;
assign addr[58693]= 618347408;
assign addr[58694]= 470399716;
assign addr[58695]= 320065829;
assign addr[58696]= 168108346;
assign addr[58697]= 15298099;
assign addr[58698]= -137589750;
assign addr[58699]= -289779648;
assign addr[58700]= -440499581;
assign addr[58701]= -588984994;
assign addr[58702]= -734482665;
assign addr[58703]= -876254528;
assign addr[58704]= -1013581418;
assign addr[58705]= -1145766716;
assign addr[58706]= -1272139887;
assign addr[58707]= -1392059879;
assign addr[58708]= -1504918373;
assign addr[58709]= -1610142873;
assign addr[58710]= -1707199606;
assign addr[58711]= -1795596234;
assign addr[58712]= -1874884346;
assign addr[58713]= -1944661739;
assign addr[58714]= -2004574453;
assign addr[58715]= -2054318569;
assign addr[58716]= -2093641749;
assign addr[58717]= -2122344521;
assign addr[58718]= -2140281282;
assign addr[58719]= -2147361045;
assign addr[58720]= -2143547897;
assign addr[58721]= -2128861181;
assign addr[58722]= -2103375398;
assign addr[58723]= -2067219829;
assign addr[58724]= -2020577882;
assign addr[58725]= -1963686155;
assign addr[58726]= -1896833245;
assign addr[58727]= -1820358275;
assign addr[58728]= -1734649179;
assign addr[58729]= -1640140734;
assign addr[58730]= -1537312353;
assign addr[58731]= -1426685652;
assign addr[58732]= -1308821808;
assign addr[58733]= -1184318708;
assign addr[58734]= -1053807919;
assign addr[58735]= -917951481;
assign addr[58736]= -777438554;
assign addr[58737]= -632981917;
assign addr[58738]= -485314355;
assign addr[58739]= -335184940;
assign addr[58740]= -183355234;
assign addr[58741]= -30595422;
assign addr[58742]= 122319591;
assign addr[58743]= 274614114;
assign addr[58744]= 425515602;
assign addr[58745]= 574258580;
assign addr[58746]= 720088517;
assign addr[58747]= 862265664;
assign addr[58748]= 1000068799;
assign addr[58749]= 1132798888;
assign addr[58750]= 1259782632;
assign addr[58751]= 1380375881;
assign addr[58752]= 1493966902;
assign addr[58753]= 1599979481;
assign addr[58754]= 1697875851;
assign addr[58755]= 1787159411;
assign addr[58756]= 1867377253;
assign addr[58757]= 1938122457;
assign addr[58758]= 1999036154;
assign addr[58759]= 2049809346;
assign addr[58760]= 2090184478;
assign addr[58761]= 2119956737;
assign addr[58762]= 2138975100;
assign addr[58763]= 2147143090;
assign addr[58764]= 2144419275;
assign addr[58765]= 2130817471;
assign addr[58766]= 2106406677;
assign addr[58767]= 2071310720;
assign addr[58768]= 2025707632;
assign addr[58769]= 1969828744;
assign addr[58770]= 1903957513;
assign addr[58771]= 1828428082;
assign addr[58772]= 1743623590;
assign addr[58773]= 1649974225;
assign addr[58774]= 1547955041;
assign addr[58775]= 1438083551;
assign addr[58776]= 1320917099;
assign addr[58777]= 1197050035;
assign addr[58778]= 1067110699;
assign addr[58779]= 931758235;
assign addr[58780]= 791679244;
assign addr[58781]= 647584304;
assign addr[58782]= 500204365;
assign addr[58783]= 350287041;
assign addr[58784]= 198592817;
assign addr[58785]= 45891193;
assign addr[58786]= -107043224;
assign addr[58787]= -259434643;
assign addr[58788]= -410510029;
assign addr[58789]= -559503022;
assign addr[58790]= -705657826;
assign addr[58791]= -848233042;
assign addr[58792]= -986505429;
assign addr[58793]= -1119773573;
assign addr[58794]= -1247361445;
assign addr[58795]= -1368621831;
assign addr[58796]= -1482939614;
assign addr[58797]= -1589734894;
assign addr[58798]= -1688465931;
assign addr[58799]= -1778631892;
assign addr[58800]= -1859775393;
assign addr[58801]= -1931484818;
assign addr[58802]= -1993396407;
assign addr[58803]= -2045196100;
assign addr[58804]= -2086621133;
assign addr[58805]= -2117461370;
assign addr[58806]= -2137560369;
assign addr[58807]= -2146816171;
assign addr[58808]= -2145181827;
assign addr[58809]= -2132665626;
assign addr[58810]= -2109331059;
assign addr[58811]= -2075296495;
assign addr[58812]= -2030734582;
assign addr[58813]= -1975871368;
assign addr[58814]= -1910985158;
assign addr[58815]= -1836405100;
assign addr[58816]= -1752509516;
assign addr[58817]= -1659723983;
assign addr[58818]= -1558519173;
assign addr[58819]= -1449408469;
assign addr[58820]= -1332945355;
assign addr[58821]= -1209720613;
assign addr[58822]= -1080359326;
assign addr[58823]= -945517704;
assign addr[58824]= -805879757;
assign addr[58825]= -662153826;
assign addr[58826]= -515068990;
assign addr[58827]= -365371365;
assign addr[58828]= -213820322;
assign addr[58829]= -61184634;
assign addr[58830]= 91761426;
assign addr[58831]= 244242007;
assign addr[58832]= 395483624;
assign addr[58833]= 544719071;
assign addr[58834]= 691191324;
assign addr[58835]= 834157373;
assign addr[58836]= 972891995;
assign addr[58837]= 1106691431;
assign addr[58838]= 1234876957;
assign addr[58839]= 1356798326;
assign addr[58840]= 1471837070;
assign addr[58841]= 1579409630;
assign addr[58842]= 1678970324;
assign addr[58843]= 1770014111;
assign addr[58844]= 1852079154;
assign addr[58845]= 1924749160;
assign addr[58846]= 1987655498;
assign addr[58847]= 2040479063;
assign addr[58848]= 2082951896;
assign addr[58849]= 2114858546;
assign addr[58850]= 2136037160;
assign addr[58851]= 2146380306;
assign addr[58852]= 2145835515;
assign addr[58853]= 2134405552;
assign addr[58854]= 2112148396;
assign addr[58855]= 2079176953;
assign addr[58856]= 2035658475;
assign addr[58857]= 1981813720;
assign addr[58858]= 1917915825;
assign addr[58859]= 1844288924;
assign addr[58860]= 1761306505;
assign addr[58861]= 1669389513;
assign addr[58862]= 1569004214;
assign addr[58863]= 1460659832;
assign addr[58864]= 1344905966;
assign addr[58865]= 1222329801;
assign addr[58866]= 1093553126;
assign addr[58867]= 959229189;
assign addr[58868]= 820039373;
assign addr[58869]= 676689746;
assign addr[58870]= 529907477;
assign addr[58871]= 380437148;
assign addr[58872]= 229036977;
assign addr[58873]= 76474970;
assign addr[58874]= -76474970;
assign addr[58875]= -229036977;
assign addr[58876]= -380437148;
assign addr[58877]= -529907477;
assign addr[58878]= -676689746;
assign addr[58879]= -820039373;
assign addr[58880]= -959229189;
assign addr[58881]= -1093553126;
assign addr[58882]= -1222329801;
assign addr[58883]= -1344905966;
assign addr[58884]= -1460659832;
assign addr[58885]= -1569004214;
assign addr[58886]= -1669389513;
assign addr[58887]= -1761306505;
assign addr[58888]= -1844288924;
assign addr[58889]= -1917915825;
assign addr[58890]= -1981813720;
assign addr[58891]= -2035658475;
assign addr[58892]= -2079176953;
assign addr[58893]= -2112148396;
assign addr[58894]= -2134405552;
assign addr[58895]= -2145835515;
assign addr[58896]= -2146380306;
assign addr[58897]= -2136037160;
assign addr[58898]= -2114858546;
assign addr[58899]= -2082951896;
assign addr[58900]= -2040479063;
assign addr[58901]= -1987655498;
assign addr[58902]= -1924749160;
assign addr[58903]= -1852079154;
assign addr[58904]= -1770014111;
assign addr[58905]= -1678970324;
assign addr[58906]= -1579409630;
assign addr[58907]= -1471837070;
assign addr[58908]= -1356798326;
assign addr[58909]= -1234876957;
assign addr[58910]= -1106691431;
assign addr[58911]= -972891995;
assign addr[58912]= -834157373;
assign addr[58913]= -691191324;
assign addr[58914]= -544719071;
assign addr[58915]= -395483624;
assign addr[58916]= -244242007;
assign addr[58917]= -91761426;
assign addr[58918]= 61184634;
assign addr[58919]= 213820322;
assign addr[58920]= 365371365;
assign addr[58921]= 515068990;
assign addr[58922]= 662153826;
assign addr[58923]= 805879757;
assign addr[58924]= 945517704;
assign addr[58925]= 1080359326;
assign addr[58926]= 1209720613;
assign addr[58927]= 1332945355;
assign addr[58928]= 1449408469;
assign addr[58929]= 1558519173;
assign addr[58930]= 1659723983;
assign addr[58931]= 1752509516;
assign addr[58932]= 1836405100;
assign addr[58933]= 1910985158;
assign addr[58934]= 1975871368;
assign addr[58935]= 2030734582;
assign addr[58936]= 2075296495;
assign addr[58937]= 2109331059;
assign addr[58938]= 2132665626;
assign addr[58939]= 2145181827;
assign addr[58940]= 2146816171;
assign addr[58941]= 2137560369;
assign addr[58942]= 2117461370;
assign addr[58943]= 2086621133;
assign addr[58944]= 2045196100;
assign addr[58945]= 1993396407;
assign addr[58946]= 1931484818;
assign addr[58947]= 1859775393;
assign addr[58948]= 1778631892;
assign addr[58949]= 1688465931;
assign addr[58950]= 1589734894;
assign addr[58951]= 1482939614;
assign addr[58952]= 1368621831;
assign addr[58953]= 1247361445;
assign addr[58954]= 1119773573;
assign addr[58955]= 986505429;
assign addr[58956]= 848233042;
assign addr[58957]= 705657826;
assign addr[58958]= 559503022;
assign addr[58959]= 410510029;
assign addr[58960]= 259434643;
assign addr[58961]= 107043224;
assign addr[58962]= -45891193;
assign addr[58963]= -198592817;
assign addr[58964]= -350287041;
assign addr[58965]= -500204365;
assign addr[58966]= -647584304;
assign addr[58967]= -791679244;
assign addr[58968]= -931758235;
assign addr[58969]= -1067110699;
assign addr[58970]= -1197050035;
assign addr[58971]= -1320917099;
assign addr[58972]= -1438083551;
assign addr[58973]= -1547955041;
assign addr[58974]= -1649974225;
assign addr[58975]= -1743623590;
assign addr[58976]= -1828428082;
assign addr[58977]= -1903957513;
assign addr[58978]= -1969828744;
assign addr[58979]= -2025707632;
assign addr[58980]= -2071310720;
assign addr[58981]= -2106406677;
assign addr[58982]= -2130817471;
assign addr[58983]= -2144419275;
assign addr[58984]= -2147143090;
assign addr[58985]= -2138975100;
assign addr[58986]= -2119956737;
assign addr[58987]= -2090184478;
assign addr[58988]= -2049809346;
assign addr[58989]= -1999036154;
assign addr[58990]= -1938122457;
assign addr[58991]= -1867377253;
assign addr[58992]= -1787159411;
assign addr[58993]= -1697875851;
assign addr[58994]= -1599979481;
assign addr[58995]= -1493966902;
assign addr[58996]= -1380375881;
assign addr[58997]= -1259782632;
assign addr[58998]= -1132798888;
assign addr[58999]= -1000068799;
assign addr[59000]= -862265664;
assign addr[59001]= -720088517;
assign addr[59002]= -574258580;
assign addr[59003]= -425515602;
assign addr[59004]= -274614114;
assign addr[59005]= -122319591;
assign addr[59006]= 30595422;
assign addr[59007]= 183355234;
assign addr[59008]= 335184940;
assign addr[59009]= 485314355;
assign addr[59010]= 632981917;
assign addr[59011]= 777438554;
assign addr[59012]= 917951481;
assign addr[59013]= 1053807919;
assign addr[59014]= 1184318708;
assign addr[59015]= 1308821808;
assign addr[59016]= 1426685652;
assign addr[59017]= 1537312353;
assign addr[59018]= 1640140734;
assign addr[59019]= 1734649179;
assign addr[59020]= 1820358275;
assign addr[59021]= 1896833245;
assign addr[59022]= 1963686155;
assign addr[59023]= 2020577882;
assign addr[59024]= 2067219829;
assign addr[59025]= 2103375398;
assign addr[59026]= 2128861181;
assign addr[59027]= 2143547897;
assign addr[59028]= 2147361045;
assign addr[59029]= 2140281282;
assign addr[59030]= 2122344521;
assign addr[59031]= 2093641749;
assign addr[59032]= 2054318569;
assign addr[59033]= 2004574453;
assign addr[59034]= 1944661739;
assign addr[59035]= 1874884346;
assign addr[59036]= 1795596234;
assign addr[59037]= 1707199606;
assign addr[59038]= 1610142873;
assign addr[59039]= 1504918373;
assign addr[59040]= 1392059879;
assign addr[59041]= 1272139887;
assign addr[59042]= 1145766716;
assign addr[59043]= 1013581418;
assign addr[59044]= 876254528;
assign addr[59045]= 734482665;
assign addr[59046]= 588984994;
assign addr[59047]= 440499581;
assign addr[59048]= 289779648;
assign addr[59049]= 137589750;
assign addr[59050]= -15298099;
assign addr[59051]= -168108346;
assign addr[59052]= -320065829;
assign addr[59053]= -470399716;
assign addr[59054]= -618347408;
assign addr[59055]= -763158411;
assign addr[59056]= -904098143;
assign addr[59057]= -1040451659;
assign addr[59058]= -1171527280;
assign addr[59059]= -1296660098;
assign addr[59060]= -1415215352;
assign addr[59061]= -1526591649;
assign addr[59062]= -1630224009;
assign addr[59063]= -1725586737;
assign addr[59064]= -1812196087;
assign addr[59065]= -1889612716;
assign addr[59066]= -1957443913;
assign addr[59067]= -2015345591;
assign addr[59068]= -2063024031;
assign addr[59069]= -2100237377;
assign addr[59070]= -2126796855;
assign addr[59071]= -2142567738;
assign addr[59072]= -2147470025;
assign addr[59073]= -2141478848;
assign addr[59074]= -2124624598;
assign addr[59075]= -2096992772;
assign addr[59076]= -2058723538;
assign addr[59077]= -2010011024;
assign addr[59078]= -1951102334;
assign addr[59079]= -1882296293;
assign addr[59080]= -1803941934;
assign addr[59081]= -1716436725;
assign addr[59082]= -1620224553;
assign addr[59083]= -1515793473;
assign addr[59084]= -1403673233;
assign addr[59085]= -1284432584;
assign addr[59086]= -1158676398;
assign addr[59087]= -1027042599;
assign addr[59088]= -890198924;
assign addr[59089]= -748839539;
assign addr[59090]= -603681519;
assign addr[59091]= -455461206;
assign addr[59092]= -304930476;
assign addr[59093]= -152852926;
assign addr[59094]= 0;
assign addr[59095]= 152852926;
assign addr[59096]= 304930476;
assign addr[59097]= 455461206;
assign addr[59098]= 603681519;
assign addr[59099]= 748839539;
assign addr[59100]= 890198924;
assign addr[59101]= 1027042599;
assign addr[59102]= 1158676398;
assign addr[59103]= 1284432584;
assign addr[59104]= 1403673233;
assign addr[59105]= 1515793473;
assign addr[59106]= 1620224553;
assign addr[59107]= 1716436725;
assign addr[59108]= 1803941934;
assign addr[59109]= 1882296293;
assign addr[59110]= 1951102334;
assign addr[59111]= 2010011024;
assign addr[59112]= 2058723538;
assign addr[59113]= 2096992772;
assign addr[59114]= 2124624598;
assign addr[59115]= 2141478848;
assign addr[59116]= 2147470025;
assign addr[59117]= 2142567738;
assign addr[59118]= 2126796855;
assign addr[59119]= 2100237377;
assign addr[59120]= 2063024031;
assign addr[59121]= 2015345591;
assign addr[59122]= 1957443913;
assign addr[59123]= 1889612716;
assign addr[59124]= 1812196087;
assign addr[59125]= 1725586737;
assign addr[59126]= 1630224009;
assign addr[59127]= 1526591649;
assign addr[59128]= 1415215352;
assign addr[59129]= 1296660098;
assign addr[59130]= 1171527280;
assign addr[59131]= 1040451659;
assign addr[59132]= 904098143;
assign addr[59133]= 763158411;
assign addr[59134]= 618347408;
assign addr[59135]= 470399716;
assign addr[59136]= 320065829;
assign addr[59137]= 168108346;
assign addr[59138]= 15298099;
assign addr[59139]= -137589750;
assign addr[59140]= -289779648;
assign addr[59141]= -440499581;
assign addr[59142]= -588984994;
assign addr[59143]= -734482665;
assign addr[59144]= -876254528;
assign addr[59145]= -1013581418;
assign addr[59146]= -1145766716;
assign addr[59147]= -1272139887;
assign addr[59148]= -1392059879;
assign addr[59149]= -1504918373;
assign addr[59150]= -1610142873;
assign addr[59151]= -1707199606;
assign addr[59152]= -1795596234;
assign addr[59153]= -1874884346;
assign addr[59154]= -1944661739;
assign addr[59155]= -2004574453;
assign addr[59156]= -2054318569;
assign addr[59157]= -2093641749;
assign addr[59158]= -2122344521;
assign addr[59159]= -2140281282;
assign addr[59160]= -2147361045;
assign addr[59161]= -2143547897;
assign addr[59162]= -2128861181;
assign addr[59163]= -2103375398;
assign addr[59164]= -2067219829;
assign addr[59165]= -2020577882;
assign addr[59166]= -1963686155;
assign addr[59167]= -1896833245;
assign addr[59168]= -1820358275;
assign addr[59169]= -1734649179;
assign addr[59170]= -1640140734;
assign addr[59171]= -1537312353;
assign addr[59172]= -1426685652;
assign addr[59173]= -1308821808;
assign addr[59174]= -1184318708;
assign addr[59175]= -1053807919;
assign addr[59176]= -917951481;
assign addr[59177]= -777438554;
assign addr[59178]= -632981917;
assign addr[59179]= -485314355;
assign addr[59180]= -335184940;
assign addr[59181]= -183355234;
assign addr[59182]= -30595422;
assign addr[59183]= 122319591;
assign addr[59184]= 274614114;
assign addr[59185]= 425515602;
assign addr[59186]= 574258580;
assign addr[59187]= 720088517;
assign addr[59188]= 862265664;
assign addr[59189]= 1000068799;
assign addr[59190]= 1132798888;
assign addr[59191]= 1259782632;
assign addr[59192]= 1380375881;
assign addr[59193]= 1493966902;
assign addr[59194]= 1599979481;
assign addr[59195]= 1697875851;
assign addr[59196]= 1787159411;
assign addr[59197]= 1867377253;
assign addr[59198]= 1938122457;
assign addr[59199]= 1999036154;
assign addr[59200]= 2049809346;
assign addr[59201]= 2090184478;
assign addr[59202]= 2119956737;
assign addr[59203]= 2138975100;
assign addr[59204]= 2147143090;
assign addr[59205]= 2144419275;
assign addr[59206]= 2130817471;
assign addr[59207]= 2106406677;
assign addr[59208]= 2071310720;
assign addr[59209]= 2025707632;
assign addr[59210]= 1969828744;
assign addr[59211]= 1903957513;
assign addr[59212]= 1828428082;
assign addr[59213]= 1743623590;
assign addr[59214]= 1649974225;
assign addr[59215]= 1547955041;
assign addr[59216]= 1438083551;
assign addr[59217]= 1320917099;
assign addr[59218]= 1197050035;
assign addr[59219]= 1067110699;
assign addr[59220]= 931758235;
assign addr[59221]= 791679244;
assign addr[59222]= 647584304;
assign addr[59223]= 500204365;
assign addr[59224]= 350287041;
assign addr[59225]= 198592817;
assign addr[59226]= 45891193;
assign addr[59227]= -107043224;
assign addr[59228]= -259434643;
assign addr[59229]= -410510029;
assign addr[59230]= -559503022;
assign addr[59231]= -705657826;
assign addr[59232]= -848233042;
assign addr[59233]= -986505429;
assign addr[59234]= -1119773573;
assign addr[59235]= -1247361445;
assign addr[59236]= -1368621831;
assign addr[59237]= -1482939614;
assign addr[59238]= -1589734894;
assign addr[59239]= -1688465931;
assign addr[59240]= -1778631892;
assign addr[59241]= -1859775393;
assign addr[59242]= -1931484818;
assign addr[59243]= -1993396407;
assign addr[59244]= -2045196100;
assign addr[59245]= -2086621133;
assign addr[59246]= -2117461370;
assign addr[59247]= -2137560369;
assign addr[59248]= -2146816171;
assign addr[59249]= -2145181827;
assign addr[59250]= -2132665626;
assign addr[59251]= -2109331059;
assign addr[59252]= -2075296495;
assign addr[59253]= -2030734582;
assign addr[59254]= -1975871368;
assign addr[59255]= -1910985158;
assign addr[59256]= -1836405100;
assign addr[59257]= -1752509516;
assign addr[59258]= -1659723983;
assign addr[59259]= -1558519173;
assign addr[59260]= -1449408469;
assign addr[59261]= -1332945355;
assign addr[59262]= -1209720613;
assign addr[59263]= -1080359326;
assign addr[59264]= -945517704;
assign addr[59265]= -805879757;
assign addr[59266]= -662153826;
assign addr[59267]= -515068990;
assign addr[59268]= -365371365;
assign addr[59269]= -213820322;
assign addr[59270]= -61184634;
assign addr[59271]= 91761426;
assign addr[59272]= 244242007;
assign addr[59273]= 395483624;
assign addr[59274]= 544719071;
assign addr[59275]= 691191324;
assign addr[59276]= 834157373;
assign addr[59277]= 972891995;
assign addr[59278]= 1106691431;
assign addr[59279]= 1234876957;
assign addr[59280]= 1356798326;
assign addr[59281]= 1471837070;
assign addr[59282]= 1579409630;
assign addr[59283]= 1678970324;
assign addr[59284]= 1770014111;
assign addr[59285]= 1852079154;
assign addr[59286]= 1924749160;
assign addr[59287]= 1987655498;
assign addr[59288]= 2040479063;
assign addr[59289]= 2082951896;
assign addr[59290]= 2114858546;
assign addr[59291]= 2136037160;
assign addr[59292]= 2146380306;
assign addr[59293]= 2145835515;
assign addr[59294]= 2134405552;
assign addr[59295]= 2112148396;
assign addr[59296]= 2079176953;
assign addr[59297]= 2035658475;
assign addr[59298]= 1981813720;
assign addr[59299]= 1917915825;
assign addr[59300]= 1844288924;
assign addr[59301]= 1761306505;
assign addr[59302]= 1669389513;
assign addr[59303]= 1569004214;
assign addr[59304]= 1460659832;
assign addr[59305]= 1344905966;
assign addr[59306]= 1222329801;
assign addr[59307]= 1093553126;
assign addr[59308]= 959229189;
assign addr[59309]= 820039373;
assign addr[59310]= 676689746;
assign addr[59311]= 529907477;
assign addr[59312]= 380437148;
assign addr[59313]= 229036977;
assign addr[59314]= 76474970;
assign addr[59315]= -76474970;
assign addr[59316]= -229036977;
assign addr[59317]= -380437148;
assign addr[59318]= -529907477;
assign addr[59319]= -676689746;
assign addr[59320]= -820039373;
assign addr[59321]= -959229189;
assign addr[59322]= -1093553126;
assign addr[59323]= -1222329801;
assign addr[59324]= -1344905966;
assign addr[59325]= -1460659832;
assign addr[59326]= -1569004214;
assign addr[59327]= -1669389513;
assign addr[59328]= -1761306505;
assign addr[59329]= -1844288924;
assign addr[59330]= -1917915825;
assign addr[59331]= -1981813720;
assign addr[59332]= -2035658475;
assign addr[59333]= -2079176953;
assign addr[59334]= -2112148396;
assign addr[59335]= -2134405552;
assign addr[59336]= -2145835515;
assign addr[59337]= -2146380306;
assign addr[59338]= -2136037160;
assign addr[59339]= -2114858546;
assign addr[59340]= -2082951896;
assign addr[59341]= -2040479063;
assign addr[59342]= -1987655498;
assign addr[59343]= -1924749160;
assign addr[59344]= -1852079154;
assign addr[59345]= -1770014111;
assign addr[59346]= -1678970324;
assign addr[59347]= -1579409630;
assign addr[59348]= -1471837070;
assign addr[59349]= -1356798326;
assign addr[59350]= -1234876957;
assign addr[59351]= -1106691431;
assign addr[59352]= -972891995;
assign addr[59353]= -834157373;
assign addr[59354]= -691191324;
assign addr[59355]= -544719071;
assign addr[59356]= -395483624;
assign addr[59357]= -244242007;
assign addr[59358]= -91761426;
assign addr[59359]= 61184634;
assign addr[59360]= 213820322;
assign addr[59361]= 365371365;
assign addr[59362]= 515068990;
assign addr[59363]= 662153826;
assign addr[59364]= 805879757;
assign addr[59365]= 945517704;
assign addr[59366]= 1080359326;
assign addr[59367]= 1209720613;
assign addr[59368]= 1332945355;
assign addr[59369]= 1449408469;
assign addr[59370]= 1558519173;
assign addr[59371]= 1659723983;
assign addr[59372]= 1752509516;
assign addr[59373]= 1836405100;
assign addr[59374]= 1910985158;
assign addr[59375]= 1975871368;
assign addr[59376]= 2030734582;
assign addr[59377]= 2075296495;
assign addr[59378]= 2109331059;
assign addr[59379]= 2132665626;
assign addr[59380]= 2145181827;
assign addr[59381]= 2146816171;
assign addr[59382]= 2137560369;
assign addr[59383]= 2117461370;
assign addr[59384]= 2086621133;
assign addr[59385]= 2045196100;
assign addr[59386]= 1993396407;
assign addr[59387]= 1931484818;
assign addr[59388]= 1859775393;
assign addr[59389]= 1778631892;
assign addr[59390]= 1688465931;
assign addr[59391]= 1589734894;
assign addr[59392]= 1482939614;
assign addr[59393]= 1368621831;
assign addr[59394]= 1247361445;
assign addr[59395]= 1119773573;
assign addr[59396]= 986505429;
assign addr[59397]= 848233042;
assign addr[59398]= 705657826;
assign addr[59399]= 559503022;
assign addr[59400]= 410510029;
assign addr[59401]= 259434643;
assign addr[59402]= 107043224;
assign addr[59403]= -45891193;
assign addr[59404]= -198592817;
assign addr[59405]= -350287041;
assign addr[59406]= -500204365;
assign addr[59407]= -647584304;
assign addr[59408]= -791679244;
assign addr[59409]= -931758235;
assign addr[59410]= -1067110699;
assign addr[59411]= -1197050035;
assign addr[59412]= -1320917099;
assign addr[59413]= -1438083551;
assign addr[59414]= -1547955041;
assign addr[59415]= -1649974225;
assign addr[59416]= -1743623590;
assign addr[59417]= -1828428082;
assign addr[59418]= -1903957513;
assign addr[59419]= -1969828744;
assign addr[59420]= -2025707632;
assign addr[59421]= -2071310720;
assign addr[59422]= -2106406677;
assign addr[59423]= -2130817471;
assign addr[59424]= -2144419275;
assign addr[59425]= -2147143090;
assign addr[59426]= -2138975100;
assign addr[59427]= -2119956737;
assign addr[59428]= -2090184478;
assign addr[59429]= -2049809346;
assign addr[59430]= -1999036154;
assign addr[59431]= -1938122457;
assign addr[59432]= -1867377253;
assign addr[59433]= -1787159411;
assign addr[59434]= -1697875851;
assign addr[59435]= -1599979481;
assign addr[59436]= -1493966902;
assign addr[59437]= -1380375881;
assign addr[59438]= -1259782632;
assign addr[59439]= -1132798888;
assign addr[59440]= -1000068799;
assign addr[59441]= -862265664;
assign addr[59442]= -720088517;
assign addr[59443]= -574258580;
assign addr[59444]= -425515602;
assign addr[59445]= -274614114;
assign addr[59446]= -122319591;
assign addr[59447]= 30595422;
assign addr[59448]= 183355234;
assign addr[59449]= 335184940;
assign addr[59450]= 485314355;
assign addr[59451]= 632981917;
assign addr[59452]= 777438554;
assign addr[59453]= 917951481;
assign addr[59454]= 1053807919;
assign addr[59455]= 1184318708;
assign addr[59456]= 1308821808;
assign addr[59457]= 1426685652;
assign addr[59458]= 1537312353;
assign addr[59459]= 1640140734;
assign addr[59460]= 1734649179;
assign addr[59461]= 1820358275;
assign addr[59462]= 1896833245;
assign addr[59463]= 1963686155;
assign addr[59464]= 2020577882;
assign addr[59465]= 2067219829;
assign addr[59466]= 2103375398;
assign addr[59467]= 2128861181;
assign addr[59468]= 2143547897;
assign addr[59469]= 2147361045;
assign addr[59470]= 2140281282;
assign addr[59471]= 2122344521;
assign addr[59472]= 2093641749;
assign addr[59473]= 2054318569;
assign addr[59474]= 2004574453;
assign addr[59475]= 1944661739;
assign addr[59476]= 1874884346;
assign addr[59477]= 1795596234;
assign addr[59478]= 1707199606;
assign addr[59479]= 1610142873;
assign addr[59480]= 1504918373;
assign addr[59481]= 1392059879;
assign addr[59482]= 1272139887;
assign addr[59483]= 1145766716;
assign addr[59484]= 1013581418;
assign addr[59485]= 876254528;
assign addr[59486]= 734482665;
assign addr[59487]= 588984994;
assign addr[59488]= 440499581;
assign addr[59489]= 289779648;
assign addr[59490]= 137589750;
assign addr[59491]= -15298099;
assign addr[59492]= -168108346;
assign addr[59493]= -320065829;
assign addr[59494]= -470399716;
assign addr[59495]= -618347408;
assign addr[59496]= -763158411;
assign addr[59497]= -904098143;
assign addr[59498]= -1040451659;
assign addr[59499]= -1171527280;
assign addr[59500]= -1296660098;
assign addr[59501]= -1415215352;
assign addr[59502]= -1526591649;
assign addr[59503]= -1630224009;
assign addr[59504]= -1725586737;
assign addr[59505]= -1812196087;
assign addr[59506]= -1889612716;
assign addr[59507]= -1957443913;
assign addr[59508]= -2015345591;
assign addr[59509]= -2063024031;
assign addr[59510]= -2100237377;
assign addr[59511]= -2126796855;
assign addr[59512]= -2142567738;
assign addr[59513]= -2147470025;
assign addr[59514]= -2141478848;
assign addr[59515]= -2124624598;
assign addr[59516]= -2096992772;
assign addr[59517]= -2058723538;
assign addr[59518]= -2010011024;
assign addr[59519]= -1951102334;
assign addr[59520]= -1882296293;
assign addr[59521]= -1803941934;
assign addr[59522]= -1716436725;
assign addr[59523]= -1620224553;
assign addr[59524]= -1515793473;
assign addr[59525]= -1403673233;
assign addr[59526]= -1284432584;
assign addr[59527]= -1158676398;
assign addr[59528]= -1027042599;
assign addr[59529]= -890198924;
assign addr[59530]= -748839539;
assign addr[59531]= -603681519;
assign addr[59532]= -455461206;
assign addr[59533]= -304930476;
assign addr[59534]= -152852926;
assign addr[59535]= 0;
assign addr[59536]= 152852926;
assign addr[59537]= 304930476;
assign addr[59538]= 455461206;
assign addr[59539]= 603681519;
assign addr[59540]= 748839539;
assign addr[59541]= 890198924;
assign addr[59542]= 1027042599;
assign addr[59543]= 1158676398;
assign addr[59544]= 1284432584;
assign addr[59545]= 1403673233;
assign addr[59546]= 1515793473;
assign addr[59547]= 1620224553;
assign addr[59548]= 1716436725;
assign addr[59549]= 1803941934;
assign addr[59550]= 1882296293;
assign addr[59551]= 1951102334;
assign addr[59552]= 2010011024;
assign addr[59553]= 2058723538;
assign addr[59554]= 2096992772;
assign addr[59555]= 2124624598;
assign addr[59556]= 2141478848;
assign addr[59557]= 2147470025;
assign addr[59558]= 2142567738;
assign addr[59559]= 2126796855;
assign addr[59560]= 2100237377;
assign addr[59561]= 2063024031;
assign addr[59562]= 2015345591;
assign addr[59563]= 1957443913;
assign addr[59564]= 1889612716;
assign addr[59565]= 1812196087;
assign addr[59566]= 1725586737;
assign addr[59567]= 1630224009;
assign addr[59568]= 1526591649;
assign addr[59569]= 1415215352;
assign addr[59570]= 1296660098;
assign addr[59571]= 1171527280;
assign addr[59572]= 1040451659;
assign addr[59573]= 904098143;
assign addr[59574]= 763158411;
assign addr[59575]= 618347408;
assign addr[59576]= 470399716;
assign addr[59577]= 320065829;
assign addr[59578]= 168108346;
assign addr[59579]= 15298099;
assign addr[59580]= -137589750;
assign addr[59581]= -289779648;
assign addr[59582]= -440499581;
assign addr[59583]= -588984994;
assign addr[59584]= -734482665;
assign addr[59585]= -876254528;
assign addr[59586]= -1013581418;
assign addr[59587]= -1145766716;
assign addr[59588]= -1272139887;
assign addr[59589]= -1392059879;
assign addr[59590]= -1504918373;
assign addr[59591]= -1610142873;
assign addr[59592]= -1707199606;
assign addr[59593]= -1795596234;
assign addr[59594]= -1874884346;
assign addr[59595]= -1944661739;
assign addr[59596]= -2004574453;
assign addr[59597]= -2054318569;
assign addr[59598]= -2093641749;
assign addr[59599]= -2122344521;
assign addr[59600]= -2140281282;
assign addr[59601]= -2147361045;
assign addr[59602]= -2143547897;
assign addr[59603]= -2128861181;
assign addr[59604]= -2103375398;
assign addr[59605]= -2067219829;
assign addr[59606]= -2020577882;
assign addr[59607]= -1963686155;
assign addr[59608]= -1896833245;
assign addr[59609]= -1820358275;
assign addr[59610]= -1734649179;
assign addr[59611]= -1640140734;
assign addr[59612]= -1537312353;
assign addr[59613]= -1426685652;
assign addr[59614]= -1308821808;
assign addr[59615]= -1184318708;
assign addr[59616]= -1053807919;
assign addr[59617]= -917951481;
assign addr[59618]= -777438554;
assign addr[59619]= -632981917;
assign addr[59620]= -485314355;
assign addr[59621]= -335184940;
assign addr[59622]= -183355234;
assign addr[59623]= -30595422;
assign addr[59624]= 122319591;
assign addr[59625]= 274614114;
assign addr[59626]= 425515602;
assign addr[59627]= 574258580;
assign addr[59628]= 720088517;
assign addr[59629]= 862265664;
assign addr[59630]= 1000068799;
assign addr[59631]= 1132798888;
assign addr[59632]= 1259782632;
assign addr[59633]= 1380375881;
assign addr[59634]= 1493966902;
assign addr[59635]= 1599979481;
assign addr[59636]= 1697875851;
assign addr[59637]= 1787159411;
assign addr[59638]= 1867377253;
assign addr[59639]= 1938122457;
assign addr[59640]= 1999036154;
assign addr[59641]= 2049809346;
assign addr[59642]= 2090184478;
assign addr[59643]= 2119956737;
assign addr[59644]= 2138975100;
assign addr[59645]= 2147143090;
assign addr[59646]= 2144419275;
assign addr[59647]= 2130817471;
assign addr[59648]= 2106406677;
assign addr[59649]= 2071310720;
assign addr[59650]= 2025707632;
assign addr[59651]= 1969828744;
assign addr[59652]= 1903957513;
assign addr[59653]= 1828428082;
assign addr[59654]= 1743623590;
assign addr[59655]= 1649974225;
assign addr[59656]= 1547955041;
assign addr[59657]= 1438083551;
assign addr[59658]= 1320917099;
assign addr[59659]= 1197050035;
assign addr[59660]= 1067110699;
assign addr[59661]= 931758235;
assign addr[59662]= 791679244;
assign addr[59663]= 647584304;
assign addr[59664]= 500204365;
assign addr[59665]= 350287041;
assign addr[59666]= 198592817;
assign addr[59667]= 45891193;
assign addr[59668]= -107043224;
assign addr[59669]= -259434643;
assign addr[59670]= -410510029;
assign addr[59671]= -559503022;
assign addr[59672]= -705657826;
assign addr[59673]= -848233042;
assign addr[59674]= -986505429;
assign addr[59675]= -1119773573;
assign addr[59676]= -1247361445;
assign addr[59677]= -1368621831;
assign addr[59678]= -1482939614;
assign addr[59679]= -1589734894;
assign addr[59680]= -1688465931;
assign addr[59681]= -1778631892;
assign addr[59682]= -1859775393;
assign addr[59683]= -1931484818;
assign addr[59684]= -1993396407;
assign addr[59685]= -2045196100;
assign addr[59686]= -2086621133;
assign addr[59687]= -2117461370;
assign addr[59688]= -2137560369;
assign addr[59689]= -2146816171;
assign addr[59690]= -2145181827;
assign addr[59691]= -2132665626;
assign addr[59692]= -2109331059;
assign addr[59693]= -2075296495;
assign addr[59694]= -2030734582;
assign addr[59695]= -1975871368;
assign addr[59696]= -1910985158;
assign addr[59697]= -1836405100;
assign addr[59698]= -1752509516;
assign addr[59699]= -1659723983;
assign addr[59700]= -1558519173;
assign addr[59701]= -1449408469;
assign addr[59702]= -1332945355;
assign addr[59703]= -1209720613;
assign addr[59704]= -1080359326;
assign addr[59705]= -945517704;
assign addr[59706]= -805879757;
assign addr[59707]= -662153826;
assign addr[59708]= -515068990;
assign addr[59709]= -365371365;
assign addr[59710]= -213820322;
assign addr[59711]= -61184634;
assign addr[59712]= 91761426;
assign addr[59713]= 244242007;
assign addr[59714]= 395483624;
assign addr[59715]= 544719071;
assign addr[59716]= 691191324;
assign addr[59717]= 834157373;
assign addr[59718]= 972891995;
assign addr[59719]= 1106691431;
assign addr[59720]= 1234876957;
assign addr[59721]= 1356798326;
assign addr[59722]= 1471837070;
assign addr[59723]= 1579409630;
assign addr[59724]= 1678970324;
assign addr[59725]= 1770014111;
assign addr[59726]= 1852079154;
assign addr[59727]= 1924749160;
assign addr[59728]= 1987655498;
assign addr[59729]= 2040479063;
assign addr[59730]= 2082951896;
assign addr[59731]= 2114858546;
assign addr[59732]= 2136037160;
assign addr[59733]= 2146380306;
assign addr[59734]= 2145835515;
assign addr[59735]= 2134405552;
assign addr[59736]= 2112148396;
assign addr[59737]= 2079176953;
assign addr[59738]= 2035658475;
assign addr[59739]= 1981813720;
assign addr[59740]= 1917915825;
assign addr[59741]= 1844288924;
assign addr[59742]= 1761306505;
assign addr[59743]= 1669389513;
assign addr[59744]= 1569004214;
assign addr[59745]= 1460659832;
assign addr[59746]= 1344905966;
assign addr[59747]= 1222329801;
assign addr[59748]= 1093553126;
assign addr[59749]= 959229189;
assign addr[59750]= 820039373;
assign addr[59751]= 676689746;
assign addr[59752]= 529907477;
assign addr[59753]= 380437148;
assign addr[59754]= 229036977;
assign addr[59755]= 76474970;
assign addr[59756]= -76474970;
assign addr[59757]= -229036977;
assign addr[59758]= -380437148;
assign addr[59759]= -529907477;
assign addr[59760]= -676689746;
assign addr[59761]= -820039373;
assign addr[59762]= -959229189;
assign addr[59763]= -1093553126;
assign addr[59764]= -1222329801;
assign addr[59765]= -1344905966;
assign addr[59766]= -1460659832;
assign addr[59767]= -1569004214;
assign addr[59768]= -1669389513;
assign addr[59769]= -1761306505;
assign addr[59770]= -1844288924;
assign addr[59771]= -1917915825;
assign addr[59772]= -1981813720;
assign addr[59773]= -2035658475;
assign addr[59774]= -2079176953;
assign addr[59775]= -2112148396;
assign addr[59776]= -2134405552;
assign addr[59777]= -2145835515;
assign addr[59778]= -2146380306;
assign addr[59779]= -2136037160;
assign addr[59780]= -2114858546;
assign addr[59781]= -2082951896;
assign addr[59782]= -2040479063;
assign addr[59783]= -1987655498;
assign addr[59784]= -1924749160;
assign addr[59785]= -1852079154;
assign addr[59786]= -1770014111;
assign addr[59787]= -1678970324;
assign addr[59788]= -1579409630;
assign addr[59789]= -1471837070;
assign addr[59790]= -1356798326;
assign addr[59791]= -1234876957;
assign addr[59792]= -1106691431;
assign addr[59793]= -972891995;
assign addr[59794]= -834157373;
assign addr[59795]= -691191324;
assign addr[59796]= -544719071;
assign addr[59797]= -395483624;
assign addr[59798]= -244242007;
assign addr[59799]= -91761426;
assign addr[59800]= 61184634;
assign addr[59801]= 213820322;
assign addr[59802]= 365371365;
assign addr[59803]= 515068990;
assign addr[59804]= 662153826;
assign addr[59805]= 805879757;
assign addr[59806]= 945517704;
assign addr[59807]= 1080359326;
assign addr[59808]= 1209720613;
assign addr[59809]= 1332945355;
assign addr[59810]= 1449408469;
assign addr[59811]= 1558519173;
assign addr[59812]= 1659723983;
assign addr[59813]= 1752509516;
assign addr[59814]= 1836405100;
assign addr[59815]= 1910985158;
assign addr[59816]= 1975871368;
assign addr[59817]= 2030734582;
assign addr[59818]= 2075296495;
assign addr[59819]= 2109331059;
assign addr[59820]= 2132665626;
assign addr[59821]= 2145181827;
assign addr[59822]= 2146816171;
assign addr[59823]= 2137560369;
assign addr[59824]= 2117461370;
assign addr[59825]= 2086621133;
assign addr[59826]= 2045196100;
assign addr[59827]= 1993396407;
assign addr[59828]= 1931484818;
assign addr[59829]= 1859775393;
assign addr[59830]= 1778631892;
assign addr[59831]= 1688465931;
assign addr[59832]= 1589734894;
assign addr[59833]= 1482939614;
assign addr[59834]= 1368621831;
assign addr[59835]= 1247361445;
assign addr[59836]= 1119773573;
assign addr[59837]= 986505429;
assign addr[59838]= 848233042;
assign addr[59839]= 705657826;
assign addr[59840]= 559503022;
assign addr[59841]= 410510029;
assign addr[59842]= 259434643;
assign addr[59843]= 107043224;
assign addr[59844]= -45891193;
assign addr[59845]= -198592817;
assign addr[59846]= -350287041;
assign addr[59847]= -500204365;
assign addr[59848]= -647584304;
assign addr[59849]= -791679244;
assign addr[59850]= -931758235;
assign addr[59851]= -1067110699;
assign addr[59852]= -1197050035;
assign addr[59853]= -1320917099;
assign addr[59854]= -1438083551;
assign addr[59855]= -1547955041;
assign addr[59856]= -1649974225;
assign addr[59857]= -1743623590;
assign addr[59858]= -1828428082;
assign addr[59859]= -1903957513;
assign addr[59860]= -1969828744;
assign addr[59861]= -2025707632;
assign addr[59862]= -2071310720;
assign addr[59863]= -2106406677;
assign addr[59864]= -2130817471;
assign addr[59865]= -2144419275;
assign addr[59866]= -2147143090;
assign addr[59867]= -2138975100;
assign addr[59868]= -2119956737;
assign addr[59869]= -2090184478;
assign addr[59870]= -2049809346;
assign addr[59871]= -1999036154;
assign addr[59872]= -1938122457;
assign addr[59873]= -1867377253;
assign addr[59874]= -1787159411;
assign addr[59875]= -1697875851;
assign addr[59876]= -1599979481;
assign addr[59877]= -1493966902;
assign addr[59878]= -1380375881;
assign addr[59879]= -1259782632;
assign addr[59880]= -1132798888;
assign addr[59881]= -1000068799;
assign addr[59882]= -862265664;
assign addr[59883]= -720088517;
assign addr[59884]= -574258580;
assign addr[59885]= -425515602;
assign addr[59886]= -274614114;
assign addr[59887]= -122319591;
assign addr[59888]= 30595422;
assign addr[59889]= 183355234;
assign addr[59890]= 335184940;
assign addr[59891]= 485314355;
assign addr[59892]= 632981917;
assign addr[59893]= 777438554;
assign addr[59894]= 917951481;
assign addr[59895]= 1053807919;
assign addr[59896]= 1184318708;
assign addr[59897]= 1308821808;
assign addr[59898]= 1426685652;
assign addr[59899]= 1537312353;
assign addr[59900]= 1640140734;
assign addr[59901]= 1734649179;
assign addr[59902]= 1820358275;
assign addr[59903]= 1896833245;
assign addr[59904]= 1963686155;
assign addr[59905]= 2020577882;
assign addr[59906]= 2067219829;
assign addr[59907]= 2103375398;
assign addr[59908]= 2128861181;
assign addr[59909]= 2143547897;
assign addr[59910]= 2147361045;
assign addr[59911]= 2140281282;
assign addr[59912]= 2122344521;
assign addr[59913]= 2093641749;
assign addr[59914]= 2054318569;
assign addr[59915]= 2004574453;
assign addr[59916]= 1944661739;
assign addr[59917]= 1874884346;
assign addr[59918]= 1795596234;
assign addr[59919]= 1707199606;
assign addr[59920]= 1610142873;
assign addr[59921]= 1504918373;
assign addr[59922]= 1392059879;
assign addr[59923]= 1272139887;
assign addr[59924]= 1145766716;
assign addr[59925]= 1013581418;
assign addr[59926]= 876254528;
assign addr[59927]= 734482665;
assign addr[59928]= 588984994;
assign addr[59929]= 440499581;
assign addr[59930]= 289779648;
assign addr[59931]= 137589750;
assign addr[59932]= -15298099;
assign addr[59933]= -168108346;
assign addr[59934]= -320065829;
assign addr[59935]= -470399716;
assign addr[59936]= -618347408;
assign addr[59937]= -763158411;
assign addr[59938]= -904098143;
assign addr[59939]= -1040451659;
assign addr[59940]= -1171527280;
assign addr[59941]= -1296660098;
assign addr[59942]= -1415215352;
assign addr[59943]= -1526591649;
assign addr[59944]= -1630224009;
assign addr[59945]= -1725586737;
assign addr[59946]= -1812196087;
assign addr[59947]= -1889612716;
assign addr[59948]= -1957443913;
assign addr[59949]= -2015345591;
assign addr[59950]= -2063024031;
assign addr[59951]= -2100237377;
assign addr[59952]= -2126796855;
assign addr[59953]= -2142567738;
assign addr[59954]= -2147470025;
assign addr[59955]= -2141478848;
assign addr[59956]= -2124624598;
assign addr[59957]= -2096992772;
assign addr[59958]= -2058723538;
assign addr[59959]= -2010011024;
assign addr[59960]= -1951102334;
assign addr[59961]= -1882296293;
assign addr[59962]= -1803941934;
assign addr[59963]= -1716436725;
assign addr[59964]= -1620224553;
assign addr[59965]= -1515793473;
assign addr[59966]= -1403673233;
assign addr[59967]= -1284432584;
assign addr[59968]= -1158676398;
assign addr[59969]= -1027042599;
assign addr[59970]= -890198924;
assign addr[59971]= -748839539;
assign addr[59972]= -603681519;
assign addr[59973]= -455461206;
assign addr[59974]= -304930476;
assign addr[59975]= -152852926;
assign addr[59976]= 0;
assign addr[59977]= 152852926;
assign addr[59978]= 304930476;
assign addr[59979]= 455461206;
assign addr[59980]= 603681519;
assign addr[59981]= 748839539;
assign addr[59982]= 890198924;
assign addr[59983]= 1027042599;
assign addr[59984]= 1158676398;
assign addr[59985]= 1284432584;
assign addr[59986]= 1403673233;
assign addr[59987]= 1515793473;
assign addr[59988]= 1620224553;
assign addr[59989]= 1716436725;
assign addr[59990]= 1803941934;
assign addr[59991]= 1882296293;
assign addr[59992]= 1951102334;
assign addr[59993]= 2010011024;
assign addr[59994]= 2058723538;
assign addr[59995]= 2096992772;
assign addr[59996]= 2124624598;
assign addr[59997]= 2141478848;
assign addr[59998]= 2147470025;
assign addr[59999]= 2142567738;
assign addr[60000]= 2126796855;
assign addr[60001]= 2100237377;
assign addr[60002]= 2063024031;
assign addr[60003]= 2015345591;
assign addr[60004]= 1957443913;
assign addr[60005]= 1889612716;
assign addr[60006]= 1812196087;
assign addr[60007]= 1725586737;
assign addr[60008]= 1630224009;
assign addr[60009]= 1526591649;
assign addr[60010]= 1415215352;
assign addr[60011]= 1296660098;
assign addr[60012]= 1171527280;
assign addr[60013]= 1040451659;
assign addr[60014]= 904098143;
assign addr[60015]= 763158411;
assign addr[60016]= 618347408;
assign addr[60017]= 470399716;
assign addr[60018]= 320065829;
assign addr[60019]= 168108346;
assign addr[60020]= 15298099;
assign addr[60021]= -137589750;
assign addr[60022]= -289779648;
assign addr[60023]= -440499581;
assign addr[60024]= -588984994;
assign addr[60025]= -734482665;
assign addr[60026]= -876254528;
assign addr[60027]= -1013581418;
assign addr[60028]= -1145766716;
assign addr[60029]= -1272139887;
assign addr[60030]= -1392059879;
assign addr[60031]= -1504918373;
assign addr[60032]= -1610142873;
assign addr[60033]= -1707199606;
assign addr[60034]= -1795596234;
assign addr[60035]= -1874884346;
assign addr[60036]= -1944661739;
assign addr[60037]= -2004574453;
assign addr[60038]= -2054318569;
assign addr[60039]= -2093641749;
assign addr[60040]= -2122344521;
assign addr[60041]= -2140281282;
assign addr[60042]= -2147361045;
assign addr[60043]= -2143547897;
assign addr[60044]= -2128861181;
assign addr[60045]= -2103375398;
assign addr[60046]= -2067219829;
assign addr[60047]= -2020577882;
assign addr[60048]= -1963686155;
assign addr[60049]= -1896833245;
assign addr[60050]= -1820358275;
assign addr[60051]= -1734649179;
assign addr[60052]= -1640140734;
assign addr[60053]= -1537312353;
assign addr[60054]= -1426685652;
assign addr[60055]= -1308821808;
assign addr[60056]= -1184318708;
assign addr[60057]= -1053807919;
assign addr[60058]= -917951481;
assign addr[60059]= -777438554;
assign addr[60060]= -632981917;
assign addr[60061]= -485314355;
assign addr[60062]= -335184940;
assign addr[60063]= -183355234;
assign addr[60064]= -30595422;
assign addr[60065]= 122319591;
assign addr[60066]= 274614114;
assign addr[60067]= 425515602;
assign addr[60068]= 574258580;
assign addr[60069]= 720088517;
assign addr[60070]= 862265664;
assign addr[60071]= 1000068799;
assign addr[60072]= 1132798888;
assign addr[60073]= 1259782632;
assign addr[60074]= 1380375881;
assign addr[60075]= 1493966902;
assign addr[60076]= 1599979481;
assign addr[60077]= 1697875851;
assign addr[60078]= 1787159411;
assign addr[60079]= 1867377253;
assign addr[60080]= 1938122457;
assign addr[60081]= 1999036154;
assign addr[60082]= 2049809346;
assign addr[60083]= 2090184478;
assign addr[60084]= 2119956737;
assign addr[60085]= 2138975100;
assign addr[60086]= 2147143090;
assign addr[60087]= 2144419275;
assign addr[60088]= 2130817471;
assign addr[60089]= 2106406677;
assign addr[60090]= 2071310720;
assign addr[60091]= 2025707632;
assign addr[60092]= 1969828744;
assign addr[60093]= 1903957513;
assign addr[60094]= 1828428082;
assign addr[60095]= 1743623590;
assign addr[60096]= 1649974225;
assign addr[60097]= 1547955041;
assign addr[60098]= 1438083551;
assign addr[60099]= 1320917099;
assign addr[60100]= 1197050035;
assign addr[60101]= 1067110699;
assign addr[60102]= 931758235;
assign addr[60103]= 791679244;
assign addr[60104]= 647584304;
assign addr[60105]= 500204365;
assign addr[60106]= 350287041;
assign addr[60107]= 198592817;
assign addr[60108]= 45891193;
assign addr[60109]= -107043224;
assign addr[60110]= -259434643;
assign addr[60111]= -410510029;
assign addr[60112]= -559503022;
assign addr[60113]= -705657826;
assign addr[60114]= -848233042;
assign addr[60115]= -986505429;
assign addr[60116]= -1119773573;
assign addr[60117]= -1247361445;
assign addr[60118]= -1368621831;
assign addr[60119]= -1482939614;
assign addr[60120]= -1589734894;
assign addr[60121]= -1688465931;
assign addr[60122]= -1778631892;
assign addr[60123]= -1859775393;
assign addr[60124]= -1931484818;
assign addr[60125]= -1993396407;
assign addr[60126]= -2045196100;
assign addr[60127]= -2086621133;
assign addr[60128]= -2117461370;
assign addr[60129]= -2137560369;
assign addr[60130]= -2146816171;
assign addr[60131]= -2145181827;
assign addr[60132]= -2132665626;
assign addr[60133]= -2109331059;
assign addr[60134]= -2075296495;
assign addr[60135]= -2030734582;
assign addr[60136]= -1975871368;
assign addr[60137]= -1910985158;
assign addr[60138]= -1836405100;
assign addr[60139]= -1752509516;
assign addr[60140]= -1659723983;
assign addr[60141]= -1558519173;
assign addr[60142]= -1449408469;
assign addr[60143]= -1332945355;
assign addr[60144]= -1209720613;
assign addr[60145]= -1080359326;
assign addr[60146]= -945517704;
assign addr[60147]= -805879757;
assign addr[60148]= -662153826;
assign addr[60149]= -515068990;
assign addr[60150]= -365371365;
assign addr[60151]= -213820322;
assign addr[60152]= -61184634;
assign addr[60153]= 91761426;
assign addr[60154]= 244242007;
assign addr[60155]= 395483624;
assign addr[60156]= 544719071;
assign addr[60157]= 691191324;
assign addr[60158]= 834157373;
assign addr[60159]= 972891995;
assign addr[60160]= 1106691431;
assign addr[60161]= 1234876957;
assign addr[60162]= 1356798326;
assign addr[60163]= 1471837070;
assign addr[60164]= 1579409630;
assign addr[60165]= 1678970324;
assign addr[60166]= 1770014111;
assign addr[60167]= 1852079154;
assign addr[60168]= 1924749160;
assign addr[60169]= 1987655498;
assign addr[60170]= 2040479063;
assign addr[60171]= 2082951896;
assign addr[60172]= 2114858546;
assign addr[60173]= 2136037160;
assign addr[60174]= 2146380306;
assign addr[60175]= 2145835515;
assign addr[60176]= 2134405552;
assign addr[60177]= 2112148396;
assign addr[60178]= 2079176953;
assign addr[60179]= 2035658475;
assign addr[60180]= 1981813720;
assign addr[60181]= 1917915825;
assign addr[60182]= 1844288924;
assign addr[60183]= 1761306505;
assign addr[60184]= 1669389513;
assign addr[60185]= 1569004214;
assign addr[60186]= 1460659832;
assign addr[60187]= 1344905966;
assign addr[60188]= 1222329801;
assign addr[60189]= 1093553126;
assign addr[60190]= 959229189;
assign addr[60191]= 820039373;
assign addr[60192]= 676689746;
assign addr[60193]= 529907477;
assign addr[60194]= 380437148;
assign addr[60195]= 229036977;
assign addr[60196]= 76474970;
assign addr[60197]= -76474970;
assign addr[60198]= -229036977;
assign addr[60199]= -380437148;
assign addr[60200]= -529907477;
assign addr[60201]= -676689746;
assign addr[60202]= -820039373;
assign addr[60203]= -959229189;
assign addr[60204]= -1093553126;
assign addr[60205]= -1222329801;
assign addr[60206]= -1344905966;
assign addr[60207]= -1460659832;
assign addr[60208]= -1569004214;
assign addr[60209]= -1669389513;
assign addr[60210]= -1761306505;
assign addr[60211]= -1844288924;
assign addr[60212]= -1917915825;
assign addr[60213]= -1981813720;
assign addr[60214]= -2035658475;
assign addr[60215]= -2079176953;
assign addr[60216]= -2112148396;
assign addr[60217]= -2134405552;
assign addr[60218]= -2145835515;
assign addr[60219]= -2146380306;
assign addr[60220]= -2136037160;
assign addr[60221]= -2114858546;
assign addr[60222]= -2082951896;
assign addr[60223]= -2040479063;
assign addr[60224]= -1987655498;
assign addr[60225]= -1924749160;
assign addr[60226]= -1852079154;
assign addr[60227]= -1770014111;
assign addr[60228]= -1678970324;
assign addr[60229]= -1579409630;
assign addr[60230]= -1471837070;
assign addr[60231]= -1356798326;
assign addr[60232]= -1234876957;
assign addr[60233]= -1106691431;
assign addr[60234]= -972891995;
assign addr[60235]= -834157373;
assign addr[60236]= -691191324;
assign addr[60237]= -544719071;
assign addr[60238]= -395483624;
assign addr[60239]= -244242007;
assign addr[60240]= -91761426;
assign addr[60241]= 61184634;
assign addr[60242]= 213820322;
assign addr[60243]= 365371365;
assign addr[60244]= 515068990;
assign addr[60245]= 662153826;
assign addr[60246]= 805879757;
assign addr[60247]= 945517704;
assign addr[60248]= 1080359326;
assign addr[60249]= 1209720613;
assign addr[60250]= 1332945355;
assign addr[60251]= 1449408469;
assign addr[60252]= 1558519173;
assign addr[60253]= 1659723983;
assign addr[60254]= 1752509516;
assign addr[60255]= 1836405100;
assign addr[60256]= 1910985158;
assign addr[60257]= 1975871368;
assign addr[60258]= 2030734582;
assign addr[60259]= 2075296495;
assign addr[60260]= 2109331059;
assign addr[60261]= 2132665626;
assign addr[60262]= 2145181827;
assign addr[60263]= 2146816171;
assign addr[60264]= 2137560369;
assign addr[60265]= 2117461370;
assign addr[60266]= 2086621133;
assign addr[60267]= 2045196100;
assign addr[60268]= 1993396407;
assign addr[60269]= 1931484818;
assign addr[60270]= 1859775393;
assign addr[60271]= 1778631892;
assign addr[60272]= 1688465931;
assign addr[60273]= 1589734894;
assign addr[60274]= 1482939614;
assign addr[60275]= 1368621831;
assign addr[60276]= 1247361445;
assign addr[60277]= 1119773573;
assign addr[60278]= 986505429;
assign addr[60279]= 848233042;
assign addr[60280]= 705657826;
assign addr[60281]= 559503022;
assign addr[60282]= 410510029;
assign addr[60283]= 259434643;
assign addr[60284]= 107043224;
assign addr[60285]= -45891193;
assign addr[60286]= -198592817;
assign addr[60287]= -350287041;
assign addr[60288]= -500204365;
assign addr[60289]= -647584304;
assign addr[60290]= -791679244;
assign addr[60291]= -931758235;
assign addr[60292]= -1067110699;
assign addr[60293]= -1197050035;
assign addr[60294]= -1320917099;
assign addr[60295]= -1438083551;
assign addr[60296]= -1547955041;
assign addr[60297]= -1649974225;
assign addr[60298]= -1743623590;
assign addr[60299]= -1828428082;
assign addr[60300]= -1903957513;
assign addr[60301]= -1969828744;
assign addr[60302]= -2025707632;
assign addr[60303]= -2071310720;
assign addr[60304]= -2106406677;
assign addr[60305]= -2130817471;
assign addr[60306]= -2144419275;
assign addr[60307]= -2147143090;
assign addr[60308]= -2138975100;
assign addr[60309]= -2119956737;
assign addr[60310]= -2090184478;
assign addr[60311]= -2049809346;
assign addr[60312]= -1999036154;
assign addr[60313]= -1938122457;
assign addr[60314]= -1867377253;
assign addr[60315]= -1787159411;
assign addr[60316]= -1697875851;
assign addr[60317]= -1599979481;
assign addr[60318]= -1493966902;
assign addr[60319]= -1380375881;
assign addr[60320]= -1259782632;
assign addr[60321]= -1132798888;
assign addr[60322]= -1000068799;
assign addr[60323]= -862265664;
assign addr[60324]= -720088517;
assign addr[60325]= -574258580;
assign addr[60326]= -425515602;
assign addr[60327]= -274614114;
assign addr[60328]= -122319591;
assign addr[60329]= 30595422;
assign addr[60330]= 183355234;
assign addr[60331]= 335184940;
assign addr[60332]= 485314355;
assign addr[60333]= 632981917;
assign addr[60334]= 777438554;
assign addr[60335]= 917951481;
assign addr[60336]= 1053807919;
assign addr[60337]= 1184318708;
assign addr[60338]= 1308821808;
assign addr[60339]= 1426685652;
assign addr[60340]= 1537312353;
assign addr[60341]= 1640140734;
assign addr[60342]= 1734649179;
assign addr[60343]= 1820358275;
assign addr[60344]= 1896833245;
assign addr[60345]= 1963686155;
assign addr[60346]= 2020577882;
assign addr[60347]= 2067219829;
assign addr[60348]= 2103375398;
assign addr[60349]= 2128861181;
assign addr[60350]= 2143547897;
assign addr[60351]= 2147361045;
assign addr[60352]= 2140281282;
assign addr[60353]= 2122344521;
assign addr[60354]= 2093641749;
assign addr[60355]= 2054318569;
assign addr[60356]= 2004574453;
assign addr[60357]= 1944661739;
assign addr[60358]= 1874884346;
assign addr[60359]= 1795596234;
assign addr[60360]= 1707199606;
assign addr[60361]= 1610142873;
assign addr[60362]= 1504918373;
assign addr[60363]= 1392059879;
assign addr[60364]= 1272139887;
assign addr[60365]= 1145766716;
assign addr[60366]= 1013581418;
assign addr[60367]= 876254528;
assign addr[60368]= 734482665;
assign addr[60369]= 588984994;
assign addr[60370]= 440499581;
assign addr[60371]= 289779648;
assign addr[60372]= 137589750;
assign addr[60373]= -15298099;
assign addr[60374]= -168108346;
assign addr[60375]= -320065829;
assign addr[60376]= -470399716;
assign addr[60377]= -618347408;
assign addr[60378]= -763158411;
assign addr[60379]= -904098143;
assign addr[60380]= -1040451659;
assign addr[60381]= -1171527280;
assign addr[60382]= -1296660098;
assign addr[60383]= -1415215352;
assign addr[60384]= -1526591649;
assign addr[60385]= -1630224009;
assign addr[60386]= -1725586737;
assign addr[60387]= -1812196087;
assign addr[60388]= -1889612716;
assign addr[60389]= -1957443913;
assign addr[60390]= -2015345591;
assign addr[60391]= -2063024031;
assign addr[60392]= -2100237377;
assign addr[60393]= -2126796855;
assign addr[60394]= -2142567738;
assign addr[60395]= -2147470025;
assign addr[60396]= -2141478848;
assign addr[60397]= -2124624598;
assign addr[60398]= -2096992772;
assign addr[60399]= -2058723538;
assign addr[60400]= -2010011024;
assign addr[60401]= -1951102334;
assign addr[60402]= -1882296293;
assign addr[60403]= -1803941934;
assign addr[60404]= -1716436725;
assign addr[60405]= -1620224553;
assign addr[60406]= -1515793473;
assign addr[60407]= -1403673233;
assign addr[60408]= -1284432584;
assign addr[60409]= -1158676398;
assign addr[60410]= -1027042599;
assign addr[60411]= -890198924;
assign addr[60412]= -748839539;
assign addr[60413]= -603681519;
assign addr[60414]= -455461206;
assign addr[60415]= -304930476;
assign addr[60416]= -152852926;
assign addr[60417]= 0;
assign addr[60418]= 152852926;
assign addr[60419]= 304930476;
assign addr[60420]= 455461206;
assign addr[60421]= 603681519;
assign addr[60422]= 748839539;
assign addr[60423]= 890198924;
assign addr[60424]= 1027042599;
assign addr[60425]= 1158676398;
assign addr[60426]= 1284432584;
assign addr[60427]= 1403673233;
assign addr[60428]= 1515793473;
assign addr[60429]= 1620224553;
assign addr[60430]= 1716436725;
assign addr[60431]= 1803941934;
assign addr[60432]= 1882296293;
assign addr[60433]= 1951102334;
assign addr[60434]= 2010011024;
assign addr[60435]= 2058723538;
assign addr[60436]= 2096992772;
assign addr[60437]= 2124624598;
assign addr[60438]= 2141478848;
assign addr[60439]= 2147470025;
assign addr[60440]= 2142567738;
assign addr[60441]= 2126796855;
assign addr[60442]= 2100237377;
assign addr[60443]= 2063024031;
assign addr[60444]= 2015345591;
assign addr[60445]= 1957443913;
assign addr[60446]= 1889612716;
assign addr[60447]= 1812196087;
assign addr[60448]= 1725586737;
assign addr[60449]= 1630224009;
assign addr[60450]= 1526591649;
assign addr[60451]= 1415215352;
assign addr[60452]= 1296660098;
assign addr[60453]= 1171527280;
assign addr[60454]= 1040451659;
assign addr[60455]= 904098143;
assign addr[60456]= 763158411;
assign addr[60457]= 618347408;
assign addr[60458]= 470399716;
assign addr[60459]= 320065829;
assign addr[60460]= 168108346;
assign addr[60461]= 15298099;
assign addr[60462]= -137589750;
assign addr[60463]= -289779648;
assign addr[60464]= -440499581;
assign addr[60465]= -588984994;
assign addr[60466]= -734482665;
assign addr[60467]= -876254528;
assign addr[60468]= -1013581418;
assign addr[60469]= -1145766716;
assign addr[60470]= -1272139887;
assign addr[60471]= -1392059879;
assign addr[60472]= -1504918373;
assign addr[60473]= -1610142873;
assign addr[60474]= -1707199606;
assign addr[60475]= -1795596234;
assign addr[60476]= -1874884346;
assign addr[60477]= -1944661739;
assign addr[60478]= -2004574453;
assign addr[60479]= -2054318569;
assign addr[60480]= -2093641749;
assign addr[60481]= -2122344521;
assign addr[60482]= -2140281282;
assign addr[60483]= -2147361045;
assign addr[60484]= -2143547897;
assign addr[60485]= -2128861181;
assign addr[60486]= -2103375398;
assign addr[60487]= -2067219829;
assign addr[60488]= -2020577882;
assign addr[60489]= -1963686155;
assign addr[60490]= -1896833245;
assign addr[60491]= -1820358275;
assign addr[60492]= -1734649179;
assign addr[60493]= -1640140734;
assign addr[60494]= -1537312353;
assign addr[60495]= -1426685652;
assign addr[60496]= -1308821808;
assign addr[60497]= -1184318708;
assign addr[60498]= -1053807919;
assign addr[60499]= -917951481;
assign addr[60500]= -777438554;
assign addr[60501]= -632981917;
assign addr[60502]= -485314355;
assign addr[60503]= -335184940;
assign addr[60504]= -183355234;
assign addr[60505]= -30595422;
assign addr[60506]= 122319591;
assign addr[60507]= 274614114;
assign addr[60508]= 425515602;
assign addr[60509]= 574258580;
assign addr[60510]= 720088517;
assign addr[60511]= 862265664;
assign addr[60512]= 1000068799;
assign addr[60513]= 1132798888;
assign addr[60514]= 1259782632;
assign addr[60515]= 1380375881;
assign addr[60516]= 1493966902;
assign addr[60517]= 1599979481;
assign addr[60518]= 1697875851;
assign addr[60519]= 1787159411;
assign addr[60520]= 1867377253;
assign addr[60521]= 1938122457;
assign addr[60522]= 1999036154;
assign addr[60523]= 2049809346;
assign addr[60524]= 2090184478;
assign addr[60525]= 2119956737;
assign addr[60526]= 2138975100;
assign addr[60527]= 2147143090;
assign addr[60528]= 2144419275;
assign addr[60529]= 2130817471;
assign addr[60530]= 2106406677;
assign addr[60531]= 2071310720;
assign addr[60532]= 2025707632;
assign addr[60533]= 1969828744;
assign addr[60534]= 1903957513;
assign addr[60535]= 1828428082;
assign addr[60536]= 1743623590;
assign addr[60537]= 1649974225;
assign addr[60538]= 1547955041;
assign addr[60539]= 1438083551;
assign addr[60540]= 1320917099;
assign addr[60541]= 1197050035;
assign addr[60542]= 1067110699;
assign addr[60543]= 931758235;
assign addr[60544]= 791679244;
assign addr[60545]= 647584304;
assign addr[60546]= 500204365;
assign addr[60547]= 350287041;
assign addr[60548]= 198592817;
assign addr[60549]= 45891193;
assign addr[60550]= -107043224;
assign addr[60551]= -259434643;
assign addr[60552]= -410510029;
assign addr[60553]= -559503022;
assign addr[60554]= -705657826;
assign addr[60555]= -848233042;
assign addr[60556]= -986505429;
assign addr[60557]= -1119773573;
assign addr[60558]= -1247361445;
assign addr[60559]= -1368621831;
assign addr[60560]= -1482939614;
assign addr[60561]= -1589734894;
assign addr[60562]= -1688465931;
assign addr[60563]= -1778631892;
assign addr[60564]= -1859775393;
assign addr[60565]= -1931484818;
assign addr[60566]= -1993396407;
assign addr[60567]= -2045196100;
assign addr[60568]= -2086621133;
assign addr[60569]= -2117461370;
assign addr[60570]= -2137560369;
assign addr[60571]= -2146816171;
assign addr[60572]= -2145181827;
assign addr[60573]= -2132665626;
assign addr[60574]= -2109331059;
assign addr[60575]= -2075296495;
assign addr[60576]= -2030734582;
assign addr[60577]= -1975871368;
assign addr[60578]= -1910985158;
assign addr[60579]= -1836405100;
assign addr[60580]= -1752509516;
assign addr[60581]= -1659723983;
assign addr[60582]= -1558519173;
assign addr[60583]= -1449408469;
assign addr[60584]= -1332945355;
assign addr[60585]= -1209720613;
assign addr[60586]= -1080359326;
assign addr[60587]= -945517704;
assign addr[60588]= -805879757;
assign addr[60589]= -662153826;
assign addr[60590]= -515068990;
assign addr[60591]= -365371365;
assign addr[60592]= -213820322;
assign addr[60593]= -61184634;
assign addr[60594]= 91761426;
assign addr[60595]= 244242007;
assign addr[60596]= 395483624;
assign addr[60597]= 544719071;
assign addr[60598]= 691191324;
assign addr[60599]= 834157373;
assign addr[60600]= 972891995;
assign addr[60601]= 1106691431;
assign addr[60602]= 1234876957;
assign addr[60603]= 1356798326;
assign addr[60604]= 1471837070;
assign addr[60605]= 1579409630;
assign addr[60606]= 1678970324;
assign addr[60607]= 1770014111;
assign addr[60608]= 1852079154;
assign addr[60609]= 1924749160;
assign addr[60610]= 1987655498;
assign addr[60611]= 2040479063;
assign addr[60612]= 2082951896;
assign addr[60613]= 2114858546;
assign addr[60614]= 2136037160;
assign addr[60615]= 2146380306;
assign addr[60616]= 2145835515;
assign addr[60617]= 2134405552;
assign addr[60618]= 2112148396;
assign addr[60619]= 2079176953;
assign addr[60620]= 2035658475;
assign addr[60621]= 1981813720;
assign addr[60622]= 1917915825;
assign addr[60623]= 1844288924;
assign addr[60624]= 1761306505;
assign addr[60625]= 1669389513;
assign addr[60626]= 1569004214;
assign addr[60627]= 1460659832;
assign addr[60628]= 1344905966;
assign addr[60629]= 1222329801;
assign addr[60630]= 1093553126;
assign addr[60631]= 959229189;
assign addr[60632]= 820039373;
assign addr[60633]= 676689746;
assign addr[60634]= 529907477;
assign addr[60635]= 380437148;
assign addr[60636]= 229036977;
assign addr[60637]= 76474970;
assign addr[60638]= -76474970;
assign addr[60639]= -229036977;
assign addr[60640]= -380437148;
assign addr[60641]= -529907477;
assign addr[60642]= -676689746;
assign addr[60643]= -820039373;
assign addr[60644]= -959229189;
assign addr[60645]= -1093553126;
assign addr[60646]= -1222329801;
assign addr[60647]= -1344905966;
assign addr[60648]= -1460659832;
assign addr[60649]= -1569004214;
assign addr[60650]= -1669389513;
assign addr[60651]= -1761306505;
assign addr[60652]= -1844288924;
assign addr[60653]= -1917915825;
assign addr[60654]= -1981813720;
assign addr[60655]= -2035658475;
assign addr[60656]= -2079176953;
assign addr[60657]= -2112148396;
assign addr[60658]= -2134405552;
assign addr[60659]= -2145835515;
assign addr[60660]= -2146380306;
assign addr[60661]= -2136037160;
assign addr[60662]= -2114858546;
assign addr[60663]= -2082951896;
assign addr[60664]= -2040479063;
assign addr[60665]= -1987655498;
assign addr[60666]= -1924749160;
assign addr[60667]= -1852079154;
assign addr[60668]= -1770014111;
assign addr[60669]= -1678970324;
assign addr[60670]= -1579409630;
assign addr[60671]= -1471837070;
assign addr[60672]= -1356798326;
assign addr[60673]= -1234876957;
assign addr[60674]= -1106691431;
assign addr[60675]= -972891995;
assign addr[60676]= -834157373;
assign addr[60677]= -691191324;
assign addr[60678]= -544719071;
assign addr[60679]= -395483624;
assign addr[60680]= -244242007;
assign addr[60681]= -91761426;
assign addr[60682]= 61184634;
assign addr[60683]= 213820322;
assign addr[60684]= 365371365;
assign addr[60685]= 515068990;
assign addr[60686]= 662153826;
assign addr[60687]= 805879757;
assign addr[60688]= 945517704;
assign addr[60689]= 1080359326;
assign addr[60690]= 1209720613;
assign addr[60691]= 1332945355;
assign addr[60692]= 1449408469;
assign addr[60693]= 1558519173;
assign addr[60694]= 1659723983;
assign addr[60695]= 1752509516;
assign addr[60696]= 1836405100;
assign addr[60697]= 1910985158;
assign addr[60698]= 1975871368;
assign addr[60699]= 2030734582;
assign addr[60700]= 2075296495;
assign addr[60701]= 2109331059;
assign addr[60702]= 2132665626;
assign addr[60703]= 2145181827;
assign addr[60704]= 2146816171;
assign addr[60705]= 2137560369;
assign addr[60706]= 2117461370;
assign addr[60707]= 2086621133;
assign addr[60708]= 2045196100;
assign addr[60709]= 1993396407;
assign addr[60710]= 1931484818;
assign addr[60711]= 1859775393;
assign addr[60712]= 1778631892;
assign addr[60713]= 1688465931;
assign addr[60714]= 1589734894;
assign addr[60715]= 1482939614;
assign addr[60716]= 1368621831;
assign addr[60717]= 1247361445;
assign addr[60718]= 1119773573;
assign addr[60719]= 986505429;
assign addr[60720]= 848233042;
assign addr[60721]= 705657826;
assign addr[60722]= 559503022;
assign addr[60723]= 410510029;
assign addr[60724]= 259434643;
assign addr[60725]= 107043224;
assign addr[60726]= -45891193;
assign addr[60727]= -198592817;
assign addr[60728]= -350287041;
assign addr[60729]= -500204365;
assign addr[60730]= -647584304;
assign addr[60731]= -791679244;
assign addr[60732]= -931758235;
assign addr[60733]= -1067110699;
assign addr[60734]= -1197050035;
assign addr[60735]= -1320917099;
assign addr[60736]= -1438083551;
assign addr[60737]= -1547955041;
assign addr[60738]= -1649974225;
assign addr[60739]= -1743623590;
assign addr[60740]= -1828428082;
assign addr[60741]= -1903957513;
assign addr[60742]= -1969828744;
assign addr[60743]= -2025707632;
assign addr[60744]= -2071310720;
assign addr[60745]= -2106406677;
assign addr[60746]= -2130817471;
assign addr[60747]= -2144419275;
assign addr[60748]= -2147143090;
assign addr[60749]= -2138975100;
assign addr[60750]= -2119956737;
assign addr[60751]= -2090184478;
assign addr[60752]= -2049809346;
assign addr[60753]= -1999036154;
assign addr[60754]= -1938122457;
assign addr[60755]= -1867377253;
assign addr[60756]= -1787159411;
assign addr[60757]= -1697875851;
assign addr[60758]= -1599979481;
assign addr[60759]= -1493966902;
assign addr[60760]= -1380375881;
assign addr[60761]= -1259782632;
assign addr[60762]= -1132798888;
assign addr[60763]= -1000068799;
assign addr[60764]= -862265664;
assign addr[60765]= -720088517;
assign addr[60766]= -574258580;
assign addr[60767]= -425515602;
assign addr[60768]= -274614114;
assign addr[60769]= -122319591;
assign addr[60770]= 30595422;
assign addr[60771]= 183355234;
assign addr[60772]= 335184940;
assign addr[60773]= 485314355;
assign addr[60774]= 632981917;
assign addr[60775]= 777438554;
assign addr[60776]= 917951481;
assign addr[60777]= 1053807919;
assign addr[60778]= 1184318708;
assign addr[60779]= 1308821808;
assign addr[60780]= 1426685652;
assign addr[60781]= 1537312353;
assign addr[60782]= 1640140734;
assign addr[60783]= 1734649179;
assign addr[60784]= 1820358275;
assign addr[60785]= 1896833245;
assign addr[60786]= 1963686155;
assign addr[60787]= 2020577882;
assign addr[60788]= 2067219829;
assign addr[60789]= 2103375398;
assign addr[60790]= 2128861181;
assign addr[60791]= 2143547897;
assign addr[60792]= 2147361045;
assign addr[60793]= 2140281282;
assign addr[60794]= 2122344521;
assign addr[60795]= 2093641749;
assign addr[60796]= 2054318569;
assign addr[60797]= 2004574453;
assign addr[60798]= 1944661739;
assign addr[60799]= 1874884346;
assign addr[60800]= 1795596234;
assign addr[60801]= 1707199606;
assign addr[60802]= 1610142873;
assign addr[60803]= 1504918373;
assign addr[60804]= 1392059879;
assign addr[60805]= 1272139887;
assign addr[60806]= 1145766716;
assign addr[60807]= 1013581418;
assign addr[60808]= 876254528;
assign addr[60809]= 734482665;
assign addr[60810]= 588984994;
assign addr[60811]= 440499581;
assign addr[60812]= 289779648;
assign addr[60813]= 137589750;
assign addr[60814]= -15298099;
assign addr[60815]= -168108346;
assign addr[60816]= -320065829;
assign addr[60817]= -470399716;
assign addr[60818]= -618347408;
assign addr[60819]= -763158411;
assign addr[60820]= -904098143;
assign addr[60821]= -1040451659;
assign addr[60822]= -1171527280;
assign addr[60823]= -1296660098;
assign addr[60824]= -1415215352;
assign addr[60825]= -1526591649;
assign addr[60826]= -1630224009;
assign addr[60827]= -1725586737;
assign addr[60828]= -1812196087;
assign addr[60829]= -1889612716;
assign addr[60830]= -1957443913;
assign addr[60831]= -2015345591;
assign addr[60832]= -2063024031;
assign addr[60833]= -2100237377;
assign addr[60834]= -2126796855;
assign addr[60835]= -2142567738;
assign addr[60836]= -2147470025;
assign addr[60837]= -2141478848;
assign addr[60838]= -2124624598;
assign addr[60839]= -2096992772;
assign addr[60840]= -2058723538;
assign addr[60841]= -2010011024;
assign addr[60842]= -1951102334;
assign addr[60843]= -1882296293;
assign addr[60844]= -1803941934;
assign addr[60845]= -1716436725;
assign addr[60846]= -1620224553;
assign addr[60847]= -1515793473;
assign addr[60848]= -1403673233;
assign addr[60849]= -1284432584;
assign addr[60850]= -1158676398;
assign addr[60851]= -1027042599;
assign addr[60852]= -890198924;
assign addr[60853]= -748839539;
assign addr[60854]= -603681519;
assign addr[60855]= -455461206;
assign addr[60856]= -304930476;
assign addr[60857]= -152852926;
assign addr[60858]= 0;
assign addr[60859]= 152852926;
assign addr[60860]= 304930476;
assign addr[60861]= 455461206;
assign addr[60862]= 603681519;
assign addr[60863]= 748839539;
assign addr[60864]= 890198924;
assign addr[60865]= 1027042599;
assign addr[60866]= 1158676398;
assign addr[60867]= 1284432584;
assign addr[60868]= 1403673233;
assign addr[60869]= 1515793473;
assign addr[60870]= 1620224553;
assign addr[60871]= 1716436725;
assign addr[60872]= 1803941934;
assign addr[60873]= 1882296293;
assign addr[60874]= 1951102334;
assign addr[60875]= 2010011024;
assign addr[60876]= 2058723538;
assign addr[60877]= 2096992772;
assign addr[60878]= 2124624598;
assign addr[60879]= 2141478848;
assign addr[60880]= 2147470025;
assign addr[60881]= 2142567738;
assign addr[60882]= 2126796855;
assign addr[60883]= 2100237377;
assign addr[60884]= 2063024031;
assign addr[60885]= 2015345591;
assign addr[60886]= 1957443913;
assign addr[60887]= 1889612716;
assign addr[60888]= 1812196087;
assign addr[60889]= 1725586737;
assign addr[60890]= 1630224009;
assign addr[60891]= 1526591649;
assign addr[60892]= 1415215352;
assign addr[60893]= 1296660098;
assign addr[60894]= 1171527280;
assign addr[60895]= 1040451659;
assign addr[60896]= 904098143;
assign addr[60897]= 763158411;
assign addr[60898]= 618347408;
assign addr[60899]= 470399716;
assign addr[60900]= 320065829;
assign addr[60901]= 168108346;
assign addr[60902]= 15298099;
assign addr[60903]= -137589750;
assign addr[60904]= -289779648;
assign addr[60905]= -440499581;
assign addr[60906]= -588984994;
assign addr[60907]= -734482665;
assign addr[60908]= -876254528;
assign addr[60909]= -1013581418;
assign addr[60910]= -1145766716;
assign addr[60911]= -1272139887;
assign addr[60912]= -1392059879;
assign addr[60913]= -1504918373;
assign addr[60914]= -1610142873;
assign addr[60915]= -1707199606;
assign addr[60916]= -1795596234;
assign addr[60917]= -1874884346;
assign addr[60918]= -1944661739;
assign addr[60919]= -2004574453;
assign addr[60920]= -2054318569;
assign addr[60921]= -2093641749;
assign addr[60922]= -2122344521;
assign addr[60923]= -2140281282;
assign addr[60924]= -2147361045;
assign addr[60925]= -2143547897;
assign addr[60926]= -2128861181;
assign addr[60927]= -2103375398;
assign addr[60928]= -2067219829;
assign addr[60929]= -2020577882;
assign addr[60930]= -1963686155;
assign addr[60931]= -1896833245;
assign addr[60932]= -1820358275;
assign addr[60933]= -1734649179;
assign addr[60934]= -1640140734;
assign addr[60935]= -1537312353;
assign addr[60936]= -1426685652;
assign addr[60937]= -1308821808;
assign addr[60938]= -1184318708;
assign addr[60939]= -1053807919;
assign addr[60940]= -917951481;
assign addr[60941]= -777438554;
assign addr[60942]= -632981917;
assign addr[60943]= -485314355;
assign addr[60944]= -335184940;
assign addr[60945]= -183355234;
assign addr[60946]= -30595422;
assign addr[60947]= 122319591;
assign addr[60948]= 274614114;
assign addr[60949]= 425515602;
assign addr[60950]= 574258580;
assign addr[60951]= 720088517;
assign addr[60952]= 862265664;
assign addr[60953]= 1000068799;
assign addr[60954]= 1132798888;
assign addr[60955]= 1259782632;
assign addr[60956]= 1380375881;
assign addr[60957]= 1493966902;
assign addr[60958]= 1599979481;
assign addr[60959]= 1697875851;
assign addr[60960]= 1787159411;
assign addr[60961]= 1867377253;
assign addr[60962]= 1938122457;
assign addr[60963]= 1999036154;
assign addr[60964]= 2049809346;
assign addr[60965]= 2090184478;
assign addr[60966]= 2119956737;
assign addr[60967]= 2138975100;
assign addr[60968]= 2147143090;
assign addr[60969]= 2144419275;
assign addr[60970]= 2130817471;
assign addr[60971]= 2106406677;
assign addr[60972]= 2071310720;
assign addr[60973]= 2025707632;
assign addr[60974]= 1969828744;
assign addr[60975]= 1903957513;
assign addr[60976]= 1828428082;
assign addr[60977]= 1743623590;
assign addr[60978]= 1649974225;
assign addr[60979]= 1547955041;
assign addr[60980]= 1438083551;
assign addr[60981]= 1320917099;
assign addr[60982]= 1197050035;
assign addr[60983]= 1067110699;
assign addr[60984]= 931758235;
assign addr[60985]= 791679244;
assign addr[60986]= 647584304;
assign addr[60987]= 500204365;
assign addr[60988]= 350287041;
assign addr[60989]= 198592817;
assign addr[60990]= 45891193;
assign addr[60991]= -107043224;
assign addr[60992]= -259434643;
assign addr[60993]= -410510029;
assign addr[60994]= -559503022;
assign addr[60995]= -705657826;
assign addr[60996]= -848233042;
assign addr[60997]= -986505429;
assign addr[60998]= -1119773573;
assign addr[60999]= -1247361445;
assign addr[61000]= -1368621831;
assign addr[61001]= -1482939614;
assign addr[61002]= -1589734894;
assign addr[61003]= -1688465931;
assign addr[61004]= -1778631892;
assign addr[61005]= -1859775393;
assign addr[61006]= -1931484818;
assign addr[61007]= -1993396407;
assign addr[61008]= -2045196100;
assign addr[61009]= -2086621133;
assign addr[61010]= -2117461370;
assign addr[61011]= -2137560369;
assign addr[61012]= -2146816171;
assign addr[61013]= -2145181827;
assign addr[61014]= -2132665626;
assign addr[61015]= -2109331059;
assign addr[61016]= -2075296495;
assign addr[61017]= -2030734582;
assign addr[61018]= -1975871368;
assign addr[61019]= -1910985158;
assign addr[61020]= -1836405100;
assign addr[61021]= -1752509516;
assign addr[61022]= -1659723983;
assign addr[61023]= -1558519173;
assign addr[61024]= -1449408469;
assign addr[61025]= -1332945355;
assign addr[61026]= -1209720613;
assign addr[61027]= -1080359326;
assign addr[61028]= -945517704;
assign addr[61029]= -805879757;
assign addr[61030]= -662153826;
assign addr[61031]= -515068990;
assign addr[61032]= -365371365;
assign addr[61033]= -213820322;
assign addr[61034]= -61184634;
assign addr[61035]= 91761426;
assign addr[61036]= 244242007;
assign addr[61037]= 395483624;
assign addr[61038]= 544719071;
assign addr[61039]= 691191324;
assign addr[61040]= 834157373;
assign addr[61041]= 972891995;
assign addr[61042]= 1106691431;
assign addr[61043]= 1234876957;
assign addr[61044]= 1356798326;
assign addr[61045]= 1471837070;
assign addr[61046]= 1579409630;
assign addr[61047]= 1678970324;
assign addr[61048]= 1770014111;
assign addr[61049]= 1852079154;
assign addr[61050]= 1924749160;
assign addr[61051]= 1987655498;
assign addr[61052]= 2040479063;
assign addr[61053]= 2082951896;
assign addr[61054]= 2114858546;
assign addr[61055]= 2136037160;
assign addr[61056]= 2146380306;
assign addr[61057]= 2145835515;
assign addr[61058]= 2134405552;
assign addr[61059]= 2112148396;
assign addr[61060]= 2079176953;
assign addr[61061]= 2035658475;
assign addr[61062]= 1981813720;
assign addr[61063]= 1917915825;
assign addr[61064]= 1844288924;
assign addr[61065]= 1761306505;
assign addr[61066]= 1669389513;
assign addr[61067]= 1569004214;
assign addr[61068]= 1460659832;
assign addr[61069]= 1344905966;
assign addr[61070]= 1222329801;
assign addr[61071]= 1093553126;
assign addr[61072]= 959229189;
assign addr[61073]= 820039373;
assign addr[61074]= 676689746;
assign addr[61075]= 529907477;
assign addr[61076]= 380437148;
assign addr[61077]= 229036977;
assign addr[61078]= 76474970;
assign addr[61079]= -76474970;
assign addr[61080]= -229036977;
assign addr[61081]= -380437148;
assign addr[61082]= -529907477;
assign addr[61083]= -676689746;
assign addr[61084]= -820039373;
assign addr[61085]= -959229189;
assign addr[61086]= -1093553126;
assign addr[61087]= -1222329801;
assign addr[61088]= -1344905966;
assign addr[61089]= -1460659832;
assign addr[61090]= -1569004214;
assign addr[61091]= -1669389513;
assign addr[61092]= -1761306505;
assign addr[61093]= -1844288924;
assign addr[61094]= -1917915825;
assign addr[61095]= -1981813720;
assign addr[61096]= -2035658475;
assign addr[61097]= -2079176953;
assign addr[61098]= -2112148396;
assign addr[61099]= -2134405552;
assign addr[61100]= -2145835515;
assign addr[61101]= -2146380306;
assign addr[61102]= -2136037160;
assign addr[61103]= -2114858546;
assign addr[61104]= -2082951896;
assign addr[61105]= -2040479063;
assign addr[61106]= -1987655498;
assign addr[61107]= -1924749160;
assign addr[61108]= -1852079154;
assign addr[61109]= -1770014111;
assign addr[61110]= -1678970324;
assign addr[61111]= -1579409630;
assign addr[61112]= -1471837070;
assign addr[61113]= -1356798326;
assign addr[61114]= -1234876957;
assign addr[61115]= -1106691431;
assign addr[61116]= -972891995;
assign addr[61117]= -834157373;
assign addr[61118]= -691191324;
assign addr[61119]= -544719071;
assign addr[61120]= -395483624;
assign addr[61121]= -244242007;
assign addr[61122]= -91761426;
assign addr[61123]= 61184634;
assign addr[61124]= 213820322;
assign addr[61125]= 365371365;
assign addr[61126]= 515068990;
assign addr[61127]= 662153826;
assign addr[61128]= 805879757;
assign addr[61129]= 945517704;
assign addr[61130]= 1080359326;
assign addr[61131]= 1209720613;
assign addr[61132]= 1332945355;
assign addr[61133]= 1449408469;
assign addr[61134]= 1558519173;
assign addr[61135]= 1659723983;
assign addr[61136]= 1752509516;
assign addr[61137]= 1836405100;
assign addr[61138]= 1910985158;
assign addr[61139]= 1975871368;
assign addr[61140]= 2030734582;
assign addr[61141]= 2075296495;
assign addr[61142]= 2109331059;
assign addr[61143]= 2132665626;
assign addr[61144]= 2145181827;
assign addr[61145]= 2146816171;
assign addr[61146]= 2137560369;
assign addr[61147]= 2117461370;
assign addr[61148]= 2086621133;
assign addr[61149]= 2045196100;
assign addr[61150]= 1993396407;
assign addr[61151]= 1931484818;
assign addr[61152]= 1859775393;
assign addr[61153]= 1778631892;
assign addr[61154]= 1688465931;
assign addr[61155]= 1589734894;
assign addr[61156]= 1482939614;
assign addr[61157]= 1368621831;
assign addr[61158]= 1247361445;
assign addr[61159]= 1119773573;
assign addr[61160]= 986505429;
assign addr[61161]= 848233042;
assign addr[61162]= 705657826;
assign addr[61163]= 559503022;
assign addr[61164]= 410510029;
assign addr[61165]= 259434643;
assign addr[61166]= 107043224;
assign addr[61167]= -45891193;
assign addr[61168]= -198592817;
assign addr[61169]= -350287041;
assign addr[61170]= -500204365;
assign addr[61171]= -647584304;
assign addr[61172]= -791679244;
assign addr[61173]= -931758235;
assign addr[61174]= -1067110699;
assign addr[61175]= -1197050035;
assign addr[61176]= -1320917099;
assign addr[61177]= -1438083551;
assign addr[61178]= -1547955041;
assign addr[61179]= -1649974225;
assign addr[61180]= -1743623590;
assign addr[61181]= -1828428082;
assign addr[61182]= -1903957513;
assign addr[61183]= -1969828744;
assign addr[61184]= -2025707632;
assign addr[61185]= -2071310720;
assign addr[61186]= -2106406677;
assign addr[61187]= -2130817471;
assign addr[61188]= -2144419275;
assign addr[61189]= -2147143090;
assign addr[61190]= -2138975100;
assign addr[61191]= -2119956737;
assign addr[61192]= -2090184478;
assign addr[61193]= -2049809346;
assign addr[61194]= -1999036154;
assign addr[61195]= -1938122457;
assign addr[61196]= -1867377253;
assign addr[61197]= -1787159411;
assign addr[61198]= -1697875851;
assign addr[61199]= -1599979481;
assign addr[61200]= -1493966902;
assign addr[61201]= -1380375881;
assign addr[61202]= -1259782632;
assign addr[61203]= -1132798888;
assign addr[61204]= -1000068799;
assign addr[61205]= -862265664;
assign addr[61206]= -720088517;
assign addr[61207]= -574258580;
assign addr[61208]= -425515602;
assign addr[61209]= -274614114;
assign addr[61210]= -122319591;
assign addr[61211]= 30595422;
assign addr[61212]= 183355234;
assign addr[61213]= 335184940;
assign addr[61214]= 485314355;
assign addr[61215]= 632981917;
assign addr[61216]= 777438554;
assign addr[61217]= 917951481;
assign addr[61218]= 1053807919;
assign addr[61219]= 1184318708;
assign addr[61220]= 1308821808;
assign addr[61221]= 1426685652;
assign addr[61222]= 1537312353;
assign addr[61223]= 1640140734;
assign addr[61224]= 1734649179;
assign addr[61225]= 1820358275;
assign addr[61226]= 1896833245;
assign addr[61227]= 1963686155;
assign addr[61228]= 2020577882;
assign addr[61229]= 2067219829;
assign addr[61230]= 2103375398;
assign addr[61231]= 2128861181;
assign addr[61232]= 2143547897;
assign addr[61233]= 2147361045;
assign addr[61234]= 2140281282;
assign addr[61235]= 2122344521;
assign addr[61236]= 2093641749;
assign addr[61237]= 2054318569;
assign addr[61238]= 2004574453;
assign addr[61239]= 1944661739;
assign addr[61240]= 1874884346;
assign addr[61241]= 1795596234;
assign addr[61242]= 1707199606;
assign addr[61243]= 1610142873;
assign addr[61244]= 1504918373;
assign addr[61245]= 1392059879;
assign addr[61246]= 1272139887;
assign addr[61247]= 1145766716;
assign addr[61248]= 1013581418;
assign addr[61249]= 876254528;
assign addr[61250]= 734482665;
assign addr[61251]= 588984994;
assign addr[61252]= 440499581;
assign addr[61253]= 289779648;
assign addr[61254]= 137589750;
assign addr[61255]= -15298099;
assign addr[61256]= -168108346;
assign addr[61257]= -320065829;
assign addr[61258]= -470399716;
assign addr[61259]= -618347408;
assign addr[61260]= -763158411;
assign addr[61261]= -904098143;
assign addr[61262]= -1040451659;
assign addr[61263]= -1171527280;
assign addr[61264]= -1296660098;
assign addr[61265]= -1415215352;
assign addr[61266]= -1526591649;
assign addr[61267]= -1630224009;
assign addr[61268]= -1725586737;
assign addr[61269]= -1812196087;
assign addr[61270]= -1889612716;
assign addr[61271]= -1957443913;
assign addr[61272]= -2015345591;
assign addr[61273]= -2063024031;
assign addr[61274]= -2100237377;
assign addr[61275]= -2126796855;
assign addr[61276]= -2142567738;
assign addr[61277]= -2147470025;
assign addr[61278]= -2141478848;
assign addr[61279]= -2124624598;
assign addr[61280]= -2096992772;
assign addr[61281]= -2058723538;
assign addr[61282]= -2010011024;
assign addr[61283]= -1951102334;
assign addr[61284]= -1882296293;
assign addr[61285]= -1803941934;
assign addr[61286]= -1716436725;
assign addr[61287]= -1620224553;
assign addr[61288]= -1515793473;
assign addr[61289]= -1403673233;
assign addr[61290]= -1284432584;
assign addr[61291]= -1158676398;
assign addr[61292]= -1027042599;
assign addr[61293]= -890198924;
assign addr[61294]= -748839539;
assign addr[61295]= -603681519;
assign addr[61296]= -455461206;
assign addr[61297]= -304930476;
assign addr[61298]= -152852926;
assign addr[61299]= 0;
assign addr[61300]= 152852926;
assign addr[61301]= 304930476;
assign addr[61302]= 455461206;
assign addr[61303]= 603681519;
assign addr[61304]= 748839539;
assign addr[61305]= 890198924;
assign addr[61306]= 1027042599;
assign addr[61307]= 1158676398;
assign addr[61308]= 1284432584;
assign addr[61309]= 1403673233;
assign addr[61310]= 1515793473;
assign addr[61311]= 1620224553;
assign addr[61312]= 1716436725;
assign addr[61313]= 1803941934;
assign addr[61314]= 1882296293;
assign addr[61315]= 1951102334;
assign addr[61316]= 2010011024;
assign addr[61317]= 2058723538;
assign addr[61318]= 2096992772;
assign addr[61319]= 2124624598;
assign addr[61320]= 2141478848;
assign addr[61321]= 2147470025;
assign addr[61322]= 2142567738;
assign addr[61323]= 2126796855;
assign addr[61324]= 2100237377;
assign addr[61325]= 2063024031;
assign addr[61326]= 2015345591;
assign addr[61327]= 1957443913;
assign addr[61328]= 1889612716;
assign addr[61329]= 1812196087;
assign addr[61330]= 1725586737;
assign addr[61331]= 1630224009;
assign addr[61332]= 1526591649;
assign addr[61333]= 1415215352;
assign addr[61334]= 1296660098;
assign addr[61335]= 1171527280;
assign addr[61336]= 1040451659;
assign addr[61337]= 904098143;
assign addr[61338]= 763158411;
assign addr[61339]= 618347408;
assign addr[61340]= 470399716;
assign addr[61341]= 320065829;
assign addr[61342]= 168108346;
assign addr[61343]= 15298099;
assign addr[61344]= -137589750;
assign addr[61345]= -289779648;
assign addr[61346]= -440499581;
assign addr[61347]= -588984994;
assign addr[61348]= -734482665;
assign addr[61349]= -876254528;
assign addr[61350]= -1013581418;
assign addr[61351]= -1145766716;
assign addr[61352]= -1272139887;
assign addr[61353]= -1392059879;
assign addr[61354]= -1504918373;
assign addr[61355]= -1610142873;
assign addr[61356]= -1707199606;
assign addr[61357]= -1795596234;
assign addr[61358]= -1874884346;
assign addr[61359]= -1944661739;
assign addr[61360]= -2004574453;
assign addr[61361]= -2054318569;
assign addr[61362]= -2093641749;
assign addr[61363]= -2122344521;
assign addr[61364]= -2140281282;
assign addr[61365]= -2147361045;
assign addr[61366]= -2143547897;
assign addr[61367]= -2128861181;
assign addr[61368]= -2103375398;
assign addr[61369]= -2067219829;
assign addr[61370]= -2020577882;
assign addr[61371]= -1963686155;
assign addr[61372]= -1896833245;
assign addr[61373]= -1820358275;
assign addr[61374]= -1734649179;
assign addr[61375]= -1640140734;
assign addr[61376]= -1537312353;
assign addr[61377]= -1426685652;
assign addr[61378]= -1308821808;
assign addr[61379]= -1184318708;
assign addr[61380]= -1053807919;
assign addr[61381]= -917951481;
assign addr[61382]= -777438554;
assign addr[61383]= -632981917;
assign addr[61384]= -485314355;
assign addr[61385]= -335184940;
assign addr[61386]= -183355234;
assign addr[61387]= -30595422;
assign addr[61388]= 122319591;
assign addr[61389]= 274614114;
assign addr[61390]= 425515602;
assign addr[61391]= 574258580;
assign addr[61392]= 720088517;
assign addr[61393]= 862265664;
assign addr[61394]= 1000068799;
assign addr[61395]= 1132798888;
assign addr[61396]= 1259782632;
assign addr[61397]= 1380375881;
assign addr[61398]= 1493966902;
assign addr[61399]= 1599979481;
assign addr[61400]= 1697875851;
assign addr[61401]= 1787159411;
assign addr[61402]= 1867377253;
assign addr[61403]= 1938122457;
assign addr[61404]= 1999036154;
assign addr[61405]= 2049809346;
assign addr[61406]= 2090184478;
assign addr[61407]= 2119956737;
assign addr[61408]= 2138975100;
assign addr[61409]= 2147143090;
assign addr[61410]= 2144419275;
assign addr[61411]= 2130817471;
assign addr[61412]= 2106406677;
assign addr[61413]= 2071310720;
assign addr[61414]= 2025707632;
assign addr[61415]= 1969828744;
assign addr[61416]= 1903957513;
assign addr[61417]= 1828428082;
assign addr[61418]= 1743623590;
assign addr[61419]= 1649974225;
assign addr[61420]= 1547955041;
assign addr[61421]= 1438083551;
assign addr[61422]= 1320917099;
assign addr[61423]= 1197050035;
assign addr[61424]= 1067110699;
assign addr[61425]= 931758235;
assign addr[61426]= 791679244;
assign addr[61427]= 647584304;
assign addr[61428]= 500204365;
assign addr[61429]= 350287041;
assign addr[61430]= 198592817;
assign addr[61431]= 45891193;
assign addr[61432]= -107043224;
assign addr[61433]= -259434643;
assign addr[61434]= -410510029;
assign addr[61435]= -559503022;
assign addr[61436]= -705657826;
assign addr[61437]= -848233042;
assign addr[61438]= -986505429;
assign addr[61439]= -1119773573;
assign addr[61440]= -1247361445;
assign addr[61441]= -1368621831;
assign addr[61442]= -1482939614;
assign addr[61443]= -1589734894;
assign addr[61444]= -1688465931;
assign addr[61445]= -1778631892;
assign addr[61446]= -1859775393;
assign addr[61447]= -1931484818;
assign addr[61448]= -1993396407;
assign addr[61449]= -2045196100;
assign addr[61450]= -2086621133;
assign addr[61451]= -2117461370;
assign addr[61452]= -2137560369;
assign addr[61453]= -2146816171;
assign addr[61454]= -2145181827;
assign addr[61455]= -2132665626;
assign addr[61456]= -2109331059;
assign addr[61457]= -2075296495;
assign addr[61458]= -2030734582;
assign addr[61459]= -1975871368;
assign addr[61460]= -1910985158;
assign addr[61461]= -1836405100;
assign addr[61462]= -1752509516;
assign addr[61463]= -1659723983;
assign addr[61464]= -1558519173;
assign addr[61465]= -1449408469;
assign addr[61466]= -1332945355;
assign addr[61467]= -1209720613;
assign addr[61468]= -1080359326;
assign addr[61469]= -945517704;
assign addr[61470]= -805879757;
assign addr[61471]= -662153826;
assign addr[61472]= -515068990;
assign addr[61473]= -365371365;
assign addr[61474]= -213820322;
assign addr[61475]= -61184634;
assign addr[61476]= 91761426;
assign addr[61477]= 244242007;
assign addr[61478]= 395483624;
assign addr[61479]= 544719071;
assign addr[61480]= 691191324;
assign addr[61481]= 834157373;
assign addr[61482]= 972891995;
assign addr[61483]= 1106691431;
assign addr[61484]= 1234876957;
assign addr[61485]= 1356798326;
assign addr[61486]= 1471837070;
assign addr[61487]= 1579409630;
assign addr[61488]= 1678970324;
assign addr[61489]= 1770014111;
assign addr[61490]= 1852079154;
assign addr[61491]= 1924749160;
assign addr[61492]= 1987655498;
assign addr[61493]= 2040479063;
assign addr[61494]= 2082951896;
assign addr[61495]= 2114858546;
assign addr[61496]= 2136037160;
assign addr[61497]= 2146380306;
assign addr[61498]= 2145835515;
assign addr[61499]= 2134405552;
assign addr[61500]= 2112148396;
assign addr[61501]= 2079176953;
assign addr[61502]= 2035658475;
assign addr[61503]= 1981813720;
assign addr[61504]= 1917915825;
assign addr[61505]= 1844288924;
assign addr[61506]= 1761306505;
assign addr[61507]= 1669389513;
assign addr[61508]= 1569004214;
assign addr[61509]= 1460659832;
assign addr[61510]= 1344905966;
assign addr[61511]= 1222329801;
assign addr[61512]= 1093553126;
assign addr[61513]= 959229189;
assign addr[61514]= 820039373;
assign addr[61515]= 676689746;
assign addr[61516]= 529907477;
assign addr[61517]= 380437148;
assign addr[61518]= 229036977;
assign addr[61519]= 76474970;
assign addr[61520]= -76474970;
assign addr[61521]= -229036977;
assign addr[61522]= -380437148;
assign addr[61523]= -529907477;
assign addr[61524]= -676689746;
assign addr[61525]= -820039373;
assign addr[61526]= -959229189;
assign addr[61527]= -1093553126;
assign addr[61528]= -1222329801;
assign addr[61529]= -1344905966;
assign addr[61530]= -1460659832;
assign addr[61531]= -1569004214;
assign addr[61532]= -1669389513;
assign addr[61533]= -1761306505;
assign addr[61534]= -1844288924;
assign addr[61535]= -1917915825;
assign addr[61536]= -1981813720;
assign addr[61537]= -2035658475;
assign addr[61538]= -2079176953;
assign addr[61539]= -2112148396;
assign addr[61540]= -2134405552;
assign addr[61541]= -2145835515;
assign addr[61542]= -2146380306;
assign addr[61543]= -2136037160;
assign addr[61544]= -2114858546;
assign addr[61545]= -2082951896;
assign addr[61546]= -2040479063;
assign addr[61547]= -1987655498;
assign addr[61548]= -1924749160;
assign addr[61549]= -1852079154;
assign addr[61550]= -1770014111;
assign addr[61551]= -1678970324;
assign addr[61552]= -1579409630;
assign addr[61553]= -1471837070;
assign addr[61554]= -1356798326;
assign addr[61555]= -1234876957;
assign addr[61556]= -1106691431;
assign addr[61557]= -972891995;
assign addr[61558]= -834157373;
assign addr[61559]= -691191324;
assign addr[61560]= -544719071;
assign addr[61561]= -395483624;
assign addr[61562]= -244242007;
assign addr[61563]= -91761426;
assign addr[61564]= 61184634;
assign addr[61565]= 213820322;
assign addr[61566]= 365371365;
assign addr[61567]= 515068990;
assign addr[61568]= 662153826;
assign addr[61569]= 805879757;
assign addr[61570]= 945517704;
assign addr[61571]= 1080359326;
assign addr[61572]= 1209720613;
assign addr[61573]= 1332945355;
assign addr[61574]= 1449408469;
assign addr[61575]= 1558519173;
assign addr[61576]= 1659723983;
assign addr[61577]= 1752509516;
assign addr[61578]= 1836405100;
assign addr[61579]= 1910985158;
assign addr[61580]= 1975871368;
assign addr[61581]= 2030734582;
assign addr[61582]= 2075296495;
assign addr[61583]= 2109331059;
assign addr[61584]= 2132665626;
assign addr[61585]= 2145181827;
assign addr[61586]= 2146816171;
assign addr[61587]= 2137560369;
assign addr[61588]= 2117461370;
assign addr[61589]= 2086621133;
assign addr[61590]= 2045196100;
assign addr[61591]= 1993396407;
assign addr[61592]= 1931484818;
assign addr[61593]= 1859775393;
assign addr[61594]= 1778631892;
assign addr[61595]= 1688465931;
assign addr[61596]= 1589734894;
assign addr[61597]= 1482939614;
assign addr[61598]= 1368621831;
assign addr[61599]= 1247361445;
assign addr[61600]= 1119773573;
assign addr[61601]= 986505429;
assign addr[61602]= 848233042;
assign addr[61603]= 705657826;
assign addr[61604]= 559503022;
assign addr[61605]= 410510029;
assign addr[61606]= 259434643;
assign addr[61607]= 107043224;
assign addr[61608]= -45891193;
assign addr[61609]= -198592817;
assign addr[61610]= -350287041;
assign addr[61611]= -500204365;
assign addr[61612]= -647584304;
assign addr[61613]= -791679244;
assign addr[61614]= -931758235;
assign addr[61615]= -1067110699;
assign addr[61616]= -1197050035;
assign addr[61617]= -1320917099;
assign addr[61618]= -1438083551;
assign addr[61619]= -1547955041;
assign addr[61620]= -1649974225;
assign addr[61621]= -1743623590;
assign addr[61622]= -1828428082;
assign addr[61623]= -1903957513;
assign addr[61624]= -1969828744;
assign addr[61625]= -2025707632;
assign addr[61626]= -2071310720;
assign addr[61627]= -2106406677;
assign addr[61628]= -2130817471;
assign addr[61629]= -2144419275;
assign addr[61630]= -2147143090;
assign addr[61631]= -2138975100;
assign addr[61632]= -2119956737;
assign addr[61633]= -2090184478;
assign addr[61634]= -2049809346;
assign addr[61635]= -1999036154;
assign addr[61636]= -1938122457;
assign addr[61637]= -1867377253;
assign addr[61638]= -1787159411;
assign addr[61639]= -1697875851;
assign addr[61640]= -1599979481;
assign addr[61641]= -1493966902;
assign addr[61642]= -1380375881;
assign addr[61643]= -1259782632;
assign addr[61644]= -1132798888;
assign addr[61645]= -1000068799;
assign addr[61646]= -862265664;
assign addr[61647]= -720088517;
assign addr[61648]= -574258580;
assign addr[61649]= -425515602;
assign addr[61650]= -274614114;
assign addr[61651]= -122319591;
assign addr[61652]= 30595422;
assign addr[61653]= 183355234;
assign addr[61654]= 335184940;
assign addr[61655]= 485314355;
assign addr[61656]= 632981917;
assign addr[61657]= 777438554;
assign addr[61658]= 917951481;
assign addr[61659]= 1053807919;
assign addr[61660]= 1184318708;
assign addr[61661]= 1308821808;
assign addr[61662]= 1426685652;
assign addr[61663]= 1537312353;
assign addr[61664]= 1640140734;
assign addr[61665]= 1734649179;
assign addr[61666]= 1820358275;
assign addr[61667]= 1896833245;
assign addr[61668]= 1963686155;
assign addr[61669]= 2020577882;
assign addr[61670]= 2067219829;
assign addr[61671]= 2103375398;
assign addr[61672]= 2128861181;
assign addr[61673]= 2143547897;
assign addr[61674]= 2147361045;
assign addr[61675]= 2140281282;
assign addr[61676]= 2122344521;
assign addr[61677]= 2093641749;
assign addr[61678]= 2054318569;
assign addr[61679]= 2004574453;
assign addr[61680]= 1944661739;
assign addr[61681]= 1874884346;
assign addr[61682]= 1795596234;
assign addr[61683]= 1707199606;
assign addr[61684]= 1610142873;
assign addr[61685]= 1504918373;
assign addr[61686]= 1392059879;
assign addr[61687]= 1272139887;
assign addr[61688]= 1145766716;
assign addr[61689]= 1013581418;
assign addr[61690]= 876254528;
assign addr[61691]= 734482665;
assign addr[61692]= 588984994;
assign addr[61693]= 440499581;
assign addr[61694]= 289779648;
assign addr[61695]= 137589750;
assign addr[61696]= -15298099;
assign addr[61697]= -168108346;
assign addr[61698]= -320065829;
assign addr[61699]= -470399716;
assign addr[61700]= -618347408;
assign addr[61701]= -763158411;
assign addr[61702]= -904098143;
assign addr[61703]= -1040451659;
assign addr[61704]= -1171527280;
assign addr[61705]= -1296660098;
assign addr[61706]= -1415215352;
assign addr[61707]= -1526591649;
assign addr[61708]= -1630224009;
assign addr[61709]= -1725586737;
assign addr[61710]= -1812196087;
assign addr[61711]= -1889612716;
assign addr[61712]= -1957443913;
assign addr[61713]= -2015345591;
assign addr[61714]= -2063024031;
assign addr[61715]= -2100237377;
assign addr[61716]= -2126796855;
assign addr[61717]= -2142567738;
assign addr[61718]= -2147470025;
assign addr[61719]= -2141478848;
assign addr[61720]= -2124624598;
assign addr[61721]= -2096992772;
assign addr[61722]= -2058723538;
assign addr[61723]= -2010011024;
assign addr[61724]= -1951102334;
assign addr[61725]= -1882296293;
assign addr[61726]= -1803941934;
assign addr[61727]= -1716436725;
assign addr[61728]= -1620224553;
assign addr[61729]= -1515793473;
assign addr[61730]= -1403673233;
assign addr[61731]= -1284432584;
assign addr[61732]= -1158676398;
assign addr[61733]= -1027042599;
assign addr[61734]= -890198924;
assign addr[61735]= -748839539;
assign addr[61736]= -603681519;
assign addr[61737]= -455461206;
assign addr[61738]= -304930476;
assign addr[61739]= -152852926;
assign addr[61740]= 0;
assign addr[61741]= 152852926;
assign addr[61742]= 304930476;
assign addr[61743]= 455461206;
assign addr[61744]= 603681519;
assign addr[61745]= 748839539;
assign addr[61746]= 890198924;
assign addr[61747]= 1027042599;
assign addr[61748]= 1158676398;
assign addr[61749]= 1284432584;
assign addr[61750]= 1403673233;
assign addr[61751]= 1515793473;
assign addr[61752]= 1620224553;
assign addr[61753]= 1716436725;
assign addr[61754]= 1803941934;
assign addr[61755]= 1882296293;
assign addr[61756]= 1951102334;
assign addr[61757]= 2010011024;
assign addr[61758]= 2058723538;
assign addr[61759]= 2096992772;
assign addr[61760]= 2124624598;
assign addr[61761]= 2141478848;
assign addr[61762]= 2147470025;
assign addr[61763]= 2142567738;
assign addr[61764]= 2126796855;
assign addr[61765]= 2100237377;
assign addr[61766]= 2063024031;
assign addr[61767]= 2015345591;
assign addr[61768]= 1957443913;
assign addr[61769]= 1889612716;
assign addr[61770]= 1812196087;
assign addr[61771]= 1725586737;
assign addr[61772]= 1630224009;
assign addr[61773]= 1526591649;
assign addr[61774]= 1415215352;
assign addr[61775]= 1296660098;
assign addr[61776]= 1171527280;
assign addr[61777]= 1040451659;
assign addr[61778]= 904098143;
assign addr[61779]= 763158411;
assign addr[61780]= 618347408;
assign addr[61781]= 470399716;
assign addr[61782]= 320065829;
assign addr[61783]= 168108346;
assign addr[61784]= 15298099;
assign addr[61785]= -137589750;
assign addr[61786]= -289779648;
assign addr[61787]= -440499581;
assign addr[61788]= -588984994;
assign addr[61789]= -734482665;
assign addr[61790]= -876254528;
assign addr[61791]= -1013581418;
assign addr[61792]= -1145766716;
assign addr[61793]= -1272139887;
assign addr[61794]= -1392059879;
assign addr[61795]= -1504918373;
assign addr[61796]= -1610142873;
assign addr[61797]= -1707199606;
assign addr[61798]= -1795596234;
assign addr[61799]= -1874884346;
assign addr[61800]= -1944661739;
assign addr[61801]= -2004574453;
assign addr[61802]= -2054318569;
assign addr[61803]= -2093641749;
assign addr[61804]= -2122344521;
assign addr[61805]= -2140281282;
assign addr[61806]= -2147361045;
assign addr[61807]= -2143547897;
assign addr[61808]= -2128861181;
assign addr[61809]= -2103375398;
assign addr[61810]= -2067219829;
assign addr[61811]= -2020577882;
assign addr[61812]= -1963686155;
assign addr[61813]= -1896833245;
assign addr[61814]= -1820358275;
assign addr[61815]= -1734649179;
assign addr[61816]= -1640140734;
assign addr[61817]= -1537312353;
assign addr[61818]= -1426685652;
assign addr[61819]= -1308821808;
assign addr[61820]= -1184318708;
assign addr[61821]= -1053807919;
assign addr[61822]= -917951481;
assign addr[61823]= -777438554;
assign addr[61824]= -632981917;
assign addr[61825]= -485314355;
assign addr[61826]= -335184940;
assign addr[61827]= -183355234;
assign addr[61828]= -30595422;
assign addr[61829]= 122319591;
assign addr[61830]= 274614114;
assign addr[61831]= 425515602;
assign addr[61832]= 574258580;
assign addr[61833]= 720088517;
assign addr[61834]= 862265664;
assign addr[61835]= 1000068799;
assign addr[61836]= 1132798888;
assign addr[61837]= 1259782632;
assign addr[61838]= 1380375881;
assign addr[61839]= 1493966902;
assign addr[61840]= 1599979481;
assign addr[61841]= 1697875851;
assign addr[61842]= 1787159411;
assign addr[61843]= 1867377253;
assign addr[61844]= 1938122457;
assign addr[61845]= 1999036154;
assign addr[61846]= 2049809346;
assign addr[61847]= 2090184478;
assign addr[61848]= 2119956737;
assign addr[61849]= 2138975100;
assign addr[61850]= 2147143090;
assign addr[61851]= 2144419275;
assign addr[61852]= 2130817471;
assign addr[61853]= 2106406677;
assign addr[61854]= 2071310720;
assign addr[61855]= 2025707632;
assign addr[61856]= 1969828744;
assign addr[61857]= 1903957513;
assign addr[61858]= 1828428082;
assign addr[61859]= 1743623590;
assign addr[61860]= 1649974225;
assign addr[61861]= 1547955041;
assign addr[61862]= 1438083551;
assign addr[61863]= 1320917099;
assign addr[61864]= 1197050035;
assign addr[61865]= 1067110699;
assign addr[61866]= 931758235;
assign addr[61867]= 791679244;
assign addr[61868]= 647584304;
assign addr[61869]= 500204365;
assign addr[61870]= 350287041;
assign addr[61871]= 198592817;
assign addr[61872]= 45891193;
assign addr[61873]= -107043224;
assign addr[61874]= -259434643;
assign addr[61875]= -410510029;
assign addr[61876]= -559503022;
assign addr[61877]= -705657826;
assign addr[61878]= -848233042;
assign addr[61879]= -986505429;
assign addr[61880]= -1119773573;
assign addr[61881]= -1247361445;
assign addr[61882]= -1368621831;
assign addr[61883]= -1482939614;
assign addr[61884]= -1589734894;
assign addr[61885]= -1688465931;
assign addr[61886]= -1778631892;
assign addr[61887]= -1859775393;
assign addr[61888]= -1931484818;
assign addr[61889]= -1993396407;
assign addr[61890]= -2045196100;
assign addr[61891]= -2086621133;
assign addr[61892]= -2117461370;
assign addr[61893]= -2137560369;
assign addr[61894]= -2146816171;
assign addr[61895]= -2145181827;
assign addr[61896]= -2132665626;
assign addr[61897]= -2109331059;
assign addr[61898]= -2075296495;
assign addr[61899]= -2030734582;
assign addr[61900]= -1975871368;
assign addr[61901]= -1910985158;
assign addr[61902]= -1836405100;
assign addr[61903]= -1752509516;
assign addr[61904]= -1659723983;
assign addr[61905]= -1558519173;
assign addr[61906]= -1449408469;
assign addr[61907]= -1332945355;
assign addr[61908]= -1209720613;
assign addr[61909]= -1080359326;
assign addr[61910]= -945517704;
assign addr[61911]= -805879757;
assign addr[61912]= -662153826;
assign addr[61913]= -515068990;
assign addr[61914]= -365371365;
assign addr[61915]= -213820322;
assign addr[61916]= -61184634;
assign addr[61917]= 91761426;
assign addr[61918]= 244242007;
assign addr[61919]= 395483624;
assign addr[61920]= 544719071;
assign addr[61921]= 691191324;
assign addr[61922]= 834157373;
assign addr[61923]= 972891995;
assign addr[61924]= 1106691431;
assign addr[61925]= 1234876957;
assign addr[61926]= 1356798326;
assign addr[61927]= 1471837070;
assign addr[61928]= 1579409630;
assign addr[61929]= 1678970324;
assign addr[61930]= 1770014111;
assign addr[61931]= 1852079154;
assign addr[61932]= 1924749160;
assign addr[61933]= 1987655498;
assign addr[61934]= 2040479063;
assign addr[61935]= 2082951896;
assign addr[61936]= 2114858546;
assign addr[61937]= 2136037160;
assign addr[61938]= 2146380306;
assign addr[61939]= 2145835515;
assign addr[61940]= 2134405552;
assign addr[61941]= 2112148396;
assign addr[61942]= 2079176953;
assign addr[61943]= 2035658475;
assign addr[61944]= 1981813720;
assign addr[61945]= 1917915825;
assign addr[61946]= 1844288924;
assign addr[61947]= 1761306505;
assign addr[61948]= 1669389513;
assign addr[61949]= 1569004214;
assign addr[61950]= 1460659832;
assign addr[61951]= 1344905966;
assign addr[61952]= 1222329801;
assign addr[61953]= 1093553126;
assign addr[61954]= 959229189;
assign addr[61955]= 820039373;
assign addr[61956]= 676689746;
assign addr[61957]= 529907477;
assign addr[61958]= 380437148;
assign addr[61959]= 229036977;
assign addr[61960]= 76474970;
assign addr[61961]= -76474970;
assign addr[61962]= -229036977;
assign addr[61963]= -380437148;
assign addr[61964]= -529907477;
assign addr[61965]= -676689746;
assign addr[61966]= -820039373;
assign addr[61967]= -959229189;
assign addr[61968]= -1093553126;
assign addr[61969]= -1222329801;
assign addr[61970]= -1344905966;
assign addr[61971]= -1460659832;
assign addr[61972]= -1569004214;
assign addr[61973]= -1669389513;
assign addr[61974]= -1761306505;
assign addr[61975]= -1844288924;
assign addr[61976]= -1917915825;
assign addr[61977]= -1981813720;
assign addr[61978]= -2035658475;
assign addr[61979]= -2079176953;
assign addr[61980]= -2112148396;
assign addr[61981]= -2134405552;
assign addr[61982]= -2145835515;
assign addr[61983]= -2146380306;
assign addr[61984]= -2136037160;
assign addr[61985]= -2114858546;
assign addr[61986]= -2082951896;
assign addr[61987]= -2040479063;
assign addr[61988]= -1987655498;
assign addr[61989]= -1924749160;
assign addr[61990]= -1852079154;
assign addr[61991]= -1770014111;
assign addr[61992]= -1678970324;
assign addr[61993]= -1579409630;
assign addr[61994]= -1471837070;
assign addr[61995]= -1356798326;
assign addr[61996]= -1234876957;
assign addr[61997]= -1106691431;
assign addr[61998]= -972891995;
assign addr[61999]= -834157373;
assign addr[62000]= -691191324;
assign addr[62001]= -544719071;
assign addr[62002]= -395483624;
assign addr[62003]= -244242007;
assign addr[62004]= -91761426;
assign addr[62005]= 61184634;
assign addr[62006]= 213820322;
assign addr[62007]= 365371365;
assign addr[62008]= 515068990;
assign addr[62009]= 662153826;
assign addr[62010]= 805879757;
assign addr[62011]= 945517704;
assign addr[62012]= 1080359326;
assign addr[62013]= 1209720613;
assign addr[62014]= 1332945355;
assign addr[62015]= 1449408469;
assign addr[62016]= 1558519173;
assign addr[62017]= 1659723983;
assign addr[62018]= 1752509516;
assign addr[62019]= 1836405100;
assign addr[62020]= 1910985158;
assign addr[62021]= 1975871368;
assign addr[62022]= 2030734582;
assign addr[62023]= 2075296495;
assign addr[62024]= 2109331059;
assign addr[62025]= 2132665626;
assign addr[62026]= 2145181827;
assign addr[62027]= 2146816171;
assign addr[62028]= 2137560369;
assign addr[62029]= 2117461370;
assign addr[62030]= 2086621133;
assign addr[62031]= 2045196100;
assign addr[62032]= 1993396407;
assign addr[62033]= 1931484818;
assign addr[62034]= 1859775393;
assign addr[62035]= 1778631892;
assign addr[62036]= 1688465931;
assign addr[62037]= 1589734894;
assign addr[62038]= 1482939614;
assign addr[62039]= 1368621831;
assign addr[62040]= 1247361445;
assign addr[62041]= 1119773573;
assign addr[62042]= 986505429;
assign addr[62043]= 848233042;
assign addr[62044]= 705657826;
assign addr[62045]= 559503022;
assign addr[62046]= 410510029;
assign addr[62047]= 259434643;
assign addr[62048]= 107043224;
assign addr[62049]= -45891193;
assign addr[62050]= -198592817;
assign addr[62051]= -350287041;
assign addr[62052]= -500204365;
assign addr[62053]= -647584304;
assign addr[62054]= -791679244;
assign addr[62055]= -931758235;
assign addr[62056]= -1067110699;
assign addr[62057]= -1197050035;
assign addr[62058]= -1320917099;
assign addr[62059]= -1438083551;
assign addr[62060]= -1547955041;
assign addr[62061]= -1649974225;
assign addr[62062]= -1743623590;
assign addr[62063]= -1828428082;
assign addr[62064]= -1903957513;
assign addr[62065]= -1969828744;
assign addr[62066]= -2025707632;
assign addr[62067]= -2071310720;
assign addr[62068]= -2106406677;
assign addr[62069]= -2130817471;
assign addr[62070]= -2144419275;
assign addr[62071]= -2147143090;
assign addr[62072]= -2138975100;
assign addr[62073]= -2119956737;
assign addr[62074]= -2090184478;
assign addr[62075]= -2049809346;
assign addr[62076]= -1999036154;
assign addr[62077]= -1938122457;
assign addr[62078]= -1867377253;
assign addr[62079]= -1787159411;
assign addr[62080]= -1697875851;
assign addr[62081]= -1599979481;
assign addr[62082]= -1493966902;
assign addr[62083]= -1380375881;
assign addr[62084]= -1259782632;
assign addr[62085]= -1132798888;
assign addr[62086]= -1000068799;
assign addr[62087]= -862265664;
assign addr[62088]= -720088517;
assign addr[62089]= -574258580;
assign addr[62090]= -425515602;
assign addr[62091]= -274614114;
assign addr[62092]= -122319591;
assign addr[62093]= 30595422;
assign addr[62094]= 183355234;
assign addr[62095]= 335184940;
assign addr[62096]= 485314355;
assign addr[62097]= 632981917;
assign addr[62098]= 777438554;
assign addr[62099]= 917951481;
assign addr[62100]= 1053807919;
assign addr[62101]= 1184318708;
assign addr[62102]= 1308821808;
assign addr[62103]= 1426685652;
assign addr[62104]= 1537312353;
assign addr[62105]= 1640140734;
assign addr[62106]= 1734649179;
assign addr[62107]= 1820358275;
assign addr[62108]= 1896833245;
assign addr[62109]= 1963686155;
assign addr[62110]= 2020577882;
assign addr[62111]= 2067219829;
assign addr[62112]= 2103375398;
assign addr[62113]= 2128861181;
assign addr[62114]= 2143547897;
assign addr[62115]= 2147361045;
assign addr[62116]= 2140281282;
assign addr[62117]= 2122344521;
assign addr[62118]= 2093641749;
assign addr[62119]= 2054318569;
assign addr[62120]= 2004574453;
assign addr[62121]= 1944661739;
assign addr[62122]= 1874884346;
assign addr[62123]= 1795596234;
assign addr[62124]= 1707199606;
assign addr[62125]= 1610142873;
assign addr[62126]= 1504918373;
assign addr[62127]= 1392059879;
assign addr[62128]= 1272139887;
assign addr[62129]= 1145766716;
assign addr[62130]= 1013581418;
assign addr[62131]= 876254528;
assign addr[62132]= 734482665;
assign addr[62133]= 588984994;
assign addr[62134]= 440499581;
assign addr[62135]= 289779648;
assign addr[62136]= 137589750;
assign addr[62137]= -15298099;
assign addr[62138]= -168108346;
assign addr[62139]= -320065829;
assign addr[62140]= -470399716;
assign addr[62141]= -618347408;
assign addr[62142]= -763158411;
assign addr[62143]= -904098143;
assign addr[62144]= -1040451659;
assign addr[62145]= -1171527280;
assign addr[62146]= -1296660098;
assign addr[62147]= -1415215352;
assign addr[62148]= -1526591649;
assign addr[62149]= -1630224009;
assign addr[62150]= -1725586737;
assign addr[62151]= -1812196087;
assign addr[62152]= -1889612716;
assign addr[62153]= -1957443913;
assign addr[62154]= -2015345591;
assign addr[62155]= -2063024031;
assign addr[62156]= -2100237377;
assign addr[62157]= -2126796855;
assign addr[62158]= -2142567738;
assign addr[62159]= -2147470025;
assign addr[62160]= -2141478848;
assign addr[62161]= -2124624598;
assign addr[62162]= -2096992772;
assign addr[62163]= -2058723538;
assign addr[62164]= -2010011024;
assign addr[62165]= -1951102334;
assign addr[62166]= -1882296293;
assign addr[62167]= -1803941934;
assign addr[62168]= -1716436725;
assign addr[62169]= -1620224553;
assign addr[62170]= -1515793473;
assign addr[62171]= -1403673233;
assign addr[62172]= -1284432584;
assign addr[62173]= -1158676398;
assign addr[62174]= -1027042599;
assign addr[62175]= -890198924;
assign addr[62176]= -748839539;
assign addr[62177]= -603681519;
assign addr[62178]= -455461206;
assign addr[62179]= -304930476;
assign addr[62180]= -152852926;
assign addr[62181]= 0;
assign addr[62182]= 152852926;
assign addr[62183]= 304930476;
assign addr[62184]= 455461206;
assign addr[62185]= 603681519;
assign addr[62186]= 748839539;
assign addr[62187]= 890198924;
assign addr[62188]= 1027042599;
assign addr[62189]= 1158676398;
assign addr[62190]= 1284432584;
assign addr[62191]= 1403673233;
assign addr[62192]= 1515793473;
assign addr[62193]= 1620224553;
assign addr[62194]= 1716436725;
assign addr[62195]= 1803941934;
assign addr[62196]= 1882296293;
assign addr[62197]= 1951102334;
assign addr[62198]= 2010011024;
assign addr[62199]= 2058723538;
assign addr[62200]= 2096992772;
assign addr[62201]= 2124624598;
assign addr[62202]= 2141478848;
assign addr[62203]= 2147470025;
assign addr[62204]= 2142567738;
assign addr[62205]= 2126796855;
assign addr[62206]= 2100237377;
assign addr[62207]= 2063024031;
assign addr[62208]= 2015345591;
assign addr[62209]= 1957443913;
assign addr[62210]= 1889612716;
assign addr[62211]= 1812196087;
assign addr[62212]= 1725586737;
assign addr[62213]= 1630224009;
assign addr[62214]= 1526591649;
assign addr[62215]= 1415215352;
assign addr[62216]= 1296660098;
assign addr[62217]= 1171527280;
assign addr[62218]= 1040451659;
assign addr[62219]= 904098143;
assign addr[62220]= 763158411;
assign addr[62221]= 618347408;
assign addr[62222]= 470399716;
assign addr[62223]= 320065829;
assign addr[62224]= 168108346;
assign addr[62225]= 15298099;
assign addr[62226]= -137589750;
assign addr[62227]= -289779648;
assign addr[62228]= -440499581;
assign addr[62229]= -588984994;
assign addr[62230]= -734482665;
assign addr[62231]= -876254528;
assign addr[62232]= -1013581418;
assign addr[62233]= -1145766716;
assign addr[62234]= -1272139887;
assign addr[62235]= -1392059879;
assign addr[62236]= -1504918373;
assign addr[62237]= -1610142873;
assign addr[62238]= -1707199606;
assign addr[62239]= -1795596234;
assign addr[62240]= -1874884346;
assign addr[62241]= -1944661739;
assign addr[62242]= -2004574453;
assign addr[62243]= -2054318569;
assign addr[62244]= -2093641749;
assign addr[62245]= -2122344521;
assign addr[62246]= -2140281282;
assign addr[62247]= -2147361045;
assign addr[62248]= -2143547897;
assign addr[62249]= -2128861181;
assign addr[62250]= -2103375398;
assign addr[62251]= -2067219829;
assign addr[62252]= -2020577882;
assign addr[62253]= -1963686155;
assign addr[62254]= -1896833245;
assign addr[62255]= -1820358275;
assign addr[62256]= -1734649179;
assign addr[62257]= -1640140734;
assign addr[62258]= -1537312353;
assign addr[62259]= -1426685652;
assign addr[62260]= -1308821808;
assign addr[62261]= -1184318708;
assign addr[62262]= -1053807919;
assign addr[62263]= -917951481;
assign addr[62264]= -777438554;
assign addr[62265]= -632981917;
assign addr[62266]= -485314355;
assign addr[62267]= -335184940;
assign addr[62268]= -183355234;
assign addr[62269]= -30595422;
assign addr[62270]= 122319591;
assign addr[62271]= 274614114;
assign addr[62272]= 425515602;
assign addr[62273]= 574258580;
assign addr[62274]= 720088517;
assign addr[62275]= 862265664;
assign addr[62276]= 1000068799;
assign addr[62277]= 1132798888;
assign addr[62278]= 1259782632;
assign addr[62279]= 1380375881;
assign addr[62280]= 1493966902;
assign addr[62281]= 1599979481;
assign addr[62282]= 1697875851;
assign addr[62283]= 1787159411;
assign addr[62284]= 1867377253;
assign addr[62285]= 1938122457;
assign addr[62286]= 1999036154;
assign addr[62287]= 2049809346;
assign addr[62288]= 2090184478;
assign addr[62289]= 2119956737;
assign addr[62290]= 2138975100;
assign addr[62291]= 2147143090;
assign addr[62292]= 2144419275;
assign addr[62293]= 2130817471;
assign addr[62294]= 2106406677;
assign addr[62295]= 2071310720;
assign addr[62296]= 2025707632;
assign addr[62297]= 1969828744;
assign addr[62298]= 1903957513;
assign addr[62299]= 1828428082;
assign addr[62300]= 1743623590;
assign addr[62301]= 1649974225;
assign addr[62302]= 1547955041;
assign addr[62303]= 1438083551;
assign addr[62304]= 1320917099;
assign addr[62305]= 1197050035;
assign addr[62306]= 1067110699;
assign addr[62307]= 931758235;
assign addr[62308]= 791679244;
assign addr[62309]= 647584304;
assign addr[62310]= 500204365;
assign addr[62311]= 350287041;
assign addr[62312]= 198592817;
assign addr[62313]= 45891193;
assign addr[62314]= -107043224;
assign addr[62315]= -259434643;
assign addr[62316]= -410510029;
assign addr[62317]= -559503022;
assign addr[62318]= -705657826;
assign addr[62319]= -848233042;
assign addr[62320]= -986505429;
assign addr[62321]= -1119773573;
assign addr[62322]= -1247361445;
assign addr[62323]= -1368621831;
assign addr[62324]= -1482939614;
assign addr[62325]= -1589734894;
assign addr[62326]= -1688465931;
assign addr[62327]= -1778631892;
assign addr[62328]= -1859775393;
assign addr[62329]= -1931484818;
assign addr[62330]= -1993396407;
assign addr[62331]= -2045196100;
assign addr[62332]= -2086621133;
assign addr[62333]= -2117461370;
assign addr[62334]= -2137560369;
assign addr[62335]= -2146816171;
assign addr[62336]= -2145181827;
assign addr[62337]= -2132665626;
assign addr[62338]= -2109331059;
assign addr[62339]= -2075296495;
assign addr[62340]= -2030734582;
assign addr[62341]= -1975871368;
assign addr[62342]= -1910985158;
assign addr[62343]= -1836405100;
assign addr[62344]= -1752509516;
assign addr[62345]= -1659723983;
assign addr[62346]= -1558519173;
assign addr[62347]= -1449408469;
assign addr[62348]= -1332945355;
assign addr[62349]= -1209720613;
assign addr[62350]= -1080359326;
assign addr[62351]= -945517704;
assign addr[62352]= -805879757;
assign addr[62353]= -662153826;
assign addr[62354]= -515068990;
assign addr[62355]= -365371365;
assign addr[62356]= -213820322;
assign addr[62357]= -61184634;
assign addr[62358]= 91761426;
assign addr[62359]= 244242007;
assign addr[62360]= 395483624;
assign addr[62361]= 544719071;
assign addr[62362]= 691191324;
assign addr[62363]= 834157373;
assign addr[62364]= 972891995;
assign addr[62365]= 1106691431;
assign addr[62366]= 1234876957;
assign addr[62367]= 1356798326;
assign addr[62368]= 1471837070;
assign addr[62369]= 1579409630;
assign addr[62370]= 1678970324;
assign addr[62371]= 1770014111;
assign addr[62372]= 1852079154;
assign addr[62373]= 1924749160;
assign addr[62374]= 1987655498;
assign addr[62375]= 2040479063;
assign addr[62376]= 2082951896;
assign addr[62377]= 2114858546;
assign addr[62378]= 2136037160;
assign addr[62379]= 2146380306;
assign addr[62380]= 2145835515;
assign addr[62381]= 2134405552;
assign addr[62382]= 2112148396;
assign addr[62383]= 2079176953;
assign addr[62384]= 2035658475;
assign addr[62385]= 1981813720;
assign addr[62386]= 1917915825;
assign addr[62387]= 1844288924;
assign addr[62388]= 1761306505;
assign addr[62389]= 1669389513;
assign addr[62390]= 1569004214;
assign addr[62391]= 1460659832;
assign addr[62392]= 1344905966;
assign addr[62393]= 1222329801;
assign addr[62394]= 1093553126;
assign addr[62395]= 959229189;
assign addr[62396]= 820039373;
assign addr[62397]= 676689746;
assign addr[62398]= 529907477;
assign addr[62399]= 380437148;
assign addr[62400]= 229036977;
assign addr[62401]= 76474970;
assign addr[62402]= -76474970;
assign addr[62403]= -229036977;
assign addr[62404]= -380437148;
assign addr[62405]= -529907477;
assign addr[62406]= -676689746;
assign addr[62407]= -820039373;
assign addr[62408]= -959229189;
assign addr[62409]= -1093553126;
assign addr[62410]= -1222329801;
assign addr[62411]= -1344905966;
assign addr[62412]= -1460659832;
assign addr[62413]= -1569004214;
assign addr[62414]= -1669389513;
assign addr[62415]= -1761306505;
assign addr[62416]= -1844288924;
assign addr[62417]= -1917915825;
assign addr[62418]= -1981813720;
assign addr[62419]= -2035658475;
assign addr[62420]= -2079176953;
assign addr[62421]= -2112148396;
assign addr[62422]= -2134405552;
assign addr[62423]= -2145835515;
assign addr[62424]= -2146380306;
assign addr[62425]= -2136037160;
assign addr[62426]= -2114858546;
assign addr[62427]= -2082951896;
assign addr[62428]= -2040479063;
assign addr[62429]= -1987655498;
assign addr[62430]= -1924749160;
assign addr[62431]= -1852079154;
assign addr[62432]= -1770014111;
assign addr[62433]= -1678970324;
assign addr[62434]= -1579409630;
assign addr[62435]= -1471837070;
assign addr[62436]= -1356798326;
assign addr[62437]= -1234876957;
assign addr[62438]= -1106691431;
assign addr[62439]= -972891995;
assign addr[62440]= -834157373;
assign addr[62441]= -691191324;
assign addr[62442]= -544719071;
assign addr[62443]= -395483624;
assign addr[62444]= -244242007;
assign addr[62445]= -91761426;
assign addr[62446]= 61184634;
assign addr[62447]= 213820322;
assign addr[62448]= 365371365;
assign addr[62449]= 515068990;
assign addr[62450]= 662153826;
assign addr[62451]= 805879757;
assign addr[62452]= 945517704;
assign addr[62453]= 1080359326;
assign addr[62454]= 1209720613;
assign addr[62455]= 1332945355;
assign addr[62456]= 1449408469;
assign addr[62457]= 1558519173;
assign addr[62458]= 1659723983;
assign addr[62459]= 1752509516;
assign addr[62460]= 1836405100;
assign addr[62461]= 1910985158;
assign addr[62462]= 1975871368;
assign addr[62463]= 2030734582;
assign addr[62464]= 2075296495;
assign addr[62465]= 2109331059;
assign addr[62466]= 2132665626;
assign addr[62467]= 2145181827;
assign addr[62468]= 2146816171;
assign addr[62469]= 2137560369;
assign addr[62470]= 2117461370;
assign addr[62471]= 2086621133;
assign addr[62472]= 2045196100;
assign addr[62473]= 1993396407;
assign addr[62474]= 1931484818;
assign addr[62475]= 1859775393;
assign addr[62476]= 1778631892;
assign addr[62477]= 1688465931;
assign addr[62478]= 1589734894;
assign addr[62479]= 1482939614;
assign addr[62480]= 1368621831;
assign addr[62481]= 1247361445;
assign addr[62482]= 1119773573;
assign addr[62483]= 986505429;
assign addr[62484]= 848233042;
assign addr[62485]= 705657826;
assign addr[62486]= 559503022;
assign addr[62487]= 410510029;
assign addr[62488]= 259434643;
assign addr[62489]= 107043224;
assign addr[62490]= -45891193;
assign addr[62491]= -198592817;
assign addr[62492]= -350287041;
assign addr[62493]= -500204365;
assign addr[62494]= -647584304;
assign addr[62495]= -791679244;
assign addr[62496]= -931758235;
assign addr[62497]= -1067110699;
assign addr[62498]= -1197050035;
assign addr[62499]= -1320917099;
assign addr[62500]= -1438083551;
assign addr[62501]= -1547955041;
assign addr[62502]= -1649974225;
assign addr[62503]= -1743623590;
assign addr[62504]= -1828428082;
assign addr[62505]= -1903957513;
assign addr[62506]= -1969828744;
assign addr[62507]= -2025707632;
assign addr[62508]= -2071310720;
assign addr[62509]= -2106406677;
assign addr[62510]= -2130817471;
assign addr[62511]= -2144419275;
assign addr[62512]= -2147143090;
assign addr[62513]= -2138975100;
assign addr[62514]= -2119956737;
assign addr[62515]= -2090184478;
assign addr[62516]= -2049809346;
assign addr[62517]= -1999036154;
assign addr[62518]= -1938122457;
assign addr[62519]= -1867377253;
assign addr[62520]= -1787159411;
assign addr[62521]= -1697875851;
assign addr[62522]= -1599979481;
assign addr[62523]= -1493966902;
assign addr[62524]= -1380375881;
assign addr[62525]= -1259782632;
assign addr[62526]= -1132798888;
assign addr[62527]= -1000068799;
assign addr[62528]= -862265664;
assign addr[62529]= -720088517;
assign addr[62530]= -574258580;
assign addr[62531]= -425515602;
assign addr[62532]= -274614114;
assign addr[62533]= -122319591;
assign addr[62534]= 30595422;
assign addr[62535]= 183355234;
assign addr[62536]= 335184940;
assign addr[62537]= 485314355;
assign addr[62538]= 632981917;
assign addr[62539]= 777438554;
assign addr[62540]= 917951481;
assign addr[62541]= 1053807919;
assign addr[62542]= 1184318708;
assign addr[62543]= 1308821808;
assign addr[62544]= 1426685652;
assign addr[62545]= 1537312353;
assign addr[62546]= 1640140734;
assign addr[62547]= 1734649179;
assign addr[62548]= 1820358275;
assign addr[62549]= 1896833245;
assign addr[62550]= 1963686155;
assign addr[62551]= 2020577882;
assign addr[62552]= 2067219829;
assign addr[62553]= 2103375398;
assign addr[62554]= 2128861181;
assign addr[62555]= 2143547897;
assign addr[62556]= 2147361045;
assign addr[62557]= 2140281282;
assign addr[62558]= 2122344521;
assign addr[62559]= 2093641749;
assign addr[62560]= 2054318569;
assign addr[62561]= 2004574453;
assign addr[62562]= 1944661739;
assign addr[62563]= 1874884346;
assign addr[62564]= 1795596234;
assign addr[62565]= 1707199606;
assign addr[62566]= 1610142873;
assign addr[62567]= 1504918373;
assign addr[62568]= 1392059879;
assign addr[62569]= 1272139887;
assign addr[62570]= 1145766716;
assign addr[62571]= 1013581418;
assign addr[62572]= 876254528;
assign addr[62573]= 734482665;
assign addr[62574]= 588984994;
assign addr[62575]= 440499581;
assign addr[62576]= 289779648;
assign addr[62577]= 137589750;
assign addr[62578]= -15298099;
assign addr[62579]= -168108346;
assign addr[62580]= -320065829;
assign addr[62581]= -470399716;
assign addr[62582]= -618347408;
assign addr[62583]= -763158411;
assign addr[62584]= -904098143;
assign addr[62585]= -1040451659;
assign addr[62586]= -1171527280;
assign addr[62587]= -1296660098;
assign addr[62588]= -1415215352;
assign addr[62589]= -1526591649;
assign addr[62590]= -1630224009;
assign addr[62591]= -1725586737;
assign addr[62592]= -1812196087;
assign addr[62593]= -1889612716;
assign addr[62594]= -1957443913;
assign addr[62595]= -2015345591;
assign addr[62596]= -2063024031;
assign addr[62597]= -2100237377;
assign addr[62598]= -2126796855;
assign addr[62599]= -2142567738;
assign addr[62600]= -2147470025;
assign addr[62601]= -2141478848;
assign addr[62602]= -2124624598;
assign addr[62603]= -2096992772;
assign addr[62604]= -2058723538;
assign addr[62605]= -2010011024;
assign addr[62606]= -1951102334;
assign addr[62607]= -1882296293;
assign addr[62608]= -1803941934;
assign addr[62609]= -1716436725;
assign addr[62610]= -1620224553;
assign addr[62611]= -1515793473;
assign addr[62612]= -1403673233;
assign addr[62613]= -1284432584;
assign addr[62614]= -1158676398;
assign addr[62615]= -1027042599;
assign addr[62616]= -890198924;
assign addr[62617]= -748839539;
assign addr[62618]= -603681519;
assign addr[62619]= -455461206;
assign addr[62620]= -304930476;
assign addr[62621]= -152852926;
assign addr[62622]= 0;
assign addr[62623]= 152852926;
assign addr[62624]= 304930476;
assign addr[62625]= 455461206;
assign addr[62626]= 603681519;
assign addr[62627]= 748839539;
assign addr[62628]= 890198924;
assign addr[62629]= 1027042599;
assign addr[62630]= 1158676398;
assign addr[62631]= 1284432584;
assign addr[62632]= 1403673233;
assign addr[62633]= 1515793473;
assign addr[62634]= 1620224553;
assign addr[62635]= 1716436725;
assign addr[62636]= 1803941934;
assign addr[62637]= 1882296293;
assign addr[62638]= 1951102334;
assign addr[62639]= 2010011024;
assign addr[62640]= 2058723538;
assign addr[62641]= 2096992772;
assign addr[62642]= 2124624598;
assign addr[62643]= 2141478848;
assign addr[62644]= 2147470025;
assign addr[62645]= 2142567738;
assign addr[62646]= 2126796855;
assign addr[62647]= 2100237377;
assign addr[62648]= 2063024031;
assign addr[62649]= 2015345591;
assign addr[62650]= 1957443913;
assign addr[62651]= 1889612716;
assign addr[62652]= 1812196087;
assign addr[62653]= 1725586737;
assign addr[62654]= 1630224009;
assign addr[62655]= 1526591649;
assign addr[62656]= 1415215352;
assign addr[62657]= 1296660098;
assign addr[62658]= 1171527280;
assign addr[62659]= 1040451659;
assign addr[62660]= 904098143;
assign addr[62661]= 763158411;
assign addr[62662]= 618347408;
assign addr[62663]= 470399716;
assign addr[62664]= 320065829;
assign addr[62665]= 168108346;
assign addr[62666]= 15298099;
assign addr[62667]= -137589750;
assign addr[62668]= -289779648;
assign addr[62669]= -440499581;
assign addr[62670]= -588984994;
assign addr[62671]= -734482665;
assign addr[62672]= -876254528;
assign addr[62673]= -1013581418;
assign addr[62674]= -1145766716;
assign addr[62675]= -1272139887;
assign addr[62676]= -1392059879;
assign addr[62677]= -1504918373;
assign addr[62678]= -1610142873;
assign addr[62679]= -1707199606;
assign addr[62680]= -1795596234;
assign addr[62681]= -1874884346;
assign addr[62682]= -1944661739;
assign addr[62683]= -2004574453;
assign addr[62684]= -2054318569;
assign addr[62685]= -2093641749;
assign addr[62686]= -2122344521;
assign addr[62687]= -2140281282;
assign addr[62688]= -2147361045;
assign addr[62689]= -2143547897;
assign addr[62690]= -2128861181;
assign addr[62691]= -2103375398;
assign addr[62692]= -2067219829;
assign addr[62693]= -2020577882;
assign addr[62694]= -1963686155;
assign addr[62695]= -1896833245;
assign addr[62696]= -1820358275;
assign addr[62697]= -1734649179;
assign addr[62698]= -1640140734;
assign addr[62699]= -1537312353;
assign addr[62700]= -1426685652;
assign addr[62701]= -1308821808;
assign addr[62702]= -1184318708;
assign addr[62703]= -1053807919;
assign addr[62704]= -917951481;
assign addr[62705]= -777438554;
assign addr[62706]= -632981917;
assign addr[62707]= -485314355;
assign addr[62708]= -335184940;
assign addr[62709]= -183355234;
assign addr[62710]= -30595422;
assign addr[62711]= 122319591;
assign addr[62712]= 274614114;
assign addr[62713]= 425515602;
assign addr[62714]= 574258580;
assign addr[62715]= 720088517;
assign addr[62716]= 862265664;
assign addr[62717]= 1000068799;
assign addr[62718]= 1132798888;
assign addr[62719]= 1259782632;
assign addr[62720]= 1380375881;
assign addr[62721]= 1493966902;
assign addr[62722]= 1599979481;
assign addr[62723]= 1697875851;
assign addr[62724]= 1787159411;
assign addr[62725]= 1867377253;
assign addr[62726]= 1938122457;
assign addr[62727]= 1999036154;
assign addr[62728]= 2049809346;
assign addr[62729]= 2090184478;
assign addr[62730]= 2119956737;
assign addr[62731]= 2138975100;
assign addr[62732]= 2147143090;
assign addr[62733]= 2144419275;
assign addr[62734]= 2130817471;
assign addr[62735]= 2106406677;
assign addr[62736]= 2071310720;
assign addr[62737]= 2025707632;
assign addr[62738]= 1969828744;
assign addr[62739]= 1903957513;
assign addr[62740]= 1828428082;
assign addr[62741]= 1743623590;
assign addr[62742]= 1649974225;
assign addr[62743]= 1547955041;
assign addr[62744]= 1438083551;
assign addr[62745]= 1320917099;
assign addr[62746]= 1197050035;
assign addr[62747]= 1067110699;
assign addr[62748]= 931758235;
assign addr[62749]= 791679244;
assign addr[62750]= 647584304;
assign addr[62751]= 500204365;
assign addr[62752]= 350287041;
assign addr[62753]= 198592817;
assign addr[62754]= 45891193;
assign addr[62755]= -107043224;
assign addr[62756]= -259434643;
assign addr[62757]= -410510029;
assign addr[62758]= -559503022;
assign addr[62759]= -705657826;
assign addr[62760]= -848233042;
assign addr[62761]= -986505429;
assign addr[62762]= -1119773573;
assign addr[62763]= -1247361445;
assign addr[62764]= -1368621831;
assign addr[62765]= -1482939614;
assign addr[62766]= -1589734894;
assign addr[62767]= -1688465931;
assign addr[62768]= -1778631892;
assign addr[62769]= -1859775393;
assign addr[62770]= -1931484818;
assign addr[62771]= -1993396407;
assign addr[62772]= -2045196100;
assign addr[62773]= -2086621133;
assign addr[62774]= -2117461370;
assign addr[62775]= -2137560369;
assign addr[62776]= -2146816171;
assign addr[62777]= -2145181827;
assign addr[62778]= -2132665626;
assign addr[62779]= -2109331059;
assign addr[62780]= -2075296495;
assign addr[62781]= -2030734582;
assign addr[62782]= -1975871368;
assign addr[62783]= -1910985158;
assign addr[62784]= -1836405100;
assign addr[62785]= -1752509516;
assign addr[62786]= -1659723983;
assign addr[62787]= -1558519173;
assign addr[62788]= -1449408469;
assign addr[62789]= -1332945355;
assign addr[62790]= -1209720613;
assign addr[62791]= -1080359326;
assign addr[62792]= -945517704;
assign addr[62793]= -805879757;
assign addr[62794]= -662153826;
assign addr[62795]= -515068990;
assign addr[62796]= -365371365;
assign addr[62797]= -213820322;
assign addr[62798]= -61184634;
assign addr[62799]= 91761426;
assign addr[62800]= 244242007;
assign addr[62801]= 395483624;
assign addr[62802]= 544719071;
assign addr[62803]= 691191324;
assign addr[62804]= 834157373;
assign addr[62805]= 972891995;
assign addr[62806]= 1106691431;
assign addr[62807]= 1234876957;
assign addr[62808]= 1356798326;
assign addr[62809]= 1471837070;
assign addr[62810]= 1579409630;
assign addr[62811]= 1678970324;
assign addr[62812]= 1770014111;
assign addr[62813]= 1852079154;
assign addr[62814]= 1924749160;
assign addr[62815]= 1987655498;
assign addr[62816]= 2040479063;
assign addr[62817]= 2082951896;
assign addr[62818]= 2114858546;
assign addr[62819]= 2136037160;
assign addr[62820]= 2146380306;
assign addr[62821]= 2145835515;
assign addr[62822]= 2134405552;
assign addr[62823]= 2112148396;
assign addr[62824]= 2079176953;
assign addr[62825]= 2035658475;
assign addr[62826]= 1981813720;
assign addr[62827]= 1917915825;
assign addr[62828]= 1844288924;
assign addr[62829]= 1761306505;
assign addr[62830]= 1669389513;
assign addr[62831]= 1569004214;
assign addr[62832]= 1460659832;
assign addr[62833]= 1344905966;
assign addr[62834]= 1222329801;
assign addr[62835]= 1093553126;
assign addr[62836]= 959229189;
assign addr[62837]= 820039373;
assign addr[62838]= 676689746;
assign addr[62839]= 529907477;
assign addr[62840]= 380437148;
assign addr[62841]= 229036977;
assign addr[62842]= 76474970;
assign addr[62843]= -76474970;
assign addr[62844]= -229036977;
assign addr[62845]= -380437148;
assign addr[62846]= -529907477;
assign addr[62847]= -676689746;
assign addr[62848]= -820039373;
assign addr[62849]= -959229189;
assign addr[62850]= -1093553126;
assign addr[62851]= -1222329801;
assign addr[62852]= -1344905966;
assign addr[62853]= -1460659832;
assign addr[62854]= -1569004214;
assign addr[62855]= -1669389513;
assign addr[62856]= -1761306505;
assign addr[62857]= -1844288924;
assign addr[62858]= -1917915825;
assign addr[62859]= -1981813720;
assign addr[62860]= -2035658475;
assign addr[62861]= -2079176953;
assign addr[62862]= -2112148396;
assign addr[62863]= -2134405552;
assign addr[62864]= -2145835515;
assign addr[62865]= -2146380306;
assign addr[62866]= -2136037160;
assign addr[62867]= -2114858546;
assign addr[62868]= -2082951896;
assign addr[62869]= -2040479063;
assign addr[62870]= -1987655498;
assign addr[62871]= -1924749160;
assign addr[62872]= -1852079154;
assign addr[62873]= -1770014111;
assign addr[62874]= -1678970324;
assign addr[62875]= -1579409630;
assign addr[62876]= -1471837070;
assign addr[62877]= -1356798326;
assign addr[62878]= -1234876957;
assign addr[62879]= -1106691431;
assign addr[62880]= -972891995;
assign addr[62881]= -834157373;
assign addr[62882]= -691191324;
assign addr[62883]= -544719071;
assign addr[62884]= -395483624;
assign addr[62885]= -244242007;
assign addr[62886]= -91761426;
assign addr[62887]= 61184634;
assign addr[62888]= 213820322;
assign addr[62889]= 365371365;
assign addr[62890]= 515068990;
assign addr[62891]= 662153826;
assign addr[62892]= 805879757;
assign addr[62893]= 945517704;
assign addr[62894]= 1080359326;
assign addr[62895]= 1209720613;
assign addr[62896]= 1332945355;
assign addr[62897]= 1449408469;
assign addr[62898]= 1558519173;
assign addr[62899]= 1659723983;
assign addr[62900]= 1752509516;
assign addr[62901]= 1836405100;
assign addr[62902]= 1910985158;
assign addr[62903]= 1975871368;
assign addr[62904]= 2030734582;
assign addr[62905]= 2075296495;
assign addr[62906]= 2109331059;
assign addr[62907]= 2132665626;
assign addr[62908]= 2145181827;
assign addr[62909]= 2146816171;
assign addr[62910]= 2137560369;
assign addr[62911]= 2117461370;
assign addr[62912]= 2086621133;
assign addr[62913]= 2045196100;
assign addr[62914]= 1993396407;
assign addr[62915]= 1931484818;
assign addr[62916]= 1859775393;
assign addr[62917]= 1778631892;
assign addr[62918]= 1688465931;
assign addr[62919]= 1589734894;
assign addr[62920]= 1482939614;
assign addr[62921]= 1368621831;
assign addr[62922]= 1247361445;
assign addr[62923]= 1119773573;
assign addr[62924]= 986505429;
assign addr[62925]= 848233042;
assign addr[62926]= 705657826;
assign addr[62927]= 559503022;
assign addr[62928]= 410510029;
assign addr[62929]= 259434643;
assign addr[62930]= 107043224;
assign addr[62931]= -45891193;
assign addr[62932]= -198592817;
assign addr[62933]= -350287041;
assign addr[62934]= -500204365;
assign addr[62935]= -647584304;
assign addr[62936]= -791679244;
assign addr[62937]= -931758235;
assign addr[62938]= -1067110699;
assign addr[62939]= -1197050035;
assign addr[62940]= -1320917099;
assign addr[62941]= -1438083551;
assign addr[62942]= -1547955041;
assign addr[62943]= -1649974225;
assign addr[62944]= -1743623590;
assign addr[62945]= -1828428082;
assign addr[62946]= -1903957513;
assign addr[62947]= -1969828744;
assign addr[62948]= -2025707632;
assign addr[62949]= -2071310720;
assign addr[62950]= -2106406677;
assign addr[62951]= -2130817471;
assign addr[62952]= -2144419275;
assign addr[62953]= -2147143090;
assign addr[62954]= -2138975100;
assign addr[62955]= -2119956737;
assign addr[62956]= -2090184478;
assign addr[62957]= -2049809346;
assign addr[62958]= -1999036154;
assign addr[62959]= -1938122457;
assign addr[62960]= -1867377253;
assign addr[62961]= -1787159411;
assign addr[62962]= -1697875851;
assign addr[62963]= -1599979481;
assign addr[62964]= -1493966902;
assign addr[62965]= -1380375881;
assign addr[62966]= -1259782632;
assign addr[62967]= -1132798888;
assign addr[62968]= -1000068799;
assign addr[62969]= -862265664;
assign addr[62970]= -720088517;
assign addr[62971]= -574258580;
assign addr[62972]= -425515602;
assign addr[62973]= -274614114;
assign addr[62974]= -122319591;
assign addr[62975]= 30595422;
assign addr[62976]= 183355234;
assign addr[62977]= 335184940;
assign addr[62978]= 485314355;
assign addr[62979]= 632981917;
assign addr[62980]= 777438554;
assign addr[62981]= 917951481;
assign addr[62982]= 1053807919;
assign addr[62983]= 1184318708;
assign addr[62984]= 1308821808;
assign addr[62985]= 1426685652;
assign addr[62986]= 1537312353;
assign addr[62987]= 1640140734;
assign addr[62988]= 1734649179;
assign addr[62989]= 1820358275;
assign addr[62990]= 1896833245;
assign addr[62991]= 1963686155;
assign addr[62992]= 2020577882;
assign addr[62993]= 2067219829;
assign addr[62994]= 2103375398;
assign addr[62995]= 2128861181;
assign addr[62996]= 2143547897;
assign addr[62997]= 2147361045;
assign addr[62998]= 2140281282;
assign addr[62999]= 2122344521;
assign addr[63000]= 2093641749;
assign addr[63001]= 2054318569;
assign addr[63002]= 2004574453;
assign addr[63003]= 1944661739;
assign addr[63004]= 1874884346;
assign addr[63005]= 1795596234;
assign addr[63006]= 1707199606;
assign addr[63007]= 1610142873;
assign addr[63008]= 1504918373;
assign addr[63009]= 1392059879;
assign addr[63010]= 1272139887;
assign addr[63011]= 1145766716;
assign addr[63012]= 1013581418;
assign addr[63013]= 876254528;
assign addr[63014]= 734482665;
assign addr[63015]= 588984994;
assign addr[63016]= 440499581;
assign addr[63017]= 289779648;
assign addr[63018]= 137589750;
assign addr[63019]= -15298099;
assign addr[63020]= -168108346;
assign addr[63021]= -320065829;
assign addr[63022]= -470399716;
assign addr[63023]= -618347408;
assign addr[63024]= -763158411;
assign addr[63025]= -904098143;
assign addr[63026]= -1040451659;
assign addr[63027]= -1171527280;
assign addr[63028]= -1296660098;
assign addr[63029]= -1415215352;
assign addr[63030]= -1526591649;
assign addr[63031]= -1630224009;
assign addr[63032]= -1725586737;
assign addr[63033]= -1812196087;
assign addr[63034]= -1889612716;
assign addr[63035]= -1957443913;
assign addr[63036]= -2015345591;
assign addr[63037]= -2063024031;
assign addr[63038]= -2100237377;
assign addr[63039]= -2126796855;
assign addr[63040]= -2142567738;
assign addr[63041]= -2147470025;
assign addr[63042]= -2141478848;
assign addr[63043]= -2124624598;
assign addr[63044]= -2096992772;
assign addr[63045]= -2058723538;
assign addr[63046]= -2010011024;
assign addr[63047]= -1951102334;
assign addr[63048]= -1882296293;
assign addr[63049]= -1803941934;
assign addr[63050]= -1716436725;
assign addr[63051]= -1620224553;
assign addr[63052]= -1515793473;
assign addr[63053]= -1403673233;
assign addr[63054]= -1284432584;
assign addr[63055]= -1158676398;
assign addr[63056]= -1027042599;
assign addr[63057]= -890198924;
assign addr[63058]= -748839539;
assign addr[63059]= -603681519;
assign addr[63060]= -455461206;
assign addr[63061]= -304930476;
assign addr[63062]= -152852926;
assign addr[63063]= 0;
assign addr[63064]= 152852926;
assign addr[63065]= 304930476;
assign addr[63066]= 455461206;
assign addr[63067]= 603681519;
assign addr[63068]= 748839539;
assign addr[63069]= 890198924;
assign addr[63070]= 1027042599;
assign addr[63071]= 1158676398;
assign addr[63072]= 1284432584;
assign addr[63073]= 1403673233;
assign addr[63074]= 1515793473;
assign addr[63075]= 1620224553;
assign addr[63076]= 1716436725;
assign addr[63077]= 1803941934;
assign addr[63078]= 1882296293;
assign addr[63079]= 1951102334;
assign addr[63080]= 2010011024;
assign addr[63081]= 2058723538;
assign addr[63082]= 2096992772;
assign addr[63083]= 2124624598;
assign addr[63084]= 2141478848;
assign addr[63085]= 2147470025;
assign addr[63086]= 2142567738;
assign addr[63087]= 2126796855;
assign addr[63088]= 2100237377;
assign addr[63089]= 2063024031;
assign addr[63090]= 2015345591;
assign addr[63091]= 1957443913;
assign addr[63092]= 1889612716;
assign addr[63093]= 1812196087;
assign addr[63094]= 1725586737;
assign addr[63095]= 1630224009;
assign addr[63096]= 1526591649;
assign addr[63097]= 1415215352;
assign addr[63098]= 1296660098;
assign addr[63099]= 1171527280;
assign addr[63100]= 1040451659;
assign addr[63101]= 904098143;
assign addr[63102]= 763158411;
assign addr[63103]= 618347408;
assign addr[63104]= 470399716;
assign addr[63105]= 320065829;
assign addr[63106]= 168108346;
assign addr[63107]= 15298099;
assign addr[63108]= -137589750;
assign addr[63109]= -289779648;
assign addr[63110]= -440499581;
assign addr[63111]= -588984994;
assign addr[63112]= -734482665;
assign addr[63113]= -876254528;
assign addr[63114]= -1013581418;
assign addr[63115]= -1145766716;
assign addr[63116]= -1272139887;
assign addr[63117]= -1392059879;
assign addr[63118]= -1504918373;
assign addr[63119]= -1610142873;
assign addr[63120]= -1707199606;
assign addr[63121]= -1795596234;
assign addr[63122]= -1874884346;
assign addr[63123]= -1944661739;
assign addr[63124]= -2004574453;
assign addr[63125]= -2054318569;
assign addr[63126]= -2093641749;
assign addr[63127]= -2122344521;
assign addr[63128]= -2140281282;
assign addr[63129]= -2147361045;
assign addr[63130]= -2143547897;
assign addr[63131]= -2128861181;
assign addr[63132]= -2103375398;
assign addr[63133]= -2067219829;
assign addr[63134]= -2020577882;
assign addr[63135]= -1963686155;
assign addr[63136]= -1896833245;
assign addr[63137]= -1820358275;
assign addr[63138]= -1734649179;
assign addr[63139]= -1640140734;
assign addr[63140]= -1537312353;
assign addr[63141]= -1426685652;
assign addr[63142]= -1308821808;
assign addr[63143]= -1184318708;
assign addr[63144]= -1053807919;
assign addr[63145]= -917951481;
assign addr[63146]= -777438554;
assign addr[63147]= -632981917;
assign addr[63148]= -485314355;
assign addr[63149]= -335184940;
assign addr[63150]= -183355234;
assign addr[63151]= -30595422;
assign addr[63152]= 122319591;
assign addr[63153]= 274614114;
assign addr[63154]= 425515602;
assign addr[63155]= 574258580;
assign addr[63156]= 720088517;
assign addr[63157]= 862265664;
assign addr[63158]= 1000068799;
assign addr[63159]= 1132798888;
assign addr[63160]= 1259782632;
assign addr[63161]= 1380375881;
assign addr[63162]= 1493966902;
assign addr[63163]= 1599979481;
assign addr[63164]= 1697875851;
assign addr[63165]= 1787159411;
assign addr[63166]= 1867377253;
assign addr[63167]= 1938122457;
assign addr[63168]= 1999036154;
assign addr[63169]= 2049809346;
assign addr[63170]= 2090184478;
assign addr[63171]= 2119956737;
assign addr[63172]= 2138975100;
assign addr[63173]= 2147143090;
assign addr[63174]= 2144419275;
assign addr[63175]= 2130817471;
assign addr[63176]= 2106406677;
assign addr[63177]= 2071310720;
assign addr[63178]= 2025707632;
assign addr[63179]= 1969828744;
assign addr[63180]= 1903957513;
assign addr[63181]= 1828428082;
assign addr[63182]= 1743623590;
assign addr[63183]= 1649974225;
assign addr[63184]= 1547955041;
assign addr[63185]= 1438083551;
assign addr[63186]= 1320917099;
assign addr[63187]= 1197050035;
assign addr[63188]= 1067110699;
assign addr[63189]= 931758235;
assign addr[63190]= 791679244;
assign addr[63191]= 647584304;
assign addr[63192]= 500204365;
assign addr[63193]= 350287041;
assign addr[63194]= 198592817;
assign addr[63195]= 45891193;
assign addr[63196]= -107043224;
assign addr[63197]= -259434643;
assign addr[63198]= -410510029;
assign addr[63199]= -559503022;
assign addr[63200]= -705657826;
assign addr[63201]= -848233042;
assign addr[63202]= -986505429;
assign addr[63203]= -1119773573;
assign addr[63204]= -1247361445;
assign addr[63205]= -1368621831;
assign addr[63206]= -1482939614;
assign addr[63207]= -1589734894;
assign addr[63208]= -1688465931;
assign addr[63209]= -1778631892;
assign addr[63210]= -1859775393;
assign addr[63211]= -1931484818;
assign addr[63212]= -1993396407;
assign addr[63213]= -2045196100;
assign addr[63214]= -2086621133;
assign addr[63215]= -2117461370;
assign addr[63216]= -2137560369;
assign addr[63217]= -2146816171;
assign addr[63218]= -2145181827;
assign addr[63219]= -2132665626;
assign addr[63220]= -2109331059;
assign addr[63221]= -2075296495;
assign addr[63222]= -2030734582;
assign addr[63223]= -1975871368;
assign addr[63224]= -1910985158;
assign addr[63225]= -1836405100;
assign addr[63226]= -1752509516;
assign addr[63227]= -1659723983;
assign addr[63228]= -1558519173;
assign addr[63229]= -1449408469;
assign addr[63230]= -1332945355;
assign addr[63231]= -1209720613;
assign addr[63232]= -1080359326;
assign addr[63233]= -945517704;
assign addr[63234]= -805879757;
assign addr[63235]= -662153826;
assign addr[63236]= -515068990;
assign addr[63237]= -365371365;
assign addr[63238]= -213820322;
assign addr[63239]= -61184634;
assign addr[63240]= 91761426;
assign addr[63241]= 244242007;
assign addr[63242]= 395483624;
assign addr[63243]= 544719071;
assign addr[63244]= 691191324;
assign addr[63245]= 834157373;
assign addr[63246]= 972891995;
assign addr[63247]= 1106691431;
assign addr[63248]= 1234876957;
assign addr[63249]= 1356798326;
assign addr[63250]= 1471837070;
assign addr[63251]= 1579409630;
assign addr[63252]= 1678970324;
assign addr[63253]= 1770014111;
assign addr[63254]= 1852079154;
assign addr[63255]= 1924749160;
assign addr[63256]= 1987655498;
assign addr[63257]= 2040479063;
assign addr[63258]= 2082951896;
assign addr[63259]= 2114858546;
assign addr[63260]= 2136037160;
assign addr[63261]= 2146380306;
assign addr[63262]= 2145835515;
assign addr[63263]= 2134405552;
assign addr[63264]= 2112148396;
assign addr[63265]= 2079176953;
assign addr[63266]= 2035658475;
assign addr[63267]= 1981813720;
assign addr[63268]= 1917915825;
assign addr[63269]= 1844288924;
assign addr[63270]= 1761306505;
assign addr[63271]= 1669389513;
assign addr[63272]= 1569004214;
assign addr[63273]= 1460659832;
assign addr[63274]= 1344905966;
assign addr[63275]= 1222329801;
assign addr[63276]= 1093553126;
assign addr[63277]= 959229189;
assign addr[63278]= 820039373;
assign addr[63279]= 676689746;
assign addr[63280]= 529907477;
assign addr[63281]= 380437148;
assign addr[63282]= 229036977;
assign addr[63283]= 76474970;
assign addr[63284]= -76474970;
assign addr[63285]= -229036977;
assign addr[63286]= -380437148;
assign addr[63287]= -529907477;
assign addr[63288]= -676689746;
assign addr[63289]= -820039373;
assign addr[63290]= -959229189;
assign addr[63291]= -1093553126;
assign addr[63292]= -1222329801;
assign addr[63293]= -1344905966;
assign addr[63294]= -1460659832;
assign addr[63295]= -1569004214;
assign addr[63296]= -1669389513;
assign addr[63297]= -1761306505;
assign addr[63298]= -1844288924;
assign addr[63299]= -1917915825;
assign addr[63300]= -1981813720;
assign addr[63301]= -2035658475;
assign addr[63302]= -2079176953;
assign addr[63303]= -2112148396;
assign addr[63304]= -2134405552;
assign addr[63305]= -2145835515;
assign addr[63306]= -2146380306;
assign addr[63307]= -2136037160;
assign addr[63308]= -2114858546;
assign addr[63309]= -2082951896;
assign addr[63310]= -2040479063;
assign addr[63311]= -1987655498;
assign addr[63312]= -1924749160;
assign addr[63313]= -1852079154;
assign addr[63314]= -1770014111;
assign addr[63315]= -1678970324;
assign addr[63316]= -1579409630;
assign addr[63317]= -1471837070;
assign addr[63318]= -1356798326;
assign addr[63319]= -1234876957;
assign addr[63320]= -1106691431;
assign addr[63321]= -972891995;
assign addr[63322]= -834157373;
assign addr[63323]= -691191324;
assign addr[63324]= -544719071;
assign addr[63325]= -395483624;
assign addr[63326]= -244242007;
assign addr[63327]= -91761426;
assign addr[63328]= 61184634;
assign addr[63329]= 213820322;
assign addr[63330]= 365371365;
assign addr[63331]= 515068990;
assign addr[63332]= 662153826;
assign addr[63333]= 805879757;
assign addr[63334]= 945517704;
assign addr[63335]= 1080359326;
assign addr[63336]= 1209720613;
assign addr[63337]= 1332945355;
assign addr[63338]= 1449408469;
assign addr[63339]= 1558519173;
assign addr[63340]= 1659723983;
assign addr[63341]= 1752509516;
assign addr[63342]= 1836405100;
assign addr[63343]= 1910985158;
assign addr[63344]= 1975871368;
assign addr[63345]= 2030734582;
assign addr[63346]= 2075296495;
assign addr[63347]= 2109331059;
assign addr[63348]= 2132665626;
assign addr[63349]= 2145181827;
assign addr[63350]= 2146816171;
assign addr[63351]= 2137560369;
assign addr[63352]= 2117461370;
assign addr[63353]= 2086621133;
assign addr[63354]= 2045196100;
assign addr[63355]= 1993396407;
assign addr[63356]= 1931484818;
assign addr[63357]= 1859775393;
assign addr[63358]= 1778631892;
assign addr[63359]= 1688465931;
assign addr[63360]= 1589734894;
assign addr[63361]= 1482939614;
assign addr[63362]= 1368621831;
assign addr[63363]= 1247361445;
assign addr[63364]= 1119773573;
assign addr[63365]= 986505429;
assign addr[63366]= 848233042;
assign addr[63367]= 705657826;
assign addr[63368]= 559503022;
assign addr[63369]= 410510029;
assign addr[63370]= 259434643;
assign addr[63371]= 107043224;
assign addr[63372]= -45891193;
assign addr[63373]= -198592817;
assign addr[63374]= -350287041;
assign addr[63375]= -500204365;
assign addr[63376]= -647584304;
assign addr[63377]= -791679244;
assign addr[63378]= -931758235;
assign addr[63379]= -1067110699;
assign addr[63380]= -1197050035;
assign addr[63381]= -1320917099;
assign addr[63382]= -1438083551;
assign addr[63383]= -1547955041;
assign addr[63384]= -1649974225;
assign addr[63385]= -1743623590;
assign addr[63386]= -1828428082;
assign addr[63387]= -1903957513;
assign addr[63388]= -1969828744;
assign addr[63389]= -2025707632;
assign addr[63390]= -2071310720;
assign addr[63391]= -2106406677;
assign addr[63392]= -2130817471;
assign addr[63393]= -2144419275;
assign addr[63394]= -2147143090;
assign addr[63395]= -2138975100;
assign addr[63396]= -2119956737;
assign addr[63397]= -2090184478;
assign addr[63398]= -2049809346;
assign addr[63399]= -1999036154;
assign addr[63400]= -1938122457;
assign addr[63401]= -1867377253;
assign addr[63402]= -1787159411;
assign addr[63403]= -1697875851;
assign addr[63404]= -1599979481;
assign addr[63405]= -1493966902;
assign addr[63406]= -1380375881;
assign addr[63407]= -1259782632;
assign addr[63408]= -1132798888;
assign addr[63409]= -1000068799;
assign addr[63410]= -862265664;
assign addr[63411]= -720088517;
assign addr[63412]= -574258580;
assign addr[63413]= -425515602;
assign addr[63414]= -274614114;
assign addr[63415]= -122319591;
assign addr[63416]= 30595422;
assign addr[63417]= 183355234;
assign addr[63418]= 335184940;
assign addr[63419]= 485314355;
assign addr[63420]= 632981917;
assign addr[63421]= 777438554;
assign addr[63422]= 917951481;
assign addr[63423]= 1053807919;
assign addr[63424]= 1184318708;
assign addr[63425]= 1308821808;
assign addr[63426]= 1426685652;
assign addr[63427]= 1537312353;
assign addr[63428]= 1640140734;
assign addr[63429]= 1734649179;
assign addr[63430]= 1820358275;
assign addr[63431]= 1896833245;
assign addr[63432]= 1963686155;
assign addr[63433]= 2020577882;
assign addr[63434]= 2067219829;
assign addr[63435]= 2103375398;
assign addr[63436]= 2128861181;
assign addr[63437]= 2143547897;
assign addr[63438]= 2147361045;
assign addr[63439]= 2140281282;
assign addr[63440]= 2122344521;
assign addr[63441]= 2093641749;
assign addr[63442]= 2054318569;
assign addr[63443]= 2004574453;
assign addr[63444]= 1944661739;
assign addr[63445]= 1874884346;
assign addr[63446]= 1795596234;
assign addr[63447]= 1707199606;
assign addr[63448]= 1610142873;
assign addr[63449]= 1504918373;
assign addr[63450]= 1392059879;
assign addr[63451]= 1272139887;
assign addr[63452]= 1145766716;
assign addr[63453]= 1013581418;
assign addr[63454]= 876254528;
assign addr[63455]= 734482665;
assign addr[63456]= 588984994;
assign addr[63457]= 440499581;
assign addr[63458]= 289779648;
assign addr[63459]= 137589750;
assign addr[63460]= -15298099;
assign addr[63461]= -168108346;
assign addr[63462]= -320065829;
assign addr[63463]= -470399716;
assign addr[63464]= -618347408;
assign addr[63465]= -763158411;
assign addr[63466]= -904098143;
assign addr[63467]= -1040451659;
assign addr[63468]= -1171527280;
assign addr[63469]= -1296660098;
assign addr[63470]= -1415215352;
assign addr[63471]= -1526591649;
assign addr[63472]= -1630224009;
assign addr[63473]= -1725586737;
assign addr[63474]= -1812196087;
assign addr[63475]= -1889612716;
assign addr[63476]= -1957443913;
assign addr[63477]= -2015345591;
assign addr[63478]= -2063024031;
assign addr[63479]= -2100237377;
assign addr[63480]= -2126796855;
assign addr[63481]= -2142567738;
assign addr[63482]= -2147470025;
assign addr[63483]= -2141478848;
assign addr[63484]= -2124624598;
assign addr[63485]= -2096992772;
assign addr[63486]= -2058723538;
assign addr[63487]= -2010011024;
assign addr[63488]= -1951102334;
assign addr[63489]= -1882296293;
assign addr[63490]= -1803941934;
assign addr[63491]= -1716436725;
assign addr[63492]= -1620224553;
assign addr[63493]= -1515793473;
assign addr[63494]= -1403673233;
assign addr[63495]= -1284432584;
assign addr[63496]= -1158676398;
assign addr[63497]= -1027042599;
assign addr[63498]= -890198924;
assign addr[63499]= -748839539;
assign addr[63500]= -603681519;
assign addr[63501]= -455461206;
assign addr[63502]= -304930476;
assign addr[63503]= -152852926;
assign addr[63504]= 0;
assign addr[63505]= 152852926;
assign addr[63506]= 304930476;
assign addr[63507]= 455461206;
assign addr[63508]= 603681519;
assign addr[63509]= 748839539;
assign addr[63510]= 890198924;
assign addr[63511]= 1027042599;
assign addr[63512]= 1158676398;
assign addr[63513]= 1284432584;
assign addr[63514]= 1403673233;
assign addr[63515]= 1515793473;
assign addr[63516]= 1620224553;
assign addr[63517]= 1716436725;
assign addr[63518]= 1803941934;
assign addr[63519]= 1882296293;
assign addr[63520]= 1951102334;
assign addr[63521]= 2010011024;
assign addr[63522]= 2058723538;
assign addr[63523]= 2096992772;
assign addr[63524]= 2124624598;
assign addr[63525]= 2141478848;
assign addr[63526]= 2147470025;
assign addr[63527]= 2142567738;
assign addr[63528]= 2126796855;
assign addr[63529]= 2100237377;
assign addr[63530]= 2063024031;
assign addr[63531]= 2015345591;
assign addr[63532]= 1957443913;
assign addr[63533]= 1889612716;
assign addr[63534]= 1812196087;
assign addr[63535]= 1725586737;
assign addr[63536]= 1630224009;
assign addr[63537]= 1526591649;
assign addr[63538]= 1415215352;
assign addr[63539]= 1296660098;
assign addr[63540]= 1171527280;
assign addr[63541]= 1040451659;
assign addr[63542]= 904098143;
assign addr[63543]= 763158411;
assign addr[63544]= 618347408;
assign addr[63545]= 470399716;
assign addr[63546]= 320065829;
assign addr[63547]= 168108346;
assign addr[63548]= 15298099;
assign addr[63549]= -137589750;
assign addr[63550]= -289779648;
assign addr[63551]= -440499581;
assign addr[63552]= -588984994;
assign addr[63553]= -734482665;
assign addr[63554]= -876254528;
assign addr[63555]= -1013581418;
assign addr[63556]= -1145766716;
assign addr[63557]= -1272139887;
assign addr[63558]= -1392059879;
assign addr[63559]= -1504918373;
assign addr[63560]= -1610142873;
assign addr[63561]= -1707199606;
assign addr[63562]= -1795596234;
assign addr[63563]= -1874884346;
assign addr[63564]= -1944661739;
assign addr[63565]= -2004574453;
assign addr[63566]= -2054318569;
assign addr[63567]= -2093641749;
assign addr[63568]= -2122344521;
assign addr[63569]= -2140281282;
assign addr[63570]= -2147361045;
assign addr[63571]= -2143547897;
assign addr[63572]= -2128861181;
assign addr[63573]= -2103375398;
assign addr[63574]= -2067219829;
assign addr[63575]= -2020577882;
assign addr[63576]= -1963686155;
assign addr[63577]= -1896833245;
assign addr[63578]= -1820358275;
assign addr[63579]= -1734649179;
assign addr[63580]= -1640140734;
assign addr[63581]= -1537312353;
assign addr[63582]= -1426685652;
assign addr[63583]= -1308821808;
assign addr[63584]= -1184318708;
assign addr[63585]= -1053807919;
assign addr[63586]= -917951481;
assign addr[63587]= -777438554;
assign addr[63588]= -632981917;
assign addr[63589]= -485314355;
assign addr[63590]= -335184940;
assign addr[63591]= -183355234;
assign addr[63592]= -30595422;
assign addr[63593]= 122319591;
assign addr[63594]= 274614114;
assign addr[63595]= 425515602;
assign addr[63596]= 574258580;
assign addr[63597]= 720088517;
assign addr[63598]= 862265664;
assign addr[63599]= 1000068799;
assign addr[63600]= 1132798888;
assign addr[63601]= 1259782632;
assign addr[63602]= 1380375881;
assign addr[63603]= 1493966902;
assign addr[63604]= 1599979481;
assign addr[63605]= 1697875851;
assign addr[63606]= 1787159411;
assign addr[63607]= 1867377253;
assign addr[63608]= 1938122457;
assign addr[63609]= 1999036154;
assign addr[63610]= 2049809346;
assign addr[63611]= 2090184478;
assign addr[63612]= 2119956737;
assign addr[63613]= 2138975100;
assign addr[63614]= 2147143090;
assign addr[63615]= 2144419275;
assign addr[63616]= 2130817471;
assign addr[63617]= 2106406677;
assign addr[63618]= 2071310720;
assign addr[63619]= 2025707632;
assign addr[63620]= 1969828744;
assign addr[63621]= 1903957513;
assign addr[63622]= 1828428082;
assign addr[63623]= 1743623590;
assign addr[63624]= 1649974225;
assign addr[63625]= 1547955041;
assign addr[63626]= 1438083551;
assign addr[63627]= 1320917099;
assign addr[63628]= 1197050035;
assign addr[63629]= 1067110699;
assign addr[63630]= 931758235;
assign addr[63631]= 791679244;
assign addr[63632]= 647584304;
assign addr[63633]= 500204365;
assign addr[63634]= 350287041;
assign addr[63635]= 198592817;
assign addr[63636]= 45891193;
assign addr[63637]= -107043224;
assign addr[63638]= -259434643;
assign addr[63639]= -410510029;
assign addr[63640]= -559503022;
assign addr[63641]= -705657826;
assign addr[63642]= -848233042;
assign addr[63643]= -986505429;
assign addr[63644]= -1119773573;
assign addr[63645]= -1247361445;
assign addr[63646]= -1368621831;
assign addr[63647]= -1482939614;
assign addr[63648]= -1589734894;
assign addr[63649]= -1688465931;
assign addr[63650]= -1778631892;
assign addr[63651]= -1859775393;
assign addr[63652]= -1931484818;
assign addr[63653]= -1993396407;
assign addr[63654]= -2045196100;
assign addr[63655]= -2086621133;
assign addr[63656]= -2117461370;
assign addr[63657]= -2137560369;
assign addr[63658]= -2146816171;
assign addr[63659]= -2145181827;
assign addr[63660]= -2132665626;
assign addr[63661]= -2109331059;
assign addr[63662]= -2075296495;
assign addr[63663]= -2030734582;
assign addr[63664]= -1975871368;
assign addr[63665]= -1910985158;
assign addr[63666]= -1836405100;
assign addr[63667]= -1752509516;
assign addr[63668]= -1659723983;
assign addr[63669]= -1558519173;
assign addr[63670]= -1449408469;
assign addr[63671]= -1332945355;
assign addr[63672]= -1209720613;
assign addr[63673]= -1080359326;
assign addr[63674]= -945517704;
assign addr[63675]= -805879757;
assign addr[63676]= -662153826;
assign addr[63677]= -515068990;
assign addr[63678]= -365371365;
assign addr[63679]= -213820322;
assign addr[63680]= -61184634;
assign addr[63681]= 91761426;
assign addr[63682]= 244242007;
assign addr[63683]= 395483624;
assign addr[63684]= 544719071;
assign addr[63685]= 691191324;
assign addr[63686]= 834157373;
assign addr[63687]= 972891995;
assign addr[63688]= 1106691431;
assign addr[63689]= 1234876957;
assign addr[63690]= 1356798326;
assign addr[63691]= 1471837070;
assign addr[63692]= 1579409630;
assign addr[63693]= 1678970324;
assign addr[63694]= 1770014111;
assign addr[63695]= 1852079154;
assign addr[63696]= 1924749160;
assign addr[63697]= 1987655498;
assign addr[63698]= 2040479063;
assign addr[63699]= 2082951896;
assign addr[63700]= 2114858546;
assign addr[63701]= 2136037160;
assign addr[63702]= 2146380306;
assign addr[63703]= 2145835515;
assign addr[63704]= 2134405552;
assign addr[63705]= 2112148396;
assign addr[63706]= 2079176953;
assign addr[63707]= 2035658475;
assign addr[63708]= 1981813720;
assign addr[63709]= 1917915825;
assign addr[63710]= 1844288924;
assign addr[63711]= 1761306505;
assign addr[63712]= 1669389513;
assign addr[63713]= 1569004214;
assign addr[63714]= 1460659832;
assign addr[63715]= 1344905966;
assign addr[63716]= 1222329801;
assign addr[63717]= 1093553126;
assign addr[63718]= 959229189;
assign addr[63719]= 820039373;
assign addr[63720]= 676689746;
assign addr[63721]= 529907477;
assign addr[63722]= 380437148;
assign addr[63723]= 229036977;
assign addr[63724]= 76474970;
assign addr[63725]= -76474970;
assign addr[63726]= -229036977;
assign addr[63727]= -380437148;
assign addr[63728]= -529907477;
assign addr[63729]= -676689746;
assign addr[63730]= -820039373;
assign addr[63731]= -959229189;
assign addr[63732]= -1093553126;
assign addr[63733]= -1222329801;
assign addr[63734]= -1344905966;
assign addr[63735]= -1460659832;
assign addr[63736]= -1569004214;
assign addr[63737]= -1669389513;
assign addr[63738]= -1761306505;
assign addr[63739]= -1844288924;
assign addr[63740]= -1917915825;
assign addr[63741]= -1981813720;
assign addr[63742]= -2035658475;
assign addr[63743]= -2079176953;
assign addr[63744]= -2112148396;
assign addr[63745]= -2134405552;
assign addr[63746]= -2145835515;
assign addr[63747]= -2146380306;
assign addr[63748]= -2136037160;
assign addr[63749]= -2114858546;
assign addr[63750]= -2082951896;
assign addr[63751]= -2040479063;
assign addr[63752]= -1987655498;
assign addr[63753]= -1924749160;
assign addr[63754]= -1852079154;
assign addr[63755]= -1770014111;
assign addr[63756]= -1678970324;
assign addr[63757]= -1579409630;
assign addr[63758]= -1471837070;
assign addr[63759]= -1356798326;
assign addr[63760]= -1234876957;
assign addr[63761]= -1106691431;
assign addr[63762]= -972891995;
assign addr[63763]= -834157373;
assign addr[63764]= -691191324;
assign addr[63765]= -544719071;
assign addr[63766]= -395483624;
assign addr[63767]= -244242007;
assign addr[63768]= -91761426;
assign addr[63769]= 61184634;
assign addr[63770]= 213820322;
assign addr[63771]= 365371365;
assign addr[63772]= 515068990;
assign addr[63773]= 662153826;
assign addr[63774]= 805879757;
assign addr[63775]= 945517704;
assign addr[63776]= 1080359326;
assign addr[63777]= 1209720613;
assign addr[63778]= 1332945355;
assign addr[63779]= 1449408469;
assign addr[63780]= 1558519173;
assign addr[63781]= 1659723983;
assign addr[63782]= 1752509516;
assign addr[63783]= 1836405100;
assign addr[63784]= 1910985158;
assign addr[63785]= 1975871368;
assign addr[63786]= 2030734582;
assign addr[63787]= 2075296495;
assign addr[63788]= 2109331059;
assign addr[63789]= 2132665626;
assign addr[63790]= 2145181827;
assign addr[63791]= 2146816171;
assign addr[63792]= 2137560369;
assign addr[63793]= 2117461370;
assign addr[63794]= 2086621133;
assign addr[63795]= 2045196100;
assign addr[63796]= 1993396407;
assign addr[63797]= 1931484818;
assign addr[63798]= 1859775393;
assign addr[63799]= 1778631892;
assign addr[63800]= 1688465931;
assign addr[63801]= 1589734894;
assign addr[63802]= 1482939614;
assign addr[63803]= 1368621831;
assign addr[63804]= 1247361445;
assign addr[63805]= 1119773573;
assign addr[63806]= 986505429;
assign addr[63807]= 848233042;
assign addr[63808]= 705657826;
assign addr[63809]= 559503022;
assign addr[63810]= 410510029;
assign addr[63811]= 259434643;
assign addr[63812]= 107043224;
assign addr[63813]= -45891193;
assign addr[63814]= -198592817;
assign addr[63815]= -350287041;
assign addr[63816]= -500204365;
assign addr[63817]= -647584304;
assign addr[63818]= -791679244;
assign addr[63819]= -931758235;
assign addr[63820]= -1067110699;
assign addr[63821]= -1197050035;
assign addr[63822]= -1320917099;
assign addr[63823]= -1438083551;
assign addr[63824]= -1547955041;
assign addr[63825]= -1649974225;
assign addr[63826]= -1743623590;
assign addr[63827]= -1828428082;
assign addr[63828]= -1903957513;
assign addr[63829]= -1969828744;
assign addr[63830]= -2025707632;
assign addr[63831]= -2071310720;
assign addr[63832]= -2106406677;
assign addr[63833]= -2130817471;
assign addr[63834]= -2144419275;
assign addr[63835]= -2147143090;
assign addr[63836]= -2138975100;
assign addr[63837]= -2119956737;
assign addr[63838]= -2090184478;
assign addr[63839]= -2049809346;
assign addr[63840]= -1999036154;
assign addr[63841]= -1938122457;
assign addr[63842]= -1867377253;
assign addr[63843]= -1787159411;
assign addr[63844]= -1697875851;
assign addr[63845]= -1599979481;
assign addr[63846]= -1493966902;
assign addr[63847]= -1380375881;
assign addr[63848]= -1259782632;
assign addr[63849]= -1132798888;
assign addr[63850]= -1000068799;
assign addr[63851]= -862265664;
assign addr[63852]= -720088517;
assign addr[63853]= -574258580;
assign addr[63854]= -425515602;
assign addr[63855]= -274614114;
assign addr[63856]= -122319591;
assign addr[63857]= 30595422;
assign addr[63858]= 183355234;
assign addr[63859]= 335184940;
assign addr[63860]= 485314355;
assign addr[63861]= 632981917;
assign addr[63862]= 777438554;
assign addr[63863]= 917951481;
assign addr[63864]= 1053807919;
assign addr[63865]= 1184318708;
assign addr[63866]= 1308821808;
assign addr[63867]= 1426685652;
assign addr[63868]= 1537312353;
assign addr[63869]= 1640140734;
assign addr[63870]= 1734649179;
assign addr[63871]= 1820358275;
assign addr[63872]= 1896833245;
assign addr[63873]= 1963686155;
assign addr[63874]= 2020577882;
assign addr[63875]= 2067219829;
assign addr[63876]= 2103375398;
assign addr[63877]= 2128861181;
assign addr[63878]= 2143547897;
assign addr[63879]= 2147361045;
assign addr[63880]= 2140281282;
assign addr[63881]= 2122344521;
assign addr[63882]= 2093641749;
assign addr[63883]= 2054318569;
assign addr[63884]= 2004574453;
assign addr[63885]= 1944661739;
assign addr[63886]= 1874884346;
assign addr[63887]= 1795596234;
assign addr[63888]= 1707199606;
assign addr[63889]= 1610142873;
assign addr[63890]= 1504918373;
assign addr[63891]= 1392059879;
assign addr[63892]= 1272139887;
assign addr[63893]= 1145766716;
assign addr[63894]= 1013581418;
assign addr[63895]= 876254528;
assign addr[63896]= 734482665;
assign addr[63897]= 588984994;
assign addr[63898]= 440499581;
assign addr[63899]= 289779648;
assign addr[63900]= 137589750;
assign addr[63901]= -15298099;
assign addr[63902]= -168108346;
assign addr[63903]= -320065829;
assign addr[63904]= -470399716;
assign addr[63905]= -618347408;
assign addr[63906]= -763158411;
assign addr[63907]= -904098143;
assign addr[63908]= -1040451659;
assign addr[63909]= -1171527280;
assign addr[63910]= -1296660098;
assign addr[63911]= -1415215352;
assign addr[63912]= -1526591649;
assign addr[63913]= -1630224009;
assign addr[63914]= -1725586737;
assign addr[63915]= -1812196087;
assign addr[63916]= -1889612716;
assign addr[63917]= -1957443913;
assign addr[63918]= -2015345591;
assign addr[63919]= -2063024031;
assign addr[63920]= -2100237377;
assign addr[63921]= -2126796855;
assign addr[63922]= -2142567738;
assign addr[63923]= -2147470025;
assign addr[63924]= -2141478848;
assign addr[63925]= -2124624598;
assign addr[63926]= -2096992772;
assign addr[63927]= -2058723538;
assign addr[63928]= -2010011024;
assign addr[63929]= -1951102334;
assign addr[63930]= -1882296293;
assign addr[63931]= -1803941934;
assign addr[63932]= -1716436725;
assign addr[63933]= -1620224553;
assign addr[63934]= -1515793473;
assign addr[63935]= -1403673233;
assign addr[63936]= -1284432584;
assign addr[63937]= -1158676398;
assign addr[63938]= -1027042599;
assign addr[63939]= -890198924;
assign addr[63940]= -748839539;
assign addr[63941]= -603681519;
assign addr[63942]= -455461206;
assign addr[63943]= -304930476;
assign addr[63944]= -152852926;
assign addr[63945]= 0;
assign addr[63946]= 152852926;
assign addr[63947]= 304930476;
assign addr[63948]= 455461206;
assign addr[63949]= 603681519;
assign addr[63950]= 748839539;
assign addr[63951]= 890198924;
assign addr[63952]= 1027042599;
assign addr[63953]= 1158676398;
assign addr[63954]= 1284432584;
assign addr[63955]= 1403673233;
assign addr[63956]= 1515793473;
assign addr[63957]= 1620224553;
assign addr[63958]= 1716436725;
assign addr[63959]= 1803941934;
assign addr[63960]= 1882296293;
assign addr[63961]= 1951102334;
assign addr[63962]= 2010011024;
assign addr[63963]= 2058723538;
assign addr[63964]= 2096992772;
assign addr[63965]= 2124624598;
assign addr[63966]= 2141478848;
assign addr[63967]= 2147470025;
assign addr[63968]= 2142567738;
assign addr[63969]= 2126796855;
assign addr[63970]= 2100237377;
assign addr[63971]= 2063024031;
assign addr[63972]= 2015345591;
assign addr[63973]= 1957443913;
assign addr[63974]= 1889612716;
assign addr[63975]= 1812196087;
assign addr[63976]= 1725586737;
assign addr[63977]= 1630224009;
assign addr[63978]= 1526591649;
assign addr[63979]= 1415215352;
assign addr[63980]= 1296660098;
assign addr[63981]= 1171527280;
assign addr[63982]= 1040451659;
assign addr[63983]= 904098143;
assign addr[63984]= 763158411;
assign addr[63985]= 618347408;
assign addr[63986]= 470399716;
assign addr[63987]= 320065829;
assign addr[63988]= 168108346;
assign addr[63989]= 15298099;
assign addr[63990]= -137589750;
assign addr[63991]= -289779648;
assign addr[63992]= -440499581;
assign addr[63993]= -588984994;
assign addr[63994]= -734482665;
assign addr[63995]= -876254528;
assign addr[63996]= -1013581418;
assign addr[63997]= -1145766716;
assign addr[63998]= -1272139887;
assign addr[63999]= -1392059879;
assign addr[64000]= -1504918373;
assign addr[64001]= -1610142873;
assign addr[64002]= -1707199606;
assign addr[64003]= -1795596234;
assign addr[64004]= -1874884346;
assign addr[64005]= -1944661739;
assign addr[64006]= -2004574453;
assign addr[64007]= -2054318569;
assign addr[64008]= -2093641749;
assign addr[64009]= -2122344521;
assign addr[64010]= -2140281282;
assign addr[64011]= -2147361045;
assign addr[64012]= -2143547897;
assign addr[64013]= -2128861181;
assign addr[64014]= -2103375398;
assign addr[64015]= -2067219829;
assign addr[64016]= -2020577882;
assign addr[64017]= -1963686155;
assign addr[64018]= -1896833245;
assign addr[64019]= -1820358275;
assign addr[64020]= -1734649179;
assign addr[64021]= -1640140734;
assign addr[64022]= -1537312353;
assign addr[64023]= -1426685652;
assign addr[64024]= -1308821808;
assign addr[64025]= -1184318708;
assign addr[64026]= -1053807919;
assign addr[64027]= -917951481;
assign addr[64028]= -777438554;
assign addr[64029]= -632981917;
assign addr[64030]= -485314355;
assign addr[64031]= -335184940;
assign addr[64032]= -183355234;
assign addr[64033]= -30595422;
assign addr[64034]= 122319591;
assign addr[64035]= 274614114;
assign addr[64036]= 425515602;
assign addr[64037]= 574258580;
assign addr[64038]= 720088517;
assign addr[64039]= 862265664;
assign addr[64040]= 1000068799;
assign addr[64041]= 1132798888;
assign addr[64042]= 1259782632;
assign addr[64043]= 1380375881;
assign addr[64044]= 1493966902;
assign addr[64045]= 1599979481;
assign addr[64046]= 1697875851;
assign addr[64047]= 1787159411;
assign addr[64048]= 1867377253;
assign addr[64049]= 1938122457;
assign addr[64050]= 1999036154;
assign addr[64051]= 2049809346;
assign addr[64052]= 2090184478;
assign addr[64053]= 2119956737;
assign addr[64054]= 2138975100;
assign addr[64055]= 2147143090;
assign addr[64056]= 2144419275;
assign addr[64057]= 2130817471;
assign addr[64058]= 2106406677;
assign addr[64059]= 2071310720;
assign addr[64060]= 2025707632;
assign addr[64061]= 1969828744;
assign addr[64062]= 1903957513;
assign addr[64063]= 1828428082;
assign addr[64064]= 1743623590;
assign addr[64065]= 1649974225;
assign addr[64066]= 1547955041;
assign addr[64067]= 1438083551;
assign addr[64068]= 1320917099;
assign addr[64069]= 1197050035;
assign addr[64070]= 1067110699;
assign addr[64071]= 931758235;
assign addr[64072]= 791679244;
assign addr[64073]= 647584304;
assign addr[64074]= 500204365;
assign addr[64075]= 350287041;
assign addr[64076]= 198592817;
assign addr[64077]= 45891193;
assign addr[64078]= -107043224;
assign addr[64079]= -259434643;
assign addr[64080]= -410510029;
assign addr[64081]= -559503022;
assign addr[64082]= -705657826;
assign addr[64083]= -848233042;
assign addr[64084]= -986505429;
assign addr[64085]= -1119773573;
assign addr[64086]= -1247361445;
assign addr[64087]= -1368621831;
assign addr[64088]= -1482939614;
assign addr[64089]= -1589734894;
assign addr[64090]= -1688465931;
assign addr[64091]= -1778631892;
assign addr[64092]= -1859775393;
assign addr[64093]= -1931484818;
assign addr[64094]= -1993396407;
assign addr[64095]= -2045196100;
assign addr[64096]= -2086621133;
assign addr[64097]= -2117461370;
assign addr[64098]= -2137560369;
assign addr[64099]= -2146816171;
assign addr[64100]= -2145181827;
assign addr[64101]= -2132665626;
assign addr[64102]= -2109331059;
assign addr[64103]= -2075296495;
assign addr[64104]= -2030734582;
assign addr[64105]= -1975871368;
assign addr[64106]= -1910985158;
assign addr[64107]= -1836405100;
assign addr[64108]= -1752509516;
assign addr[64109]= -1659723983;
assign addr[64110]= -1558519173;
assign addr[64111]= -1449408469;
assign addr[64112]= -1332945355;
assign addr[64113]= -1209720613;
assign addr[64114]= -1080359326;
assign addr[64115]= -945517704;
assign addr[64116]= -805879757;
assign addr[64117]= -662153826;
assign addr[64118]= -515068990;
assign addr[64119]= -365371365;
assign addr[64120]= -213820322;
assign addr[64121]= -61184634;
assign addr[64122]= 91761426;
assign addr[64123]= 244242007;
assign addr[64124]= 395483624;
assign addr[64125]= 544719071;
assign addr[64126]= 691191324;
assign addr[64127]= 834157373;
assign addr[64128]= 972891995;
assign addr[64129]= 1106691431;
assign addr[64130]= 1234876957;
assign addr[64131]= 1356798326;
assign addr[64132]= 1471837070;
assign addr[64133]= 1579409630;
assign addr[64134]= 1678970324;
assign addr[64135]= 1770014111;
assign addr[64136]= 1852079154;
assign addr[64137]= 1924749160;
assign addr[64138]= 1987655498;
assign addr[64139]= 2040479063;
assign addr[64140]= 2082951896;
assign addr[64141]= 2114858546;
assign addr[64142]= 2136037160;
assign addr[64143]= 2146380306;
assign addr[64144]= 2145835515;
assign addr[64145]= 2134405552;
assign addr[64146]= 2112148396;
assign addr[64147]= 2079176953;
assign addr[64148]= 2035658475;
assign addr[64149]= 1981813720;
assign addr[64150]= 1917915825;
assign addr[64151]= 1844288924;
assign addr[64152]= 1761306505;
assign addr[64153]= 1669389513;
assign addr[64154]= 1569004214;
assign addr[64155]= 1460659832;
assign addr[64156]= 1344905966;
assign addr[64157]= 1222329801;
assign addr[64158]= 1093553126;
assign addr[64159]= 959229189;
assign addr[64160]= 820039373;
assign addr[64161]= 676689746;
assign addr[64162]= 529907477;
assign addr[64163]= 380437148;
assign addr[64164]= 229036977;
assign addr[64165]= 76474970;
assign addr[64166]= -76474970;
assign addr[64167]= -229036977;
assign addr[64168]= -380437148;
assign addr[64169]= -529907477;
assign addr[64170]= -676689746;
assign addr[64171]= -820039373;
assign addr[64172]= -959229189;
assign addr[64173]= -1093553126;
assign addr[64174]= -1222329801;
assign addr[64175]= -1344905966;
assign addr[64176]= -1460659832;
assign addr[64177]= -1569004214;
assign addr[64178]= -1669389513;
assign addr[64179]= -1761306505;
assign addr[64180]= -1844288924;
assign addr[64181]= -1917915825;
assign addr[64182]= -1981813720;
assign addr[64183]= -2035658475;
assign addr[64184]= -2079176953;
assign addr[64185]= -2112148396;
assign addr[64186]= -2134405552;
assign addr[64187]= -2145835515;
assign addr[64188]= -2146380306;
assign addr[64189]= -2136037160;
assign addr[64190]= -2114858546;
assign addr[64191]= -2082951896;
assign addr[64192]= -2040479063;
assign addr[64193]= -1987655498;
assign addr[64194]= -1924749160;
assign addr[64195]= -1852079154;
assign addr[64196]= -1770014111;
assign addr[64197]= -1678970324;
assign addr[64198]= -1579409630;
assign addr[64199]= -1471837070;
assign addr[64200]= -1356798326;
assign addr[64201]= -1234876957;
assign addr[64202]= -1106691431;
assign addr[64203]= -972891995;
assign addr[64204]= -834157373;
assign addr[64205]= -691191324;
assign addr[64206]= -544719071;
assign addr[64207]= -395483624;
assign addr[64208]= -244242007;
assign addr[64209]= -91761426;
assign addr[64210]= 61184634;
assign addr[64211]= 213820322;
assign addr[64212]= 365371365;
assign addr[64213]= 515068990;
assign addr[64214]= 662153826;
assign addr[64215]= 805879757;
assign addr[64216]= 945517704;
assign addr[64217]= 1080359326;
assign addr[64218]= 1209720613;
assign addr[64219]= 1332945355;
assign addr[64220]= 1449408469;
assign addr[64221]= 1558519173;
assign addr[64222]= 1659723983;
assign addr[64223]= 1752509516;
assign addr[64224]= 1836405100;
assign addr[64225]= 1910985158;
assign addr[64226]= 1975871368;
assign addr[64227]= 2030734582;
assign addr[64228]= 2075296495;
assign addr[64229]= 2109331059;
assign addr[64230]= 2132665626;
assign addr[64231]= 2145181827;
assign addr[64232]= 2146816171;
assign addr[64233]= 2137560369;
assign addr[64234]= 2117461370;
assign addr[64235]= 2086621133;
assign addr[64236]= 2045196100;
assign addr[64237]= 1993396407;
assign addr[64238]= 1931484818;
assign addr[64239]= 1859775393;
assign addr[64240]= 1778631892;
assign addr[64241]= 1688465931;
assign addr[64242]= 1589734894;
assign addr[64243]= 1482939614;
assign addr[64244]= 1368621831;
assign addr[64245]= 1247361445;
assign addr[64246]= 1119773573;
assign addr[64247]= 986505429;
assign addr[64248]= 848233042;
assign addr[64249]= 705657826;
assign addr[64250]= 559503022;
assign addr[64251]= 410510029;
assign addr[64252]= 259434643;
assign addr[64253]= 107043224;
assign addr[64254]= -45891193;
assign addr[64255]= -198592817;
assign addr[64256]= -350287041;
assign addr[64257]= -500204365;
assign addr[64258]= -647584304;
assign addr[64259]= -791679244;
assign addr[64260]= -931758235;
assign addr[64261]= -1067110699;
assign addr[64262]= -1197050035;
assign addr[64263]= -1320917099;
assign addr[64264]= -1438083551;
assign addr[64265]= -1547955041;
assign addr[64266]= -1649974225;
assign addr[64267]= -1743623590;
assign addr[64268]= -1828428082;
assign addr[64269]= -1903957513;
assign addr[64270]= -1969828744;
assign addr[64271]= -2025707632;
assign addr[64272]= -2071310720;
assign addr[64273]= -2106406677;
assign addr[64274]= -2130817471;
assign addr[64275]= -2144419275;
assign addr[64276]= -2147143090;
assign addr[64277]= -2138975100;
assign addr[64278]= -2119956737;
assign addr[64279]= -2090184478;
assign addr[64280]= -2049809346;
assign addr[64281]= -1999036154;
assign addr[64282]= -1938122457;
assign addr[64283]= -1867377253;
assign addr[64284]= -1787159411;
assign addr[64285]= -1697875851;
assign addr[64286]= -1599979481;
assign addr[64287]= -1493966902;
assign addr[64288]= -1380375881;
assign addr[64289]= -1259782632;
assign addr[64290]= -1132798888;
assign addr[64291]= -1000068799;
assign addr[64292]= -862265664;
assign addr[64293]= -720088517;
assign addr[64294]= -574258580;
assign addr[64295]= -425515602;
assign addr[64296]= -274614114;
assign addr[64297]= -122319591;
assign addr[64298]= 30595422;
assign addr[64299]= 183355234;
assign addr[64300]= 335184940;
assign addr[64301]= 485314355;
assign addr[64302]= 632981917;
assign addr[64303]= 777438554;
assign addr[64304]= 917951481;
assign addr[64305]= 1053807919;
assign addr[64306]= 1184318708;
assign addr[64307]= 1308821808;
assign addr[64308]= 1426685652;
assign addr[64309]= 1537312353;
assign addr[64310]= 1640140734;
assign addr[64311]= 1734649179;
assign addr[64312]= 1820358275;
assign addr[64313]= 1896833245;
assign addr[64314]= 1963686155;
assign addr[64315]= 2020577882;
assign addr[64316]= 2067219829;
assign addr[64317]= 2103375398;
assign addr[64318]= 2128861181;
assign addr[64319]= 2143547897;
assign addr[64320]= 2147361045;
assign addr[64321]= 2140281282;
assign addr[64322]= 2122344521;
assign addr[64323]= 2093641749;
assign addr[64324]= 2054318569;
assign addr[64325]= 2004574453;
assign addr[64326]= 1944661739;
assign addr[64327]= 1874884346;
assign addr[64328]= 1795596234;
assign addr[64329]= 1707199606;
assign addr[64330]= 1610142873;
assign addr[64331]= 1504918373;
assign addr[64332]= 1392059879;
assign addr[64333]= 1272139887;
assign addr[64334]= 1145766716;
assign addr[64335]= 1013581418;
assign addr[64336]= 876254528;
assign addr[64337]= 734482665;
assign addr[64338]= 588984994;
assign addr[64339]= 440499581;
assign addr[64340]= 289779648;
assign addr[64341]= 137589750;
assign addr[64342]= -15298099;
assign addr[64343]= -168108346;
assign addr[64344]= -320065829;
assign addr[64345]= -470399716;
assign addr[64346]= -618347408;
assign addr[64347]= -763158411;
assign addr[64348]= -904098143;
assign addr[64349]= -1040451659;
assign addr[64350]= -1171527280;
assign addr[64351]= -1296660098;
assign addr[64352]= -1415215352;
assign addr[64353]= -1526591649;
assign addr[64354]= -1630224009;
assign addr[64355]= -1725586737;
assign addr[64356]= -1812196087;
assign addr[64357]= -1889612716;
assign addr[64358]= -1957443913;
assign addr[64359]= -2015345591;
assign addr[64360]= -2063024031;
assign addr[64361]= -2100237377;
assign addr[64362]= -2126796855;
assign addr[64363]= -2142567738;
assign addr[64364]= -2147470025;
assign addr[64365]= -2141478848;
assign addr[64366]= -2124624598;
assign addr[64367]= -2096992772;
assign addr[64368]= -2058723538;
assign addr[64369]= -2010011024;
assign addr[64370]= -1951102334;
assign addr[64371]= -1882296293;
assign addr[64372]= -1803941934;
assign addr[64373]= -1716436725;
assign addr[64374]= -1620224553;
assign addr[64375]= -1515793473;
assign addr[64376]= -1403673233;
assign addr[64377]= -1284432584;
assign addr[64378]= -1158676398;
assign addr[64379]= -1027042599;
assign addr[64380]= -890198924;
assign addr[64381]= -748839539;
assign addr[64382]= -603681519;
assign addr[64383]= -455461206;
assign addr[64384]= -304930476;
assign addr[64385]= -152852926;
assign addr[64386]= 0;
assign addr[64387]= 152852926;
assign addr[64388]= 304930476;
assign addr[64389]= 455461206;
assign addr[64390]= 603681519;
assign addr[64391]= 748839539;
assign addr[64392]= 890198924;
assign addr[64393]= 1027042599;
assign addr[64394]= 1158676398;
assign addr[64395]= 1284432584;
assign addr[64396]= 1403673233;
assign addr[64397]= 1515793473;
assign addr[64398]= 1620224553;
assign addr[64399]= 1716436725;
assign addr[64400]= 1803941934;
assign addr[64401]= 1882296293;
assign addr[64402]= 1951102334;
assign addr[64403]= 2010011024;
assign addr[64404]= 2058723538;
assign addr[64405]= 2096992772;
assign addr[64406]= 2124624598;
assign addr[64407]= 2141478848;
assign addr[64408]= 2147470025;
assign addr[64409]= 2142567738;
assign addr[64410]= 2126796855;
assign addr[64411]= 2100237377;
assign addr[64412]= 2063024031;
assign addr[64413]= 2015345591;
assign addr[64414]= 1957443913;
assign addr[64415]= 1889612716;
assign addr[64416]= 1812196087;
assign addr[64417]= 1725586737;
assign addr[64418]= 1630224009;
assign addr[64419]= 1526591649;
assign addr[64420]= 1415215352;
assign addr[64421]= 1296660098;
assign addr[64422]= 1171527280;
assign addr[64423]= 1040451659;
assign addr[64424]= 904098143;
assign addr[64425]= 763158411;
assign addr[64426]= 618347408;
assign addr[64427]= 470399716;
assign addr[64428]= 320065829;
assign addr[64429]= 168108346;
assign addr[64430]= 15298099;
assign addr[64431]= -137589750;
assign addr[64432]= -289779648;
assign addr[64433]= -440499581;
assign addr[64434]= -588984994;
assign addr[64435]= -734482665;
assign addr[64436]= -876254528;
assign addr[64437]= -1013581418;
assign addr[64438]= -1145766716;
assign addr[64439]= -1272139887;
assign addr[64440]= -1392059879;
assign addr[64441]= -1504918373;
assign addr[64442]= -1610142873;
assign addr[64443]= -1707199606;
assign addr[64444]= -1795596234;
assign addr[64445]= -1874884346;
assign addr[64446]= -1944661739;
assign addr[64447]= -2004574453;
assign addr[64448]= -2054318569;
assign addr[64449]= -2093641749;
assign addr[64450]= -2122344521;
assign addr[64451]= -2140281282;
assign addr[64452]= -2147361045;
assign addr[64453]= -2143547897;
assign addr[64454]= -2128861181;
assign addr[64455]= -2103375398;
assign addr[64456]= -2067219829;
assign addr[64457]= -2020577882;
assign addr[64458]= -1963686155;
assign addr[64459]= -1896833245;
assign addr[64460]= -1820358275;
assign addr[64461]= -1734649179;
assign addr[64462]= -1640140734;
assign addr[64463]= -1537312353;
assign addr[64464]= -1426685652;
assign addr[64465]= -1308821808;
assign addr[64466]= -1184318708;
assign addr[64467]= -1053807919;
assign addr[64468]= -917951481;
assign addr[64469]= -777438554;
assign addr[64470]= -632981917;
assign addr[64471]= -485314355;
assign addr[64472]= -335184940;
assign addr[64473]= -183355234;
assign addr[64474]= -30595422;
assign addr[64475]= 122319591;
assign addr[64476]= 274614114;
assign addr[64477]= 425515602;
assign addr[64478]= 574258580;
assign addr[64479]= 720088517;
assign addr[64480]= 862265664;
assign addr[64481]= 1000068799;
assign addr[64482]= 1132798888;
assign addr[64483]= 1259782632;
assign addr[64484]= 1380375881;
assign addr[64485]= 1493966902;
assign addr[64486]= 1599979481;
assign addr[64487]= 1697875851;
assign addr[64488]= 1787159411;
assign addr[64489]= 1867377253;
assign addr[64490]= 1938122457;
assign addr[64491]= 1999036154;
assign addr[64492]= 2049809346;
assign addr[64493]= 2090184478;
assign addr[64494]= 2119956737;
assign addr[64495]= 2138975100;
assign addr[64496]= 2147143090;
assign addr[64497]= 2144419275;
assign addr[64498]= 2130817471;
assign addr[64499]= 2106406677;
assign addr[64500]= 2071310720;
assign addr[64501]= 2025707632;
assign addr[64502]= 1969828744;
assign addr[64503]= 1903957513;
assign addr[64504]= 1828428082;
assign addr[64505]= 1743623590;
assign addr[64506]= 1649974225;
assign addr[64507]= 1547955041;
assign addr[64508]= 1438083551;
assign addr[64509]= 1320917099;
assign addr[64510]= 1197050035;
assign addr[64511]= 1067110699;
assign addr[64512]= 931758235;
assign addr[64513]= 791679244;
assign addr[64514]= 647584304;
assign addr[64515]= 500204365;
assign addr[64516]= 350287041;
assign addr[64517]= 198592817;
assign addr[64518]= 45891193;
assign addr[64519]= -107043224;
assign addr[64520]= -259434643;
assign addr[64521]= -410510029;
assign addr[64522]= -559503022;
assign addr[64523]= -705657826;
assign addr[64524]= -848233042;
assign addr[64525]= -986505429;
assign addr[64526]= -1119773573;
assign addr[64527]= -1247361445;
assign addr[64528]= -1368621831;
assign addr[64529]= -1482939614;
assign addr[64530]= -1589734894;
assign addr[64531]= -1688465931;
assign addr[64532]= -1778631892;
assign addr[64533]= -1859775393;
assign addr[64534]= -1931484818;
assign addr[64535]= -1993396407;
assign addr[64536]= -2045196100;
assign addr[64537]= -2086621133;
assign addr[64538]= -2117461370;
assign addr[64539]= -2137560369;
assign addr[64540]= -2146816171;
assign addr[64541]= -2145181827;
assign addr[64542]= -2132665626;
assign addr[64543]= -2109331059;
assign addr[64544]= -2075296495;
assign addr[64545]= -2030734582;
assign addr[64546]= -1975871368;
assign addr[64547]= -1910985158;
assign addr[64548]= -1836405100;
assign addr[64549]= -1752509516;
assign addr[64550]= -1659723983;
assign addr[64551]= -1558519173;
assign addr[64552]= -1449408469;
assign addr[64553]= -1332945355;
assign addr[64554]= -1209720613;
assign addr[64555]= -1080359326;
assign addr[64556]= -945517704;
assign addr[64557]= -805879757;
assign addr[64558]= -662153826;
assign addr[64559]= -515068990;
assign addr[64560]= -365371365;
assign addr[64561]= -213820322;
assign addr[64562]= -61184634;
assign addr[64563]= 91761426;
assign addr[64564]= 244242007;
assign addr[64565]= 395483624;
assign addr[64566]= 544719071;
assign addr[64567]= 691191324;
assign addr[64568]= 834157373;
assign addr[64569]= 972891995;
assign addr[64570]= 1106691431;
assign addr[64571]= 1234876957;
assign addr[64572]= 1356798326;
assign addr[64573]= 1471837070;
assign addr[64574]= 1579409630;
assign addr[64575]= 1678970324;
assign addr[64576]= 1770014111;
assign addr[64577]= 1852079154;
assign addr[64578]= 1924749160;
assign addr[64579]= 1987655498;
assign addr[64580]= 2040479063;
assign addr[64581]= 2082951896;
assign addr[64582]= 2114858546;
assign addr[64583]= 2136037160;
assign addr[64584]= 2146380306;
assign addr[64585]= 2145835515;
assign addr[64586]= 2134405552;
assign addr[64587]= 2112148396;
assign addr[64588]= 2079176953;
assign addr[64589]= 2035658475;
assign addr[64590]= 1981813720;
assign addr[64591]= 1917915825;
assign addr[64592]= 1844288924;
assign addr[64593]= 1761306505;
assign addr[64594]= 1669389513;
assign addr[64595]= 1569004214;
assign addr[64596]= 1460659832;
assign addr[64597]= 1344905966;
assign addr[64598]= 1222329801;
assign addr[64599]= 1093553126;
assign addr[64600]= 959229189;
assign addr[64601]= 820039373;
assign addr[64602]= 676689746;
assign addr[64603]= 529907477;
assign addr[64604]= 380437148;
assign addr[64605]= 229036977;
assign addr[64606]= 76474970;
assign addr[64607]= -76474970;
assign addr[64608]= -229036977;
assign addr[64609]= -380437148;
assign addr[64610]= -529907477;
assign addr[64611]= -676689746;
assign addr[64612]= -820039373;
assign addr[64613]= -959229189;
assign addr[64614]= -1093553126;
assign addr[64615]= -1222329801;
assign addr[64616]= -1344905966;
assign addr[64617]= -1460659832;
assign addr[64618]= -1569004214;
assign addr[64619]= -1669389513;
assign addr[64620]= -1761306505;
assign addr[64621]= -1844288924;
assign addr[64622]= -1917915825;
assign addr[64623]= -1981813720;
assign addr[64624]= -2035658475;
assign addr[64625]= -2079176953;
assign addr[64626]= -2112148396;
assign addr[64627]= -2134405552;
assign addr[64628]= -2145835515;
assign addr[64629]= -2146380306;
assign addr[64630]= -2136037160;
assign addr[64631]= -2114858546;
assign addr[64632]= -2082951896;
assign addr[64633]= -2040479063;
assign addr[64634]= -1987655498;
assign addr[64635]= -1924749160;
assign addr[64636]= -1852079154;
assign addr[64637]= -1770014111;
assign addr[64638]= -1678970324;
assign addr[64639]= -1579409630;
assign addr[64640]= -1471837070;
assign addr[64641]= -1356798326;
assign addr[64642]= -1234876957;
assign addr[64643]= -1106691431;
assign addr[64644]= -972891995;
assign addr[64645]= -834157373;
assign addr[64646]= -691191324;
assign addr[64647]= -544719071;
assign addr[64648]= -395483624;
assign addr[64649]= -244242007;
assign addr[64650]= -91761426;
assign addr[64651]= 61184634;
assign addr[64652]= 213820322;
assign addr[64653]= 365371365;
assign addr[64654]= 515068990;
assign addr[64655]= 662153826;
assign addr[64656]= 805879757;
assign addr[64657]= 945517704;
assign addr[64658]= 1080359326;
assign addr[64659]= 1209720613;
assign addr[64660]= 1332945355;
assign addr[64661]= 1449408469;
assign addr[64662]= 1558519173;
assign addr[64663]= 1659723983;
assign addr[64664]= 1752509516;
assign addr[64665]= 1836405100;
assign addr[64666]= 1910985158;
assign addr[64667]= 1975871368;
assign addr[64668]= 2030734582;
assign addr[64669]= 2075296495;
assign addr[64670]= 2109331059;
assign addr[64671]= 2132665626;
assign addr[64672]= 2145181827;
assign addr[64673]= 2146816171;
assign addr[64674]= 2137560369;
assign addr[64675]= 2117461370;
assign addr[64676]= 2086621133;
assign addr[64677]= 2045196100;
assign addr[64678]= 1993396407;
assign addr[64679]= 1931484818;
assign addr[64680]= 1859775393;
assign addr[64681]= 1778631892;
assign addr[64682]= 1688465931;
assign addr[64683]= 1589734894;
assign addr[64684]= 1482939614;
assign addr[64685]= 1368621831;
assign addr[64686]= 1247361445;
assign addr[64687]= 1119773573;
assign addr[64688]= 986505429;
assign addr[64689]= 848233042;
assign addr[64690]= 705657826;
assign addr[64691]= 559503022;
assign addr[64692]= 410510029;
assign addr[64693]= 259434643;
assign addr[64694]= 107043224;
assign addr[64695]= -45891193;
assign addr[64696]= -198592817;
assign addr[64697]= -350287041;
assign addr[64698]= -500204365;
assign addr[64699]= -647584304;
assign addr[64700]= -791679244;
assign addr[64701]= -931758235;
assign addr[64702]= -1067110699;
assign addr[64703]= -1197050035;
assign addr[64704]= -1320917099;
assign addr[64705]= -1438083551;
assign addr[64706]= -1547955041;
assign addr[64707]= -1649974225;
assign addr[64708]= -1743623590;
assign addr[64709]= -1828428082;
assign addr[64710]= -1903957513;
assign addr[64711]= -1969828744;
assign addr[64712]= -2025707632;
assign addr[64713]= -2071310720;
assign addr[64714]= -2106406677;
assign addr[64715]= -2130817471;
assign addr[64716]= -2144419275;
assign addr[64717]= -2147143090;
assign addr[64718]= -2138975100;
assign addr[64719]= -2119956737;
assign addr[64720]= -2090184478;
assign addr[64721]= -2049809346;
assign addr[64722]= -1999036154;
assign addr[64723]= -1938122457;
assign addr[64724]= -1867377253;
assign addr[64725]= -1787159411;
assign addr[64726]= -1697875851;
assign addr[64727]= -1599979481;
assign addr[64728]= -1493966902;
assign addr[64729]= -1380375881;
assign addr[64730]= -1259782632;
assign addr[64731]= -1132798888;
assign addr[64732]= -1000068799;
assign addr[64733]= -862265664;
assign addr[64734]= -720088517;
assign addr[64735]= -574258580;
assign addr[64736]= -425515602;
assign addr[64737]= -274614114;
assign addr[64738]= -122319591;
assign addr[64739]= 30595422;
assign addr[64740]= 183355234;
assign addr[64741]= 335184940;
assign addr[64742]= 485314355;
assign addr[64743]= 632981917;
assign addr[64744]= 777438554;
assign addr[64745]= 917951481;
assign addr[64746]= 1053807919;
assign addr[64747]= 1184318708;
assign addr[64748]= 1308821808;
assign addr[64749]= 1426685652;
assign addr[64750]= 1537312353;
assign addr[64751]= 1640140734;
assign addr[64752]= 1734649179;
assign addr[64753]= 1820358275;
assign addr[64754]= 1896833245;
assign addr[64755]= 1963686155;
assign addr[64756]= 2020577882;
assign addr[64757]= 2067219829;
assign addr[64758]= 2103375398;
assign addr[64759]= 2128861181;
assign addr[64760]= 2143547897;
assign addr[64761]= 2147361045;
assign addr[64762]= 2140281282;
assign addr[64763]= 2122344521;
assign addr[64764]= 2093641749;
assign addr[64765]= 2054318569;
assign addr[64766]= 2004574453;
assign addr[64767]= 1944661739;
assign addr[64768]= 1874884346;
assign addr[64769]= 1795596234;
assign addr[64770]= 1707199606;
assign addr[64771]= 1610142873;
assign addr[64772]= 1504918373;
assign addr[64773]= 1392059879;
assign addr[64774]= 1272139887;
assign addr[64775]= 1145766716;
assign addr[64776]= 1013581418;
assign addr[64777]= 876254528;
assign addr[64778]= 734482665;
assign addr[64779]= 588984994;
assign addr[64780]= 440499581;
assign addr[64781]= 289779648;
assign addr[64782]= 137589750;
assign addr[64783]= -15298099;
assign addr[64784]= -168108346;
assign addr[64785]= -320065829;
assign addr[64786]= -470399716;
assign addr[64787]= -618347408;
assign addr[64788]= -763158411;
assign addr[64789]= -904098143;
assign addr[64790]= -1040451659;
assign addr[64791]= -1171527280;
assign addr[64792]= -1296660098;
assign addr[64793]= -1415215352;
assign addr[64794]= -1526591649;
assign addr[64795]= -1630224009;
assign addr[64796]= -1725586737;
assign addr[64797]= -1812196087;
assign addr[64798]= -1889612716;
assign addr[64799]= -1957443913;
assign addr[64800]= -2015345591;
assign addr[64801]= -2063024031;
assign addr[64802]= -2100237377;
assign addr[64803]= -2126796855;
assign addr[64804]= -2142567738;
assign addr[64805]= -2147470025;
assign addr[64806]= -2141478848;
assign addr[64807]= -2124624598;
assign addr[64808]= -2096992772;
assign addr[64809]= -2058723538;
assign addr[64810]= -2010011024;
assign addr[64811]= -1951102334;
assign addr[64812]= -1882296293;
assign addr[64813]= -1803941934;
assign addr[64814]= -1716436725;
assign addr[64815]= -1620224553;
assign addr[64816]= -1515793473;
assign addr[64817]= -1403673233;
assign addr[64818]= -1284432584;
assign addr[64819]= -1158676398;
assign addr[64820]= -1027042599;
assign addr[64821]= -890198924;
assign addr[64822]= -748839539;
assign addr[64823]= -603681519;
assign addr[64824]= -455461206;
assign addr[64825]= -304930476;
assign addr[64826]= -152852926;
assign addr[64827]= 0;
assign addr[64828]= 152852926;
assign addr[64829]= 304930476;
assign addr[64830]= 455461206;
assign addr[64831]= 603681519;
assign addr[64832]= 748839539;
assign addr[64833]= 890198924;
assign addr[64834]= 1027042599;
assign addr[64835]= 1158676398;
assign addr[64836]= 1284432584;
assign addr[64837]= 1403673233;
assign addr[64838]= 1515793473;
assign addr[64839]= 1620224553;
assign addr[64840]= 1716436725;
assign addr[64841]= 1803941934;
assign addr[64842]= 1882296293;
assign addr[64843]= 1951102334;
assign addr[64844]= 2010011024;
assign addr[64845]= 2058723538;
assign addr[64846]= 2096992772;
assign addr[64847]= 2124624598;
assign addr[64848]= 2141478848;
assign addr[64849]= 2147470025;
assign addr[64850]= 2142567738;
assign addr[64851]= 2126796855;
assign addr[64852]= 2100237377;
assign addr[64853]= 2063024031;
assign addr[64854]= 2015345591;
assign addr[64855]= 1957443913;
assign addr[64856]= 1889612716;
assign addr[64857]= 1812196087;
assign addr[64858]= 1725586737;
assign addr[64859]= 1630224009;
assign addr[64860]= 1526591649;
assign addr[64861]= 1415215352;
assign addr[64862]= 1296660098;
assign addr[64863]= 1171527280;
assign addr[64864]= 1040451659;
assign addr[64865]= 904098143;
assign addr[64866]= 763158411;
assign addr[64867]= 618347408;
assign addr[64868]= 470399716;
assign addr[64869]= 320065829;
assign addr[64870]= 168108346;
assign addr[64871]= 15298099;
assign addr[64872]= -137589750;
assign addr[64873]= -289779648;
assign addr[64874]= -440499581;
assign addr[64875]= -588984994;
assign addr[64876]= -734482665;
assign addr[64877]= -876254528;
assign addr[64878]= -1013581418;
assign addr[64879]= -1145766716;
assign addr[64880]= -1272139887;
assign addr[64881]= -1392059879;
assign addr[64882]= -1504918373;
assign addr[64883]= -1610142873;
assign addr[64884]= -1707199606;
assign addr[64885]= -1795596234;
assign addr[64886]= -1874884346;
assign addr[64887]= -1944661739;
assign addr[64888]= -2004574453;
assign addr[64889]= -2054318569;
assign addr[64890]= -2093641749;
assign addr[64891]= -2122344521;
assign addr[64892]= -2140281282;
assign addr[64893]= -2147361045;
assign addr[64894]= -2143547897;
assign addr[64895]= -2128861181;
assign addr[64896]= -2103375398;
assign addr[64897]= -2067219829;
assign addr[64898]= -2020577882;
assign addr[64899]= -1963686155;
assign addr[64900]= -1896833245;
assign addr[64901]= -1820358275;
assign addr[64902]= -1734649179;
assign addr[64903]= -1640140734;
assign addr[64904]= -1537312353;
assign addr[64905]= -1426685652;
assign addr[64906]= -1308821808;
assign addr[64907]= -1184318708;
assign addr[64908]= -1053807919;
assign addr[64909]= -917951481;
assign addr[64910]= -777438554;
assign addr[64911]= -632981917;
assign addr[64912]= -485314355;
assign addr[64913]= -335184940;
assign addr[64914]= -183355234;
assign addr[64915]= -30595422;
assign addr[64916]= 122319591;
assign addr[64917]= 274614114;
assign addr[64918]= 425515602;
assign addr[64919]= 574258580;
assign addr[64920]= 720088517;
assign addr[64921]= 862265664;
assign addr[64922]= 1000068799;
assign addr[64923]= 1132798888;
assign addr[64924]= 1259782632;
assign addr[64925]= 1380375881;
assign addr[64926]= 1493966902;
assign addr[64927]= 1599979481;
assign addr[64928]= 1697875851;
assign addr[64929]= 1787159411;
assign addr[64930]= 1867377253;
assign addr[64931]= 1938122457;
assign addr[64932]= 1999036154;
assign addr[64933]= 2049809346;
assign addr[64934]= 2090184478;
assign addr[64935]= 2119956737;
assign addr[64936]= 2138975100;
assign addr[64937]= 2147143090;
assign addr[64938]= 2144419275;
assign addr[64939]= 2130817471;
assign addr[64940]= 2106406677;
assign addr[64941]= 2071310720;
assign addr[64942]= 2025707632;
assign addr[64943]= 1969828744;
assign addr[64944]= 1903957513;
assign addr[64945]= 1828428082;
assign addr[64946]= 1743623590;
assign addr[64947]= 1649974225;
assign addr[64948]= 1547955041;
assign addr[64949]= 1438083551;
assign addr[64950]= 1320917099;
assign addr[64951]= 1197050035;
assign addr[64952]= 1067110699;
assign addr[64953]= 931758235;
assign addr[64954]= 791679244;
assign addr[64955]= 647584304;
assign addr[64956]= 500204365;
assign addr[64957]= 350287041;
assign addr[64958]= 198592817;
assign addr[64959]= 45891193;
assign addr[64960]= -107043224;
assign addr[64961]= -259434643;
assign addr[64962]= -410510029;
assign addr[64963]= -559503022;
assign addr[64964]= -705657826;
assign addr[64965]= -848233042;
assign addr[64966]= -986505429;
assign addr[64967]= -1119773573;
assign addr[64968]= -1247361445;
assign addr[64969]= -1368621831;
assign addr[64970]= -1482939614;
assign addr[64971]= -1589734894;
assign addr[64972]= -1688465931;
assign addr[64973]= -1778631892;
assign addr[64974]= -1859775393;
assign addr[64975]= -1931484818;
assign addr[64976]= -1993396407;
assign addr[64977]= -2045196100;
assign addr[64978]= -2086621133;
assign addr[64979]= -2117461370;
assign addr[64980]= -2137560369;
assign addr[64981]= -2146816171;
assign addr[64982]= -2145181827;
assign addr[64983]= -2132665626;
assign addr[64984]= -2109331059;
assign addr[64985]= -2075296495;
assign addr[64986]= -2030734582;
assign addr[64987]= -1975871368;
assign addr[64988]= -1910985158;
assign addr[64989]= -1836405100;
assign addr[64990]= -1752509516;
assign addr[64991]= -1659723983;
assign addr[64992]= -1558519173;
assign addr[64993]= -1449408469;
assign addr[64994]= -1332945355;
assign addr[64995]= -1209720613;
assign addr[64996]= -1080359326;
assign addr[64997]= -945517704;
assign addr[64998]= -805879757;
assign addr[64999]= -662153826;
assign addr[65000]= -515068990;
assign addr[65001]= -365371365;
assign addr[65002]= -213820322;
assign addr[65003]= -61184634;
assign addr[65004]= 91761426;
assign addr[65005]= 244242007;
assign addr[65006]= 395483624;
assign addr[65007]= 544719071;
assign addr[65008]= 691191324;
assign addr[65009]= 834157373;
assign addr[65010]= 972891995;
assign addr[65011]= 1106691431;
assign addr[65012]= 1234876957;
assign addr[65013]= 1356798326;
assign addr[65014]= 1471837070;
assign addr[65015]= 1579409630;
assign addr[65016]= 1678970324;
assign addr[65017]= 1770014111;
assign addr[65018]= 1852079154;
assign addr[65019]= 1924749160;
assign addr[65020]= 1987655498;
assign addr[65021]= 2040479063;
assign addr[65022]= 2082951896;
assign addr[65023]= 2114858546;
assign addr[65024]= 2136037160;
assign addr[65025]= 2146380306;
assign addr[65026]= 2145835515;
assign addr[65027]= 2134405552;
assign addr[65028]= 2112148396;
assign addr[65029]= 2079176953;
assign addr[65030]= 2035658475;
assign addr[65031]= 1981813720;
assign addr[65032]= 1917915825;
assign addr[65033]= 1844288924;
assign addr[65034]= 1761306505;
assign addr[65035]= 1669389513;
assign addr[65036]= 1569004214;
assign addr[65037]= 1460659832;
assign addr[65038]= 1344905966;
assign addr[65039]= 1222329801;
assign addr[65040]= 1093553126;
assign addr[65041]= 959229189;
assign addr[65042]= 820039373;
assign addr[65043]= 676689746;
assign addr[65044]= 529907477;
assign addr[65045]= 380437148;
assign addr[65046]= 229036977;
assign addr[65047]= 76474970;
assign addr[65048]= -76474970;
assign addr[65049]= -229036977;
assign addr[65050]= -380437148;
assign addr[65051]= -529907477;
assign addr[65052]= -676689746;
assign addr[65053]= -820039373;
assign addr[65054]= -959229189;
assign addr[65055]= -1093553126;
assign addr[65056]= -1222329801;
assign addr[65057]= -1344905966;
assign addr[65058]= -1460659832;
assign addr[65059]= -1569004214;
assign addr[65060]= -1669389513;
assign addr[65061]= -1761306505;
assign addr[65062]= -1844288924;
assign addr[65063]= -1917915825;
assign addr[65064]= -1981813720;
assign addr[65065]= -2035658475;
assign addr[65066]= -2079176953;
assign addr[65067]= -2112148396;
assign addr[65068]= -2134405552;
assign addr[65069]= -2145835515;
assign addr[65070]= -2146380306;
assign addr[65071]= -2136037160;
assign addr[65072]= -2114858546;
assign addr[65073]= -2082951896;
assign addr[65074]= -2040479063;
assign addr[65075]= -1987655498;
assign addr[65076]= -1924749160;
assign addr[65077]= -1852079154;
assign addr[65078]= -1770014111;
assign addr[65079]= -1678970324;
assign addr[65080]= -1579409630;
assign addr[65081]= -1471837070;
assign addr[65082]= -1356798326;
assign addr[65083]= -1234876957;
assign addr[65084]= -1106691431;
assign addr[65085]= -972891995;
assign addr[65086]= -834157373;
assign addr[65087]= -691191324;
assign addr[65088]= -544719071;
assign addr[65089]= -395483624;
assign addr[65090]= -244242007;
assign addr[65091]= -91761426;
assign addr[65092]= 61184634;
assign addr[65093]= 213820322;
assign addr[65094]= 365371365;
assign addr[65095]= 515068990;
assign addr[65096]= 662153826;
assign addr[65097]= 805879757;
assign addr[65098]= 945517704;
assign addr[65099]= 1080359326;
assign addr[65100]= 1209720613;
assign addr[65101]= 1332945355;
assign addr[65102]= 1449408469;
assign addr[65103]= 1558519173;
assign addr[65104]= 1659723983;
assign addr[65105]= 1752509516;
assign addr[65106]= 1836405100;
assign addr[65107]= 1910985158;
assign addr[65108]= 1975871368;
assign addr[65109]= 2030734582;
assign addr[65110]= 2075296495;
assign addr[65111]= 2109331059;
assign addr[65112]= 2132665626;
assign addr[65113]= 2145181827;
assign addr[65114]= 2146816171;
assign addr[65115]= 2137560369;
assign addr[65116]= 2117461370;
assign addr[65117]= 2086621133;
assign addr[65118]= 2045196100;
assign addr[65119]= 1993396407;
assign addr[65120]= 1931484818;
assign addr[65121]= 1859775393;
assign addr[65122]= 1778631892;
assign addr[65123]= 1688465931;
assign addr[65124]= 1589734894;
assign addr[65125]= 1482939614;
assign addr[65126]= 1368621831;
assign addr[65127]= 1247361445;
assign addr[65128]= 1119773573;
assign addr[65129]= 986505429;
assign addr[65130]= 848233042;
assign addr[65131]= 705657826;
assign addr[65132]= 559503022;
assign addr[65133]= 410510029;
assign addr[65134]= 259434643;
assign addr[65135]= 107043224;
assign addr[65136]= -45891193;
assign addr[65137]= -198592817;
assign addr[65138]= -350287041;
assign addr[65139]= -500204365;
assign addr[65140]= -647584304;
assign addr[65141]= -791679244;
assign addr[65142]= -931758235;
assign addr[65143]= -1067110699;
assign addr[65144]= -1197050035;
assign addr[65145]= -1320917099;
assign addr[65146]= -1438083551;
assign addr[65147]= -1547955041;
assign addr[65148]= -1649974225;
assign addr[65149]= -1743623590;
assign addr[65150]= -1828428082;
assign addr[65151]= -1903957513;
assign addr[65152]= -1969828744;
assign addr[65153]= -2025707632;
assign addr[65154]= -2071310720;
assign addr[65155]= -2106406677;
assign addr[65156]= -2130817471;
assign addr[65157]= -2144419275;
assign addr[65158]= -2147143090;
assign addr[65159]= -2138975100;
assign addr[65160]= -2119956737;
assign addr[65161]= -2090184478;
assign addr[65162]= -2049809346;
assign addr[65163]= -1999036154;
assign addr[65164]= -1938122457;
assign addr[65165]= -1867377253;
assign addr[65166]= -1787159411;
assign addr[65167]= -1697875851;
assign addr[65168]= -1599979481;
assign addr[65169]= -1493966902;
assign addr[65170]= -1380375881;
assign addr[65171]= -1259782632;
assign addr[65172]= -1132798888;
assign addr[65173]= -1000068799;
assign addr[65174]= -862265664;
assign addr[65175]= -720088517;
assign addr[65176]= -574258580;
assign addr[65177]= -425515602;
assign addr[65178]= -274614114;
assign addr[65179]= -122319591;
assign addr[65180]= 30595422;
assign addr[65181]= 183355234;
assign addr[65182]= 335184940;
assign addr[65183]= 485314355;
assign addr[65184]= 632981917;
assign addr[65185]= 777438554;
assign addr[65186]= 917951481;
assign addr[65187]= 1053807919;
assign addr[65188]= 1184318708;
assign addr[65189]= 1308821808;
assign addr[65190]= 1426685652;
assign addr[65191]= 1537312353;
assign addr[65192]= 1640140734;
assign addr[65193]= 1734649179;
assign addr[65194]= 1820358275;
assign addr[65195]= 1896833245;
assign addr[65196]= 1963686155;
assign addr[65197]= 2020577882;
assign addr[65198]= 2067219829;
assign addr[65199]= 2103375398;
assign addr[65200]= 2128861181;
assign addr[65201]= 2143547897;
assign addr[65202]= 2147361045;
assign addr[65203]= 2140281282;
assign addr[65204]= 2122344521;
assign addr[65205]= 2093641749;
assign addr[65206]= 2054318569;
assign addr[65207]= 2004574453;
assign addr[65208]= 1944661739;
assign addr[65209]= 1874884346;
assign addr[65210]= 1795596234;
assign addr[65211]= 1707199606;
assign addr[65212]= 1610142873;
assign addr[65213]= 1504918373;
assign addr[65214]= 1392059879;
assign addr[65215]= 1272139887;
assign addr[65216]= 1145766716;
assign addr[65217]= 1013581418;
assign addr[65218]= 876254528;
assign addr[65219]= 734482665;
assign addr[65220]= 588984994;
assign addr[65221]= 440499581;
assign addr[65222]= 289779648;
assign addr[65223]= 137589750;
assign addr[65224]= -15298099;
assign addr[65225]= -168108346;
assign addr[65226]= -320065829;
assign addr[65227]= -470399716;
assign addr[65228]= -618347408;
assign addr[65229]= -763158411;
assign addr[65230]= -904098143;
assign addr[65231]= -1040451659;
assign addr[65232]= -1171527280;
assign addr[65233]= -1296660098;
assign addr[65234]= -1415215352;
assign addr[65235]= -1526591649;
assign addr[65236]= -1630224009;
assign addr[65237]= -1725586737;
assign addr[65238]= -1812196087;
assign addr[65239]= -1889612716;
assign addr[65240]= -1957443913;
assign addr[65241]= -2015345591;
assign addr[65242]= -2063024031;
assign addr[65243]= -2100237377;
assign addr[65244]= -2126796855;
assign addr[65245]= -2142567738;
assign addr[65246]= -2147470025;
assign addr[65247]= -2141478848;
assign addr[65248]= -2124624598;
assign addr[65249]= -2096992772;
assign addr[65250]= -2058723538;
assign addr[65251]= -2010011024;
assign addr[65252]= -1951102334;
assign addr[65253]= -1882296293;
assign addr[65254]= -1803941934;
assign addr[65255]= -1716436725;
assign addr[65256]= -1620224553;
assign addr[65257]= -1515793473;
assign addr[65258]= -1403673233;
assign addr[65259]= -1284432584;
assign addr[65260]= -1158676398;
assign addr[65261]= -1027042599;
assign addr[65262]= -890198924;
assign addr[65263]= -748839539;
assign addr[65264]= -603681519;
assign addr[65265]= -455461206;
assign addr[65266]= -304930476;
assign addr[65267]= -152852926;
assign addr[65268]= 0;
assign addr[65269]= 152852926;
assign addr[65270]= 304930476;
assign addr[65271]= 455461206;
assign addr[65272]= 603681519;
assign addr[65273]= 748839539;
assign addr[65274]= 890198924;
assign addr[65275]= 1027042599;
assign addr[65276]= 1158676398;
assign addr[65277]= 1284432584;
assign addr[65278]= 1403673233;
assign addr[65279]= 1515793473;
assign addr[65280]= 1620224553;
assign addr[65281]= 1716436725;
assign addr[65282]= 1803941934;
assign addr[65283]= 1882296293;
assign addr[65284]= 1951102334;
assign addr[65285]= 2010011024;
assign addr[65286]= 2058723538;
assign addr[65287]= 2096992772;
assign addr[65288]= 2124624598;
assign addr[65289]= 2141478848;
assign addr[65290]= 2147470025;
assign addr[65291]= 2142567738;
assign addr[65292]= 2126796855;
assign addr[65293]= 2100237377;
assign addr[65294]= 2063024031;
assign addr[65295]= 2015345591;
assign addr[65296]= 1957443913;
assign addr[65297]= 1889612716;
assign addr[65298]= 1812196087;
assign addr[65299]= 1725586737;
assign addr[65300]= 1630224009;
assign addr[65301]= 1526591649;
assign addr[65302]= 1415215352;
assign addr[65303]= 1296660098;
assign addr[65304]= 1171527280;
assign addr[65305]= 1040451659;
assign addr[65306]= 904098143;
assign addr[65307]= 763158411;
assign addr[65308]= 618347408;
assign addr[65309]= 470399716;
assign addr[65310]= 320065829;
assign addr[65311]= 168108346;
assign addr[65312]= 15298099;
assign addr[65313]= -137589750;
assign addr[65314]= -289779648;
assign addr[65315]= -440499581;
assign addr[65316]= -588984994;
assign addr[65317]= -734482665;
assign addr[65318]= -876254528;
assign addr[65319]= -1013581418;
assign addr[65320]= -1145766716;
assign addr[65321]= -1272139887;
assign addr[65322]= -1392059879;
assign addr[65323]= -1504918373;
assign addr[65324]= -1610142873;
assign addr[65325]= -1707199606;
assign addr[65326]= -1795596234;
assign addr[65327]= -1874884346;
assign addr[65328]= -1944661739;
assign addr[65329]= -2004574453;
assign addr[65330]= -2054318569;
assign addr[65331]= -2093641749;
assign addr[65332]= -2122344521;
assign addr[65333]= -2140281282;
assign addr[65334]= -2147361045;
assign addr[65335]= -2143547897;
assign addr[65336]= -2128861181;
assign addr[65337]= -2103375398;
assign addr[65338]= -2067219829;
assign addr[65339]= -2020577882;
assign addr[65340]= -1963686155;
assign addr[65341]= -1896833245;
assign addr[65342]= -1820358275;
assign addr[65343]= -1734649179;
assign addr[65344]= -1640140734;
assign addr[65345]= -1537312353;
assign addr[65346]= -1426685652;
assign addr[65347]= -1308821808;
assign addr[65348]= -1184318708;
assign addr[65349]= -1053807919;
assign addr[65350]= -917951481;
assign addr[65351]= -777438554;
assign addr[65352]= -632981917;
assign addr[65353]= -485314355;
assign addr[65354]= -335184940;
assign addr[65355]= -183355234;
assign addr[65356]= -30595422;
assign addr[65357]= 122319591;
assign addr[65358]= 274614114;
assign addr[65359]= 425515602;
assign addr[65360]= 574258580;
assign addr[65361]= 720088517;
assign addr[65362]= 862265664;
assign addr[65363]= 1000068799;
assign addr[65364]= 1132798888;
assign addr[65365]= 1259782632;
assign addr[65366]= 1380375881;
assign addr[65367]= 1493966902;
assign addr[65368]= 1599979481;
assign addr[65369]= 1697875851;
assign addr[65370]= 1787159411;
assign addr[65371]= 1867377253;
assign addr[65372]= 1938122457;
assign addr[65373]= 1999036154;
assign addr[65374]= 2049809346;
assign addr[65375]= 2090184478;
assign addr[65376]= 2119956737;
assign addr[65377]= 2138975100;
assign addr[65378]= 2147143090;
assign addr[65379]= 2144419275;
assign addr[65380]= 2130817471;
assign addr[65381]= 2106406677;
assign addr[65382]= 2071310720;
assign addr[65383]= 2025707632;
assign addr[65384]= 1969828744;
assign addr[65385]= 1903957513;
assign addr[65386]= 1828428082;
assign addr[65387]= 1743623590;
assign addr[65388]= 1649974225;
assign addr[65389]= 1547955041;
assign addr[65390]= 1438083551;
assign addr[65391]= 1320917099;
assign addr[65392]= 1197050035;
assign addr[65393]= 1067110699;
assign addr[65394]= 931758235;
assign addr[65395]= 791679244;
assign addr[65396]= 647584304;
assign addr[65397]= 500204365;
assign addr[65398]= 350287041;
assign addr[65399]= 198592817;
assign addr[65400]= 45891193;
assign addr[65401]= -107043224;
assign addr[65402]= -259434643;
assign addr[65403]= -410510029;
assign addr[65404]= -559503022;
assign addr[65405]= -705657826;
assign addr[65406]= -848233042;
assign addr[65407]= -986505429;
assign addr[65408]= -1119773573;
assign addr[65409]= -1247361445;
assign addr[65410]= -1368621831;
assign addr[65411]= -1482939614;
assign addr[65412]= -1589734894;
assign addr[65413]= -1688465931;
assign addr[65414]= -1778631892;
assign addr[65415]= -1859775393;
assign addr[65416]= -1931484818;
assign addr[65417]= -1993396407;
assign addr[65418]= -2045196100;
assign addr[65419]= -2086621133;
assign addr[65420]= -2117461370;
assign addr[65421]= -2137560369;
assign addr[65422]= -2146816171;
assign addr[65423]= -2145181827;
assign addr[65424]= -2132665626;
assign addr[65425]= -2109331059;
assign addr[65426]= -2075296495;
assign addr[65427]= -2030734582;
assign addr[65428]= -1975871368;
assign addr[65429]= -1910985158;
assign addr[65430]= -1836405100;
assign addr[65431]= -1752509516;
assign addr[65432]= -1659723983;
assign addr[65433]= -1558519173;
assign addr[65434]= -1449408469;
assign addr[65435]= -1332945355;
assign addr[65436]= -1209720613;
assign addr[65437]= -1080359326;
assign addr[65438]= -945517704;
assign addr[65439]= -805879757;
assign addr[65440]= -662153826;
assign addr[65441]= -515068990;
assign addr[65442]= -365371365;
assign addr[65443]= -213820322;
assign addr[65444]= -61184634;
assign addr[65445]= 91761426;
assign addr[65446]= 244242007;
assign addr[65447]= 395483624;
assign addr[65448]= 544719071;
assign addr[65449]= 691191324;
assign addr[65450]= 834157373;
assign addr[65451]= 972891995;
assign addr[65452]= 1106691431;
assign addr[65453]= 1234876957;
assign addr[65454]= 1356798326;
assign addr[65455]= 1471837070;
assign addr[65456]= 1579409630;
assign addr[65457]= 1678970324;
assign addr[65458]= 1770014111;
assign addr[65459]= 1852079154;
assign addr[65460]= 1924749160;
assign addr[65461]= 1987655498;
assign addr[65462]= 2040479063;
assign addr[65463]= 2082951896;
assign addr[65464]= 2114858546;
assign addr[65465]= 2136037160;
assign addr[65466]= 2146380306;
assign addr[65467]= 2145835515;
assign addr[65468]= 2134405552;
assign addr[65469]= 2112148396;
assign addr[65470]= 2079176953;
assign addr[65471]= 2035658475;
assign addr[65472]= 1981813720;
assign addr[65473]= 1917915825;
assign addr[65474]= 1844288924;
assign addr[65475]= 1761306505;
assign addr[65476]= 1669389513;
assign addr[65477]= 1569004214;
assign addr[65478]= 1460659832;
assign addr[65479]= 1344905966;
assign addr[65480]= 1222329801;
assign addr[65481]= 1093553126;
assign addr[65482]= 959229189;
assign addr[65483]= 820039373;
assign addr[65484]= 676689746;
assign addr[65485]= 529907477;
assign addr[65486]= 380437148;
assign addr[65487]= 229036977;
assign addr[65488]= 76474970;
assign addr[65489]= -76474970;
assign addr[65490]= -229036977;
assign addr[65491]= -380437148;
assign addr[65492]= -529907477;
assign addr[65493]= -676689746;
assign addr[65494]= -820039373;
assign addr[65495]= -959229189;
assign addr[65496]= -1093553126;
assign addr[65497]= -1222329801;
assign addr[65498]= -1344905966;
assign addr[65499]= -1460659832;
assign addr[65500]= -1569004214;
assign addr[65501]= -1669389513;
assign addr[65502]= -1761306505;
assign addr[65503]= -1844288924;
assign addr[65504]= -1917915825;
assign addr[65505]= -1981813720;
assign addr[65506]= -2035658475;
assign addr[65507]= -2079176953;
assign addr[65508]= -2112148396;
assign addr[65509]= -2134405552;
assign addr[65510]= -2145835515;
assign addr[65511]= -2146380306;
assign addr[65512]= -2136037160;
assign addr[65513]= -2114858546;
assign addr[65514]= -2082951896;
assign addr[65515]= -2040479063;
assign addr[65516]= -1987655498;
assign addr[65517]= -1924749160;
assign addr[65518]= -1852079154;
assign addr[65519]= -1770014111;
assign addr[65520]= -1678970324;
assign addr[65521]= -1579409630;
assign addr[65522]= -1471837070;
assign addr[65523]= -1356798326;
assign addr[65524]= -1234876957;
assign addr[65525]= -1106691431;
assign addr[65526]= -972891995;
assign addr[65527]= -834157373;
assign addr[65528]= -691191324;
assign addr[65529]= -544719071;
assign addr[65530]= -395483624;
assign addr[65531]= -244242007;
assign addr[65532]= -91761426;
assign addr[65533]= 61184634;
assign addr[65534]= 213820322;
assign addr[65535]= 365371365;
endmodule